
module FIFOTop ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, ClkW, Reseter
 );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(n195), .WriteReq(n194), .ClkR(ClkR), .ClkW(ClkW), .Reset(n193) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({n228, n227, n226, 
        n225, n224, n223, n222, n221, n220, n219, n218, n217, n216, n215, n214, 
        n213, n212, n211, n210, n209, n208, n207, n206, n205, n204, n203, n202, 
        n201, n200, n199, n198, n197}), .AddrR(SM_ReadAddr), .AddrW(
        SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), .ChipEna(1'b1), .Read(n196), 
        .Write(SM_MemWriteCmd), .Reset(n193) );
  CKBXD0 U2 ( .I(Reseter), .Z(n193) );
  DEL2 U3 ( .I(n6), .Z(n228) );
  DEL4 U4 ( .I(Din[31]), .Z(n1) );
  DEL4 U5 ( .I(n1), .Z(n2) );
  DEL4 U6 ( .I(n2), .Z(n3) );
  DEL4 U7 ( .I(n3), .Z(n4) );
  DEL4 U8 ( .I(n4), .Z(n5) );
  DEL4 U9 ( .I(n5), .Z(n6) );
  DEL2 U10 ( .I(n12), .Z(n227) );
  DEL4 U11 ( .I(Din[30]), .Z(n7) );
  DEL4 U12 ( .I(n7), .Z(n8) );
  DEL4 U13 ( .I(n8), .Z(n9) );
  DEL4 U14 ( .I(n9), .Z(n10) );
  DEL4 U15 ( .I(n10), .Z(n11) );
  DEL4 U16 ( .I(n11), .Z(n12) );
  DEL2 U17 ( .I(n18), .Z(n226) );
  DEL4 U18 ( .I(Din[29]), .Z(n13) );
  DEL4 U19 ( .I(n13), .Z(n14) );
  DEL4 U20 ( .I(n14), .Z(n15) );
  DEL4 U21 ( .I(n15), .Z(n16) );
  DEL4 U22 ( .I(n16), .Z(n17) );
  DEL4 U23 ( .I(n17), .Z(n18) );
  DEL2 U24 ( .I(n24), .Z(n225) );
  DEL4 U25 ( .I(Din[28]), .Z(n19) );
  DEL4 U26 ( .I(n19), .Z(n20) );
  DEL4 U27 ( .I(n20), .Z(n21) );
  DEL4 U28 ( .I(n21), .Z(n22) );
  DEL4 U29 ( .I(n22), .Z(n23) );
  DEL4 U30 ( .I(n23), .Z(n24) );
  DEL2 U31 ( .I(n30), .Z(n224) );
  DEL4 U32 ( .I(Din[27]), .Z(n25) );
  DEL4 U33 ( .I(n25), .Z(n26) );
  DEL4 U34 ( .I(n26), .Z(n27) );
  DEL4 U35 ( .I(n27), .Z(n28) );
  DEL4 U36 ( .I(n28), .Z(n29) );
  DEL4 U37 ( .I(n29), .Z(n30) );
  DEL2 U38 ( .I(n36), .Z(n223) );
  DEL4 U39 ( .I(Din[26]), .Z(n31) );
  DEL4 U40 ( .I(n31), .Z(n32) );
  DEL4 U41 ( .I(n32), .Z(n33) );
  DEL4 U42 ( .I(n33), .Z(n34) );
  DEL4 U43 ( .I(n34), .Z(n35) );
  DEL4 U44 ( .I(n35), .Z(n36) );
  DEL2 U45 ( .I(n42), .Z(n222) );
  DEL4 U46 ( .I(Din[25]), .Z(n37) );
  DEL4 U47 ( .I(n37), .Z(n38) );
  DEL4 U48 ( .I(n38), .Z(n39) );
  DEL4 U49 ( .I(n39), .Z(n40) );
  DEL4 U50 ( .I(n40), .Z(n41) );
  DEL4 U51 ( .I(n41), .Z(n42) );
  DEL2 U52 ( .I(n48), .Z(n221) );
  DEL4 U53 ( .I(Din[24]), .Z(n43) );
  DEL4 U54 ( .I(n43), .Z(n44) );
  DEL4 U55 ( .I(n44), .Z(n45) );
  DEL4 U56 ( .I(n45), .Z(n46) );
  DEL4 U57 ( .I(n46), .Z(n47) );
  DEL4 U58 ( .I(n47), .Z(n48) );
  DEL2 U59 ( .I(n54), .Z(n220) );
  DEL4 U60 ( .I(Din[23]), .Z(n49) );
  DEL4 U61 ( .I(n49), .Z(n50) );
  DEL4 U62 ( .I(n50), .Z(n51) );
  DEL4 U63 ( .I(n51), .Z(n52) );
  DEL4 U64 ( .I(n52), .Z(n53) );
  DEL4 U65 ( .I(n53), .Z(n54) );
  DEL2 U66 ( .I(n60), .Z(n219) );
  DEL4 U67 ( .I(Din[22]), .Z(n55) );
  DEL4 U68 ( .I(n55), .Z(n56) );
  DEL4 U69 ( .I(n56), .Z(n57) );
  DEL4 U70 ( .I(n57), .Z(n58) );
  DEL4 U71 ( .I(n58), .Z(n59) );
  DEL4 U72 ( .I(n59), .Z(n60) );
  DEL2 U73 ( .I(n66), .Z(n218) );
  DEL4 U74 ( .I(Din[21]), .Z(n61) );
  DEL4 U75 ( .I(n61), .Z(n62) );
  DEL4 U76 ( .I(n62), .Z(n63) );
  DEL4 U77 ( .I(n63), .Z(n64) );
  DEL4 U78 ( .I(n64), .Z(n65) );
  DEL4 U79 ( .I(n65), .Z(n66) );
  DEL2 U80 ( .I(n72), .Z(n217) );
  DEL4 U81 ( .I(Din[20]), .Z(n67) );
  DEL4 U82 ( .I(n67), .Z(n68) );
  DEL4 U83 ( .I(n68), .Z(n69) );
  DEL4 U84 ( .I(n69), .Z(n70) );
  DEL4 U85 ( .I(n70), .Z(n71) );
  DEL4 U86 ( .I(n71), .Z(n72) );
  DEL2 U87 ( .I(n78), .Z(n216) );
  DEL4 U88 ( .I(Din[19]), .Z(n73) );
  DEL4 U89 ( .I(n73), .Z(n74) );
  DEL4 U90 ( .I(n74), .Z(n75) );
  DEL4 U91 ( .I(n75), .Z(n76) );
  DEL4 U92 ( .I(n76), .Z(n77) );
  DEL4 U93 ( .I(n77), .Z(n78) );
  DEL2 U94 ( .I(n84), .Z(n215) );
  DEL4 U95 ( .I(Din[18]), .Z(n79) );
  DEL4 U96 ( .I(n79), .Z(n80) );
  DEL4 U97 ( .I(n80), .Z(n81) );
  DEL4 U98 ( .I(n81), .Z(n82) );
  DEL4 U99 ( .I(n82), .Z(n83) );
  DEL4 U100 ( .I(n83), .Z(n84) );
  DEL2 U101 ( .I(n90), .Z(n214) );
  DEL4 U102 ( .I(Din[17]), .Z(n85) );
  DEL4 U103 ( .I(n85), .Z(n86) );
  DEL4 U104 ( .I(n86), .Z(n87) );
  DEL4 U105 ( .I(n87), .Z(n88) );
  DEL4 U106 ( .I(n88), .Z(n89) );
  DEL4 U107 ( .I(n89), .Z(n90) );
  DEL2 U108 ( .I(n96), .Z(n213) );
  DEL4 U109 ( .I(Din[16]), .Z(n91) );
  DEL4 U110 ( .I(n91), .Z(n92) );
  DEL4 U111 ( .I(n92), .Z(n93) );
  DEL4 U112 ( .I(n93), .Z(n94) );
  DEL4 U113 ( .I(n94), .Z(n95) );
  DEL4 U114 ( .I(n95), .Z(n96) );
  DEL2 U115 ( .I(n102), .Z(n212) );
  DEL4 U116 ( .I(Din[15]), .Z(n97) );
  DEL4 U117 ( .I(n97), .Z(n98) );
  DEL4 U118 ( .I(n98), .Z(n99) );
  DEL4 U119 ( .I(n99), .Z(n100) );
  DEL4 U120 ( .I(n100), .Z(n101) );
  DEL4 U121 ( .I(n101), .Z(n102) );
  DEL2 U122 ( .I(n108), .Z(n211) );
  DEL4 U123 ( .I(Din[14]), .Z(n103) );
  DEL4 U124 ( .I(n103), .Z(n104) );
  DEL4 U125 ( .I(n104), .Z(n105) );
  DEL4 U126 ( .I(n105), .Z(n106) );
  DEL4 U127 ( .I(n106), .Z(n107) );
  DEL4 U128 ( .I(n107), .Z(n108) );
  DEL2 U129 ( .I(n114), .Z(n210) );
  DEL4 U130 ( .I(Din[13]), .Z(n109) );
  DEL4 U131 ( .I(n109), .Z(n110) );
  DEL4 U132 ( .I(n110), .Z(n111) );
  DEL4 U133 ( .I(n111), .Z(n112) );
  DEL4 U134 ( .I(n112), .Z(n113) );
  DEL4 U135 ( .I(n113), .Z(n114) );
  DEL2 U136 ( .I(n120), .Z(n209) );
  DEL4 U137 ( .I(Din[12]), .Z(n115) );
  DEL4 U138 ( .I(n115), .Z(n116) );
  DEL4 U139 ( .I(n116), .Z(n117) );
  DEL4 U140 ( .I(n117), .Z(n118) );
  DEL4 U141 ( .I(n118), .Z(n119) );
  DEL4 U142 ( .I(n119), .Z(n120) );
  DEL2 U143 ( .I(n126), .Z(n208) );
  DEL4 U144 ( .I(Din[11]), .Z(n121) );
  DEL4 U145 ( .I(n121), .Z(n122) );
  DEL4 U146 ( .I(n122), .Z(n123) );
  DEL4 U147 ( .I(n123), .Z(n124) );
  DEL4 U148 ( .I(n124), .Z(n125) );
  DEL4 U149 ( .I(n125), .Z(n126) );
  DEL2 U150 ( .I(n132), .Z(n207) );
  DEL4 U151 ( .I(Din[10]), .Z(n127) );
  DEL4 U152 ( .I(n127), .Z(n128) );
  DEL4 U153 ( .I(n128), .Z(n129) );
  DEL4 U154 ( .I(n129), .Z(n130) );
  DEL4 U155 ( .I(n130), .Z(n131) );
  DEL4 U156 ( .I(n131), .Z(n132) );
  DEL2 U157 ( .I(n138), .Z(n206) );
  DEL4 U158 ( .I(Din[9]), .Z(n133) );
  DEL4 U159 ( .I(n133), .Z(n134) );
  DEL4 U160 ( .I(n134), .Z(n135) );
  DEL4 U161 ( .I(n135), .Z(n136) );
  DEL4 U162 ( .I(n136), .Z(n137) );
  DEL4 U163 ( .I(n137), .Z(n138) );
  DEL2 U164 ( .I(n144), .Z(n205) );
  DEL4 U165 ( .I(Din[8]), .Z(n139) );
  DEL4 U166 ( .I(n139), .Z(n140) );
  DEL4 U167 ( .I(n140), .Z(n141) );
  DEL4 U168 ( .I(n141), .Z(n142) );
  DEL4 U169 ( .I(n142), .Z(n143) );
  DEL4 U170 ( .I(n143), .Z(n144) );
  DEL2 U171 ( .I(n150), .Z(n204) );
  DEL4 U172 ( .I(Din[7]), .Z(n145) );
  DEL4 U173 ( .I(n145), .Z(n146) );
  DEL4 U174 ( .I(n146), .Z(n147) );
  DEL4 U175 ( .I(n147), .Z(n148) );
  DEL4 U176 ( .I(n148), .Z(n149) );
  DEL4 U177 ( .I(n149), .Z(n150) );
  DEL2 U178 ( .I(n156), .Z(n203) );
  DEL4 U179 ( .I(Din[6]), .Z(n151) );
  DEL4 U180 ( .I(n151), .Z(n152) );
  DEL4 U181 ( .I(n152), .Z(n153) );
  DEL4 U182 ( .I(n153), .Z(n154) );
  DEL4 U183 ( .I(n154), .Z(n155) );
  DEL4 U184 ( .I(n155), .Z(n156) );
  DEL2 U185 ( .I(n162), .Z(n202) );
  DEL4 U186 ( .I(Din[5]), .Z(n157) );
  DEL4 U187 ( .I(n157), .Z(n158) );
  DEL4 U188 ( .I(n158), .Z(n159) );
  DEL4 U189 ( .I(n159), .Z(n160) );
  DEL4 U190 ( .I(n160), .Z(n161) );
  DEL4 U191 ( .I(n161), .Z(n162) );
  DEL2 U192 ( .I(n168), .Z(n201) );
  DEL4 U193 ( .I(Din[4]), .Z(n163) );
  DEL4 U194 ( .I(n163), .Z(n164) );
  DEL4 U195 ( .I(n164), .Z(n165) );
  DEL4 U196 ( .I(n165), .Z(n166) );
  DEL4 U197 ( .I(n166), .Z(n167) );
  DEL4 U198 ( .I(n167), .Z(n168) );
  DEL2 U199 ( .I(n174), .Z(n200) );
  DEL4 U200 ( .I(Din[3]), .Z(n169) );
  DEL4 U201 ( .I(n169), .Z(n170) );
  DEL4 U202 ( .I(n170), .Z(n171) );
  DEL4 U203 ( .I(n171), .Z(n172) );
  DEL4 U204 ( .I(n172), .Z(n173) );
  DEL4 U205 ( .I(n173), .Z(n174) );
  DEL2 U206 ( .I(n180), .Z(n199) );
  DEL4 U207 ( .I(Din[2]), .Z(n175) );
  DEL4 U208 ( .I(n175), .Z(n176) );
  DEL4 U209 ( .I(n176), .Z(n177) );
  DEL4 U210 ( .I(n177), .Z(n178) );
  DEL4 U211 ( .I(n178), .Z(n179) );
  DEL4 U212 ( .I(n179), .Z(n180) );
  DEL2 U213 ( .I(n186), .Z(n198) );
  DEL4 U214 ( .I(Din[1]), .Z(n181) );
  DEL4 U215 ( .I(n181), .Z(n182) );
  DEL4 U216 ( .I(n182), .Z(n183) );
  DEL4 U217 ( .I(n183), .Z(n184) );
  DEL4 U218 ( .I(n184), .Z(n185) );
  DEL4 U219 ( .I(n185), .Z(n186) );
  DEL2 U220 ( .I(n192), .Z(n197) );
  DEL4 U221 ( .I(Din[0]), .Z(n187) );
  DEL4 U222 ( .I(n187), .Z(n188) );
  DEL4 U223 ( .I(n188), .Z(n189) );
  DEL4 U224 ( .I(n189), .Z(n190) );
  DEL4 U225 ( .I(n190), .Z(n191) );
  DEL4 U226 ( .I(n191), .Z(n192) );
  DEL4 U227 ( .I(ReadIn), .Z(n195) );
  DEL4 U228 ( .I(WriteIn), .Z(n194) );
  BUFFD1 U229 ( .I(SM_MemReadCmd), .Z(n196) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n277, n278, n279, n280, StateClockRaw, StateClock, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N217, N219, N220, N221, N445, N447, N448, N449,
         n6, n8, n9, n10, n11, n12, n13, n14, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n123, n124, n125, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, \add_384/carry[2] , \add_384/carry[3] ,
         \add_384/carry[4] , \add_303/carry[2] , \add_303/carry[3] ,
         \add_303/carry[4] , n1, n2, n3, n4, n5, n7, n15, n16, n63, n81, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n126, n127, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n246,
         n247, n248, n249, n251, n253, n254, n260, n261, n262, n263, n272,
         n273, n274, n275, n276;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [4:0] OldReadAr;
  wire   [4:0] OldWriteAr;
  assign ReadAddr[0] = N217;
  assign WriteAddr[0] = N445;
  assign WriteAddr[1] = \add_384/carry[2] ;
  assign ReadAddr[1] = \add_303/carry[2] ;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  OA21D1 U110 ( .A1(CurState[2]), .A2(n42), .B(n83), .Z(n30) );
  FIFOStateM_AWid5_DW01_inc_0 r105 ( .A({WriteAddr[4:2], \add_384/carry[2] , 
        N445}), .SUM({N76, N75, N74, N73, N72}) );
  FIFOStateM_AWid5_DW01_inc_1 r104 ( .A({ReadAddr[4], n209, n213, 
        \add_303/carry[2] , N217}), .SUM({N51, N50, N49, N48, N47}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n119), .CPN(StateClock), .CDN(n272), .QN(
        n103) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n126), .CPN(StateClock), .CDN(n272), .QN(
        n23) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n148), .CPN(StateClock), .CDN(n272), .QN(
        n20) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n152), .CPN(StateClock), .CDN(n272), .QN(n14) );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n156), .CPN(StateClock), .CDN(n272), .Q(
        OldWriteAr[4]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n160), .CPN(StateClock), .CDN(n273), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n164), .CPN(StateClock), .CDN(n272), .Q(
        OldReadAr[3]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n168), .CPN(StateClock), .CDN(n272), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n172), .CPN(StateClock), .CDN(n272), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n176), .CPN(StateClock), .CDN(n272), .Q(
        OldReadAr[4]) );
  DFNCND1 \NextState_reg[1]  ( .D(n180), .CPN(StateClock), .CDN(n273), .Q(
        NextState[1]), .QN(n125) );
  DFNCND1 \NextState_reg[2]  ( .D(n184), .CPN(StateClock), .CDN(n273), .Q(
        NextState[2]), .QN(n124) );
  DFNCND1 \NextState_reg[0]  ( .D(n188), .CPN(StateClock), .CDN(n273), .Q(
        NextState[0]), .QN(n123) );
  DFNCND1 ReadCmdr_reg ( .D(n192), .CPN(StateClock), .CDN(n273), .Q(n279) );
  DFNCND1 WriteCmdr_reg ( .D(n196), .CPN(StateClock), .CDN(n273), .Q(n280) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n273), 
        .Q(CurState[0]) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n273), 
        .Q(CurState[1]) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n144), 
        .Q(CurState[2]), .QN(n261) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n200), .E(N56), .CP(StateClock), .CDN(n144), 
        .QN(n275) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N52), .E(N56), .CP(StateClock), .CDN(n144), 
        .QN(n274) );
  EDFCND1 \ReadAr_reg[4]  ( .D(n205), .E(N56), .CP(StateClock), .CDN(n144), 
        .Q(ReadAddr[4]), .QN(n276) );
  EDFCND1 \ReadAr_reg[3]  ( .D(n206), .E(N56), .CP(StateClock), .CDN(n144), 
        .Q(ReadAddr[3]) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n210), .E(N56), .CP(StateClock), .CDN(n144), 
        .Q(ReadAddr[2]) );
  EDFCND1 \WriteAr_reg[1]  ( .D(n216), .E(n238), .CP(StateClock), .CDN(n144), 
        .Q(\add_384/carry[2] ), .QN(n21) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n221), .E(n238), .CP(StateClock), .CDN(n144), 
        .Q(N445), .QN(n24) );
  EDFCND1 \WriteAr_reg[4]  ( .D(n226), .E(n238), .CP(StateClock), .CDN(n144), 
        .Q(WriteAddr[4]) );
  EDFCND1 \WriteAr_reg[3]  ( .D(n230), .E(n238), .CP(StateClock), .CDN(n144), 
        .Q(WriteAddr[3]), .QN(n17) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n234), .E(n238), .CP(StateClock), .CDN(n144), 
        .Q(WriteAddr[2]), .QN(n22) );
  DFND1 FullFIFOr_reg ( .D(n1), .CPN(StateClock), .Q(n278) );
  DFND1 EmptyFIFOr_reg ( .D(n5), .CPN(StateClock), .Q(n277) );
  DEL3 U3 ( .I(n2), .Z(n1) );
  DEL4 U4 ( .I(n3), .Z(n2) );
  DEL4 U5 ( .I(n4), .Z(n3) );
  DEL4 U6 ( .I(n129), .Z(n4) );
  OAI31D4 U7 ( .A1(n8), .A2(Reset), .A3(ReadReq), .B(n9), .ZN(n129) );
  DEL3 U8 ( .I(n7), .Z(n5) );
  DEL4 U9 ( .I(n15), .Z(n7) );
  DEL4 U10 ( .I(n16), .Z(n15) );
  DEL4 U11 ( .I(n128), .Z(n16) );
  OAI31D4 U12 ( .A1(n6), .A2(WriteReq), .A3(Reset), .B(n63), .ZN(n128) );
  AO22D0 U13 ( .A1(n110), .A2(N74), .B1(n53), .B2(ReadAddr[2]), .Z(N79) );
  AO22D0 U14 ( .A1(n110), .A2(N75), .B1(n53), .B2(ReadAddr[3]), .Z(N80) );
  IOA22D0 U15 ( .B1(n239), .B2(n276), .A1(n110), .A2(N76), .ZN(N81) );
  OAI22D2 U16 ( .A1(n239), .A2(n225), .B1(n29), .B2(n82), .ZN(N77) );
  OAI22D0 U17 ( .A1(n239), .A2(n220), .B1(n29), .B2(n80), .ZN(N78) );
  OAI32D1 U18 ( .A1(n26), .A2(n27), .A3(n28), .B1(n29), .B2(n25), .ZN(n139) );
  OAI32D1 U19 ( .A1(n99), .A2(n100), .A3(n98), .B1(n101), .B2(n102), .ZN(n143)
         );
  OAI21D1 U20 ( .A1(n37), .A2(n123), .B(n38), .ZN(n140) );
  OAI22D0 U21 ( .A1(n37), .A2(n124), .B1(n50), .B2(n51), .ZN(n141) );
  DEL2 U22 ( .I(n125), .Z(n182) );
  MOAI22D1 U23 ( .A1(n276), .A2(n13), .B1(n13), .B2(OldReadAr[4]), .ZN(n133)
         );
  MOAI22D1 U24 ( .A1(n17), .A2(n18), .B1(n18), .B2(OldWriteAr[3]), .ZN(n134)
         );
  MOAI22D1 U25 ( .A1(n22), .A2(n18), .B1(n18), .B2(OldWriteAr[2]), .ZN(n136)
         );
  AO22D0 U26 ( .A1(ReadAddr[3]), .A2(n12), .B1(n13), .B2(OldReadAr[3]), .Z(
        n130) );
  AO22D0 U27 ( .A1(ReadAddr[2]), .A2(n12), .B1(n13), .B2(OldReadAr[2]), .Z(
        n132) );
  AO22D0 U28 ( .A1(WriteAddr[4]), .A2(n19), .B1(n18), .B2(OldWriteAr[4]), .Z(
        n137) );
  OAI22D0 U29 ( .A1(n12), .A2(n14), .B1(n275), .B2(n13), .ZN(n131) );
  OAI22D0 U30 ( .A1(n19), .A2(n20), .B1(n21), .B2(n18), .ZN(n135) );
  OAI22D0 U31 ( .A1(n19), .A2(n23), .B1(n24), .B2(n18), .ZN(n138) );
  OAI22D0 U32 ( .A1(n12), .A2(n103), .B1(n274), .B2(n13), .ZN(n145) );
  CKND2D0 U33 ( .A1(n260), .A2(n277), .ZN(n63) );
  AN2D1 U34 ( .A1(n261), .A2(n262), .Z(n81) );
  DEL4 U35 ( .I(n114), .Z(WriteCmd) );
  DEL4 U36 ( .I(n115), .Z(n114) );
  DEL4 U37 ( .I(n116), .Z(n115) );
  DEL4 U38 ( .I(n117), .Z(n116) );
  DEL4 U39 ( .I(n118), .Z(n117) );
  DEL4 U40 ( .I(n280), .Z(n118) );
  DEL3 U41 ( .I(n120), .Z(n119) );
  DEL4 U42 ( .I(n121), .Z(n120) );
  DEL4 U43 ( .I(n122), .Z(n121) );
  DEL4 U44 ( .I(n145), .Z(n122) );
  DEL3 U45 ( .I(n127), .Z(n126) );
  DEL4 U46 ( .I(n146), .Z(n127) );
  DEL4 U47 ( .I(n147), .Z(n146) );
  DEL4 U48 ( .I(n138), .Z(n147) );
  DEL3 U49 ( .I(n149), .Z(n148) );
  DEL4 U50 ( .I(n150), .Z(n149) );
  DEL4 U51 ( .I(n151), .Z(n150) );
  DEL4 U52 ( .I(n135), .Z(n151) );
  DEL3 U53 ( .I(n153), .Z(n152) );
  DEL4 U54 ( .I(n154), .Z(n153) );
  DEL4 U55 ( .I(n155), .Z(n154) );
  DEL4 U56 ( .I(n131), .Z(n155) );
  DEL3 U57 ( .I(n157), .Z(n156) );
  DEL4 U58 ( .I(n158), .Z(n157) );
  DEL4 U59 ( .I(n159), .Z(n158) );
  DEL4 U60 ( .I(n137), .Z(n159) );
  DEL3 U61 ( .I(n161), .Z(n160) );
  DEL4 U62 ( .I(n162), .Z(n161) );
  DEL4 U63 ( .I(n163), .Z(n162) );
  DEL4 U64 ( .I(n132), .Z(n163) );
  DEL3 U65 ( .I(n165), .Z(n164) );
  DEL4 U66 ( .I(n166), .Z(n165) );
  DEL4 U67 ( .I(n167), .Z(n166) );
  DEL4 U68 ( .I(n130), .Z(n167) );
  DEL3 U69 ( .I(n169), .Z(n168) );
  DEL4 U70 ( .I(n170), .Z(n169) );
  DEL4 U71 ( .I(n171), .Z(n170) );
  DEL4 U72 ( .I(n136), .Z(n171) );
  DEL3 U73 ( .I(n173), .Z(n172) );
  DEL4 U74 ( .I(n174), .Z(n173) );
  DEL4 U75 ( .I(n175), .Z(n174) );
  DEL4 U76 ( .I(n134), .Z(n175) );
  DEL3 U77 ( .I(n177), .Z(n176) );
  DEL4 U78 ( .I(n178), .Z(n177) );
  DEL4 U79 ( .I(n179), .Z(n178) );
  DEL4 U80 ( .I(n133), .Z(n179) );
  OAI22D0 U81 ( .A1(n37), .A2(n182), .B1(n50), .B2(n58), .ZN(n142) );
  DEL4 U82 ( .I(n181), .Z(n180) );
  DEL4 U83 ( .I(n183), .Z(n181) );
  DEL4 U84 ( .I(n142), .Z(n183) );
  DEL3 U85 ( .I(n185), .Z(n184) );
  DEL4 U86 ( .I(n186), .Z(n185) );
  DEL4 U87 ( .I(n187), .Z(n186) );
  DEL4 U88 ( .I(n141), .Z(n187) );
  DEL3 U89 ( .I(n189), .Z(n188) );
  DEL4 U90 ( .I(n190), .Z(n189) );
  DEL4 U91 ( .I(n191), .Z(n190) );
  DEL4 U92 ( .I(n140), .Z(n191) );
  DEL4 U93 ( .I(n193), .Z(n192) );
  DEL4 U94 ( .I(n194), .Z(n193) );
  DEL4 U95 ( .I(n195), .Z(n194) );
  DEL4 U96 ( .I(n143), .Z(n195) );
  DEL4 U97 ( .I(n197), .Z(n196) );
  DEL4 U98 ( .I(n198), .Z(n197) );
  DEL4 U99 ( .I(n199), .Z(n198) );
  DEL4 U100 ( .I(n139), .Z(n199) );
  DEL2 U101 ( .I(N53), .Z(n200) );
  NR2D0 U102 ( .A1(n70), .A2(n101), .ZN(N53) );
  DEL4 U103 ( .I(n275), .Z(n201) );
  DEL4 U104 ( .I(n201), .Z(n202) );
  DEL4 U105 ( .I(n274), .Z(n203) );
  DEL4 U106 ( .I(n203), .Z(n204) );
  DEL2 U107 ( .I(N57), .Z(n205) );
  INR2D0 U108 ( .A1(N51), .B1(n101), .ZN(N57) );
  DEL2 U109 ( .I(n207), .Z(n206) );
  INR2D0 U111 ( .A1(N50), .B1(n101), .ZN(N55) );
  DEL4 U112 ( .I(n208), .Z(n207) );
  DEL4 U113 ( .I(N55), .Z(n208) );
  DEL4 U114 ( .I(ReadAddr[3]), .Z(n209) );
  DEL2 U115 ( .I(n211), .Z(n210) );
  INR2D0 U116 ( .A1(N49), .B1(n101), .ZN(N54) );
  DEL4 U117 ( .I(n212), .Z(n211) );
  DEL4 U118 ( .I(N54), .Z(n212) );
  DEL4 U119 ( .I(ReadAddr[2]), .Z(n213) );
  DEL1 U120 ( .I(n11), .Z(n214) );
  ND2D0 U121 ( .A1(n240), .A2(n101), .ZN(N56) );
  DEL4 U122 ( .I(n214), .Z(n215) );
  NR3D0 U123 ( .A1(CurState[1]), .A2(CurState[2]), .A3(CurState[0]), .ZN(n11)
         );
  DEL2 U124 ( .I(n217), .Z(n216) );
  DEL4 U125 ( .I(n218), .Z(n217) );
  DEL4 U126 ( .I(n219), .Z(n218) );
  DEL4 U127 ( .I(N78), .Z(n219) );
  DEL4 U128 ( .I(n202), .Z(n220) );
  DEL2 U129 ( .I(n222), .Z(n221) );
  DEL4 U130 ( .I(n223), .Z(n222) );
  DEL4 U131 ( .I(n224), .Z(n223) );
  DEL4 U132 ( .I(N77), .Z(n224) );
  DEL4 U133 ( .I(n204), .Z(n225) );
  DEL2 U134 ( .I(n227), .Z(n226) );
  DEL4 U135 ( .I(n228), .Z(n227) );
  DEL4 U136 ( .I(n229), .Z(n228) );
  DEL4 U137 ( .I(N81), .Z(n229) );
  DEL2 U138 ( .I(n231), .Z(n230) );
  DEL4 U139 ( .I(n232), .Z(n231) );
  DEL4 U140 ( .I(n233), .Z(n232) );
  DEL4 U141 ( .I(N80), .Z(n233) );
  DEL2 U142 ( .I(n235), .Z(n234) );
  DEL4 U143 ( .I(n236), .Z(n235) );
  DEL4 U144 ( .I(n237), .Z(n236) );
  DEL4 U145 ( .I(N79), .Z(n237) );
  DEL1 U146 ( .I(n242), .Z(n238) );
  BUFFD0 U147 ( .I(n8), .Z(n239) );
  DEL4 U148 ( .I(n241), .Z(n240) );
  DEL4 U149 ( .I(n6), .Z(n241) );
  CKNXD0 U150 ( .I(n215), .ZN(n6) );
  INVD0 U151 ( .I(CurState[1]), .ZN(n42) );
  DEL4 U152 ( .I(n243), .Z(n242) );
  DEL4 U153 ( .I(n244), .Z(n243) );
  DEL4 U154 ( .I(N82), .Z(n244) );
  ND3D8 U155 ( .A1(n239), .A2(n240), .A3(n29), .ZN(N82) );
  DEL2 U156 ( .I(n246), .Z(ReadCmd) );
  DEL4 U157 ( .I(n247), .Z(n246) );
  DEL4 U158 ( .I(n248), .Z(n247) );
  DEL4 U159 ( .I(n279), .Z(n248) );
  DEL4 U160 ( .I(n254), .Z(n249) );
  CKNXD16 U161 ( .I(n249), .ZN(EmptyFIFO) );
  DEL4 U162 ( .I(n253), .Z(n251) );
  CKNXD16 U163 ( .I(n251), .ZN(FullFIFO) );
  CKND0 U164 ( .CLK(n278), .CN(n253) );
  CKND0 U165 ( .CLK(n277), .CN(n254) );
  OAI21D0 U166 ( .A1(n10), .A2(Reset), .B(n278), .ZN(n9) );
  CKND0 U167 ( .CLK(Reset), .CN(n262) );
  CKND0 U168 ( .CLK(CurState[0]), .CN(n263) );
  CKND2D0 U169 ( .A1(n263), .A2(n81), .ZN(n260) );
  INVD1 U170 ( .I(N48), .ZN(n70) );
  INVD1 U171 ( .I(n53), .ZN(n8) );
  INVD1 U172 ( .I(n13), .ZN(n12) );
  INVD1 U173 ( .I(n18), .ZN(n19) );
  INVD1 U174 ( .I(Reset), .ZN(n272) );
  INVD1 U175 ( .I(Reset), .ZN(n273) );
  AOI221D0 U176 ( .A1(CurState[0]), .A2(n54), .B1(n62), .B2(n263), .C(n41), 
        .ZN(n61) );
  OAI31D0 U177 ( .A1(n71), .A2(n47), .A3(n45), .B(n72), .ZN(n62) );
  INVD1 U178 ( .I(n73), .ZN(n72) );
  IND3D1 U179 ( .A1(n46), .B1(n49), .B2(n48), .ZN(n71) );
  ND3D1 U180 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n54) );
  XNR2D1 U181 ( .A1(n274), .A2(n82), .ZN(n74) );
  XNR2D1 U182 ( .A1(n275), .A2(n80), .ZN(n75) );
  NR3D0 U183 ( .A1(n77), .A2(n78), .A3(n79), .ZN(n76) );
  AN2D1 U184 ( .A1(n55), .A2(CurState[0]), .Z(n41) );
  XNR2D1 U185 ( .A1(n17), .A2(N50), .ZN(n67) );
  XNR2D1 U186 ( .A1(n276), .A2(N76), .ZN(n79) );
  XNR2D1 U187 ( .A1(n22), .A2(N49), .ZN(n68) );
  INVD1 U188 ( .I(n225), .ZN(N217) );
  INVD1 U189 ( .I(n220), .ZN(\add_303/carry[2] ) );
  ND3D1 U190 ( .A1(n25), .A2(n26), .A3(WriteReq), .ZN(n18) );
  ND3D1 U191 ( .A1(n102), .A2(n99), .A3(ReadReq), .ZN(n13) );
  NR3D0 U192 ( .A1(n42), .A2(n263), .A3(n261), .ZN(n53) );
  INVD1 U193 ( .I(n102), .ZN(n100) );
  INVD1 U194 ( .I(WriteReq), .ZN(n28) );
  INVD1 U195 ( .I(n25), .ZN(n27) );
  ND2D1 U196 ( .A1(n30), .A2(n8), .ZN(n102) );
  ND2D1 U197 ( .A1(n30), .A2(n6), .ZN(n25) );
  INVD1 U198 ( .I(n37), .ZN(n50) );
  ND3D1 U199 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n26) );
  XNR2D1 U200 ( .A1(n24), .A2(n23), .ZN(n31) );
  XNR2D1 U201 ( .A1(n21), .A2(n20), .ZN(n32) );
  NR3D0 U202 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n33) );
  ND3D1 U203 ( .A1(n104), .A2(n105), .A3(n106), .ZN(n99) );
  XNR2D1 U204 ( .A1(n274), .A2(n103), .ZN(n104) );
  XNR2D1 U205 ( .A1(n275), .A2(n14), .ZN(n105) );
  NR3D0 U206 ( .A1(n107), .A2(n108), .A3(n109), .ZN(n106) );
  INVD1 U207 ( .I(n29), .ZN(n110) );
  INR2D1 U208 ( .A1(N47), .B1(n101), .ZN(N52) );
  ND3D1 U209 ( .A1(n48), .A2(n261), .A3(n49), .ZN(n44) );
  XNR2D1 U210 ( .A1(n21), .A2(\add_303/carry[2] ), .ZN(n93) );
  XNR2D1 U211 ( .A1(n24), .A2(N47), .ZN(n69) );
  XNR2D1 U212 ( .A1(n24), .A2(N217), .ZN(n95) );
  ND3D1 U213 ( .A1(n84), .A2(n85), .A3(n86), .ZN(n57) );
  XNR2D1 U214 ( .A1(n21), .A2(\add_303/carry[2] ), .ZN(n84) );
  NR3D0 U215 ( .A1(n87), .A2(n88), .A3(n89), .ZN(n86) );
  XNR2D1 U216 ( .A1(N449), .A2(ReadAddr[4]), .ZN(n85) );
  INVD1 U217 ( .I(N73), .ZN(n80) );
  XOR2D1 U218 ( .A1(\add_303/carry[2] ), .A2(n21), .Z(n47) );
  INVD1 U219 ( .I(ReadReq), .ZN(n98) );
  INVD1 U220 ( .I(Reset), .ZN(n144) );
  AOI21D1 U221 ( .A1(CurState[0]), .A2(n52), .B(n53), .ZN(n51) );
  OAI32D1 U222 ( .A1(n54), .A2(n55), .A3(n42), .B1(n56), .B2(n261), .ZN(n52)
         );
  INVD1 U223 ( .I(n57), .ZN(n56) );
  OAI211D1 U224 ( .A1(CurState[0]), .A2(n39), .B(n40), .C(n37), .ZN(n38) );
  NR4D0 U225 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n39) );
  OAI21D1 U226 ( .A1(n41), .A2(n42), .B(n261), .ZN(n40) );
  AOI21D1 U227 ( .A1(CurState[2]), .A2(CurState[0]), .B(n11), .ZN(n10) );
  NR3D0 U228 ( .A1(n59), .A2(n11), .A3(n60), .ZN(n58) );
  AOI21D1 U229 ( .A1(n73), .A2(n57), .B(n83), .ZN(n59) );
  NR3D0 U230 ( .A1(n42), .A2(CurState[2]), .A3(n61), .ZN(n60) );
  XOR2D1 U231 ( .A1(N221), .A2(WriteAddr[4]), .Z(n45) );
  AN3D1 U232 ( .A1(n64), .A2(n65), .A3(n66), .Z(n55) );
  XNR2D1 U233 ( .A1(n21), .A2(n70), .ZN(n64) );
  NR3D0 U234 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n66) );
  XNR2D1 U235 ( .A1(WriteAddr[4]), .A2(N51), .ZN(n65) );
  OAI211D1 U236 ( .A1(CurState[1]), .A2(n263), .B(n30), .C(n96), .ZN(n37) );
  AOI21D1 U237 ( .A1(WriteReq), .A2(n11), .B(n97), .ZN(n96) );
  AOI21D1 U238 ( .A1(CurState[0]), .A2(n98), .B(n261), .ZN(n97) );
  ND2D1 U239 ( .A1(ReadCmd), .A2(n240), .ZN(n101) );
  ND2D1 U240 ( .A1(n280), .A2(n239), .ZN(n29) );
  XNR2D1 U241 ( .A1(N219), .A2(WriteAddr[2]), .ZN(n49) );
  ND3D1 U242 ( .A1(CurState[0]), .A2(n42), .A3(CurState[2]), .ZN(n83) );
  ND3D1 U243 ( .A1(n90), .A2(n91), .A3(n92), .ZN(n73) );
  XNR2D1 U244 ( .A1(ReadAddr[4]), .A2(WriteAddr[4]), .ZN(n90) );
  XNR2D1 U245 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n91) );
  NR3D0 U246 ( .A1(n93), .A2(n94), .A3(n95), .ZN(n92) );
  XNR2D1 U247 ( .A1(N220), .A2(WriteAddr[3]), .ZN(n48) );
  INVD1 U248 ( .I(N72), .ZN(n82) );
  XOR2D1 U249 ( .A1(N217), .A2(N445), .Z(n46) );
  XNR2D1 U250 ( .A1(n17), .A2(ReadAddr[3]), .ZN(n94) );
  XOR2D1 U251 ( .A1(ReadAddr[3]), .A2(N75), .Z(n77) );
  XNR2D1 U252 ( .A1(n274), .A2(N445), .ZN(n89) );
  XOR2D1 U253 ( .A1(ReadAddr[3]), .A2(N448), .Z(n87) );
  XOR2D1 U254 ( .A1(ReadAddr[3]), .A2(OldReadAr[3]), .Z(n107) );
  XOR2D1 U255 ( .A1(ReadAddr[2]), .A2(N74), .Z(n78) );
  XOR2D1 U256 ( .A1(ReadAddr[2]), .A2(N447), .Z(n88) );
  XOR2D1 U257 ( .A1(WriteAddr[4]), .A2(OldWriteAr[4]), .Z(n36) );
  XOR2D1 U258 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .Z(n108) );
  XNR2D1 U259 ( .A1(n17), .A2(OldWriteAr[3]), .ZN(n34) );
  XNR2D1 U260 ( .A1(n22), .A2(OldWriteAr[2]), .ZN(n35) );
  XNR2D1 U261 ( .A1(n276), .A2(OldReadAr[4]), .ZN(n109) );
  ND2D1 U262 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  CKXOR2D0 U263 ( .A1(ReadAddr[4]), .A2(\add_303/carry[4] ), .Z(N221) );
  AN2D0 U264 ( .A1(ReadAddr[3]), .A2(\add_303/carry[3] ), .Z(
        \add_303/carry[4] ) );
  CKXOR2D0 U265 ( .A1(\add_303/carry[3] ), .A2(ReadAddr[3]), .Z(N220) );
  AN2D0 U266 ( .A1(ReadAddr[2]), .A2(\add_303/carry[2] ), .Z(
        \add_303/carry[3] ) );
  CKXOR2D0 U267 ( .A1(\add_303/carry[2] ), .A2(ReadAddr[2]), .Z(N219) );
  CKXOR2D0 U268 ( .A1(WriteAddr[4]), .A2(\add_384/carry[4] ), .Z(N449) );
  AN2D0 U269 ( .A1(WriteAddr[3]), .A2(\add_384/carry[3] ), .Z(
        \add_384/carry[4] ) );
  CKXOR2D0 U270 ( .A1(\add_384/carry[3] ), .A2(WriteAddr[3]), .Z(N448) );
  AN2D0 U271 ( .A1(WriteAddr[2]), .A2(\add_384/carry[2] ), .Z(
        \add_384/carry[3] ) );
  CKXOR2D0 U272 ( .A1(\add_384/carry[2] ), .A2(WriteAddr[2]), .Z(N447) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N79, N80, N81, N82, N83, ClockR, ClockW,
         Dreadyr, \Storage[31][32] , \Storage[31][31] , \Storage[31][30] ,
         \Storage[31][29] , \Storage[31][28] , \Storage[31][27] ,
         \Storage[31][26] , \Storage[31][25] , \Storage[31][24] ,
         \Storage[31][23] , \Storage[31][22] , \Storage[31][21] ,
         \Storage[31][20] , \Storage[31][19] , \Storage[31][18] ,
         \Storage[31][17] , \Storage[31][16] , \Storage[31][15] ,
         \Storage[31][14] , \Storage[31][13] , \Storage[31][12] ,
         \Storage[31][11] , \Storage[31][10] , \Storage[31][9] ,
         \Storage[31][8] , \Storage[31][7] , \Storage[31][6] ,
         \Storage[31][5] , \Storage[31][4] , \Storage[31][3] ,
         \Storage[31][2] , \Storage[31][1] , \Storage[31][0] ,
         \Storage[30][32] , \Storage[30][31] , \Storage[30][30] ,
         \Storage[30][29] , \Storage[30][28] , \Storage[30][27] ,
         \Storage[30][26] , \Storage[30][25] , \Storage[30][24] ,
         \Storage[30][23] , \Storage[30][22] , \Storage[30][21] ,
         \Storage[30][20] , \Storage[30][19] , \Storage[30][18] ,
         \Storage[30][17] , \Storage[30][16] , \Storage[30][15] ,
         \Storage[30][14] , \Storage[30][13] , \Storage[30][12] ,
         \Storage[30][11] , \Storage[30][10] , \Storage[30][9] ,
         \Storage[30][8] , \Storage[30][7] , \Storage[30][6] ,
         \Storage[30][5] , \Storage[30][4] , \Storage[30][3] ,
         \Storage[30][2] , \Storage[30][1] , \Storage[30][0] ,
         \Storage[29][32] , \Storage[29][31] , \Storage[29][30] ,
         \Storage[29][29] , \Storage[29][28] , \Storage[29][27] ,
         \Storage[29][26] , \Storage[29][25] , \Storage[29][24] ,
         \Storage[29][23] , \Storage[29][22] , \Storage[29][21] ,
         \Storage[29][20] , \Storage[29][19] , \Storage[29][18] ,
         \Storage[29][17] , \Storage[29][16] , \Storage[29][15] ,
         \Storage[29][14] , \Storage[29][13] , \Storage[29][12] ,
         \Storage[29][11] , \Storage[29][10] , \Storage[29][9] ,
         \Storage[29][8] , \Storage[29][7] , \Storage[29][6] ,
         \Storage[29][5] , \Storage[29][4] , \Storage[29][3] ,
         \Storage[29][2] , \Storage[29][1] , \Storage[29][0] ,
         \Storage[28][32] , \Storage[28][31] , \Storage[28][30] ,
         \Storage[28][29] , \Storage[28][28] , \Storage[28][27] ,
         \Storage[28][26] , \Storage[28][25] , \Storage[28][24] ,
         \Storage[28][23] , \Storage[28][22] , \Storage[28][21] ,
         \Storage[28][20] , \Storage[28][19] , \Storage[28][18] ,
         \Storage[28][17] , \Storage[28][16] , \Storage[28][15] ,
         \Storage[28][14] , \Storage[28][13] , \Storage[28][12] ,
         \Storage[28][11] , \Storage[28][10] , \Storage[28][9] ,
         \Storage[28][8] , \Storage[28][7] , \Storage[28][6] ,
         \Storage[28][5] , \Storage[28][4] , \Storage[28][3] ,
         \Storage[28][2] , \Storage[28][1] , \Storage[28][0] ,
         \Storage[27][32] , \Storage[27][31] , \Storage[27][30] ,
         \Storage[27][29] , \Storage[27][28] , \Storage[27][27] ,
         \Storage[27][26] , \Storage[27][25] , \Storage[27][24] ,
         \Storage[27][23] , \Storage[27][22] , \Storage[27][21] ,
         \Storage[27][20] , \Storage[27][19] , \Storage[27][18] ,
         \Storage[27][17] , \Storage[27][16] , \Storage[27][15] ,
         \Storage[27][14] , \Storage[27][13] , \Storage[27][12] ,
         \Storage[27][11] , \Storage[27][10] , \Storage[27][9] ,
         \Storage[27][8] , \Storage[27][7] , \Storage[27][6] ,
         \Storage[27][5] , \Storage[27][4] , \Storage[27][3] ,
         \Storage[27][2] , \Storage[27][1] , \Storage[27][0] ,
         \Storage[26][32] , \Storage[26][31] , \Storage[26][30] ,
         \Storage[26][29] , \Storage[26][28] , \Storage[26][27] ,
         \Storage[26][26] , \Storage[26][25] , \Storage[26][24] ,
         \Storage[26][23] , \Storage[26][22] , \Storage[26][21] ,
         \Storage[26][20] , \Storage[26][19] , \Storage[26][18] ,
         \Storage[26][17] , \Storage[26][16] , \Storage[26][15] ,
         \Storage[26][14] , \Storage[26][13] , \Storage[26][12] ,
         \Storage[26][11] , \Storage[26][10] , \Storage[26][9] ,
         \Storage[26][8] , \Storage[26][7] , \Storage[26][6] ,
         \Storage[26][5] , \Storage[26][4] , \Storage[26][3] ,
         \Storage[26][2] , \Storage[26][1] , \Storage[26][0] ,
         \Storage[25][32] , \Storage[25][31] , \Storage[25][30] ,
         \Storage[25][29] , \Storage[25][28] , \Storage[25][27] ,
         \Storage[25][26] , \Storage[25][25] , \Storage[25][24] ,
         \Storage[25][23] , \Storage[25][22] , \Storage[25][21] ,
         \Storage[25][20] , \Storage[25][19] , \Storage[25][18] ,
         \Storage[25][17] , \Storage[25][16] , \Storage[25][15] ,
         \Storage[25][14] , \Storage[25][13] , \Storage[25][12] ,
         \Storage[25][11] , \Storage[25][10] , \Storage[25][9] ,
         \Storage[25][8] , \Storage[25][7] , \Storage[25][6] ,
         \Storage[25][5] , \Storage[25][4] , \Storage[25][3] ,
         \Storage[25][2] , \Storage[25][1] , \Storage[25][0] ,
         \Storage[24][32] , \Storage[24][31] , \Storage[24][30] ,
         \Storage[24][29] , \Storage[24][28] , \Storage[24][27] ,
         \Storage[24][26] , \Storage[24][25] , \Storage[24][24] ,
         \Storage[24][23] , \Storage[24][22] , \Storage[24][21] ,
         \Storage[24][20] , \Storage[24][19] , \Storage[24][18] ,
         \Storage[24][17] , \Storage[24][16] , \Storage[24][15] ,
         \Storage[24][14] , \Storage[24][13] , \Storage[24][12] ,
         \Storage[24][11] , \Storage[24][10] , \Storage[24][9] ,
         \Storage[24][8] , \Storage[24][7] , \Storage[24][6] ,
         \Storage[24][5] , \Storage[24][4] , \Storage[24][3] ,
         \Storage[24][2] , \Storage[24][1] , \Storage[24][0] ,
         \Storage[23][32] , \Storage[23][31] , \Storage[23][30] ,
         \Storage[23][29] , \Storage[23][28] , \Storage[23][27] ,
         \Storage[23][26] , \Storage[23][25] , \Storage[23][24] ,
         \Storage[23][23] , \Storage[23][22] , \Storage[23][21] ,
         \Storage[23][20] , \Storage[23][19] , \Storage[23][18] ,
         \Storage[23][17] , \Storage[23][16] , \Storage[23][15] ,
         \Storage[23][14] , \Storage[23][13] , \Storage[23][12] ,
         \Storage[23][11] , \Storage[23][10] , \Storage[23][9] ,
         \Storage[23][8] , \Storage[23][7] , \Storage[23][6] ,
         \Storage[23][5] , \Storage[23][4] , \Storage[23][3] ,
         \Storage[23][2] , \Storage[23][1] , \Storage[23][0] ,
         \Storage[22][32] , \Storage[22][31] , \Storage[22][30] ,
         \Storage[22][29] , \Storage[22][28] , \Storage[22][27] ,
         \Storage[22][26] , \Storage[22][25] , \Storage[22][24] ,
         \Storage[22][23] , \Storage[22][22] , \Storage[22][21] ,
         \Storage[22][20] , \Storage[22][19] , \Storage[22][18] ,
         \Storage[22][17] , \Storage[22][16] , \Storage[22][15] ,
         \Storage[22][14] , \Storage[22][13] , \Storage[22][12] ,
         \Storage[22][11] , \Storage[22][10] , \Storage[22][9] ,
         \Storage[22][8] , \Storage[22][7] , \Storage[22][6] ,
         \Storage[22][5] , \Storage[22][4] , \Storage[22][3] ,
         \Storage[22][2] , \Storage[22][1] , \Storage[22][0] ,
         \Storage[21][32] , \Storage[21][31] , \Storage[21][30] ,
         \Storage[21][29] , \Storage[21][28] , \Storage[21][27] ,
         \Storage[21][26] , \Storage[21][25] , \Storage[21][24] ,
         \Storage[21][23] , \Storage[21][22] , \Storage[21][21] ,
         \Storage[21][20] , \Storage[21][19] , \Storage[21][18] ,
         \Storage[21][17] , \Storage[21][16] , \Storage[21][15] ,
         \Storage[21][14] , \Storage[21][13] , \Storage[21][12] ,
         \Storage[21][11] , \Storage[21][10] , \Storage[21][9] ,
         \Storage[21][8] , \Storage[21][7] , \Storage[21][6] ,
         \Storage[21][5] , \Storage[21][4] , \Storage[21][3] ,
         \Storage[21][2] , \Storage[21][1] , \Storage[21][0] ,
         \Storage[20][32] , \Storage[20][31] , \Storage[20][30] ,
         \Storage[20][29] , \Storage[20][28] , \Storage[20][27] ,
         \Storage[20][26] , \Storage[20][25] , \Storage[20][24] ,
         \Storage[20][23] , \Storage[20][22] , \Storage[20][21] ,
         \Storage[20][20] , \Storage[20][19] , \Storage[20][18] ,
         \Storage[20][17] , \Storage[20][16] , \Storage[20][15] ,
         \Storage[20][14] , \Storage[20][13] , \Storage[20][12] ,
         \Storage[20][11] , \Storage[20][10] , \Storage[20][9] ,
         \Storage[20][8] , \Storage[20][7] , \Storage[20][6] ,
         \Storage[20][5] , \Storage[20][4] , \Storage[20][3] ,
         \Storage[20][2] , \Storage[20][1] , \Storage[20][0] ,
         \Storage[19][32] , \Storage[19][31] , \Storage[19][30] ,
         \Storage[19][29] , \Storage[19][28] , \Storage[19][27] ,
         \Storage[19][26] , \Storage[19][25] , \Storage[19][24] ,
         \Storage[19][23] , \Storage[19][22] , \Storage[19][21] ,
         \Storage[19][20] , \Storage[19][19] , \Storage[19][18] ,
         \Storage[19][17] , \Storage[19][16] , \Storage[19][15] ,
         \Storage[19][14] , \Storage[19][13] , \Storage[19][12] ,
         \Storage[19][11] , \Storage[19][10] , \Storage[19][9] ,
         \Storage[19][8] , \Storage[19][7] , \Storage[19][6] ,
         \Storage[19][5] , \Storage[19][4] , \Storage[19][3] ,
         \Storage[19][2] , \Storage[19][1] , \Storage[19][0] ,
         \Storage[18][32] , \Storage[18][31] , \Storage[18][30] ,
         \Storage[18][29] , \Storage[18][28] , \Storage[18][27] ,
         \Storage[18][26] , \Storage[18][25] , \Storage[18][24] ,
         \Storage[18][23] , \Storage[18][22] , \Storage[18][21] ,
         \Storage[18][20] , \Storage[18][19] , \Storage[18][18] ,
         \Storage[18][17] , \Storage[18][16] , \Storage[18][15] ,
         \Storage[18][14] , \Storage[18][13] , \Storage[18][12] ,
         \Storage[18][11] , \Storage[18][10] , \Storage[18][9] ,
         \Storage[18][8] , \Storage[18][7] , \Storage[18][6] ,
         \Storage[18][5] , \Storage[18][4] , \Storage[18][3] ,
         \Storage[18][2] , \Storage[18][1] , \Storage[18][0] ,
         \Storage[17][32] , \Storage[17][31] , \Storage[17][30] ,
         \Storage[17][29] , \Storage[17][28] , \Storage[17][27] ,
         \Storage[17][26] , \Storage[17][25] , \Storage[17][24] ,
         \Storage[17][23] , \Storage[17][22] , \Storage[17][21] ,
         \Storage[17][20] , \Storage[17][19] , \Storage[17][18] ,
         \Storage[17][17] , \Storage[17][16] , \Storage[17][15] ,
         \Storage[17][14] , \Storage[17][13] , \Storage[17][12] ,
         \Storage[17][11] , \Storage[17][10] , \Storage[17][9] ,
         \Storage[17][8] , \Storage[17][7] , \Storage[17][6] ,
         \Storage[17][5] , \Storage[17][4] , \Storage[17][3] ,
         \Storage[17][2] , \Storage[17][1] , \Storage[17][0] ,
         \Storage[16][32] , \Storage[16][31] , \Storage[16][30] ,
         \Storage[16][29] , \Storage[16][28] , \Storage[16][27] ,
         \Storage[16][26] , \Storage[16][25] , \Storage[16][24] ,
         \Storage[16][23] , \Storage[16][22] , \Storage[16][21] ,
         \Storage[16][20] , \Storage[16][19] , \Storage[16][18] ,
         \Storage[16][17] , \Storage[16][16] , \Storage[16][15] ,
         \Storage[16][14] , \Storage[16][13] , \Storage[16][12] ,
         \Storage[16][11] , \Storage[16][10] , \Storage[16][9] ,
         \Storage[16][8] , \Storage[16][7] , \Storage[16][6] ,
         \Storage[16][5] , \Storage[16][4] , \Storage[16][3] ,
         \Storage[16][2] , \Storage[16][1] , \Storage[16][0] ,
         \Storage[15][32] , \Storage[15][31] , \Storage[15][30] ,
         \Storage[15][29] , \Storage[15][28] , \Storage[15][27] ,
         \Storage[15][26] , \Storage[15][25] , \Storage[15][24] ,
         \Storage[15][23] , \Storage[15][22] , \Storage[15][21] ,
         \Storage[15][20] , \Storage[15][19] , \Storage[15][18] ,
         \Storage[15][17] , \Storage[15][16] , \Storage[15][15] ,
         \Storage[15][14] , \Storage[15][13] , \Storage[15][12] ,
         \Storage[15][11] , \Storage[15][10] , \Storage[15][9] ,
         \Storage[15][8] , \Storage[15][7] , \Storage[15][6] ,
         \Storage[15][5] , \Storage[15][4] , \Storage[15][3] ,
         \Storage[15][2] , \Storage[15][1] , \Storage[15][0] ,
         \Storage[14][32] , \Storage[14][31] , \Storage[14][30] ,
         \Storage[14][29] , \Storage[14][28] , \Storage[14][27] ,
         \Storage[14][26] , \Storage[14][25] , \Storage[14][24] ,
         \Storage[14][23] , \Storage[14][22] , \Storage[14][21] ,
         \Storage[14][20] , \Storage[14][19] , \Storage[14][18] ,
         \Storage[14][17] , \Storage[14][16] , \Storage[14][15] ,
         \Storage[14][14] , \Storage[14][13] , \Storage[14][12] ,
         \Storage[14][11] , \Storage[14][10] , \Storage[14][9] ,
         \Storage[14][8] , \Storage[14][7] , \Storage[14][6] ,
         \Storage[14][5] , \Storage[14][4] , \Storage[14][3] ,
         \Storage[14][2] , \Storage[14][1] , \Storage[14][0] ,
         \Storage[13][32] , \Storage[13][31] , \Storage[13][30] ,
         \Storage[13][29] , \Storage[13][28] , \Storage[13][27] ,
         \Storage[13][26] , \Storage[13][25] , \Storage[13][24] ,
         \Storage[13][23] , \Storage[13][22] , \Storage[13][21] ,
         \Storage[13][20] , \Storage[13][19] , \Storage[13][18] ,
         \Storage[13][17] , \Storage[13][16] , \Storage[13][15] ,
         \Storage[13][14] , \Storage[13][13] , \Storage[13][12] ,
         \Storage[13][11] , \Storage[13][10] , \Storage[13][9] ,
         \Storage[13][8] , \Storage[13][7] , \Storage[13][6] ,
         \Storage[13][5] , \Storage[13][4] , \Storage[13][3] ,
         \Storage[13][2] , \Storage[13][1] , \Storage[13][0] ,
         \Storage[12][32] , \Storage[12][31] , \Storage[12][30] ,
         \Storage[12][29] , \Storage[12][28] , \Storage[12][27] ,
         \Storage[12][26] , \Storage[12][25] , \Storage[12][24] ,
         \Storage[12][23] , \Storage[12][22] , \Storage[12][21] ,
         \Storage[12][20] , \Storage[12][19] , \Storage[12][18] ,
         \Storage[12][17] , \Storage[12][16] , \Storage[12][15] ,
         \Storage[12][14] , \Storage[12][13] , \Storage[12][12] ,
         \Storage[12][11] , \Storage[12][10] , \Storage[12][9] ,
         \Storage[12][8] , \Storage[12][7] , \Storage[12][6] ,
         \Storage[12][5] , \Storage[12][4] , \Storage[12][3] ,
         \Storage[12][2] , \Storage[12][1] , \Storage[12][0] ,
         \Storage[11][32] , \Storage[11][31] , \Storage[11][30] ,
         \Storage[11][29] , \Storage[11][28] , \Storage[11][27] ,
         \Storage[11][26] , \Storage[11][25] , \Storage[11][24] ,
         \Storage[11][23] , \Storage[11][22] , \Storage[11][21] ,
         \Storage[11][20] , \Storage[11][19] , \Storage[11][18] ,
         \Storage[11][17] , \Storage[11][16] , \Storage[11][15] ,
         \Storage[11][14] , \Storage[11][13] , \Storage[11][12] ,
         \Storage[11][11] , \Storage[11][10] , \Storage[11][9] ,
         \Storage[11][8] , \Storage[11][7] , \Storage[11][6] ,
         \Storage[11][5] , \Storage[11][4] , \Storage[11][3] ,
         \Storage[11][2] , \Storage[11][1] , \Storage[11][0] ,
         \Storage[10][32] , \Storage[10][31] , \Storage[10][30] ,
         \Storage[10][29] , \Storage[10][28] , \Storage[10][27] ,
         \Storage[10][26] , \Storage[10][25] , \Storage[10][24] ,
         \Storage[10][23] , \Storage[10][22] , \Storage[10][21] ,
         \Storage[10][20] , \Storage[10][19] , \Storage[10][18] ,
         \Storage[10][17] , \Storage[10][16] , \Storage[10][15] ,
         \Storage[10][14] , \Storage[10][13] , \Storage[10][12] ,
         \Storage[10][11] , \Storage[10][10] , \Storage[10][9] ,
         \Storage[10][8] , \Storage[10][7] , \Storage[10][6] ,
         \Storage[10][5] , \Storage[10][4] , \Storage[10][3] ,
         \Storage[10][2] , \Storage[10][1] , \Storage[10][0] ,
         \Storage[9][32] , \Storage[9][31] , \Storage[9][30] ,
         \Storage[9][29] , \Storage[9][28] , \Storage[9][27] ,
         \Storage[9][26] , \Storage[9][25] , \Storage[9][24] ,
         \Storage[9][23] , \Storage[9][22] , \Storage[9][21] ,
         \Storage[9][20] , \Storage[9][19] , \Storage[9][18] ,
         \Storage[9][17] , \Storage[9][16] , \Storage[9][15] ,
         \Storage[9][14] , \Storage[9][13] , \Storage[9][12] ,
         \Storage[9][11] , \Storage[9][10] , \Storage[9][9] , \Storage[9][8] ,
         \Storage[9][7] , \Storage[9][6] , \Storage[9][5] , \Storage[9][4] ,
         \Storage[9][3] , \Storage[9][2] , \Storage[9][1] , \Storage[9][0] ,
         \Storage[8][32] , \Storage[8][31] , \Storage[8][30] ,
         \Storage[8][29] , \Storage[8][28] , \Storage[8][27] ,
         \Storage[8][26] , \Storage[8][25] , \Storage[8][24] ,
         \Storage[8][23] , \Storage[8][22] , \Storage[8][21] ,
         \Storage[8][20] , \Storage[8][19] , \Storage[8][18] ,
         \Storage[8][17] , \Storage[8][16] , \Storage[8][15] ,
         \Storage[8][14] , \Storage[8][13] , \Storage[8][12] ,
         \Storage[8][11] , \Storage[8][10] , \Storage[8][9] , \Storage[8][8] ,
         \Storage[8][7] , \Storage[8][6] , \Storage[8][5] , \Storage[8][4] ,
         \Storage[8][3] , \Storage[8][2] , \Storage[8][1] , \Storage[8][0] ,
         \Storage[7][32] , \Storage[7][31] , \Storage[7][30] ,
         \Storage[7][29] , \Storage[7][28] , \Storage[7][27] ,
         \Storage[7][26] , \Storage[7][25] , \Storage[7][24] ,
         \Storage[7][23] , \Storage[7][22] , \Storage[7][21] ,
         \Storage[7][20] , \Storage[7][19] , \Storage[7][18] ,
         \Storage[7][17] , \Storage[7][16] , \Storage[7][15] ,
         \Storage[7][14] , \Storage[7][13] , \Storage[7][12] ,
         \Storage[7][11] , \Storage[7][10] , \Storage[7][9] , \Storage[7][8] ,
         \Storage[7][7] , \Storage[7][6] , \Storage[7][5] , \Storage[7][4] ,
         \Storage[7][3] , \Storage[7][2] , \Storage[7][1] , \Storage[7][0] ,
         \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899;
  wire   [31:0] DataOr;
  assign N79 = AddrR[0];
  assign N80 = AddrR[1];
  assign N81 = AddrR[2];
  assign N82 = AddrR[3];
  assign N83 = AddrR[4];

  XNR4D1 U25 ( .A1(n884), .A2(n882), .A3(n888), .A4(n886), .ZN(n88) );
  XOR4D1 U26 ( .A1(n892), .A2(n890), .A3(n896), .A4(n894), .Z(n87) );
  XOR4D1 U27 ( .A1(n874), .A2(n872), .A3(n898), .A4(n876), .Z(n84) );
  XOR4D1 U28 ( .A1(n864), .A2(n862), .A3(DataI[22]), .A4(n878), .Z(n81) );
  XNR4D1 U29 ( .A1(n850), .A2(n842), .A3(DataI[9]), .A4(n852), .ZN(n78) );
  XOR4D1 U33 ( .A1(n41), .A2(n157), .A3(n94), .A4(n133), .Z(n92) );
  XNR4D1 U34 ( .A1(n181), .A2(n189), .A3(n165), .A4(n173), .ZN(n94) );
  XNR4D1 U39 ( .A1(n54), .A2(N32), .A3(n113), .A4(n58), .ZN(n100) );
  XOR4D1 U40 ( .A1(n129), .A2(n117), .A3(n145), .A4(n137), .Z(n99) );
  XNR4D1 U41 ( .A1(n185), .A2(n177), .A3(n201), .A4(n193), .ZN(n96) );
  XNR4D1 U42 ( .A1(n50), .A2(n109), .A3(n46), .A4(n42), .ZN(n90) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n830), .E(n713), .CP(n781), .CDN(n661), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(n713), .CP(n781), .CDN(
        n660), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(n712), .CP(n781), .CDN(
        n660), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(n713), .CP(n781), .CDN(
        n660), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(n712), .CP(n782), .CDN(
        n660), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(n890), .E(n713), .CP(n782), .CDN(n660), 
        .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(n712), .CP(n782), .CDN(
        n660), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(n713), .CP(n782), .CDN(
        n660), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(n712), .CP(n782), .CDN(
        n660), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(n882), .E(n713), .CP(n782), .CDN(n660), 
        .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(n712), .CP(n782), .CDN(
        n660), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(n712), .CP(n782), .CDN(
        n660), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(n712), .CP(n782), .CDN(
        n659), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(n712), .CP(n782), .CDN(
        n659), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(n872), .E(n712), .CP(n783), .CDN(n659), 
        .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(n712), .CP(n783), .CDN(
        n659), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(n712), .CP(n783), .CDN(
        n659), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(n712), .CP(n783), .CDN(
        n659), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(n712), .CP(n783), .CDN(
        n659), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(n862), .E(n712), .CP(n783), .CDN(n659), 
        .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(n713), .CP(n783), .CDN(
        n659), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(n713), .CP(n783), .CDN(
        n659), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(n713), .CP(n783), .CDN(
        n659), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(n713), .CP(n783), .CDN(n658), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(n713), .CP(n784), .CDN(n658), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(n713), .CP(n784), .CDN(n658), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(DataI[6]), .E(n713), .CP(n784), .CDN(n658), .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(DataI[5]), .E(n713), .CP(n784), .CDN(n658), .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(n713), .CP(n784), .CDN(n658), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(n842), .E(n713), .CP(n784), .CDN(n658), 
        .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(n712), .CP(n784), .CDN(n658), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(n712), .CP(n784), .CDN(n658), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(n836), .E(n713), .CP(n784), .CDN(n658), 
        .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n829), .E(n721), .CP(n794), .CDN(n649), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(n721), .CP(n794), .CDN(
        n648), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(DataI[30]), .E(n720), .CP(n795), .CDN(
        n648), .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(n721), .CP(n795), .CDN(
        n648), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(n720), .CP(n795), .CDN(
        n648), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(n721), .CP(n795), .CDN(
        n648), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(DataI[26]), .E(n720), .CP(n795), .CDN(
        n648), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(DataI[25]), .E(n721), .CP(n795), .CDN(
        n648), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(n720), .CP(n795), .CDN(
        n648), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(n721), .CP(n795), .CDN(
        n648), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n880), .E(n720), .CP(n795), .CDN(n648), 
        .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(DataI[21]), .E(n720), .CP(n795), .CDN(
        n648), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(DataI[18]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(DataI[14]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(n720), .CP(n796), .CDN(
        n647), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n860), .E(n721), .CP(n796), .CDN(n647), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(DataI[11]), .E(n721), .CP(n796), .CDN(
        n647), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(n721), .CP(n797), .CDN(
        n647), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n854), .E(n721), .CP(n797), .CDN(n646), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(DataI[8]), .E(n721), .CP(n797), .CDN(n646), .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(n721), .CP(n797), .CDN(n646), .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n848), .E(n721), .CP(n797), .CDN(n646), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(DataI[5]), .E(n721), .CP(n797), .CDN(n646), .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n844), .E(n721), .CP(n797), .CDN(n646), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(n721), .CP(n797), .CDN(n646), .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n840), .E(n720), .CP(n797), .CDN(n646), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(n720), .CP(n797), .CDN(n646), .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n836), .E(n721), .CP(n798), .CDN(n646), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(n829), .E(n729), .CP(n805), .CDN(n638), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n898), .E(n729), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n896), .E(n728), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n894), .E(n729), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n892), .E(n728), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(n729), .CP(n805), .CDN(
        n637), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n888), .E(n728), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n886), .E(n729), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n884), .E(n728), .CP(n805), .CDN(n637), 
        .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(n729), .CP(n805), .CDN(
        n637), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n880), .E(n728), .CP(n806), .CDN(n637), 
        .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n878), .E(n728), .CP(n806), .CDN(n637), 
        .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n876), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n874), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(n728), .CP(n806), .CDN(
        n636), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n870), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n868), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n866), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n864), .E(n728), .CP(n806), .CDN(n636), 
        .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(DataI[13]), .E(n728), .CP(n806), .CDN(
        n636), .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n860), .E(n729), .CP(n816), .CDN(n636), 
        .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n858), .E(n729), .CP(n783), .CDN(n636), 
        .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n856), .E(n729), .CP(n774), .CDN(n636), 
        .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n854), .E(n729), .CP(n823), .CDN(n635), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n852), .E(n729), .CP(n819), .CDN(n635), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n850), .E(n729), .CP(n825), .CDN(n635), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n848), .E(n729), .CP(n826), .CDN(n635), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n846), .E(n729), .CP(n824), .CDN(n635), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n844), .E(n729), .CP(n807), .CDN(n635), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(DataI[3]), .E(n729), .CP(n793), .CDN(n635), .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n840), .E(n728), .CP(n809), .CDN(n635), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n838), .E(n728), .CP(n819), .CDN(n635), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n836), .E(n729), .CP(n824), .CDN(n635), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n829), .E(n737), .CP(ClockW), .CDN(n627), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n898), .E(n737), .CP(n785), .CDN(n626), 
        .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n896), .E(n736), .CP(n773), .CDN(n626), 
        .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(DataI[29]), .E(n737), .CP(n816), .CDN(
        n626), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(DataI[28]), .E(n736), .CP(n815), .CDN(
        n626), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n890), .E(n737), .CP(n814), .CDN(n626), 
        .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n888), .E(n736), .CP(n811), .CDN(n626), 
        .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(DataI[25]), .E(n737), .CP(n812), .CDN(
        n626), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(DataI[24]), .E(n736), .CP(n804), .CDN(
        n626), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n882), .E(n737), .CP(n808), .CDN(n626), 
        .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n880), .E(n736), .CP(n807), .CDN(n626), 
        .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(DataI[21]), .E(n736), .CP(n811), .CDN(
        n626), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(DataI[20]), .E(n736), .CP(n819), .CDN(
        n625), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(DataI[19]), .E(n736), .CP(n818), .CDN(
        n625), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n872), .E(n736), .CP(n817), .CDN(n625), 
        .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n870), .E(n736), .CP(n820), .CDN(n625), 
        .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(DataI[16]), .E(n736), .CP(n822), .CDN(
        n625), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(DataI[15]), .E(n736), .CP(n803), .CDN(
        n625), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(DataI[14]), .E(n736), .CP(n792), .CDN(
        n625), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n862), .E(n736), .CP(n826), .CDN(n625), 
        .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n860), .E(n737), .CP(n775), .CDN(n625), 
        .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(DataI[11]), .E(n737), .CP(n776), .CDN(
        n625), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(DataI[10]), .E(n737), .CP(n817), .CDN(
        n625), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n854), .E(n737), .CP(n787), .CDN(n624), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(DataI[8]), .E(n737), .CP(n802), .CDN(n624), .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(DataI[7]), .E(n737), .CP(ClockW), .CDN(
        n624), .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n848), .E(n737), .CP(n783), .CDN(n624), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(DataI[5]), .E(n737), .CP(n790), .CDN(n624), .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n844), .E(n737), .CP(n798), .CDN(n624), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n842), .E(n737), .CP(n787), .CDN(n624), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n840), .E(n736), .CP(n788), .CDN(n624), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(DataI[1]), .E(n736), .CP(n789), .CDN(n624), .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n836), .E(n737), .CP(n790), .CDN(n624), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n829), .E(n745), .CP(n796), .CDN(n615), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(n745), .CP(n779), .CDN(
        n614), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(n744), .CP(n780), .CDN(
        n614), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n745), .CP(n775), .CDN(
        n614), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(n744), .CP(n776), .CDN(
        n614), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(n745), .CP(n774), .CDN(
        n614), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(n744), .CP(n811), .CDN(
        n614), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(n745), .CP(n822), .CDN(
        n614), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(n744), .CP(n820), .CDN(
        n614), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(n745), .CP(n801), .CDN(
        n614), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n880), .E(n744), .CP(n800), .CDN(n614), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(n744), .CP(n807), .CDN(
        n614), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n744), .CP(n791), .CDN(
        n613), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(n744), .CP(n806), .CDN(
        n613), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(n744), .CP(n777), .CDN(
        n613), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n744), .CP(ClockW), .CDN(
        n613), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(n744), .CP(n785), .CDN(
        n613), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n744), .CP(n818), .CDN(
        n613), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(n744), .CP(n819), .CDN(
        n613), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(n744), .CP(n810), .CDN(
        n613), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n860), .E(n745), .CP(n807), .CDN(n613), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(n745), .CP(n808), .CDN(
        n613), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n745), .CP(n825), .CDN(
        n613), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n854), .E(n745), .CP(n781), .CDN(n612), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(n745), .CP(ClockW), .CDN(
        n612), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(n745), .CP(n822), .CDN(n612), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n848), .E(n745), .CP(n817), .CDN(n612), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(n745), .CP(n811), .CDN(n612), .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n844), .E(n745), .CP(n810), .CDN(n612), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(n745), .CP(n809), .CDN(n612), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n840), .E(n744), .CP(n783), .CDN(n612), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n744), .CP(n808), .CDN(n612), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n836), .E(n745), .CP(n807), .CDN(n612), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n830), .E(n753), .CP(n812), .CDN(n603), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n898), .E(n753), .CP(n785), .CDN(n595), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n896), .E(n752), .CP(n789), .CDN(n602), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n894), .E(n753), .CP(n781), .CDN(n668), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n892), .E(n752), .CP(n773), .CDN(n586), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n890), .E(n753), .CP(n772), .CDN(n587), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n888), .E(n752), .CP(ClockW), .CDN(n598), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n886), .E(n753), .CP(n786), .CDN(n599), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n884), .E(n752), .CP(n797), .CDN(n602), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n882), .E(n753), .CP(n805), .CDN(n668), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n752), .CP(n812), .CDN(
        n592), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n878), .E(n752), .CP(n789), .CDN(n586), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n876), .E(n752), .CP(n802), .CDN(n602), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n874), .E(n752), .CP(n805), .CDN(n602), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n872), .E(n752), .CP(n824), .CDN(n602), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n870), .E(n752), .CP(n813), .CDN(n602), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n868), .E(n752), .CP(n809), .CDN(n602), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n866), .E(n752), .CP(n773), .CDN(n602), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n864), .E(n752), .CP(n808), .CDN(n602), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n862), .E(n752), .CP(n807), .CDN(n602), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n753), .CP(n772), .CDN(
        n602), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n858), .E(n753), .CP(n817), .CDN(n602), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n856), .E(n753), .CP(n783), .CDN(n602), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(n753), .CP(n819), .CDN(n601), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n852), .E(n753), .CP(n823), .CDN(n601), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n850), .E(n753), .CP(n774), .CDN(n601), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(n753), .CP(n776), .CDN(n601), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n846), .E(n753), .CP(n819), .CDN(n601), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n753), .CP(n779), .CDN(n601), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n842), .E(n753), .CP(n806), .CDN(n601), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(n752), .CP(n787), .CDN(n601), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n838), .E(n752), .CP(n781), .CDN(n601), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n753), .CP(n826), .CDN(n601), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n830), .E(n761), .CP(n802), .CDN(n592), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n898), .E(n761), .CP(n795), .CDN(n591), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n896), .E(n760), .CP(n797), .CDN(n591), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n894), .E(n761), .CP(n820), .CDN(n591), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n892), .E(n760), .CP(n798), .CDN(n591), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n890), .E(n761), .CP(n820), .CDN(n591), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n888), .E(n760), .CP(n819), .CDN(n591), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n886), .E(n761), .CP(n795), .CDN(n591), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n884), .E(n760), .CP(n812), .CDN(n591), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n882), .E(n761), .CP(n800), .CDN(n591), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n760), .CP(n823), .CDN(
        n591), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n878), .E(n760), .CP(n818), .CDN(n591), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n876), .E(n760), .CP(ClockW), .CDN(n590), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n874), .E(n760), .CP(n790), .CDN(n590), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n872), .E(n760), .CP(n804), .CDN(n590), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n870), .E(n760), .CP(n809), .CDN(n590), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n868), .E(n760), .CP(n788), .CDN(n590), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n866), .E(n760), .CP(n812), .CDN(n590), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n864), .E(n760), .CP(n791), .CDN(n590), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n862), .E(n760), .CP(n819), .CDN(n590), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n761), .CP(n809), .CDN(
        n590), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n858), .E(n761), .CP(n817), .CDN(n590), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n856), .E(n761), .CP(n826), .CDN(n590), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n761), .CP(n786), .CDN(n589), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n852), .E(n761), .CP(n808), .CDN(n589), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n850), .E(n761), .CP(n774), .CDN(n589), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n761), .CP(n823), .CDN(n589), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n846), .E(n761), .CP(n824), .CDN(n589), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n761), .CP(n825), .CDN(n589), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n842), .E(n761), .CP(n826), .CDN(n589), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n760), .CP(n825), .CDN(n589), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n838), .E(n760), .CP(n792), .CDN(n589), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n761), .CP(n772), .CDN(n589), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n830), .E(n769), .CP(n814), .CDN(n581), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n898), .E(n769), .CP(n812), .CDN(n580), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n896), .E(n768), .CP(n819), .CDN(n580), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n894), .E(n769), .CP(n818), .CDN(n580), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n892), .E(n768), .CP(n817), .CDN(n580), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n890), .E(n769), .CP(n822), .CDN(n580), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n888), .E(n768), .CP(n821), .CDN(n580), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n886), .E(n769), .CP(n820), .CDN(n580), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n884), .E(n768), .CP(n816), .CDN(n580), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n882), .E(n769), .CP(n815), .CDN(n580), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n768), .CP(n816), .CDN(
        n580), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n878), .E(n768), .CP(n773), .CDN(n580), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n876), .E(n768), .CP(n811), .CDN(n579), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n874), .E(n768), .CP(n781), .CDN(n579), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n872), .E(n768), .CP(n793), .CDN(n579), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n870), .E(n768), .CP(n813), .CDN(n579), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n868), .E(n768), .CP(n789), .CDN(n579), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n866), .E(n768), .CP(n800), .CDN(n579), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n864), .E(n768), .CP(n779), .CDN(n579), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n862), .E(n768), .CP(n776), .CDN(n579), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n769), .CP(n798), .CDN(
        n579), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n858), .E(n769), .CP(n808), .CDN(n579), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n856), .E(n769), .CP(n772), .CDN(n579), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n769), .CP(n778), .CDN(n578), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n852), .E(n769), .CP(n797), .CDN(n578), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n850), .E(n769), .CP(n773), .CDN(n578), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n769), .CP(n799), .CDN(n578), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n846), .E(n769), .CP(n809), .CDN(n578), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n769), .CP(n786), .CDN(n578), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n842), .E(n769), .CP(n773), .CDN(n578), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n768), .CP(n823), .CDN(n578), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n838), .E(n768), .CP(ClockW), .CDN(n578), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n769), .CP(n821), .CDN(n578), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n829), .E(n709), .CP(n775), .CDN(n667), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(n709), .CP(n775), .CDN(
        n666), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(n708), .CP(n775), .CDN(
        n666), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(n709), .CP(n775), .CDN(
        n666), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(n708), .CP(n775), .CDN(
        n666), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(n709), .CP(n775), .CDN(
        n666), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(n708), .CP(n775), .CDN(
        n666), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(n709), .CP(n775), .CDN(
        n666), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(n708), .CP(n775), .CDN(
        n666), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(n709), .CP(n775), .CDN(
        n666), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(n880), .E(n708), .CP(n776), .CDN(n666), 
        .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(n708), .CP(n776), .CDN(
        n666), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(n708), .CP(n776), .CDN(
        n665), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(n860), .E(n709), .CP(n777), .CDN(n665), 
        .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(n709), .CP(n777), .CDN(
        n665), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(n709), .CP(n777), .CDN(
        n665), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(n854), .E(n709), .CP(n777), .CDN(n664), 
        .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(n709), .CP(n777), .CDN(n664), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(n709), .CP(n777), .CDN(n664), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n848), .E(n709), .CP(n777), .CDN(n664), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(n709), .CP(n777), .CDN(n664), .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(n844), .E(n709), .CP(n777), .CDN(n664), 
        .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(n709), .CP(n777), .CDN(n664), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(n840), .E(n708), .CP(n778), .CDN(n664), 
        .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(n708), .CP(n778), .CDN(n664), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(n836), .E(n709), .CP(n778), .CDN(n664), 
        .Q(\Storage[31][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(n829), .E(n711), .CP(n778), .CDN(n664), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(n711), .CP(n778), .CDN(
        n663), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n710), .CP(n778), .CDN(
        n663), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(n711), .CP(n778), .CDN(
        n663), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(n710), .CP(n778), .CDN(
        n663), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(n711), .CP(n778), .CDN(
        n663), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n710), .CP(n778), .CDN(
        n663), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n711), .CP(n779), .CDN(
        n663), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(n710), .CP(n779), .CDN(
        n663), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(n711), .CP(n779), .CDN(
        n663), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(n880), .E(n710), .CP(n779), .CDN(n663), 
        .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n710), .CP(n779), .CDN(
        n663), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(n710), .CP(n779), .CDN(
        n662), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(n710), .CP(n779), .CDN(
        n662), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n710), .CP(n779), .CDN(
        n662), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(n710), .CP(n779), .CDN(
        n662), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(n710), .CP(n779), .CDN(
        n662), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(n710), .CP(n780), .CDN(
        n662), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n710), .CP(n780), .CDN(
        n662), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(n710), .CP(n780), .CDN(
        n662), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(n860), .E(n711), .CP(n780), .CDN(n662), 
        .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n711), .CP(n780), .CDN(
        n662), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(n711), .CP(n780), .CDN(
        n662), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(n854), .E(n711), .CP(n780), .CDN(n661), 
        .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n711), .CP(n780), .CDN(n661), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(n711), .CP(n780), .CDN(n661), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n848), .E(n711), .CP(n780), .CDN(n661), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(DataI[5]), .E(n711), .CP(n781), .CDN(n661), .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(n844), .E(n711), .CP(n781), .CDN(n661), 
        .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(n711), .CP(n781), .CDN(n661), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(n840), .E(n710), .CP(n781), .CDN(n661), 
        .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(n710), .CP(n781), .CDN(n661), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(n836), .E(n711), .CP(n781), .CDN(n661), 
        .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(n830), .E(n715), .CP(n784), .CDN(n658), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(n715), .CP(n785), .CDN(
        n657), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(DataI[30]), .E(n714), .CP(n785), .CDN(
        n657), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(DataI[29]), .E(n715), .CP(n785), .CDN(
        n657), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(n714), .CP(n785), .CDN(
        n657), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(n715), .CP(n785), .CDN(
        n657), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(DataI[26]), .E(n714), .CP(n785), .CDN(
        n657), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(DataI[25]), .E(n715), .CP(n785), .CDN(
        n657), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(n714), .CP(n785), .CDN(
        n657), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(n715), .CP(n785), .CDN(
        n657), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n880), .E(n714), .CP(n785), .CDN(n657), 
        .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(DataI[21]), .E(n714), .CP(n786), .CDN(
        n657), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(DataI[18]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(DataI[17]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(DataI[15]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(DataI[14]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(n714), .CP(n786), .CDN(
        n656), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n860), .E(n715), .CP(n786), .CDN(n656), 
        .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(DataI[11]), .E(n715), .CP(n787), .CDN(
        n656), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(DataI[10]), .E(n715), .CP(n787), .CDN(
        n656), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n854), .E(n715), .CP(n787), .CDN(n655), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(DataI[8]), .E(n715), .CP(n787), .CDN(n655), .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(DataI[7]), .E(n715), .CP(n787), .CDN(n655), .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n848), .E(n715), .CP(n787), .CDN(n655), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(DataI[5]), .E(n715), .CP(n787), .CDN(n655), .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n844), .E(n715), .CP(n787), .CDN(n655), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(DataI[3]), .E(n715), .CP(n787), .CDN(n655), .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n840), .E(n714), .CP(n787), .CDN(n655), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(DataI[1]), .E(n714), .CP(n788), .CDN(n655), .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n836), .E(n715), .CP(n788), .CDN(n655), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n829), .E(n717), .CP(n788), .CDN(n655), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(n717), .CP(n788), .CDN(
        n654), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(n716), .CP(n788), .CDN(
        n654), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(DataI[29]), .E(n717), .CP(n788), .CDN(
        n654), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(n716), .CP(n788), .CDN(
        n654), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(n717), .CP(n788), .CDN(
        n654), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(n716), .CP(n788), .CDN(
        n654), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(n717), .CP(n788), .CDN(
        n654), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(n716), .CP(n789), .CDN(
        n654), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(n717), .CP(n789), .CDN(
        n654), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n880), .E(n716), .CP(n789), .CDN(n654), 
        .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(n716), .CP(n789), .CDN(
        n654), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(DataI[17]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(DataI[15]), .E(n716), .CP(n789), .CDN(
        n653), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(DataI[14]), .E(n716), .CP(n790), .CDN(
        n653), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(n716), .CP(n790), .CDN(
        n653), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n860), .E(n717), .CP(n790), .CDN(n653), 
        .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(n717), .CP(n790), .CDN(
        n653), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(DataI[10]), .E(n717), .CP(n790), .CDN(
        n653), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n854), .E(n717), .CP(n790), .CDN(n652), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(n717), .CP(n790), .CDN(n652), .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(DataI[7]), .E(n717), .CP(n790), .CDN(n652), .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n848), .E(n717), .CP(n790), .CDN(n652), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(n717), .CP(n790), .CDN(n652), .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n844), .E(n717), .CP(n791), .CDN(n652), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(DataI[3]), .E(n717), .CP(n791), .CDN(n652), .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n840), .E(n716), .CP(n791), .CDN(n652), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(DataI[1]), .E(n716), .CP(n791), .CDN(n652), .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n836), .E(n717), .CP(n791), .CDN(n652), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(n830), .E(n719), .CP(n791), .CDN(n652), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(n719), .CP(n791), .CDN(
        n651), .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(DataI[30]), .E(n718), .CP(n791), .CDN(
        n651), .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(DataI[29]), .E(n719), .CP(n791), .CDN(
        n651), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(n718), .CP(n791), .CDN(
        n651), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(n719), .CP(n792), .CDN(
        n651), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(DataI[26]), .E(n718), .CP(n792), .CDN(
        n651), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(DataI[25]), .E(n719), .CP(n792), .CDN(
        n651), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(n718), .CP(n792), .CDN(
        n651), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(n719), .CP(n792), .CDN(
        n651), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n880), .E(n718), .CP(n792), .CDN(n651), 
        .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(DataI[21]), .E(n718), .CP(n792), .CDN(
        n651), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(n718), .CP(n792), .CDN(
        n650), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(n718), .CP(n792), .CDN(
        n650), .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(DataI[18]), .E(n718), .CP(n792), .CDN(
        n650), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(DataI[17]), .E(n718), .CP(n793), .CDN(
        n650), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(n718), .CP(n793), .CDN(
        n650), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(DataI[15]), .E(n718), .CP(n793), .CDN(
        n650), .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(DataI[14]), .E(n718), .CP(n793), .CDN(
        n650), .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(n718), .CP(n793), .CDN(
        n650), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n860), .E(n719), .CP(n793), .CDN(n650), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(DataI[11]), .E(n719), .CP(n793), .CDN(
        n650), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(DataI[10]), .E(n719), .CP(n793), .CDN(
        n650), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n854), .E(n719), .CP(n793), .CDN(n649), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(DataI[8]), .E(n719), .CP(n793), .CDN(n649), .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(DataI[7]), .E(n719), .CP(n794), .CDN(n649), .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n848), .E(n719), .CP(n794), .CDN(n649), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(DataI[5]), .E(n719), .CP(n794), .CDN(n649), .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n844), .E(n719), .CP(n794), .CDN(n649), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(DataI[3]), .E(n719), .CP(n794), .CDN(n649), .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n840), .E(n718), .CP(n794), .CDN(n649), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(n718), .CP(n794), .CDN(n649), .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n836), .E(n719), .CP(n794), .CDN(n649), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(n829), .E(n723), .CP(n798), .CDN(n646), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(DataI[31]), .E(n723), .CP(n798), .CDN(
        n645), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(DataI[30]), .E(n722), .CP(n798), .CDN(
        n645), .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(DataI[29]), .E(n723), .CP(n798), .CDN(
        n645), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(DataI[28]), .E(n722), .CP(n798), .CDN(
        n645), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(DataI[27]), .E(n723), .CP(n798), .CDN(
        n645), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(DataI[26]), .E(n722), .CP(n798), .CDN(
        n645), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(DataI[25]), .E(n723), .CP(n798), .CDN(
        n645), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(DataI[24]), .E(n722), .CP(n798), .CDN(
        n645), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(DataI[23]), .E(n723), .CP(n799), .CDN(
        n645), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n880), .E(n722), .CP(n799), .CDN(n645), 
        .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(DataI[21]), .E(n722), .CP(n799), .CDN(
        n645), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(DataI[20]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(DataI[19]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(DataI[18]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(DataI[17]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(DataI[16]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(DataI[15]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(DataI[14]), .E(n722), .CP(n799), .CDN(
        n644), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(DataI[13]), .E(n722), .CP(n800), .CDN(
        n644), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n860), .E(n723), .CP(n800), .CDN(n644), 
        .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(DataI[11]), .E(n723), .CP(n800), .CDN(
        n644), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(DataI[10]), .E(n723), .CP(n800), .CDN(
        n644), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n854), .E(n723), .CP(n800), .CDN(n643), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(DataI[8]), .E(n723), .CP(n800), .CDN(n643), .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(DataI[7]), .E(n723), .CP(n800), .CDN(n643), .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n848), .E(n723), .CP(n800), .CDN(n643), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(DataI[5]), .E(n723), .CP(n800), .CDN(n643), .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n844), .E(n723), .CP(n800), .CDN(n643), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(DataI[3]), .E(n723), .CP(n801), .CDN(n643), .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n840), .E(n722), .CP(n801), .CDN(n643), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(DataI[1]), .E(n722), .CP(n801), .CDN(n643), .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n836), .E(n723), .CP(n801), .CDN(n643), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n830), .E(n725), .CP(n801), .CDN(n643), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(DataI[31]), .E(n725), .CP(n801), .CDN(
        n642), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(DataI[30]), .E(n724), .CP(n801), .CDN(
        n642), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(DataI[29]), .E(n725), .CP(n801), .CDN(
        n642), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(DataI[28]), .E(n724), .CP(n801), .CDN(
        n642), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(DataI[27]), .E(n725), .CP(n801), .CDN(
        n642), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(DataI[26]), .E(n724), .CP(n802), .CDN(
        n642), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(DataI[25]), .E(n725), .CP(n802), .CDN(
        n642), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(DataI[24]), .E(n724), .CP(n802), .CDN(
        n642), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(DataI[23]), .E(n725), .CP(n802), .CDN(
        n642), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n880), .E(n724), .CP(n802), .CDN(n642), 
        .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(DataI[21]), .E(n724), .CP(n802), .CDN(
        n642), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(DataI[20]), .E(n724), .CP(n802), .CDN(
        n641), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(DataI[19]), .E(n724), .CP(n802), .CDN(
        n641), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(DataI[18]), .E(n724), .CP(n802), .CDN(
        n641), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(DataI[17]), .E(n724), .CP(n802), .CDN(
        n641), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(DataI[16]), .E(n724), .CP(n803), .CDN(
        n641), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(DataI[15]), .E(n724), .CP(n803), .CDN(
        n641), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(DataI[14]), .E(n724), .CP(n803), .CDN(
        n641), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(DataI[13]), .E(n724), .CP(n803), .CDN(
        n641), .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n860), .E(n725), .CP(n803), .CDN(n641), 
        .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(DataI[11]), .E(n725), .CP(n803), .CDN(
        n641), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(DataI[10]), .E(n725), .CP(n803), .CDN(
        n641), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n854), .E(n725), .CP(n803), .CDN(n640), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(DataI[8]), .E(n725), .CP(n803), .CDN(n640), .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(DataI[7]), .E(n725), .CP(n803), .CDN(n640), .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n848), .E(n725), .CP(n781), .CDN(n640), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(DataI[5]), .E(n725), .CP(n820), .CDN(n640), .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n844), .E(n725), .CP(n808), .CDN(n640), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(DataI[3]), .E(n725), .CP(n818), .CDN(n640), .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n840), .E(n724), .CP(n807), .CDN(n640), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(DataI[1]), .E(n724), .CP(n813), .CDN(n640), .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n836), .E(n725), .CP(n811), .CDN(n640), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(n829), .E(n727), .CP(n814), .CDN(n640), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n898), .E(n727), .CP(ClockW), .CDN(n639), 
        .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n896), .E(n726), .CP(n779), .CDN(n639), 
        .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(DataI[29]), .E(n727), .CP(n799), .CDN(
        n639), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(DataI[28]), .E(n726), .CP(n800), .CDN(
        n639), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(DataI[27]), .E(n727), .CP(n801), .CDN(
        n639), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n888), .E(n726), .CP(n802), .CDN(n639), 
        .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(DataI[25]), .E(n727), .CP(n810), .CDN(
        n639), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(DataI[24]), .E(n726), .CP(n812), .CDN(
        n639), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(DataI[23]), .E(n727), .CP(n811), .CDN(
        n639), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(DataI[22]), .E(n726), .CP(n815), .CDN(
        n639), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(DataI[21]), .E(n726), .CP(n816), .CDN(
        n639), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(DataI[20]), .E(n726), .CP(n814), .CDN(
        n609), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(DataI[19]), .E(n726), .CP(n800), .CDN(
        n668), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(DataI[18]), .E(n726), .CP(n793), .CDN(
        n668), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n870), .E(n726), .CP(n794), .CDN(n668), 
        .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(DataI[16]), .E(n726), .CP(n795), .CDN(
        n668), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(DataI[15]), .E(n726), .CP(n796), .CDN(
        n668), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(DataI[14]), .E(n726), .CP(n797), .CDN(
        n668), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(DataI[13]), .E(n726), .CP(n798), .CDN(
        n668), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(DataI[12]), .E(n727), .CP(n806), .CDN(
        n610), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(DataI[11]), .E(n727), .CP(n790), .CDN(
        n613), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(DataI[10]), .E(n727), .CP(n787), .CDN(
        n614), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(DataI[9]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(DataI[8]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(DataI[7]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(DataI[6]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(DataI[5]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(DataI[4]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(DataI[3]), .E(n727), .CP(n804), .CDN(n638), .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(DataI[2]), .E(n726), .CP(n804), .CDN(n638), .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(DataI[1]), .E(n726), .CP(n804), .CDN(n638), .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n836), .E(n727), .CP(n804), .CDN(n638), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(n829), .E(n731), .CP(n778), .CDN(n635), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(n731), .CP(n823), .CDN(
        n634), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(n730), .CP(n818), .CDN(
        n634), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(DataI[29]), .E(n731), .CP(n772), .CDN(
        n634), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(n730), .CP(n773), .CDN(
        n634), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(n731), .CP(n816), .CDN(
        n634), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(n730), .CP(n815), .CDN(
        n634), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(n731), .CP(n792), .CDN(
        n634), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(n730), .CP(n805), .CDN(
        n634), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(n731), .CP(n806), .CDN(
        n634), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n880), .E(n730), .CP(n814), .CDN(n634), 
        .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(n730), .CP(n807), .CDN(
        n634), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(DataI[20]), .E(n730), .CP(n808), .CDN(
        n633), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(n730), .CP(n820), .CDN(
        n633), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(n730), .CP(n821), .CDN(
        n633), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(DataI[17]), .E(n730), .CP(n822), .CDN(
        n633), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(n730), .CP(n817), .CDN(
        n633), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(DataI[15]), .E(n730), .CP(n784), .CDN(
        n633), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(n730), .CP(n818), .CDN(
        n633), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(n730), .CP(n804), .CDN(
        n633), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n860), .E(n731), .CP(n802), .CDN(n633), 
        .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(n731), .CP(n785), .CDN(
        n633), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(DataI[10]), .E(n731), .CP(n779), .CDN(
        n633), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n854), .E(n731), .CP(n780), .CDN(n632), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(n731), .CP(n777), .CDN(n632), .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(DataI[7]), .E(n731), .CP(n778), .CDN(n632), .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n848), .E(n731), .CP(n775), .CDN(n632), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(DataI[5]), .E(n731), .CP(n802), .CDN(n632), .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n844), .E(n731), .CP(n799), .CDN(n632), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(DataI[3]), .E(n731), .CP(n800), .CDN(n632), .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n840), .E(n730), .CP(n799), .CDN(n632), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(DataI[1]), .E(n730), .CP(n803), .CDN(n632), .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n836), .E(n731), .CP(n803), .CDN(n632), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(n829), .E(n733), .CP(n819), .CDN(n632), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(DataI[31]), .E(n733), .CP(n774), .CDN(
        n631), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(DataI[30]), .E(n732), .CP(n809), .CDN(
        n631), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(n733), .CP(n810), .CDN(
        n631), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(DataI[28]), .E(n732), .CP(n792), .CDN(
        n631), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(DataI[27]), .E(n733), .CP(n810), .CDN(
        n631), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(DataI[26]), .E(n732), .CP(n785), .CDN(
        n631), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(DataI[25]), .E(n733), .CP(n817), .CDN(
        n631), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(DataI[24]), .E(n732), .CP(n821), .CDN(
        n631), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(DataI[23]), .E(n733), .CP(n775), .CDN(
        n631), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n880), .E(n732), .CP(n797), .CDN(n631), 
        .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(DataI[21]), .E(n732), .CP(n780), .CDN(
        n631), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(n732), .CP(ClockW), .CDN(
        n630), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(DataI[19]), .E(n732), .CP(n786), .CDN(
        n630), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(DataI[18]), .E(n732), .CP(n776), .CDN(
        n630), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(n732), .CP(n791), .CDN(
        n630), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(DataI[16]), .E(n732), .CP(n794), .CDN(
        n630), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(n732), .CP(n793), .CDN(
        n630), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(DataI[14]), .E(n732), .CP(n796), .CDN(
        n630), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(DataI[13]), .E(n732), .CP(n795), .CDN(
        n630), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n860), .E(n733), .CP(n798), .CDN(n630), 
        .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(DataI[11]), .E(n733), .CP(n791), .CDN(
        n630), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(n733), .CP(n785), .CDN(
        n630), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n854), .E(n733), .CP(n799), .CDN(n629), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(DataI[8]), .E(n733), .CP(n820), .CDN(n629), .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(n733), .CP(n822), .CDN(n629), .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n848), .E(n733), .CP(n821), .CDN(n629), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(DataI[5]), .E(n733), .CP(n817), .CDN(n629), .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n844), .E(n733), .CP(n806), .CDN(n629), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(n733), .CP(n809), .CDN(n629), .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n840), .E(n732), .CP(n798), .CDN(n629), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(n732), .CP(n808), .CDN(n629), .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n836), .E(n733), .CP(n807), .CDN(n629), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(n829), .E(n735), .CP(n815), .CDN(n629), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(DataI[31]), .E(n735), .CP(n779), .CDN(
        n597), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(DataI[30]), .E(n734), .CP(n817), .CDN(
        n597), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(n735), .CP(n775), .CDN(
        n597), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(DataI[28]), .E(n734), .CP(n776), .CDN(
        n597), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(DataI[27]), .E(n735), .CP(n777), .CDN(
        n597), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(DataI[26]), .E(n734), .CP(n778), .CDN(
        n597), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(DataI[25]), .E(n735), .CP(n782), .CDN(
        n668), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(DataI[24]), .E(n734), .CP(n781), .CDN(
        n597), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(DataI[23]), .E(n735), .CP(n815), .CDN(
        n668), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n880), .E(n734), .CP(n810), .CDN(n597), 
        .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(DataI[21]), .E(n734), .CP(n782), .CDN(
        n668), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(n734), .CP(n786), .CDN(
        n628), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(DataI[19]), .E(n734), .CP(n811), .CDN(
        n628), .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(DataI[18]), .E(n734), .CP(n812), .CDN(
        n628), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(n734), .CP(n813), .CDN(
        n628), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(DataI[16]), .E(n734), .CP(n814), .CDN(
        n628), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(n734), .CP(n816), .CDN(
        n628), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(DataI[14]), .E(n734), .CP(n815), .CDN(
        n628), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(DataI[13]), .E(n734), .CP(n773), .CDN(
        n628), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n860), .E(n735), .CP(n823), .CDN(n628), 
        .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(DataI[11]), .E(n735), .CP(n794), .CDN(
        n628), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(n735), .CP(n793), .CDN(
        n628), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n854), .E(n735), .CP(n795), .CDN(n627), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(DataI[8]), .E(n735), .CP(n796), .CDN(n627), .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(n735), .CP(n798), .CDN(n627), .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n848), .E(n735), .CP(n797), .CDN(n627), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(DataI[5]), .E(n735), .CP(n787), .CDN(n627), .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n844), .E(n735), .CP(n788), .CDN(n627), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(n735), .CP(n789), .CDN(n627), .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n840), .E(n734), .CP(n790), .CDN(n627), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(n734), .CP(n813), .CDN(n627), .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n836), .E(n735), .CP(n804), .CDN(n627), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(n829), .E(n738), .CP(n791), .CDN(n624), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(DataI[31]), .E(n738), .CP(n792), .CDN(
        n623), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(DataI[30]), .E(n739), .CP(n793), .CDN(
        n623), .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(DataI[29]), .E(n738), .CP(n794), .CDN(
        n623), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(DataI[28]), .E(n739), .CP(n795), .CDN(
        n623), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(DataI[27]), .E(n738), .CP(n825), .CDN(
        n623), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(DataI[26]), .E(n739), .CP(n774), .CDN(
        n623), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(DataI[25]), .E(n738), .CP(n772), .CDN(
        n623), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(DataI[24]), .E(n739), .CP(n823), .CDN(
        n623), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(DataI[23]), .E(n738), .CP(n824), .CDN(
        n623), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n880), .E(n738), .CP(n820), .CDN(n623), 
        .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(DataI[21]), .E(n738), .CP(n826), .CDN(
        n623), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(DataI[20]), .E(n738), .CP(n816), .CDN(
        n622), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(DataI[19]), .E(n738), .CP(n815), .CDN(
        n622), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(DataI[18]), .E(n738), .CP(n773), .CDN(
        n622), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(DataI[17]), .E(n738), .CP(n786), .CDN(
        n622), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(DataI[16]), .E(n738), .CP(n787), .CDN(
        n622), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(DataI[15]), .E(n738), .CP(n788), .CDN(
        n622), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(DataI[14]), .E(n738), .CP(n789), .CDN(
        n622), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(DataI[13]), .E(n738), .CP(n790), .CDN(
        n622), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n860), .E(n739), .CP(n791), .CDN(n622), 
        .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(DataI[11]), .E(n739), .CP(n792), .CDN(
        n622), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(DataI[10]), .E(n739), .CP(n793), .CDN(
        n622), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n854), .E(n739), .CP(n794), .CDN(n621), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(DataI[8]), .E(n739), .CP(n795), .CDN(n621), .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(DataI[7]), .E(n739), .CP(n807), .CDN(n621), .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n848), .E(n739), .CP(n797), .CDN(n621), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(DataI[5]), .E(n739), .CP(n810), .CDN(n621), .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n844), .E(n739), .CP(n772), .CDN(n621), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(DataI[3]), .E(n739), .CP(n822), .CDN(n621), .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n840), .E(n739), .CP(n821), .CDN(n621), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(DataI[1]), .E(n739), .CP(n778), .CDN(n621), .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n836), .E(n738), .CP(n790), .CDN(n621), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n829), .E(n741), .CP(n781), .CDN(n621), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n741), .CP(n818), .CDN(
        n620), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(n740), .CP(n782), .CDN(
        n620), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(n741), .CP(n786), .CDN(
        n620), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(n740), .CP(n773), .CDN(
        n620), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(n741), .CP(n816), .CDN(
        n620), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(n740), .CP(n815), .CDN(
        n620), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(n741), .CP(n814), .CDN(
        n620), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(n740), .CP(n812), .CDN(
        n620), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(n741), .CP(n813), .CDN(
        n620), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n880), .E(n740), .CP(n819), .CDN(n620), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n740), .CP(n817), .CDN(
        n620), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(n740), .CP(n783), .CDN(
        n619), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n740), .CP(n820), .CDN(
        n619), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n740), .CP(n775), .CDN(
        n619), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(n740), .CP(n776), .CDN(
        n619), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n740), .CP(n813), .CDN(
        n619), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(n740), .CP(n787), .CDN(
        n619), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n740), .CP(n806), .CDN(
        n619), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n740), .CP(n779), .CDN(
        n619), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n860), .E(n741), .CP(n780), .CDN(n619), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n741), .CP(n781), .CDN(
        n619), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(n741), .CP(n809), .CDN(
        n619), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n854), .E(n741), .CP(n784), .CDN(n618), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(n741), .CP(n785), .CDN(n618), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(n741), .CP(n786), .CDN(n618), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n848), .E(n741), .CP(n799), .CDN(n618), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(n741), .CP(n800), .CDN(n618), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n844), .E(n741), .CP(n796), .CDN(n618), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(n741), .CP(n797), .CDN(n618), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n840), .E(n740), .CP(n822), .CDN(n618), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(n740), .CP(n797), .CDN(n618), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n836), .E(n741), .CP(n821), .CDN(n618), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n829), .E(n743), .CP(n805), .CDN(n618), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(n743), .CP(n804), .CDN(
        n617), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(n742), .CP(n803), .CDN(
        n617), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(n743), .CP(n779), .CDN(
        n617), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n742), .CP(n800), .CDN(
        n617), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n743), .CP(n799), .CDN(
        n617), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n742), .CP(n816), .CDN(
        n617), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(n743), .CP(n803), .CDN(
        n617), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n742), .CP(n802), .CDN(
        n617), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n743), .CP(n795), .CDN(
        n617), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n880), .E(n742), .CP(n806), .CDN(n617), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n742), .CP(n787), .CDN(
        n617), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(n742), .CP(n788), .CDN(
        n616), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n742), .CP(n789), .CDN(
        n616), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(n742), .CP(n790), .CDN(
        n616), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(n742), .CP(n791), .CDN(
        n616), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(n742), .CP(n792), .CDN(
        n616), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(n742), .CP(n793), .CDN(
        n616), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(n742), .CP(n794), .CDN(
        n616), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(n742), .CP(n814), .CDN(
        n616), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n860), .E(n743), .CP(n826), .CDN(n616), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n743), .CP(n801), .CDN(
        n616), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(n743), .CP(n789), .CDN(
        n616), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n854), .E(n743), .CP(n800), .CDN(n615), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n743), .CP(n772), .CDN(n615), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(n743), .CP(n791), .CDN(n615), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n848), .E(n743), .CP(n824), .CDN(n615), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(n743), .CP(n780), .CDN(n615), .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n844), .E(n743), .CP(n810), .CDN(n615), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(n743), .CP(n796), .CDN(n615), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n840), .E(n742), .CP(n817), .CDN(n615), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(n742), .CP(n777), .CDN(n615), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n836), .E(n743), .CP(n820), .CDN(n615), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(n829), .E(n747), .CP(n813), .CDN(n612), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(n747), .CP(n819), .CDN(
        n611), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(n746), .CP(n818), .CDN(
        n611), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n894), .E(n747), .CP(n802), .CDN(n611), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n892), .E(n746), .CP(n774), .CDN(n611), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(n747), .CP(n794), .CDN(
        n611), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(n746), .CP(n781), .CDN(
        n611), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n886), .E(n747), .CP(n792), .CDN(n611), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n884), .E(n746), .CP(ClockW), .CDN(n611), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(n747), .CP(n804), .CDN(
        n611), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n880), .E(n746), .CP(ClockW), .CDN(n611), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n878), .E(n746), .CP(n774), .CDN(n611), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n876), .E(n746), .CP(n798), .CDN(n610), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n874), .E(n746), .CP(n821), .CDN(n610), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(n746), .CP(n774), .CDN(
        n610), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(n746), .CP(n825), .CDN(
        n610), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n868), .E(n746), .CP(n826), .CDN(n610), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n866), .E(n746), .CP(n774), .CDN(n610), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n864), .E(n746), .CP(n794), .CDN(n610), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(n746), .CP(n824), .CDN(
        n610), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n860), .E(n747), .CP(n822), .CDN(n610), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n858), .E(n747), .CP(n772), .CDN(n610), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n856), .E(n747), .CP(n784), .CDN(n610), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n854), .E(n747), .CP(n811), .CDN(n609), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n852), .E(n747), .CP(n812), .CDN(n609), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n850), .E(n747), .CP(n818), .CDN(n609), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n848), .E(n747), .CP(n791), .CDN(n609), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n846), .E(n747), .CP(n823), .CDN(n609), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n844), .E(n747), .CP(n772), .CDN(n609), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(n747), .CP(n773), .CDN(n609), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n840), .E(n746), .CP(n814), .CDN(n609), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n838), .E(n746), .CP(n815), .CDN(n609), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(n747), .CP(n816), .CDN(n609), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n830), .E(n749), .CP(n783), .CDN(n609), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(n749), .CP(n784), .CDN(
        n608), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(n748), .CP(n784), .CDN(
        n608), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n894), .E(n749), .CP(n808), .CDN(n608), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n892), .E(n748), .CP(n799), .CDN(n608), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(n749), .CP(n824), .CDN(
        n608), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(n748), .CP(n805), .CDN(
        n608), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n886), .E(n749), .CP(n805), .CDN(n608), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n884), .E(n748), .CP(n801), .CDN(n608), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(n749), .CP(n824), .CDN(
        n608), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n880), .E(n748), .CP(n778), .CDN(n608), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n878), .E(n748), .CP(n803), .CDN(n608), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n876), .E(n748), .CP(ClockW), .CDN(n607), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n874), .E(n748), .CP(n782), .CDN(n607), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(n748), .CP(n781), .CDN(
        n607), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(n748), .CP(n784), .CDN(
        n607), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n868), .E(n748), .CP(n783), .CDN(n607), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n866), .E(n748), .CP(n786), .CDN(n607), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n864), .E(n748), .CP(n785), .CDN(n607), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(n748), .CP(n777), .CDN(
        n607), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n860), .E(n749), .CP(n826), .CDN(n607), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n858), .E(n749), .CP(n811), .CDN(n607), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n856), .E(n749), .CP(n784), .CDN(n607), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n854), .E(n749), .CP(n826), .CDN(n606), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n852), .E(n749), .CP(n820), .CDN(n606), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n850), .E(n749), .CP(n774), .CDN(n606), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n848), .E(n749), .CP(n823), .CDN(n606), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n846), .E(n749), .CP(n824), .CDN(n606), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n844), .E(n749), .CP(n825), .CDN(n606), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(n749), .CP(n826), .CDN(n606), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n840), .E(n748), .CP(ClockW), .CDN(n606), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n838), .E(n748), .CP(n816), .CDN(n606), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(n749), .CP(n782), .CDN(n606), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(n830), .E(n751), .CP(n780), .CDN(n606), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(n751), .CP(n775), .CDN(
        n605), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(n750), .CP(n788), .CDN(
        n605), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n894), .E(n751), .CP(n786), .CDN(n605), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n892), .E(n750), .CP(n788), .CDN(n605), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n890), .E(n751), .CP(n819), .CDN(n605), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(n750), .CP(n825), .CDN(
        n605), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n886), .E(n751), .CP(n815), .CDN(n605), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n884), .E(n750), .CP(n822), .CDN(n605), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n882), .E(n751), .CP(n821), .CDN(n605), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n880), .E(n750), .CP(n772), .CDN(n605), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n878), .E(n750), .CP(n822), .CDN(n605), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n876), .E(n750), .CP(n821), .CDN(n604), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n874), .E(n750), .CP(n820), .CDN(n604), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n872), .E(n750), .CP(n819), .CDN(n604), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(n750), .CP(n818), .CDN(
        n604), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n868), .E(n750), .CP(n817), .CDN(n604), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n866), .E(n750), .CP(n803), .CDN(n604), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n864), .E(n750), .CP(n825), .CDN(n604), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n862), .E(n750), .CP(n814), .CDN(n604), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n860), .E(n751), .CP(n813), .CDN(n604), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n858), .E(n751), .CP(n812), .CDN(n604), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n856), .E(n751), .CP(n811), .CDN(n604), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n854), .E(n751), .CP(n779), .CDN(n603), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n852), .E(n751), .CP(n782), .CDN(n603), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n850), .E(n751), .CP(n809), .CDN(n603), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n848), .E(n751), .CP(n801), .CDN(n603), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n846), .E(n751), .CP(n806), .CDN(n603), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n844), .E(n751), .CP(n773), .CDN(n603), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n842), .E(n751), .CP(n815), .CDN(n603), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n840), .E(n750), .CP(n816), .CDN(n603), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n838), .E(n750), .CP(n814), .CDN(n603), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(n751), .CP(n813), .CDN(n603), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(n830), .E(n755), .CP(n825), .CDN(n601), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n898), .E(n755), .CP(n825), .CDN(n600), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n896), .E(n754), .CP(n815), .CDN(n600), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n894), .E(n755), .CP(n772), .CDN(n600), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n892), .E(n754), .CP(n811), .CDN(n600), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n890), .E(n755), .CP(n821), .CDN(n600), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n888), .E(n754), .CP(n803), .CDN(n600), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n886), .E(n755), .CP(n822), .CDN(n600), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n884), .E(n754), .CP(n785), .CDN(n600), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n882), .E(n755), .CP(n818), .CDN(n600), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(n754), .CP(n807), .CDN(
        n600), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n878), .E(n754), .CP(n810), .CDN(n600), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n876), .E(n754), .CP(n816), .CDN(n599), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n874), .E(n754), .CP(n772), .CDN(n599), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n872), .E(n754), .CP(n773), .CDN(n599), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n870), .E(n754), .CP(n804), .CDN(n599), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n868), .E(n754), .CP(n780), .CDN(n599), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n866), .E(n754), .CP(n792), .CDN(n599), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n864), .E(n754), .CP(n825), .CDN(n599), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n862), .E(n754), .CP(n802), .CDN(n599), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n755), .CP(n798), .CDN(
        n599), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n858), .E(n755), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n856), .E(n755), .CP(n814), .CDN(n599), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(n755), .CP(n822), .CDN(n598), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n852), .E(n755), .CP(n821), .CDN(n598), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n850), .E(n755), .CP(n820), .CDN(n598), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(n755), .CP(n819), .CDN(n598), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n846), .E(n755), .CP(n818), .CDN(n598), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(n755), .CP(n817), .CDN(n598), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n842), .E(n755), .CP(n809), .CDN(n598), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(n754), .CP(n774), .CDN(n598), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n838), .E(n754), .CP(n799), .CDN(n598), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n755), .CP(n805), .CDN(n598), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n830), .E(n757), .CP(n818), .CDN(n598), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n898), .E(n757), .CP(n816), .CDN(n597), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n896), .E(n756), .CP(n815), .CDN(n597), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n894), .E(n757), .CP(n813), .CDN(n597), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n892), .E(n756), .CP(n812), .CDN(n597), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n890), .E(n757), .CP(n811), .CDN(n597), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n888), .E(n756), .CP(n783), .CDN(n597), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n886), .E(n757), .CP(n796), .CDN(n597), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n884), .E(n756), .CP(n782), .CDN(n597), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n882), .E(n757), .CP(n774), .CDN(n597), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n756), .CP(n776), .CDN(
        n597), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n878), .E(n756), .CP(n775), .CDN(n597), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n876), .E(n756), .CP(n810), .CDN(n596), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n874), .E(n756), .CP(n809), .CDN(n596), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n872), .E(n756), .CP(n807), .CDN(n596), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n870), .E(n756), .CP(n814), .CDN(n596), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n868), .E(n756), .CP(n803), .CDN(n596), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n866), .E(n756), .CP(n801), .CDN(n596), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n864), .E(n756), .CP(n823), .CDN(n596), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n862), .E(n756), .CP(n820), .CDN(n596), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n757), .CP(n788), .CDN(
        n596), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n858), .E(n757), .CP(n774), .CDN(n596), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n856), .E(n757), .CP(n826), .CDN(n596), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n757), .CP(n810), .CDN(n595), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n852), .E(n757), .CP(n824), .CDN(n595), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n850), .E(n757), .CP(n811), .CDN(n595), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n757), .CP(n801), .CDN(n595), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n846), .E(n757), .CP(n791), .CDN(n595), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n757), .CP(n817), .CDN(n595), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n842), .E(n757), .CP(n811), .CDN(n595), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n756), .CP(n825), .CDN(n595), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n838), .E(n756), .CP(n778), .CDN(n595), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n757), .CP(n813), .CDN(n595), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n830), .E(n759), .CP(n826), .CDN(n595), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n898), .E(n759), .CP(n774), .CDN(n594), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n896), .E(n758), .CP(n808), .CDN(n594), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n894), .E(n759), .CP(n810), .CDN(n594), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n892), .E(n758), .CP(n825), .CDN(n594), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n890), .E(n759), .CP(n806), .CDN(n594), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n888), .E(n758), .CP(n823), .CDN(n594), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n886), .E(n759), .CP(n790), .CDN(n594), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n884), .E(n758), .CP(n780), .CDN(n594), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n882), .E(n759), .CP(n816), .CDN(n594), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n758), .CP(n815), .CDN(
        n594), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n878), .E(n758), .CP(n813), .CDN(n594), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n876), .E(n758), .CP(n788), .CDN(n593), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n874), .E(n758), .CP(n775), .CDN(n593), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n872), .E(n758), .CP(n805), .CDN(n593), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n870), .E(n758), .CP(n795), .CDN(n593), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n868), .E(n758), .CP(ClockW), .CDN(n593), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n866), .E(n758), .CP(n815), .CDN(n593), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n864), .E(n758), .CP(n813), .CDN(n593), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n862), .E(n758), .CP(n812), .CDN(n593), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n759), .CP(n811), .CDN(
        n593), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n858), .E(n759), .CP(n804), .CDN(n593), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n856), .E(n759), .CP(n808), .CDN(n593), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n759), .CP(n807), .CDN(n592), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n852), .E(n759), .CP(n806), .CDN(n592), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n850), .E(n759), .CP(n811), .CDN(n592), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n759), .CP(n804), .CDN(n592), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n846), .E(n759), .CP(n802), .CDN(n592), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n759), .CP(n821), .CDN(n592), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n842), .E(n759), .CP(n799), .CDN(n592), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n758), .CP(n778), .CDN(n592), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n838), .E(n758), .CP(n821), .CDN(n592), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n759), .CP(n809), .CDN(n592), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(n830), .E(n763), .CP(n814), .CDN(n589), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n898), .E(n763), .CP(n820), .CDN(n588), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n896), .E(n762), .CP(n808), .CDN(n588), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n894), .E(n763), .CP(n814), .CDN(n588), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n892), .E(n762), .CP(n777), .CDN(n588), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n890), .E(n763), .CP(n821), .CDN(n588), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n888), .E(n762), .CP(n807), .CDN(n588), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n886), .E(n763), .CP(n809), .CDN(n588), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n884), .E(n762), .CP(n789), .CDN(n588), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n882), .E(n763), .CP(n794), .CDN(n588), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n762), .CP(n810), .CDN(
        n588), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n878), .E(n762), .CP(n819), .CDN(n588), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n876), .E(n762), .CP(n818), .CDN(n587), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n874), .E(n762), .CP(n816), .CDN(n587), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n872), .E(n762), .CP(n815), .CDN(n587), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n870), .E(n762), .CP(n814), .CDN(n587), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n868), .E(n762), .CP(n813), .CDN(n587), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n866), .E(n762), .CP(n812), .CDN(n587), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n864), .E(n762), .CP(n811), .CDN(n587), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n862), .E(n762), .CP(n795), .CDN(n587), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n763), .CP(n822), .CDN(
        n587), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n858), .E(n763), .CP(n812), .CDN(n587), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n856), .E(n763), .CP(n804), .CDN(n587), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n763), .CP(n801), .CDN(n586), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n852), .E(n763), .CP(n826), .CDN(n586), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n850), .E(n763), .CP(n822), .CDN(n586), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n763), .CP(n810), .CDN(n586), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n846), .E(n763), .CP(n777), .CDN(n586), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n763), .CP(n810), .CDN(n586), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n842), .E(n763), .CP(n797), .CDN(n586), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n762), .CP(n817), .CDN(n586), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n838), .E(n762), .CP(n822), .CDN(n586), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n763), .CP(n823), .CDN(n586), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n830), .E(n765), .CP(n772), .CDN(n586), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n898), .E(n765), .CP(n813), .CDN(n585), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n896), .E(n764), .CP(n823), .CDN(n585), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n894), .E(n765), .CP(n824), .CDN(n585), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n892), .E(n764), .CP(n777), .CDN(n585), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n890), .E(n765), .CP(n801), .CDN(n585), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n888), .E(n764), .CP(n825), .CDN(n585), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n886), .E(n765), .CP(n820), .CDN(n585), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n884), .E(n764), .CP(n796), .CDN(n585), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n882), .E(n765), .CP(n773), .CDN(n585), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n764), .CP(n821), .CDN(
        n585), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n878), .E(n764), .CP(n818), .CDN(n585), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n876), .E(n764), .CP(n798), .CDN(n584), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n874), .E(n764), .CP(n818), .CDN(n584), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n872), .E(n764), .CP(n815), .CDN(n584), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n870), .E(n764), .CP(n824), .CDN(n584), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n868), .E(n764), .CP(n796), .CDN(n584), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n866), .E(n764), .CP(n809), .CDN(n584), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n864), .E(n764), .CP(n824), .CDN(n584), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n862), .E(n764), .CP(n808), .CDN(n584), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n765), .CP(n793), .CDN(
        n584), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n858), .E(n765), .CP(n808), .CDN(n584), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n856), .E(n765), .CP(n774), .CDN(n584), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n765), .CP(n823), .CDN(n595), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n852), .E(n765), .CP(n826), .CDN(n583), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n850), .E(n765), .CP(n788), .CDN(n583), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n765), .CP(n772), .CDN(n583), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n846), .E(n765), .CP(n816), .CDN(n600), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n765), .CP(n809), .CDN(n601), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n842), .E(n765), .CP(ClockW), .CDN(n602), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n764), .CP(n807), .CDN(n593), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n838), .E(n764), .CP(n814), .CDN(n592), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n765), .CP(n778), .CDN(n593), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(n830), .E(n767), .CP(n784), .CDN(n594), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n898), .E(n767), .CP(n817), .CDN(n583), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n896), .E(n766), .CP(ClockW), .CDN(n583), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n894), .E(n767), .CP(n822), .CDN(n583), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n892), .E(n766), .CP(n772), .CDN(n583), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n890), .E(n767), .CP(n824), .CDN(n583), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n888), .E(n766), .CP(n801), .CDN(n583), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n886), .E(n767), .CP(n783), .CDN(n583), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n884), .E(n766), .CP(n793), .CDN(n583), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n882), .E(n767), .CP(n800), .CDN(n583), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n766), .CP(n810), .CDN(
        n583), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n878), .E(n766), .CP(n812), .CDN(n583), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n876), .E(n766), .CP(n773), .CDN(n582), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n874), .E(n766), .CP(n817), .CDN(n582), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n872), .E(n766), .CP(ClockW), .CDN(n582), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n870), .E(n766), .CP(n807), .CDN(n582), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n868), .E(n766), .CP(n808), .CDN(n582), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n866), .E(n766), .CP(n805), .CDN(n582), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n864), .E(n766), .CP(n809), .CDN(n582), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n862), .E(n766), .CP(n810), .CDN(n582), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n767), .CP(n820), .CDN(
        n582), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n858), .E(n767), .CP(n821), .CDN(n582), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n856), .E(n767), .CP(n822), .CDN(n582), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n767), .CP(n773), .CDN(n581), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n852), .E(n767), .CP(n813), .CDN(n581), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n850), .E(n767), .CP(ClockW), .CDN(n581), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n767), .CP(n824), .CDN(n581), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n846), .E(n767), .CP(n810), .CDN(n581), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n767), .CP(n809), .CDN(n581), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n842), .E(n767), .CP(n780), .CDN(n581), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n766), .CP(n808), .CDN(n581), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n838), .E(n766), .CP(n807), .CDN(n581), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n836), .E(n767), .CP(n787), .CDN(n581), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(n830), .E(n771), .CP(n808), .CDN(n578), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n898), .E(n770), .CP(n784), .CDN(n577), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n896), .E(n770), .CP(n773), .CDN(n577), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n894), .E(n771), .CP(n803), .CDN(n577), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n892), .E(n770), .CP(n823), .CDN(n577), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n890), .E(n771), .CP(n774), .CDN(n577), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n888), .E(n770), .CP(n774), .CDN(n577), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n886), .E(n771), .CP(n772), .CDN(n577), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n884), .E(n770), .CP(n808), .CDN(n577), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n882), .E(n771), .CP(n821), .CDN(n577), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n770), .CP(n818), .CDN(
        n577), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n878), .E(n770), .CP(n776), .CDN(n577), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n876), .E(n770), .CP(n819), .CDN(n576), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n874), .E(n770), .CP(n814), .CDN(n576), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n872), .E(n770), .CP(n826), .CDN(n576), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n870), .E(n770), .CP(n782), .CDN(n576), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n868), .E(n770), .CP(n807), .CDN(n576), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n866), .E(n770), .CP(n812), .CDN(n576), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n864), .E(n770), .CP(n825), .CDN(n576), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n862), .E(n770), .CP(n823), .CDN(n576), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n771), .CP(n824), .CDN(
        n576), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n858), .E(n771), .CP(n777), .CDN(n576), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n856), .E(n771), .CP(n794), .CDN(n576), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n771), .CP(n805), .CDN(n575), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n852), .E(n771), .CP(n782), .CDN(n575), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n850), .E(n771), .CP(n812), .CDN(n575), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n771), .CP(n796), .CDN(n575), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n846), .E(n771), .CP(n772), .CDN(n575), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n771), .CP(n773), .CDN(n575), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n842), .E(n771), .CP(n787), .CDN(n575), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n771), .CP(n790), .CDN(n575), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n838), .E(n770), .CP(n825), .CDN(n575), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n771), .CP(n826), .CDN(n575), 
        .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n34), .CP(ClockR), .CDN(n575), .Q(Dreadyr) );
  EDFCNQD1 Parityr_reg ( .D(n38), .E(n831), .CP(ClockR), .CDN(n667), .Q(
        ParityErr) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n46), .E(n831), .CP(ClockR), .CDN(n667), .Q(
        DataOr[0]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n42), .E(n831), .CP(ClockR), .CDN(n667), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n54), .E(Read), .CP(n827), .CDN(n668), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n50), .E(Read), .CP(ClockR), .CDN(n667), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n62), .E(Read), .CP(ClockR), .CDN(n667), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n58), .E(n831), .CP(ClockR), .CDN(n668), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n113), .E(n831), .CP(ClockR), .CDN(n615), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n109), .E(Read), .CP(n827), .CDN(n667), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n121), .E(Read), .CP(ClockR), .CDN(n667), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n117), .E(n831), .CP(ClockR), .CDN(n701), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n125), .E(n831), .CP(n827), .CDN(n667), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n129), .E(n831), .CP(ClockR), .CDN(n629), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n133), .E(Read), .CP(ClockR), .CDN(n667), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n137), .E(n831), .CP(ClockR), .CDN(n665), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n141), .E(n831), .CP(n827), .CDN(n667), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n145), .E(n831), .CP(ClockR), .CDN(n666), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n149), .E(Read), .CP(ClockR), .CDN(n636), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n153), .E(Read), .CP(n827), .CDN(n668), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n157), .E(n831), .CP(n827), .CDN(n668), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n161), .E(Read), .CP(n827), .CDN(n637), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n165), .E(Read), .CP(ClockR), .CDN(n668), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n169), .E(Read), .CP(ClockR), .CDN(n664), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n173), .E(n831), .CP(n827), .CDN(n629), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n177), .E(n831), .CP(n827), .CDN(n661), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n181), .E(Read), .CP(n827), .CDN(n665), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n185), .E(Read), .CP(n827), .CDN(n668), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n189), .E(Read), .CP(n827), .CDN(n666), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n193), .E(Read), .CP(n827), .CDN(n668), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n197), .E(Read), .CP(n827), .CDN(n596), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n201), .E(Read), .CP(n827), .CDN(n580), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n205), .E(Read), .CP(n827), .CDN(n579), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n209), .E(Read), .CP(n827), .CDN(n616), .Q(
        DataOr[17]) );
  DEL3 U3 ( .I(n55), .Z(n54) );
  DEL4 U4 ( .I(n56), .Z(n55) );
  DEL4 U5 ( .I(n57), .Z(n56) );
  DEL4 U6 ( .I(N33), .Z(n57) );
  DEL3 U7 ( .I(n59), .Z(n58) );
  DEL4 U8 ( .I(n60), .Z(n59) );
  DEL4 U9 ( .I(n61), .Z(n60) );
  DEL4 U10 ( .I(N34), .Z(n61) );
  DEL3 U11 ( .I(n114), .Z(n113) );
  DEL4 U12 ( .I(n115), .Z(n114) );
  DEL4 U13 ( .I(n116), .Z(n115) );
  DEL4 U14 ( .I(N35), .Z(n116) );
  DEL3 U15 ( .I(n118), .Z(n117) );
  DEL4 U16 ( .I(n119), .Z(n118) );
  DEL4 U17 ( .I(n120), .Z(n119) );
  DEL4 U18 ( .I(N36), .Z(n120) );
  DEL3 U19 ( .I(n130), .Z(n129) );
  DEL4 U20 ( .I(n131), .Z(n130) );
  DEL4 U21 ( .I(n132), .Z(n131) );
  DEL4 U22 ( .I(N37), .Z(n132) );
  DEL3 U23 ( .I(n138), .Z(n137) );
  DEL4 U24 ( .I(n139), .Z(n138) );
  DEL4 U30 ( .I(n140), .Z(n139) );
  DEL4 U31 ( .I(N38), .Z(n140) );
  DEL3 U32 ( .I(n146), .Z(n145) );
  DEL4 U35 ( .I(n147), .Z(n146) );
  DEL4 U36 ( .I(n148), .Z(n147) );
  DEL4 U37 ( .I(N39), .Z(n148) );
  DEL3 U38 ( .I(n154), .Z(n153) );
  DEL4 U43 ( .I(n155), .Z(n154) );
  DEL4 U44 ( .I(n156), .Z(n155) );
  DEL4 U45 ( .I(N40), .Z(n156) );
  DEL3 U46 ( .I(n162), .Z(n161) );
  DEL4 U47 ( .I(n163), .Z(n162) );
  DEL4 U48 ( .I(n164), .Z(n163) );
  DEL4 U49 ( .I(N41), .Z(n164) );
  DEL3 U50 ( .I(n170), .Z(n169) );
  DEL4 U51 ( .I(n171), .Z(n170) );
  DEL4 U52 ( .I(n172), .Z(n171) );
  DEL4 U53 ( .I(N42), .Z(n172) );
  XNR3D1 U54 ( .A1(DataI[6]), .A2(n846), .A3(n77), .ZN(n1) );
  OR2D1 U55 ( .A1(n69), .A2(n70), .Z(n2) );
  OR2D1 U56 ( .A1(n67), .A2(n70), .Z(n3) );
  OR2D1 U57 ( .A1(n68), .A2(n70), .Z(n4) );
  OR2D1 U58 ( .A1(n69), .A2(n103), .Z(n5) );
  OR2D1 U59 ( .A1(n67), .A2(n103), .Z(n6) );
  OR2D1 U60 ( .A1(n75), .A2(n103), .Z(n7) );
  OR2D1 U61 ( .A1(n74), .A2(n103), .Z(n8) );
  OR2D1 U62 ( .A1(n72), .A2(n103), .Z(n9) );
  OR2D1 U63 ( .A1(n71), .A2(n103), .Z(n10) );
  OR2D1 U64 ( .A1(n69), .A2(n101), .Z(n11) );
  OR2D1 U65 ( .A1(n67), .A2(n101), .Z(n12) );
  OR2D1 U66 ( .A1(n75), .A2(n101), .Z(n13) );
  OR2D1 U67 ( .A1(n74), .A2(n101), .Z(n14) );
  OR2D1 U68 ( .A1(n72), .A2(n101), .Z(n15) );
  OR2D1 U69 ( .A1(n71), .A2(n101), .Z(n16) );
  OR2D1 U70 ( .A1(n68), .A2(n103), .Z(n17) );
  OR2D1 U71 ( .A1(n73), .A2(n103), .Z(n18) );
  OR2D1 U72 ( .A1(n68), .A2(n101), .Z(n19) );
  OR2D1 U73 ( .A1(n73), .A2(n101), .Z(n20) );
  OR2D1 U74 ( .A1(n66), .A2(n69), .Z(n21) );
  OR2D1 U75 ( .A1(n66), .A2(n67), .Z(n22) );
  OR2D1 U76 ( .A1(n66), .A2(n75), .Z(n23) );
  OR2D1 U77 ( .A1(n66), .A2(n74), .Z(n24) );
  OR2D1 U78 ( .A1(n66), .A2(n72), .Z(n25) );
  OR2D1 U79 ( .A1(n66), .A2(n71), .Z(n26) );
  OR2D1 U80 ( .A1(n66), .A2(n68), .Z(n27) );
  OR2D1 U81 ( .A1(n66), .A2(n73), .Z(n28) );
  OR2D1 U82 ( .A1(n70), .A2(n75), .Z(n29) );
  OR2D1 U83 ( .A1(n70), .A2(n74), .Z(n30) );
  OR2D1 U84 ( .A1(n70), .A2(n72), .Z(n31) );
  OR2D1 U85 ( .A1(n70), .A2(n71), .Z(n32) );
  OR2D1 U86 ( .A1(n70), .A2(n73), .Z(n33) );
  DEL3 U87 ( .I(n35), .Z(n34) );
  DEL4 U88 ( .I(n36), .Z(n35) );
  DEL4 U89 ( .I(n37), .Z(n36) );
  DEL4 U90 ( .I(n107), .Z(n37) );
  OR2D0 U91 ( .A1(n831), .A2(Dreadyr), .Z(n107) );
  DEL2 U92 ( .I(N65), .Z(n38) );
  XOR3D0 U93 ( .A1(n62), .A2(n141), .A3(n40), .Z(N65) );
  DEL4 U94 ( .I(n97), .Z(n39) );
  XOR3D0 U95 ( .A1(n169), .A2(n161), .A3(n98), .Z(n97) );
  DEL4 U96 ( .I(n89), .Z(n40) );
  XOR3D0 U97 ( .A1(n149), .A2(n90), .A3(n91), .Z(n89) );
  DEL4 U98 ( .I(n93), .Z(n41) );
  XOR3D0 U99 ( .A1(n197), .A2(n205), .A3(n95), .Z(n93) );
  MUX4D0 U100 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n574), .S1(n560), .Z(
        n540) );
  DEL3 U101 ( .I(n43), .Z(n42) );
  MUX2ND0 U102 ( .I0(n213), .I1(n214), .S(N83), .ZN(N63) );
  DEL4 U103 ( .I(n44), .Z(n43) );
  DEL4 U104 ( .I(n45), .Z(n44) );
  DEL4 U105 ( .I(N63), .Z(n45) );
  MUX4D0 U106 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n567), .S1(n553), .Z(
        n292) );
  DEL3 U107 ( .I(n47), .Z(n46) );
  MUX2ND0 U108 ( .I0(n255), .I1(n256), .S(N83), .ZN(N64) );
  DEL4 U109 ( .I(n48), .Z(n47) );
  DEL4 U110 ( .I(n49), .Z(n48) );
  DEL4 U111 ( .I(N64), .Z(n49) );
  MUX4D0 U112 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n566), .S1(n552), .Z(
        n284) );
  DEL3 U113 ( .I(n51), .Z(n50) );
  MUX2ND0 U114 ( .I0(n215), .I1(n216), .S(N83), .ZN(N62) );
  DEL4 U115 ( .I(n52), .Z(n51) );
  DEL4 U116 ( .I(n53), .Z(n52) );
  DEL4 U117 ( .I(N62), .Z(n53) );
  MUX4D0 U118 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n567), .S1(n553), .Z(
        n300) );
  MUX2ND0 U119 ( .I0(n233), .I1(n234), .S(n835), .ZN(N33) );
  MUX4D0 U120 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n574), .S1(n560), .Z(
        n532) );
  MUX2ND0 U121 ( .I0(n231), .I1(n232), .S(n835), .ZN(N34) );
  MUX4D0 U122 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n573), .S1(n559), .Z(
        n524) );
  DEL3 U123 ( .I(n63), .Z(n62) );
  MUX2ND0 U124 ( .I0(n257), .I1(n258), .S(n835), .ZN(N61) );
  DEL4 U125 ( .I(n64), .Z(n63) );
  DEL4 U126 ( .I(n65), .Z(n64) );
  DEL4 U127 ( .I(N61), .Z(n65) );
  MUX4D0 U128 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n568), .S1(n554), .Z(
        n308) );
  DEL3 U129 ( .I(n110), .Z(n109) );
  MUX2ND0 U130 ( .I0(n245), .I1(n246), .S(N83), .ZN(N60) );
  DEL4 U131 ( .I(n111), .Z(n110) );
  DEL4 U132 ( .I(n112), .Z(n111) );
  DEL4 U133 ( .I(N60), .Z(n112) );
  MUX4D0 U134 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n569), .S1(n555), .Z(
        n316) );
  MUX2ND0 U135 ( .I0(n275), .I1(n276), .S(n835), .ZN(N35) );
  MUX4D0 U136 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n572), .S1(n558), .Z(
        n516) );
  MUX2ND0 U137 ( .I0(n253), .I1(n254), .S(n835), .ZN(N36) );
  MUX4D0 U138 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n572), .S1(n558), .Z(
        n508) );
  DEL3 U139 ( .I(n122), .Z(n121) );
  MUX2ND0 U140 ( .I0(n259), .I1(n260), .S(n835), .ZN(N59) );
  DEL4 U141 ( .I(n123), .Z(n122) );
  DEL4 U142 ( .I(n124), .Z(n123) );
  DEL4 U143 ( .I(N59), .Z(n124) );
  MUX4D0 U144 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n569), .S1(n555), .Z(
        n324) );
  DEL3 U145 ( .I(n126), .Z(n125) );
  MUX2ND0 U146 ( .I0(n235), .I1(n236), .S(N83), .ZN(N58) );
  DEL4 U147 ( .I(n127), .Z(n126) );
  DEL4 U148 ( .I(n128), .Z(n127) );
  DEL4 U149 ( .I(N58), .Z(n128) );
  MUX4D0 U150 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n564), .S1(n560), .Z(
        n332) );
  MUX2ND0 U151 ( .I0(n229), .I1(n230), .S(n835), .ZN(N37) );
  MUX4D0 U152 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n571), .S1(n557), .Z(
        n500) );
  DEL3 U153 ( .I(n134), .Z(n133) );
  MUX2ND0 U154 ( .I0(n217), .I1(n218), .S(N83), .ZN(N57) );
  DEL4 U155 ( .I(n135), .Z(n134) );
  DEL4 U156 ( .I(n136), .Z(n135) );
  DEL4 U157 ( .I(N57), .Z(n136) );
  MUX4D0 U158 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n573), .S1(n559), .Z(
        n340) );
  MUX2ND0 U159 ( .I0(n227), .I1(n228), .S(n835), .ZN(N38) );
  MUX4D0 U160 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n571), .S1(n550), .Z(
        n492) );
  DEL3 U161 ( .I(n142), .Z(n141) );
  MUX2ND0 U162 ( .I0(n237), .I1(n238), .S(n835), .ZN(N56) );
  DEL4 U163 ( .I(n143), .Z(n142) );
  DEL4 U164 ( .I(n144), .Z(n143) );
  DEL4 U165 ( .I(N56), .Z(n144) );
  MUX4D0 U166 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n563), .S1(n549), .Z(
        n348) );
  MUX2ND0 U167 ( .I0(n273), .I1(n274), .S(n835), .ZN(N39) );
  MUX4D0 U168 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n562), .S1(n558), .Z(
        n484) );
  DEL3 U169 ( .I(n150), .Z(n149) );
  MUX2ND0 U170 ( .I0(n261), .I1(n262), .S(n835), .ZN(N55) );
  DEL4 U171 ( .I(n151), .Z(n150) );
  DEL4 U172 ( .I(n152), .Z(n151) );
  DEL4 U173 ( .I(N55), .Z(n152) );
  MUX4D0 U174 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n574), .S1(n559), .Z(
        n356) );
  MUX2ND0 U175 ( .I0(n243), .I1(n244), .S(n835), .ZN(N40) );
  MUX4D0 U176 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n565), .S1(n550), .Z(
        n476) );
  DEL3 U177 ( .I(n158), .Z(n157) );
  MUX2ND0 U178 ( .I0(n247), .I1(n248), .S(N83), .ZN(N54) );
  DEL4 U179 ( .I(n159), .Z(n158) );
  DEL4 U180 ( .I(n160), .Z(n159) );
  DEL4 U181 ( .I(N54), .Z(n160) );
  MUX4D0 U182 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n567), .S1(n555), .Z(
        n364) );
  MUX2ND0 U183 ( .I0(n241), .I1(n242), .S(n835), .ZN(N41) );
  MUX4D0 U184 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n563), .S1(n547), .Z(
        n468) );
  DEL3 U185 ( .I(n166), .Z(n165) );
  MUX2ND0 U186 ( .I0(n263), .I1(n264), .S(N83), .ZN(N53) );
  DEL4 U187 ( .I(n167), .Z(n166) );
  DEL4 U188 ( .I(n168), .Z(n167) );
  DEL4 U189 ( .I(N53), .Z(n168) );
  MUX4D0 U190 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n564), .S1(n557), .Z(
        n372) );
  MUX2ND0 U191 ( .I0(n271), .I1(n272), .S(n835), .ZN(N42) );
  MUX4D0 U192 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(N79), .S1(N80), .Z(
        n460) );
  DEL3 U193 ( .I(n174), .Z(n173) );
  MUX2ND0 U194 ( .I0(n219), .I1(n220), .S(N83), .ZN(N52) );
  DEL4 U195 ( .I(n175), .Z(n174) );
  DEL4 U196 ( .I(n176), .Z(n175) );
  DEL4 U197 ( .I(N52), .Z(n176) );
  MUX4D0 U198 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n567), .S1(n554), .Z(
        n380) );
  DEL3 U199 ( .I(n178), .Z(n177) );
  MUX2ND0 U200 ( .I0(n251), .I1(n252), .S(n835), .ZN(N43) );
  DEL4 U201 ( .I(n179), .Z(n178) );
  DEL4 U202 ( .I(n180), .Z(n179) );
  DEL4 U203 ( .I(N43), .Z(n180) );
  MUX4D0 U204 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n563), .S1(n549), .Z(
        n452) );
  DEL3 U205 ( .I(n182), .Z(n181) );
  MUX2ND0 U206 ( .I0(n221), .I1(n222), .S(N83), .ZN(N51) );
  DEL4 U207 ( .I(n183), .Z(n182) );
  DEL4 U208 ( .I(n184), .Z(n183) );
  DEL4 U209 ( .I(N51), .Z(n184) );
  MUX4D0 U210 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n568), .S1(n552), .Z(
        n388) );
  DEL3 U211 ( .I(n186), .Z(n185) );
  MUX2ND0 U212 ( .I0(n225), .I1(n226), .S(N83), .ZN(N44) );
  DEL4 U213 ( .I(n187), .Z(n186) );
  DEL4 U214 ( .I(n188), .Z(n187) );
  DEL4 U215 ( .I(N44), .Z(n188) );
  MUX4D0 U216 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(N79), .S1(N80), .Z(
        n444) );
  DEL3 U217 ( .I(n190), .Z(n189) );
  MUX2ND0 U218 ( .I0(n249), .I1(n250), .S(N83), .ZN(N50) );
  DEL4 U219 ( .I(n191), .Z(n190) );
  DEL4 U220 ( .I(n192), .Z(n191) );
  DEL4 U221 ( .I(N50), .Z(n192) );
  MUX4D0 U222 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n571), .S1(n553), .Z(
        n396) );
  DEL3 U223 ( .I(n194), .Z(n193) );
  MUX2ND0 U224 ( .I0(n223), .I1(n224), .S(n835), .ZN(N45) );
  DEL4 U225 ( .I(n195), .Z(n194) );
  DEL4 U226 ( .I(n196), .Z(n195) );
  DEL4 U227 ( .I(N45), .Z(n196) );
  MUX4D0 U228 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(N79), .S1(N80), .Z(
        n436) );
  DEL3 U229 ( .I(n198), .Z(n197) );
  MUX2ND0 U230 ( .I0(n265), .I1(n266), .S(N83), .ZN(N49) );
  DEL4 U231 ( .I(n199), .Z(n198) );
  DEL4 U232 ( .I(n200), .Z(n199) );
  DEL4 U233 ( .I(N49), .Z(n200) );
  MUX4D0 U234 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n564), .S1(n551), .Z(
        n404) );
  DEL3 U235 ( .I(n202), .Z(n201) );
  MUX2ND0 U236 ( .I0(n269), .I1(n270), .S(n835), .ZN(N46) );
  DEL4 U237 ( .I(n203), .Z(n202) );
  DEL4 U238 ( .I(n204), .Z(n203) );
  DEL4 U239 ( .I(N46), .Z(n204) );
  MUX4D0 U240 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n570), .S1(n556), .Z(
        n428) );
  DEL3 U241 ( .I(n206), .Z(n205) );
  MUX2ND0 U242 ( .I0(n239), .I1(n240), .S(N83), .ZN(N48) );
  DEL4 U243 ( .I(n207), .Z(n206) );
  DEL4 U244 ( .I(n208), .Z(n207) );
  DEL4 U245 ( .I(N48), .Z(n208) );
  MUX4D0 U246 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n562), .S1(n548), .Z(
        n412) );
  DEL3 U247 ( .I(n210), .Z(n209) );
  MUX2ND0 U248 ( .I0(n267), .I1(n268), .S(N83), .ZN(N47) );
  DEL4 U249 ( .I(n211), .Z(n210) );
  DEL4 U250 ( .I(n212), .Z(n211) );
  DEL4 U251 ( .I(N47), .Z(n212) );
  MUX4D0 U252 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n565), .S1(n551), .Z(
        n420) );
  AN2D1 U253 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U254 ( .I(DataI[10]), .ZN(n857) );
  INVD1 U255 ( .I(DataI[11]), .ZN(n859) );
  INVD1 U256 ( .I(DataI[13]), .ZN(n863) );
  INVD1 U257 ( .I(DataI[14]), .ZN(n865) );
  INVD1 U258 ( .I(DataI[15]), .ZN(n867) );
  INVD1 U259 ( .I(DataI[16]), .ZN(n869) );
  INVD1 U260 ( .I(DataI[17]), .ZN(n871) );
  INVD1 U261 ( .I(DataI[18]), .ZN(n873) );
  INVD1 U262 ( .I(DataI[19]), .ZN(n875) );
  INVD1 U263 ( .I(DataI[20]), .ZN(n877) );
  INVD1 U264 ( .I(DataI[21]), .ZN(n879) );
  INVD1 U265 ( .I(DataI[22]), .ZN(n881) );
  INVD1 U266 ( .I(DataI[23]), .ZN(n883) );
  INVD1 U267 ( .I(DataI[24]), .ZN(n885) );
  INVD1 U268 ( .I(DataI[25]), .ZN(n887) );
  INVD1 U269 ( .I(DataI[26]), .ZN(n889) );
  INVD1 U270 ( .I(DataI[27]), .ZN(n891) );
  INVD1 U271 ( .I(DataI[28]), .ZN(n893) );
  INVD1 U272 ( .I(DataI[29]), .ZN(n895) );
  INVD1 U273 ( .I(DataI[30]), .ZN(n897) );
  INVD1 U274 ( .I(DataI[31]), .ZN(n899) );
  INVD1 U275 ( .I(DataI[0]), .ZN(n837) );
  INVD1 U276 ( .I(DataI[1]), .ZN(n839) );
  INVD1 U277 ( .I(DataI[2]), .ZN(n841) );
  INVD1 U278 ( .I(DataI[3]), .ZN(n843) );
  INVD1 U279 ( .I(DataI[4]), .ZN(n845) );
  INVD1 U280 ( .I(DataI[5]), .ZN(n847) );
  INVD1 U281 ( .I(DataI[6]), .ZN(n849) );
  INVD1 U282 ( .I(DataI[7]), .ZN(n851) );
  INVD1 U283 ( .I(DataI[8]), .ZN(n853) );
  INVD1 U284 ( .I(DataI[9]), .ZN(n855) );
  INVD1 U285 ( .I(DataI[12]), .ZN(n861) );
  BUFFD1 U286 ( .I(n689), .Z(n581) );
  BUFFD1 U287 ( .I(n674), .Z(n582) );
  BUFFD1 U288 ( .I(n704), .Z(n583) );
  BUFFD1 U289 ( .I(n700), .Z(n584) );
  BUFFD1 U290 ( .I(n700), .Z(n585) );
  BUFFD1 U291 ( .I(n697), .Z(n586) );
  BUFFD1 U292 ( .I(n696), .Z(n587) );
  BUFFD1 U293 ( .I(n699), .Z(n588) );
  BUFFD1 U294 ( .I(n699), .Z(n589) );
  BUFFD1 U295 ( .I(n699), .Z(n590) );
  BUFFD1 U296 ( .I(n699), .Z(n591) );
  BUFFD1 U297 ( .I(n698), .Z(n592) );
  BUFFD1 U298 ( .I(n698), .Z(n593) );
  BUFFD1 U299 ( .I(n697), .Z(n594) );
  BUFFD1 U300 ( .I(n697), .Z(n595) );
  BUFFD1 U301 ( .I(n701), .Z(n596) );
  BUFFD1 U302 ( .I(n706), .Z(n597) );
  BUFFD1 U303 ( .I(n696), .Z(n598) );
  BUFFD1 U304 ( .I(n696), .Z(n599) );
  BUFFD1 U305 ( .I(n695), .Z(n600) );
  BUFFD1 U306 ( .I(n695), .Z(n601) );
  BUFFD1 U307 ( .I(n694), .Z(n602) );
  BUFFD1 U308 ( .I(n693), .Z(n603) );
  BUFFD1 U309 ( .I(n693), .Z(n604) );
  BUFFD1 U310 ( .I(n692), .Z(n605) );
  BUFFD1 U311 ( .I(n692), .Z(n606) );
  BUFFD1 U312 ( .I(n691), .Z(n607) );
  BUFFD1 U313 ( .I(n691), .Z(n608) );
  BUFFD1 U314 ( .I(n690), .Z(n609) );
  BUFFD1 U315 ( .I(n690), .Z(n610) );
  BUFFD1 U316 ( .I(n689), .Z(n611) );
  BUFFD1 U317 ( .I(n689), .Z(n612) );
  BUFFD1 U318 ( .I(n688), .Z(n613) );
  BUFFD1 U319 ( .I(n688), .Z(n614) );
  BUFFD1 U320 ( .I(n687), .Z(n615) );
  BUFFD1 U321 ( .I(n687), .Z(n616) );
  BUFFD1 U322 ( .I(n686), .Z(n617) );
  BUFFD1 U323 ( .I(n686), .Z(n618) );
  BUFFD1 U324 ( .I(n685), .Z(n619) );
  BUFFD1 U325 ( .I(n685), .Z(n620) );
  BUFFD1 U326 ( .I(n684), .Z(n621) );
  BUFFD1 U327 ( .I(n684), .Z(n622) );
  BUFFD1 U328 ( .I(n683), .Z(n623) );
  BUFFD1 U329 ( .I(n683), .Z(n624) );
  BUFFD1 U330 ( .I(n682), .Z(n625) );
  BUFFD1 U331 ( .I(n682), .Z(n626) );
  BUFFD1 U332 ( .I(n681), .Z(n627) );
  BUFFD1 U333 ( .I(n681), .Z(n628) );
  BUFFD1 U334 ( .I(n705), .Z(n629) );
  BUFFD1 U335 ( .I(n680), .Z(n630) );
  BUFFD1 U336 ( .I(n680), .Z(n631) );
  BUFFD1 U337 ( .I(n679), .Z(n632) );
  BUFFD1 U338 ( .I(n679), .Z(n633) );
  BUFFD1 U339 ( .I(n672), .Z(n634) );
  BUFFD1 U340 ( .I(n669), .Z(n635) );
  BUFFD1 U341 ( .I(n678), .Z(n636) );
  BUFFD1 U342 ( .I(n678), .Z(n637) );
  BUFFD1 U343 ( .I(n689), .Z(n638) );
  BUFFD1 U344 ( .I(n677), .Z(n639) );
  BUFFD1 U345 ( .I(n677), .Z(n640) );
  BUFFD1 U346 ( .I(n676), .Z(n641) );
  BUFFD1 U347 ( .I(n676), .Z(n642) );
  BUFFD1 U348 ( .I(n676), .Z(n643) );
  BUFFD1 U349 ( .I(n677), .Z(n644) );
  BUFFD1 U350 ( .I(n675), .Z(n645) );
  BUFFD1 U351 ( .I(n675), .Z(n646) );
  BUFFD1 U352 ( .I(n675), .Z(n647) );
  BUFFD1 U353 ( .I(n675), .Z(n648) );
  BUFFD1 U354 ( .I(n674), .Z(n649) );
  BUFFD1 U355 ( .I(n674), .Z(n650) );
  BUFFD1 U356 ( .I(n673), .Z(n651) );
  BUFFD1 U357 ( .I(n673), .Z(n652) );
  BUFFD1 U358 ( .I(n673), .Z(n653) );
  BUFFD1 U359 ( .I(n674), .Z(n654) );
  BUFFD1 U360 ( .I(n672), .Z(n655) );
  BUFFD1 U361 ( .I(n672), .Z(n656) );
  BUFFD1 U362 ( .I(n671), .Z(n657) );
  BUFFD1 U363 ( .I(n671), .Z(n658) );
  BUFFD1 U364 ( .I(n671), .Z(n659) );
  BUFFD1 U365 ( .I(n671), .Z(n660) );
  BUFFD1 U366 ( .I(n678), .Z(n661) );
  BUFFD1 U367 ( .I(n678), .Z(n662) );
  BUFFD1 U368 ( .I(n678), .Z(n663) );
  BUFFD1 U369 ( .I(n678), .Z(n664) );
  BUFFD1 U370 ( .I(n670), .Z(n665) );
  BUFFD1 U371 ( .I(n670), .Z(n666) );
  BUFFD1 U372 ( .I(n669), .Z(n667) );
  BUFFD1 U373 ( .I(n703), .Z(n575) );
  BUFFD1 U374 ( .I(n703), .Z(n576) );
  BUFFD1 U375 ( .I(n702), .Z(n577) );
  BUFFD1 U376 ( .I(n702), .Z(n578) );
  BUFFD1 U377 ( .I(n701), .Z(n579) );
  BUFFD1 U378 ( .I(n701), .Z(n580) );
  BUFFD1 U379 ( .I(n704), .Z(n700) );
  BUFFD1 U380 ( .I(n704), .Z(n699) );
  BUFFD1 U381 ( .I(n707), .Z(n698) );
  BUFFD1 U382 ( .I(n707), .Z(n697) );
  BUFFD1 U383 ( .I(n707), .Z(n696) );
  BUFFD1 U384 ( .I(n707), .Z(n695) );
  BUFFD1 U385 ( .I(n707), .Z(n694) );
  BUFFD1 U386 ( .I(n696), .Z(n693) );
  BUFFD1 U387 ( .I(n697), .Z(n692) );
  BUFFD1 U388 ( .I(n698), .Z(n691) );
  BUFFD1 U389 ( .I(n704), .Z(n690) );
  BUFFD1 U390 ( .I(n704), .Z(n689) );
  BUFFD1 U391 ( .I(n704), .Z(n688) );
  BUFFD1 U392 ( .I(n707), .Z(n687) );
  BUFFD1 U393 ( .I(n687), .Z(n686) );
  BUFFD1 U394 ( .I(n695), .Z(n685) );
  BUFFD1 U395 ( .I(n698), .Z(n684) );
  BUFFD1 U396 ( .I(n694), .Z(n683) );
  BUFFD1 U397 ( .I(n695), .Z(n682) );
  BUFFD1 U398 ( .I(n705), .Z(n681) );
  BUFFD1 U399 ( .I(n705), .Z(n680) );
  BUFFD1 U400 ( .I(n705), .Z(n679) );
  BUFFD1 U401 ( .I(n706), .Z(n678) );
  BUFFD1 U402 ( .I(n704), .Z(n677) );
  BUFFD1 U403 ( .I(n704), .Z(n676) );
  BUFFD1 U404 ( .I(n704), .Z(n675) );
  BUFFD1 U405 ( .I(n704), .Z(n674) );
  BUFFD1 U406 ( .I(n704), .Z(n673) );
  BUFFD1 U407 ( .I(n670), .Z(n672) );
  BUFFD1 U408 ( .I(n704), .Z(n671) );
  BUFFD1 U409 ( .I(n706), .Z(n670) );
  BUFFD1 U410 ( .I(n670), .Z(n669) );
  BUFFD1 U411 ( .I(n565), .Z(n566) );
  BUFFD1 U412 ( .I(n565), .Z(n567) );
  BUFFD1 U413 ( .I(n564), .Z(n568) );
  BUFFD1 U414 ( .I(n564), .Z(n569) );
  BUFFD1 U415 ( .I(n561), .Z(n570) );
  BUFFD1 U416 ( .I(n568), .Z(n571) );
  BUFFD1 U417 ( .I(n569), .Z(n572) );
  BUFFD1 U418 ( .I(n562), .Z(n573) );
  BUFFD1 U419 ( .I(n562), .Z(n574) );
  BUFFD1 U420 ( .I(n551), .Z(n552) );
  BUFFD1 U421 ( .I(n551), .Z(n553) );
  BUFFD1 U422 ( .I(n550), .Z(n554) );
  BUFFD1 U423 ( .I(n550), .Z(n555) );
  BUFFD1 U424 ( .I(n547), .Z(n556) );
  BUFFD1 U425 ( .I(n550), .Z(n557) );
  BUFFD1 U426 ( .I(n552), .Z(n558) );
  BUFFD1 U427 ( .I(n548), .Z(n559) );
  BUFFD1 U428 ( .I(n548), .Z(n560) );
  BUFFD1 U429 ( .I(n789), .Z(n806) );
  BUFFD1 U430 ( .I(n807), .Z(n805) );
  BUFFD1 U431 ( .I(n807), .Z(n804) );
  BUFFD1 U432 ( .I(n792), .Z(n803) );
  BUFFD1 U433 ( .I(n809), .Z(n802) );
  BUFFD1 U434 ( .I(n809), .Z(n801) );
  BUFFD1 U435 ( .I(n810), .Z(n800) );
  BUFFD1 U436 ( .I(n810), .Z(n799) );
  BUFFD1 U437 ( .I(n811), .Z(n798) );
  BUFFD1 U438 ( .I(n811), .Z(n797) );
  BUFFD1 U439 ( .I(n812), .Z(n796) );
  BUFFD1 U440 ( .I(n812), .Z(n795) );
  BUFFD1 U441 ( .I(n813), .Z(n794) );
  BUFFD1 U442 ( .I(n813), .Z(n793) );
  BUFFD1 U443 ( .I(n814), .Z(n792) );
  BUFFD1 U444 ( .I(n814), .Z(n791) );
  BUFFD1 U445 ( .I(n815), .Z(n790) );
  BUFFD1 U446 ( .I(n815), .Z(n789) );
  BUFFD1 U447 ( .I(n816), .Z(n788) );
  BUFFD1 U448 ( .I(n816), .Z(n787) );
  BUFFD1 U449 ( .I(n817), .Z(n786) );
  BUFFD1 U450 ( .I(n817), .Z(n785) );
  BUFFD1 U451 ( .I(n818), .Z(n784) );
  BUFFD1 U452 ( .I(n818), .Z(n783) );
  BUFFD1 U453 ( .I(n819), .Z(n782) );
  BUFFD1 U454 ( .I(n819), .Z(n781) );
  BUFFD1 U455 ( .I(n820), .Z(n780) );
  BUFFD1 U456 ( .I(n820), .Z(n779) );
  BUFFD1 U457 ( .I(n821), .Z(n778) );
  BUFFD1 U458 ( .I(n821), .Z(n777) );
  BUFFD1 U459 ( .I(n822), .Z(n776) );
  BUFFD1 U460 ( .I(n822), .Z(n775) );
  BUFFD1 U461 ( .I(n706), .Z(n668) );
  INVD1 U462 ( .I(n1), .ZN(n830) );
  INVD1 U463 ( .I(n1), .ZN(n829) );
  BUFFD1 U464 ( .I(n694), .Z(n702) );
  BUFFD1 U465 ( .I(n707), .Z(n701) );
  BUFFD1 U466 ( .I(n694), .Z(n703) );
  BUFFD1 U467 ( .I(n108), .Z(n704) );
  BUFFD1 U468 ( .I(n706), .Z(n705) );
  BUFFD1 U469 ( .I(n561), .Z(n565) );
  BUFFD1 U470 ( .I(n547), .Z(n551) );
  BUFFD1 U471 ( .I(n561), .Z(n564) );
  BUFFD1 U472 ( .I(n547), .Z(n550) );
  BUFFD1 U473 ( .I(N79), .Z(n563) );
  BUFFD1 U474 ( .I(N80), .Z(n549) );
  BUFFD1 U475 ( .I(n563), .Z(n562) );
  BUFFD1 U476 ( .I(n549), .Z(n548) );
  BUFFD1 U477 ( .I(n785), .Z(n807) );
  BUFFD1 U478 ( .I(n779), .Z(n808) );
  BUFFD1 U479 ( .I(n819), .Z(n809) );
  BUFFD1 U480 ( .I(n813), .Z(n810) );
  BUFFD1 U481 ( .I(n826), .Z(n811) );
  BUFFD1 U482 ( .I(n826), .Z(n812) );
  BUFFD1 U483 ( .I(n826), .Z(n813) );
  BUFFD1 U484 ( .I(n825), .Z(n814) );
  BUFFD1 U485 ( .I(n825), .Z(n815) );
  BUFFD1 U486 ( .I(n825), .Z(n816) );
  BUFFD1 U487 ( .I(n824), .Z(n817) );
  BUFFD1 U488 ( .I(n824), .Z(n818) );
  BUFFD1 U489 ( .I(n824), .Z(n819) );
  BUFFD1 U490 ( .I(n823), .Z(n820) );
  BUFFD1 U491 ( .I(n823), .Z(n821) );
  BUFFD1 U492 ( .I(n823), .Z(n822) );
  BUFFD1 U493 ( .I(n108), .Z(n707) );
  BUFFD1 U494 ( .I(n108), .Z(n706) );
  BUFFD1 U495 ( .I(N79), .Z(n561) );
  BUFFD1 U496 ( .I(N80), .Z(n547) );
  INVD1 U497 ( .I(n29), .ZN(n733) );
  INVD1 U498 ( .I(n29), .ZN(n732) );
  INVD1 U499 ( .I(n30), .ZN(n731) );
  INVD1 U500 ( .I(n30), .ZN(n730) );
  INVD1 U501 ( .I(n33), .ZN(n729) );
  INVD1 U502 ( .I(n33), .ZN(n728) );
  INVD1 U503 ( .I(n31), .ZN(n727) );
  INVD1 U504 ( .I(n31), .ZN(n726) );
  INVD1 U505 ( .I(n32), .ZN(n725) );
  INVD1 U506 ( .I(n32), .ZN(n724) );
  INVD1 U507 ( .I(n21), .ZN(n723) );
  INVD1 U508 ( .I(n21), .ZN(n722) );
  INVD1 U509 ( .I(n27), .ZN(n721) );
  INVD1 U510 ( .I(n27), .ZN(n720) );
  INVD1 U511 ( .I(n22), .ZN(n719) );
  INVD1 U512 ( .I(n22), .ZN(n718) );
  INVD1 U513 ( .I(n23), .ZN(n717) );
  INVD1 U514 ( .I(n23), .ZN(n716) );
  INVD1 U515 ( .I(n24), .ZN(n715) );
  INVD1 U516 ( .I(n24), .ZN(n714) );
  INVD1 U517 ( .I(n28), .ZN(n713) );
  INVD1 U518 ( .I(n28), .ZN(n712) );
  INVD1 U519 ( .I(n25), .ZN(n711) );
  INVD1 U520 ( .I(n25), .ZN(n710) );
  INVD1 U521 ( .I(n26), .ZN(n709) );
  INVD1 U522 ( .I(n26), .ZN(n708) );
  INVD1 U523 ( .I(n5), .ZN(n771) );
  INVD1 U524 ( .I(n5), .ZN(n770) );
  INVD1 U525 ( .I(n17), .ZN(n769) );
  INVD1 U526 ( .I(n17), .ZN(n768) );
  INVD1 U527 ( .I(n6), .ZN(n767) );
  INVD1 U528 ( .I(n6), .ZN(n766) );
  INVD1 U529 ( .I(n7), .ZN(n765) );
  INVD1 U530 ( .I(n7), .ZN(n764) );
  INVD1 U531 ( .I(n8), .ZN(n763) );
  INVD1 U532 ( .I(n8), .ZN(n762) );
  INVD1 U533 ( .I(n18), .ZN(n761) );
  INVD1 U534 ( .I(n18), .ZN(n760) );
  INVD1 U535 ( .I(n9), .ZN(n759) );
  INVD1 U536 ( .I(n9), .ZN(n758) );
  INVD1 U537 ( .I(n10), .ZN(n757) );
  INVD1 U538 ( .I(n10), .ZN(n756) );
  INVD1 U539 ( .I(n11), .ZN(n755) );
  INVD1 U540 ( .I(n11), .ZN(n754) );
  INVD1 U541 ( .I(n19), .ZN(n753) );
  INVD1 U542 ( .I(n19), .ZN(n752) );
  INVD1 U543 ( .I(n12), .ZN(n751) );
  INVD1 U544 ( .I(n12), .ZN(n750) );
  INVD1 U545 ( .I(n13), .ZN(n749) );
  INVD1 U546 ( .I(n13), .ZN(n748) );
  INVD1 U547 ( .I(n14), .ZN(n747) );
  INVD1 U548 ( .I(n14), .ZN(n746) );
  INVD1 U549 ( .I(n20), .ZN(n745) );
  INVD1 U550 ( .I(n20), .ZN(n744) );
  INVD1 U551 ( .I(n15), .ZN(n743) );
  INVD1 U552 ( .I(n15), .ZN(n742) );
  INVD1 U553 ( .I(n16), .ZN(n741) );
  INVD1 U554 ( .I(n16), .ZN(n740) );
  INVD1 U555 ( .I(n2), .ZN(n739) );
  INVD1 U556 ( .I(n2), .ZN(n738) );
  INVD1 U557 ( .I(n4), .ZN(n737) );
  INVD1 U558 ( .I(n4), .ZN(n736) );
  INVD1 U559 ( .I(n3), .ZN(n735) );
  INVD1 U560 ( .I(n3), .ZN(n734) );
  BUFFD1 U561 ( .I(n773), .Z(n826) );
  BUFFD1 U562 ( .I(n773), .Z(n825) );
  BUFFD1 U563 ( .I(n772), .Z(n824) );
  BUFFD1 U564 ( .I(n772), .Z(n823) );
  XOR3D1 U565 ( .A1(DataI[4]), .A2(n78), .A3(n79), .Z(n77) );
  XOR3D1 U566 ( .A1(n84), .A2(n856), .A3(n85), .Z(n83) );
  XOR3D1 U567 ( .A1(n870), .A2(n868), .A3(n86), .Z(n85) );
  XOR3D1 U568 ( .A1(n87), .A2(n866), .A3(n88), .Z(n86) );
  XOR3D1 U569 ( .A1(DataI[2]), .A2(n838), .A3(n80), .Z(n79) );
  XOR3D1 U570 ( .A1(n81), .A2(DataI[0]), .A3(n82), .Z(n80) );
  XOR3D1 U571 ( .A1(DataI[12]), .A2(n858), .A3(n83), .Z(n82) );
  BUFFD1 U572 ( .I(n834), .Z(n544) );
  BUFFD1 U573 ( .I(N83), .Z(n835) );
  BUFFD1 U574 ( .I(n833), .Z(n546) );
  BUFFD1 U575 ( .I(n834), .Z(n543) );
  BUFFD1 U576 ( .I(n833), .Z(n545) );
  INVD1 U577 ( .I(n832), .ZN(n831) );
  BUFFD1 U578 ( .I(n774), .Z(n773) );
  BUFFD1 U579 ( .I(n774), .Z(n772) );
  INVD1 U580 ( .I(n828), .ZN(n827) );
  INVD1 U581 ( .I(n875), .ZN(n874) );
  INVD1 U582 ( .I(n877), .ZN(n876) );
  INVD1 U583 ( .I(n885), .ZN(n884) );
  INVD1 U584 ( .I(n887), .ZN(n886) );
  INVD1 U585 ( .I(n893), .ZN(n892) );
  INVD1 U586 ( .I(n895), .ZN(n894) );
  INVD1 U587 ( .I(n867), .ZN(n866) );
  INVD1 U588 ( .I(n869), .ZN(n868) );
  INVD1 U589 ( .I(n873), .ZN(n872) );
  INVD1 U590 ( .I(n883), .ZN(n882) );
  INVD1 U591 ( .I(n891), .ZN(n890) );
  INVD1 U592 ( .I(n871), .ZN(n870) );
  INVD1 U593 ( .I(n889), .ZN(n888) );
  INVD1 U594 ( .I(n897), .ZN(n896) );
  INVD1 U595 ( .I(n899), .ZN(n898) );
  INVD1 U596 ( .I(n851), .ZN(n850) );
  INVD1 U597 ( .I(n853), .ZN(n852) );
  INVD1 U598 ( .I(n865), .ZN(n864) );
  INVD1 U599 ( .I(n879), .ZN(n878) );
  INVD1 U600 ( .I(n839), .ZN(n838) );
  INVD1 U601 ( .I(n847), .ZN(n846) );
  INVD1 U602 ( .I(n857), .ZN(n856) );
  INVD1 U603 ( .I(n859), .ZN(n858) );
  INVD1 U604 ( .I(n837), .ZN(n836) );
  INVD1 U605 ( .I(n843), .ZN(n842) );
  INVD1 U606 ( .I(n863), .ZN(n862) );
  INVD1 U607 ( .I(n841), .ZN(n840) );
  INVD1 U608 ( .I(n845), .ZN(n844) );
  INVD1 U609 ( .I(n849), .ZN(n848) );
  INVD1 U610 ( .I(n855), .ZN(n854) );
  INVD1 U611 ( .I(n861), .ZN(n860) );
  INVD1 U612 ( .I(n881), .ZN(n880) );
  INVD1 U613 ( .I(Reset), .ZN(n108) );
  XOR3D1 U614 ( .A1(n99), .A2(n153), .A3(n100), .Z(n98) );
  XOR3D1 U615 ( .A1(n209), .A2(n96), .A3(n39), .Z(n95) );
  XOR3D1 U616 ( .A1(n121), .A2(n125), .A3(n92), .Z(n91) );
  ND3D1 U617 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  INVD1 U618 ( .I(ClockR), .ZN(n828) );
  BUFFD1 U619 ( .I(ClockW), .Z(n774) );
  MUX4D0 U620 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n574), .S1(n560), .Z(
        n535) );
  MUX4D0 U621 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n574), .S1(n560), .Z(
        n537) );
  MUX4D0 U622 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n574), .S1(n560), .Z(
        n538) );
  MUX4D0 U623 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n574), .S1(n560), .Z(
        n539) );
  MUX4D0 U624 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n574), .S1(n560), .Z(
        n541) );
  MUX4D0 U625 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n574), .S1(n560), .Z(
        n542) );
  MUX4D0 U626 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n566), .S1(n552), .Z(
        n279) );
  MUX4D0 U627 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n566), .S1(n552), .Z(
        n281) );
  MUX4D0 U628 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n566), .S1(n552), .Z(
        n282) );
  MUX4D0 U629 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n566), .S1(n552), .Z(
        n283) );
  MUX4D0 U630 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n566), .S1(n552), .Z(n285)
         );
  MUX4D0 U631 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n566), .S1(n552), .Z(n286)
         );
  MUX4D0 U632 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n566), .S1(n552), .Z(
        n287) );
  MUX4D0 U633 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n566), .S1(n552), .Z(
        n289) );
  MUX4D0 U634 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n566), .S1(n552), .Z(
        n290) );
  MUX4D0 U635 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n567), .S1(n553), .Z(
        n291) );
  MUX4D0 U636 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n567), .S1(n553), .Z(n293)
         );
  MUX4D0 U637 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n567), .S1(n553), .Z(n294)
         );
  MUX4D0 U638 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n567), .S1(n553), .Z(
        n295) );
  MUX4D0 U639 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n567), .S1(n553), .Z(
        n297) );
  MUX4D0 U640 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n567), .S1(n553), .Z(
        n298) );
  MUX4D0 U641 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n567), .S1(n553), .Z(
        n299) );
  MUX4D0 U642 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n567), .S1(n553), .Z(n301)
         );
  MUX4D0 U643 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n567), .S1(n553), .Z(n302)
         );
  MUX4D0 U644 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n568), .S1(n554), .Z(
        n303) );
  MUX4D0 U645 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n568), .S1(n554), .Z(
        n305) );
  MUX4D0 U646 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n568), .S1(n554), .Z(
        n306) );
  MUX4D0 U647 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n568), .S1(n554), .Z(
        n307) );
  MUX4D0 U648 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n568), .S1(n554), .Z(n309)
         );
  MUX4D0 U649 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n568), .S1(n554), .Z(n310)
         );
  MUX4D0 U650 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n568), .S1(n554), .Z(
        n311) );
  MUX4D0 U651 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n568), .S1(n554), .Z(
        n313) );
  MUX4D0 U652 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n568), .S1(n554), .Z(
        n314) );
  MUX4D0 U653 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n569), .S1(n555), .Z(
        n315) );
  MUX4D0 U654 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n569), .S1(n555), .Z(n317)
         );
  MUX4D0 U655 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n569), .S1(n555), .Z(n318)
         );
  MUX4D0 U656 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n569), .S1(n555), .Z(
        n319) );
  MUX4D0 U657 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n569), .S1(n555), .Z(
        n321) );
  MUX4D0 U658 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n569), .S1(n555), .Z(
        n322) );
  MUX4D0 U659 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n569), .S1(n555), .Z(
        n323) );
  MUX4D0 U660 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n569), .S1(n555), .Z(n325)
         );
  MUX4D0 U661 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n569), .S1(n555), .Z(n326)
         );
  MUX4D0 U662 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n562), .S1(n549), .Z(
        n327) );
  MUX4D0 U663 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n565), .S1(n559), .Z(
        n329) );
  MUX4D0 U664 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n562), .S1(n548), .Z(
        n330) );
  MUX4D0 U665 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n567), .S1(n548), .Z(
        n331) );
  MUX4D0 U666 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n562), .S1(n551), .Z(n333)
         );
  MUX4D0 U667 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n566), .S1(n559), .Z(n334)
         );
  MUX4D0 U668 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n565), .S1(n550), .Z(
        n335) );
  MUX4D0 U669 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n562), .S1(n548), .Z(
        n337) );
  MUX4D0 U670 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n562), .S1(n560), .Z(
        n338) );
  MUX4D0 U671 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n562), .S1(n551), .Z(
        n339) );
  MUX4D0 U672 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n562), .S1(n548), .Z(n341)
         );
  MUX4D0 U673 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n564), .S1(n550), .Z(n342)
         );
  MUX4D0 U674 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n571), .S1(n550), .Z(
        n343) );
  MUX4D0 U675 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(N79), .S1(N80), .Z(n345)
         );
  MUX4D0 U676 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n573), .S1(n559), .Z(
        n346) );
  MUX4D0 U677 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n571), .S1(n557), .Z(
        n347) );
  MUX4D0 U678 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n572), .S1(n558), .Z(n349)
         );
  MUX4D0 U679 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n561), .S1(n547), .Z(n350)
         );
  MUX4D0 U680 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n574), .S1(n560), .Z(
        n351) );
  MUX4D0 U681 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n573), .S1(n558), .Z(
        n353) );
  MUX4D0 U682 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n573), .S1(n560), .Z(
        n354) );
  MUX4D0 U683 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n574), .S1(n559), .Z(
        n355) );
  MUX4D0 U684 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n573), .S1(n560), .Z(n357)
         );
  MUX4D0 U685 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n573), .S1(n560), .Z(n358)
         );
  MUX4D0 U686 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n574), .S1(n560), .Z(
        n359) );
  MUX4D0 U687 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n573), .S1(n559), .Z(
        n361) );
  MUX4D0 U688 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n573), .S1(n558), .Z(
        n362) );
  MUX4D0 U689 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n568), .S1(n554), .Z(
        n363) );
  MUX4D0 U690 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n569), .S1(n553), .Z(
        n365) );
  MUX4D0 U691 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n566), .S1(n552), .Z(
        n366) );
  MUX4D0 U692 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n563), .S1(n557), .Z(
        n367) );
  MUX4D0 U693 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n567), .S1(n553), .Z(
        n369) );
  MUX4D0 U694 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n571), .S1(n554), .Z(
        n370) );
  MUX4D0 U695 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n565), .S1(n557), .Z(
        n371) );
  MUX4D0 U696 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n572), .S1(n552), .Z(
        n373) );
  MUX4D0 U697 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n569), .S1(n555), .Z(
        n374) );
  MUX4D0 U698 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n566), .S1(n555), .Z(
        n375) );
  MUX4D0 U699 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n568), .S1(n552), .Z(
        n377) );
  MUX4D0 U700 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n568), .S1(n554), .Z(
        n378) );
  MUX4D0 U701 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n567), .S1(n553), .Z(
        n379) );
  MUX4D0 U702 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n566), .S1(n555), .Z(
        n381) );
  MUX4D0 U703 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n566), .S1(n555), .Z(
        n382) );
  MUX4D0 U704 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n571), .S1(n554), .Z(
        n383) );
  MUX4D0 U705 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n567), .S1(n553), .Z(
        n385) );
  MUX4D0 U706 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n567), .S1(n553), .Z(
        n386) );
  MUX4D0 U707 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n569), .S1(n552), .Z(
        n387) );
  MUX4D0 U708 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n567), .S1(n553), .Z(
        n389) );
  MUX4D0 U709 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n566), .S1(n551), .Z(
        n390) );
  MUX4D0 U710 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n568), .S1(n552), .Z(
        n391) );
  MUX4D0 U711 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n569), .S1(n554), .Z(
        n393) );
  MUX4D0 U712 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n569), .S1(n552), .Z(
        n394) );
  MUX4D0 U713 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n572), .S1(n553), .Z(
        n395) );
  MUX4D0 U714 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n564), .S1(n555), .Z(
        n397) );
  MUX4D0 U715 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n568), .S1(n554), .Z(
        n398) );
  MUX4D0 U716 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n565), .S1(n550), .Z(
        n399) );
  MUX4D0 U717 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n565), .S1(n551), .Z(
        n401) );
  MUX4D0 U718 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n562), .S1(n551), .Z(
        n402) );
  MUX4D0 U719 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n562), .S1(n548), .Z(
        n403) );
  MUX4D0 U720 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n565), .S1(n548), .Z(
        n405) );
  MUX4D0 U721 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n565), .S1(n550), .Z(
        n406) );
  MUX4D0 U722 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n562), .S1(n551), .Z(
        n407) );
  MUX4D0 U723 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n564), .S1(n548), .Z(
        n409) );
  MUX4D0 U724 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n562), .S1(n550), .Z(
        n410) );
  MUX4D0 U725 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n562), .S1(n548), .Z(
        n411) );
  MUX4D0 U726 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n564), .S1(n548), .Z(
        n413) );
  MUX4D0 U727 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n564), .S1(n550), .Z(
        n414) );
  MUX4D0 U728 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n565), .S1(n551), .Z(
        n415) );
  MUX4D0 U729 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n564), .S1(n550), .Z(
        n417) );
  MUX4D0 U730 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n565), .S1(n551), .Z(
        n418) );
  MUX4D0 U731 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n565), .S1(n550), .Z(
        n419) );
  MUX4D0 U732 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n564), .S1(n550), .Z(
        n421) );
  MUX4D0 U733 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n565), .S1(n551), .Z(
        n422) );
  MUX4D0 U734 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n570), .S1(n556), .Z(
        n423) );
  MUX4D0 U735 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n570), .S1(n556), .Z(
        n425) );
  MUX4D0 U736 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n570), .S1(n556), .Z(
        n426) );
  MUX4D0 U737 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n570), .S1(n556), .Z(
        n427) );
  MUX4D0 U738 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n570), .S1(n556), .Z(
        n429) );
  MUX4D0 U739 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n570), .S1(n556), .Z(
        n430) );
  MUX4D0 U740 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n570), .S1(n556), .Z(
        n431) );
  MUX4D0 U741 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n570), .S1(n556), .Z(
        n433) );
  MUX4D0 U742 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n570), .S1(n556), .Z(
        n434) );
  MUX4D0 U743 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(N79), .S1(N80), .Z(
        n435) );
  MUX4D0 U744 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(N79), .S1(N80), .Z(n437)
         );
  MUX4D0 U745 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n561), .S1(n547), .Z(
        n438) );
  MUX4D0 U746 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(N79), .S1(N80), .Z(
        n439) );
  MUX4D0 U747 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(N79), .S1(N80), .Z(
        n441) );
  MUX4D0 U748 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(N79), .S1(N80), .Z(
        n442) );
  MUX4D0 U749 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(N79), .S1(N80), .Z(
        n443) );
  MUX4D0 U750 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(N79), .S1(N80), .Z(n445)
         );
  MUX4D0 U751 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n563), .S1(n549), .Z(
        n446) );
  MUX4D0 U752 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n563), .S1(n549), .Z(
        n447) );
  MUX4D0 U753 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n563), .S1(n549), .Z(
        n449) );
  MUX4D0 U754 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n563), .S1(n549), .Z(
        n450) );
  MUX4D0 U755 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n563), .S1(n549), .Z(
        n451) );
  MUX4D0 U756 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n563), .S1(n549), .Z(
        n453) );
  MUX4D0 U757 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n563), .S1(n549), .Z(
        n454) );
  MUX4D0 U758 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n563), .S1(n549), .Z(
        n455) );
  MUX4D0 U759 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n563), .S1(n547), .Z(
        n457) );
  MUX4D0 U760 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n563), .S1(n549), .Z(
        n458) );
  MUX4D0 U761 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(N79), .S1(n549), .Z(
        n459) );
  MUX4D0 U762 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n561), .S1(n549), .Z(
        n461) );
  MUX4D0 U763 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(N79), .S1(n547), .Z(n462) );
  MUX4D0 U764 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n563), .S1(n547), .Z(
        n463) );
  MUX4D0 U765 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n561), .S1(n547), .Z(
        n465) );
  MUX4D0 U766 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n561), .S1(n549), .Z(
        n466) );
  MUX4D0 U767 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n563), .S1(n547), .Z(
        n467) );
  MUX4D0 U768 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n561), .S1(n549), .Z(
        n469) );
  MUX4D0 U769 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n561), .S1(n549), .Z(
        n470) );
  MUX4D0 U770 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n564), .S1(n551), .Z(
        n471) );
  MUX4D0 U771 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n565), .S1(n551), .Z(
        n473) );
  MUX4D0 U772 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n562), .S1(n548), .Z(
        n474) );
  MUX4D0 U773 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n564), .S1(n550), .Z(
        n475) );
  MUX4D0 U774 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n564), .S1(n551), .Z(
        n477) );
  MUX4D0 U775 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n562), .S1(n548), .Z(
        n478) );
  MUX4D0 U776 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n564), .S1(n550), .Z(
        n479) );
  MUX4D0 U777 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n565), .S1(n551), .Z(
        n481) );
  MUX4D0 U778 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n562), .S1(n548), .Z(
        n482) );
  MUX4D0 U779 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n564), .S1(n548), .Z(
        n483) );
  MUX4D0 U780 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n572), .S1(n558), .Z(
        n485) );
  MUX4D0 U781 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n564), .S1(n557), .Z(
        n486) );
  MUX4D0 U782 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n571), .S1(n551), .Z(
        n487) );
  MUX4D0 U783 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n572), .S1(n557), .Z(
        n489) );
  MUX4D0 U784 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n572), .S1(n558), .Z(
        n490) );
  MUX4D0 U785 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n568), .S1(n548), .Z(
        n491) );
  MUX4D0 U786 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n572), .S1(n558), .Z(
        n493) );
  MUX4D0 U787 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n569), .S1(n558), .Z(
        n494) );
  MUX4D0 U788 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n571), .S1(n557), .Z(
        n495) );
  MUX4D0 U789 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n571), .S1(n557), .Z(
        n497) );
  MUX4D0 U790 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n571), .S1(n557), .Z(
        n498) );
  MUX4D0 U791 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n571), .S1(n557), .Z(
        n499) );
  MUX4D0 U792 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n571), .S1(n557), .Z(
        n501) );
  MUX4D0 U793 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n571), .S1(n557), .Z(
        n502) );
  MUX4D0 U794 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n571), .S1(n557), .Z(
        n503) );
  MUX4D0 U795 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n571), .S1(n557), .Z(
        n505) );
  MUX4D0 U796 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n571), .S1(n557), .Z(
        n506) );
  MUX4D0 U797 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n572), .S1(n558), .Z(
        n507) );
  MUX4D0 U798 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n572), .S1(n558), .Z(
        n509) );
  MUX4D0 U799 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n572), .S1(n558), .Z(
        n510) );
  MUX4D0 U800 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n572), .S1(n558), .Z(
        n511) );
  MUX4D0 U801 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n572), .S1(n558), .Z(
        n513) );
  MUX4D0 U802 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n572), .S1(n558), .Z(
        n514) );
  MUX4D0 U803 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n572), .S1(n558), .Z(
        n515) );
  MUX4D0 U804 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n572), .S1(n558), .Z(
        n517) );
  MUX4D0 U805 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n572), .S1(n558), .Z(
        n518) );
  MUX4D0 U806 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n573), .S1(n559), .Z(
        n519) );
  MUX4D0 U807 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n573), .S1(n559), .Z(
        n521) );
  MUX4D0 U808 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n573), .S1(n559), .Z(
        n522) );
  MUX4D0 U809 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n573), .S1(n559), .Z(
        n523) );
  MUX4D0 U810 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n573), .S1(n559), .Z(
        n525) );
  MUX4D0 U811 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n573), .S1(n559), .Z(
        n526) );
  MUX4D0 U812 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n573), .S1(n559), .Z(
        n527) );
  MUX4D0 U813 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n573), .S1(n559), .Z(
        n529) );
  MUX4D0 U814 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n573), .S1(n559), .Z(
        n530) );
  MUX4D0 U815 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n574), .S1(n560), .Z(
        n531) );
  MUX4D0 U816 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n574), .S1(n560), .Z(
        n533) );
  MUX4D0 U817 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n574), .S1(n560), .Z(
        n534) );
  MUX4D0 U818 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .I2(
        \Storage[26][32] ), .I3(\Storage[27][32] ), .S0(n574), .S1(n560), .Z(
        n536) );
  MUX4D0 U819 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .I2(
        \Storage[26][0] ), .I3(\Storage[27][0] ), .S0(n566), .S1(n552), .Z(
        n280) );
  MUX4D0 U820 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .I2(
        \Storage[26][1] ), .I3(\Storage[27][1] ), .S0(n566), .S1(n552), .Z(
        n288) );
  MUX4D0 U821 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .I2(
        \Storage[26][2] ), .I3(\Storage[27][2] ), .S0(n567), .S1(n553), .Z(
        n296) );
  MUX4D0 U822 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .I2(
        \Storage[26][3] ), .I3(\Storage[27][3] ), .S0(n568), .S1(n554), .Z(
        n304) );
  MUX4D0 U823 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .I2(
        \Storage[26][4] ), .I3(\Storage[27][4] ), .S0(n568), .S1(n554), .Z(
        n312) );
  MUX4D0 U824 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .I2(
        \Storage[26][5] ), .I3(\Storage[27][5] ), .S0(n569), .S1(n555), .Z(
        n320) );
  MUX4D0 U825 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .I2(
        \Storage[26][6] ), .I3(\Storage[27][6] ), .S0(n572), .S1(n550), .Z(
        n328) );
  MUX4D0 U826 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .I2(
        \Storage[26][7] ), .I3(\Storage[27][7] ), .S0(n574), .S1(n548), .Z(
        n336) );
  MUX4D0 U827 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .I2(
        \Storage[26][8] ), .I3(\Storage[27][8] ), .S0(n574), .S1(n560), .Z(
        n344) );
  MUX4D0 U828 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .I2(
        \Storage[26][9] ), .I3(\Storage[27][9] ), .S0(n574), .S1(n559), .Z(
        n352) );
  MUX4D0 U829 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .I2(
        \Storage[26][10] ), .I3(\Storage[27][10] ), .S0(n574), .S1(n557), .Z(
        n360) );
  MUX4D0 U830 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .I2(
        \Storage[26][11] ), .I3(\Storage[27][11] ), .S0(n565), .S1(n557), .Z(
        n368) );
  MUX4D0 U831 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .I2(
        \Storage[26][12] ), .I3(\Storage[27][12] ), .S0(n566), .S1(n555), .Z(
        n376) );
  MUX4D0 U832 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .I2(
        \Storage[26][13] ), .I3(\Storage[27][13] ), .S0(n569), .S1(n554), .Z(
        n384) );
  MUX4D0 U833 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .I2(
        \Storage[26][14] ), .I3(\Storage[27][14] ), .S0(n566), .S1(n555), .Z(
        n392) );
  MUX4D0 U834 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .I2(
        \Storage[26][15] ), .I3(\Storage[27][15] ), .S0(n564), .S1(n548), .Z(
        n400) );
  MUX4D0 U835 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .I2(
        \Storage[26][16] ), .I3(\Storage[27][16] ), .S0(n562), .S1(n548), .Z(
        n408) );
  MUX4D0 U836 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .I2(
        \Storage[26][17] ), .I3(\Storage[27][17] ), .S0(n564), .S1(n550), .Z(
        n416) );
  MUX4D0 U837 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .I2(
        \Storage[26][18] ), .I3(\Storage[27][18] ), .S0(n570), .S1(n556), .Z(
        n424) );
  MUX4D0 U838 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .I2(
        \Storage[26][19] ), .I3(\Storage[27][19] ), .S0(n570), .S1(n556), .Z(
        n432) );
  MUX4D0 U839 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .I2(
        \Storage[26][20] ), .I3(\Storage[27][20] ), .S0(N79), .S1(N80), .Z(
        n440) );
  MUX4D0 U840 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .I2(
        \Storage[26][21] ), .I3(\Storage[27][21] ), .S0(n563), .S1(n549), .Z(
        n448) );
  MUX4D0 U841 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .I2(
        \Storage[26][22] ), .I3(\Storage[27][22] ), .S0(n563), .S1(n549), .Z(
        n456) );
  MUX4D0 U842 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .I2(
        \Storage[26][23] ), .I3(\Storage[27][23] ), .S0(n563), .S1(n547), .Z(
        n464) );
  MUX4D0 U843 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .I2(
        \Storage[26][24] ), .I3(\Storage[27][24] ), .S0(n565), .S1(n550), .Z(
        n472) );
  MUX4D0 U844 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .I2(
        \Storage[26][25] ), .I3(\Storage[27][25] ), .S0(n565), .S1(n551), .Z(
        n480) );
  MUX4D0 U845 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .I2(
        \Storage[26][26] ), .I3(\Storage[27][26] ), .S0(n571), .S1(n551), .Z(
        n488) );
  MUX4D0 U846 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .I2(
        \Storage[26][27] ), .I3(\Storage[27][27] ), .S0(n571), .S1(n557), .Z(
        n496) );
  MUX4D0 U847 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .I2(
        \Storage[26][28] ), .I3(\Storage[27][28] ), .S0(n571), .S1(n557), .Z(
        n504) );
  MUX4D0 U848 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .I2(
        \Storage[26][29] ), .I3(\Storage[27][29] ), .S0(n572), .S1(n558), .Z(
        n512) );
  MUX4D0 U849 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .I2(
        \Storage[26][30] ), .I3(\Storage[27][30] ), .S0(n573), .S1(n559), .Z(
        n520) );
  MUX4D0 U850 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .I2(
        \Storage[26][31] ), .I3(\Storage[27][31] ), .S0(n573), .S1(n559), .Z(
        n528) );
  MUX4ND0 U851 ( .I0(n294), .I1(n292), .I2(n293), .I3(n291), .S0(n543), .S1(
        n545), .ZN(n213) );
  MUX4ND0 U852 ( .I0(n290), .I1(n288), .I2(n289), .I3(n287), .S0(n543), .S1(
        n545), .ZN(n214) );
  MUX4ND0 U853 ( .I0(n302), .I1(n300), .I2(n301), .I3(n299), .S0(n543), .S1(
        n545), .ZN(n215) );
  MUX4ND0 U854 ( .I0(n298), .I1(n296), .I2(n297), .I3(n295), .S0(n543), .S1(
        n545), .ZN(n216) );
  MUX4ND0 U855 ( .I0(n342), .I1(n340), .I2(n341), .I3(n339), .S0(n544), .S1(
        n546), .ZN(n217) );
  MUX4ND0 U856 ( .I0(n338), .I1(n336), .I2(n337), .I3(n335), .S0(n544), .S1(
        n546), .ZN(n218) );
  MUX4ND0 U857 ( .I0(n382), .I1(n380), .I2(n381), .I3(n379), .S0(n834), .S1(
        n833), .ZN(n219) );
  MUX4ND0 U858 ( .I0(n378), .I1(n376), .I2(n377), .I3(n375), .S0(n834), .S1(
        n833), .ZN(n220) );
  MUX4ND0 U859 ( .I0(n390), .I1(n388), .I2(n389), .I3(n387), .S0(n834), .S1(
        n833), .ZN(n221) );
  MUX4ND0 U860 ( .I0(n386), .I1(n384), .I2(n385), .I3(n383), .S0(n834), .S1(
        n833), .ZN(n222) );
  MUX4ND0 U861 ( .I0(n438), .I1(n436), .I2(n437), .I3(n435), .S0(n834), .S1(
        N81), .ZN(n223) );
  MUX4ND0 U862 ( .I0(n434), .I1(n432), .I2(n433), .I3(n431), .S0(N82), .S1(N81), .ZN(n224) );
  MUX4ND0 U863 ( .I0(n446), .I1(n444), .I2(n445), .I3(n443), .S0(N82), .S1(
        n833), .ZN(n225) );
  MUX4ND0 U864 ( .I0(n442), .I1(n440), .I2(n441), .I3(n439), .S0(N82), .S1(N81), .ZN(n226) );
  MUX4ND0 U865 ( .I0(n494), .I1(n492), .I2(n493), .I3(n491), .S0(n544), .S1(
        n546), .ZN(n227) );
  MUX4ND0 U866 ( .I0(n490), .I1(n488), .I2(n489), .I3(n487), .S0(n543), .S1(
        n545), .ZN(n228) );
  MUX4ND0 U867 ( .I0(n502), .I1(n500), .I2(n501), .I3(n499), .S0(n543), .S1(
        n545), .ZN(n229) );
  MUX4ND0 U868 ( .I0(n498), .I1(n496), .I2(n497), .I3(n495), .S0(n543), .S1(
        n545), .ZN(n230) );
  MUX4ND0 U869 ( .I0(n526), .I1(n524), .I2(n525), .I3(n523), .S0(n543), .S1(
        n545), .ZN(n231) );
  MUX4ND0 U870 ( .I0(n522), .I1(n520), .I2(n521), .I3(n519), .S0(n543), .S1(
        n545), .ZN(n232) );
  MUX4ND0 U871 ( .I0(n534), .I1(n532), .I2(n533), .I3(n531), .S0(n543), .S1(
        n545), .ZN(n233) );
  MUX4ND0 U872 ( .I0(n530), .I1(n528), .I2(n529), .I3(n527), .S0(n543), .S1(
        n545), .ZN(n234) );
  MUX4ND0 U873 ( .I0(n334), .I1(n332), .I2(n333), .I3(n331), .S0(n544), .S1(
        n546), .ZN(n235) );
  MUX4ND0 U874 ( .I0(n330), .I1(n328), .I2(n329), .I3(n327), .S0(n544), .S1(
        n546), .ZN(n236) );
  MUX4ND0 U875 ( .I0(n350), .I1(n348), .I2(n349), .I3(n347), .S0(n544), .S1(
        n546), .ZN(n237) );
  MUX4ND0 U876 ( .I0(n346), .I1(n344), .I2(n345), .I3(n343), .S0(n544), .S1(
        n546), .ZN(n238) );
  MUX4ND0 U877 ( .I0(n414), .I1(n412), .I2(n413), .I3(n411), .S0(N82), .S1(N81), .ZN(n239) );
  MUX4ND0 U878 ( .I0(n410), .I1(n408), .I2(n409), .I3(n407), .S0(n834), .S1(
        n833), .ZN(n240) );
  MUX4ND0 U879 ( .I0(n470), .I1(n468), .I2(n469), .I3(n467), .S0(n544), .S1(
        n545), .ZN(n241) );
  MUX4ND0 U880 ( .I0(n466), .I1(n464), .I2(n465), .I3(n463), .S0(n544), .S1(
        n546), .ZN(n242) );
  MUX4ND0 U881 ( .I0(n478), .I1(n476), .I2(n477), .I3(n475), .S0(n544), .S1(
        n546), .ZN(n243) );
  MUX4ND0 U882 ( .I0(n474), .I1(n472), .I2(n473), .I3(n471), .S0(n543), .S1(
        n545), .ZN(n244) );
  MUX4ND0 U883 ( .I0(n318), .I1(n316), .I2(n317), .I3(n315), .S0(n544), .S1(
        n546), .ZN(n245) );
  MUX4ND0 U884 ( .I0(n314), .I1(n312), .I2(n313), .I3(n311), .S0(n544), .S1(
        n546), .ZN(n246) );
  MUX4ND0 U885 ( .I0(n366), .I1(n364), .I2(n365), .I3(n363), .S0(n834), .S1(
        n833), .ZN(n247) );
  MUX4ND0 U886 ( .I0(n362), .I1(n360), .I2(n361), .I3(n359), .S0(n834), .S1(
        n833), .ZN(n248) );
  MUX4ND0 U887 ( .I0(n398), .I1(n396), .I2(n397), .I3(n395), .S0(n834), .S1(
        n833), .ZN(n249) );
  MUX4ND0 U888 ( .I0(n394), .I1(n392), .I2(n393), .I3(n391), .S0(n834), .S1(
        n833), .ZN(n250) );
  MUX4ND0 U889 ( .I0(n454), .I1(n452), .I2(n453), .I3(n451), .S0(n834), .S1(
        n833), .ZN(n251) );
  MUX4ND0 U890 ( .I0(n450), .I1(n448), .I2(n449), .I3(n447), .S0(n834), .S1(
        n833), .ZN(n252) );
  MUX4ND0 U891 ( .I0(n510), .I1(n508), .I2(n509), .I3(n507), .S0(n543), .S1(
        n545), .ZN(n253) );
  MUX4ND0 U892 ( .I0(n506), .I1(n504), .I2(n505), .I3(n503), .S0(n543), .S1(
        n545), .ZN(n254) );
  MUX4ND0 U893 ( .I0(n286), .I1(n284), .I2(n285), .I3(n283), .S0(n543), .S1(
        n545), .ZN(n255) );
  MUX4ND0 U894 ( .I0(n282), .I1(n280), .I2(n281), .I3(n279), .S0(n543), .S1(
        n545), .ZN(n256) );
  MUX4ND0 U895 ( .I0(n310), .I1(n308), .I2(n309), .I3(n307), .S0(n544), .S1(
        n546), .ZN(n257) );
  MUX4ND0 U896 ( .I0(n306), .I1(n304), .I2(n305), .I3(n303), .S0(n544), .S1(
        n546), .ZN(n258) );
  MUX4ND0 U897 ( .I0(n326), .I1(n324), .I2(n325), .I3(n323), .S0(n544), .S1(
        n546), .ZN(n259) );
  MUX4ND0 U898 ( .I0(n322), .I1(n320), .I2(n321), .I3(n319), .S0(n544), .S1(
        n546), .ZN(n260) );
  MUX4ND0 U899 ( .I0(n358), .I1(n356), .I2(n357), .I3(n355), .S0(n834), .S1(
        n833), .ZN(n261) );
  MUX4ND0 U900 ( .I0(n354), .I1(n352), .I2(n353), .I3(n351), .S0(n834), .S1(
        n833), .ZN(n262) );
  MUX4ND0 U901 ( .I0(n374), .I1(n372), .I2(n373), .I3(n371), .S0(n834), .S1(
        n833), .ZN(n263) );
  MUX4ND0 U902 ( .I0(n370), .I1(n368), .I2(n369), .I3(n367), .S0(n834), .S1(
        n833), .ZN(n264) );
  MUX4ND0 U903 ( .I0(n406), .I1(n404), .I2(n405), .I3(n403), .S0(N82), .S1(N81), .ZN(n265) );
  MUX4ND0 U904 ( .I0(n402), .I1(n400), .I2(n401), .I3(n399), .S0(N82), .S1(N81), .ZN(n266) );
  MUX4ND0 U905 ( .I0(n422), .I1(n420), .I2(n421), .I3(n419), .S0(N82), .S1(N81), .ZN(n267) );
  MUX4ND0 U906 ( .I0(n418), .I1(n416), .I2(n417), .I3(n415), .S0(N82), .S1(N81), .ZN(n268) );
  MUX4ND0 U907 ( .I0(n430), .I1(n428), .I2(n429), .I3(n427), .S0(N82), .S1(N81), .ZN(n269) );
  MUX4ND0 U908 ( .I0(n426), .I1(n424), .I2(n425), .I3(n423), .S0(N82), .S1(N81), .ZN(n270) );
  MUX4ND0 U909 ( .I0(n462), .I1(n460), .I2(n461), .I3(n459), .S0(n544), .S1(
        n546), .ZN(n271) );
  MUX4ND0 U910 ( .I0(n458), .I1(n456), .I2(n457), .I3(n455), .S0(n544), .S1(
        n546), .ZN(n272) );
  MUX4ND0 U911 ( .I0(n486), .I1(n484), .I2(n485), .I3(n483), .S0(n544), .S1(
        n546), .ZN(n273) );
  MUX4ND0 U912 ( .I0(n482), .I1(n480), .I2(n481), .I3(n479), .S0(n543), .S1(
        n546), .ZN(n274) );
  MUX4ND0 U913 ( .I0(n518), .I1(n516), .I2(n517), .I3(n515), .S0(n543), .S1(
        n545), .ZN(n275) );
  MUX4ND0 U914 ( .I0(n514), .I1(n512), .I2(n513), .I3(n511), .S0(n543), .S1(
        n545), .ZN(n276) );
  MUX2ND0 U915 ( .I0(n277), .I1(n278), .S(n835), .ZN(N32) );
  MUX4ND0 U916 ( .I0(n542), .I1(n540), .I2(n541), .I3(n539), .S0(n544), .S1(
        n545), .ZN(n277) );
  MUX4ND0 U917 ( .I0(n538), .I1(n536), .I2(n537), .I3(n535), .S0(n543), .S1(
        n546), .ZN(n278) );
  BUFFD1 U918 ( .I(N81), .Z(n833) );
  BUFFD1 U919 ( .I(N82), .Z(n834) );
  ND3D1 U920 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U921 ( .A1(AddrW[4]), .A2(n76), .A3(Write), .ZN(n70) );
  ND3D1 U922 ( .A1(n76), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U923 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U924 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n75) );
  ND3D1 U925 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  ND3D1 U926 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n73) );
  ND3D1 U927 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U928 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n74) );
  ND3D1 U929 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  ND3D1 U930 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  INVD1 U931 ( .I(AddrW[2]), .ZN(n105) );
  INVD1 U932 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U933 ( .I(AddrW[1]), .ZN(n106) );
  INVD1 U934 ( .I(AddrW[4]), .ZN(n102) );
  INVD1 U935 ( .I(AddrW[3]), .ZN(n76) );
  INVD1 U936 ( .I(Read), .ZN(n832) );
  AN2D1 U937 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  AN2D1 U938 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U5 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U6 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n6, \carry[4] , \carry[3] , \carry[2] , n3, n4, n5;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  DEL2 U5 ( .I(n5), .Z(SUM[0]) );
  INVD0 U6 ( .I(A[0]), .ZN(n5) );
  DEL4 U7 ( .I(n3), .Z(SUM[4]) );
  DEL4 U8 ( .I(n4), .Z(n3) );
  DEL4 U9 ( .I(n6), .Z(n4) );
  XOR2D0 U10 ( .A1(\carry[4] ), .A2(A[4]), .Z(n6) );
endmodule

