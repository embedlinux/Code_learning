
module Deserializer ( ParOut, ParValid, DecoderParClk, FIFOEmpty, FIFOFull, 
        ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   ParValidDecode, SerialClk, SerRxToDecode, n2, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid5_DWid32 FIFO_U1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(n871), .WriteIn(ParValidDecode), 
        .ClkR(n870), .ClkW(DecoderParClk), .Reseter(n485) );
  DesDecoder_DWid32 DesDecoder_U1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n869) );
  SerialRx SerialRx_U1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n869) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(n4), .CP(n870), .CDN(n2), .Q(ParOut[31]) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(n31), .CP(ParOutClk), .CDN(n2), .Q(ParOut[30])
         );
  DFCNQD1 \ParBuf_reg[29]  ( .D(n58), .CP(ParOutClk), .CDN(n2), .Q(ParOut[29])
         );
  DFCNQD1 \ParBuf_reg[28]  ( .D(n85), .CP(ParOutClk), .CDN(n2), .Q(ParOut[28])
         );
  DFCNQD1 \ParBuf_reg[27]  ( .D(n112), .CP(n870), .CDN(n2), .Q(ParOut[27]) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(n139), .CP(ParOutClk), .CDN(n2), .Q(ParOut[26]) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(n166), .CP(n870), .CDN(n2), .Q(ParOut[25]) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(n193), .CP(ParOutClk), .CDN(n2), .Q(ParOut[24]) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(n586), .CP(n870), .CDN(n2), .Q(ParOut[23]) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(n595), .CP(ParOutClk), .CDN(n2), .Q(ParOut[22]) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(n477), .CP(n870), .CDN(n2), .Q(ParOut[21]) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(n220), .CP(ParOutClk), .CDN(n2), .Q(ParOut[20]) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(n247), .CP(n870), .CDN(n2), .Q(ParOut[19]) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(n629), .CP(ParOutClk), .CDN(n2), .Q(ParOut[18]) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(n638), .CP(n870), .CDN(n2), .Q(ParOut[17]) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(n479), .CP(ParOutClk), .CDN(n2), .Q(ParOut[16]) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(n274), .CP(n870), .CDN(n2), .Q(ParOut[15]) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(n301), .CP(ParOutClk), .CDN(n2), .Q(ParOut[14]) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(n672), .CP(n870), .CDN(n2), .Q(ParOut[13]) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(n681), .CP(ParOutClk), .CDN(n2), .Q(ParOut[12]) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(n481), .CP(n870), .CDN(n2), .Q(ParOut[11]) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(n328), .CP(ParOutClk), .CDN(n2), .Q(ParOut[10]) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(n355), .CP(n870), .CDN(n2), .Q(ParOut[9]) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(n715), .CP(ParOutClk), .CDN(n2), .Q(ParOut[8])
         );
  DFCNQD1 \ParBuf_reg[7]  ( .D(n724), .CP(n870), .CDN(n2), .Q(ParOut[7]) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(n733), .CP(ParOutClk), .CDN(n2), .Q(ParOut[6])
         );
  DFCNQD1 \ParBuf_reg[5]  ( .D(n483), .CP(n870), .CDN(n2), .Q(ParOut[5]) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(n382), .CP(ParOutClk), .CDN(n2), .Q(ParOut[4])
         );
  DFCNQD1 \ParBuf_reg[3]  ( .D(n409), .CP(n870), .CDN(n2), .Q(ParOut[3]) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(n767), .CP(ParOutClk), .CDN(n2), .Q(ParOut[2])
         );
  DFCNQD1 \ParBuf_reg[1]  ( .D(n776), .CP(n870), .CDN(n2), .Q(ParOut[1]) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(n785), .CP(ParOutClk), .CDN(n2), .Q(ParOut[0])
         );
  DFCNQD1 ParValidr_reg ( .D(n436), .CP(n870), .CDN(n2), .Q(ParValid) );
  INVD5 U38 ( .I(n513), .ZN(n514) );
  BUFFD0 U39 ( .I(n5), .Z(n4) );
  BUFFD0 U40 ( .I(n6), .Z(n5) );
  BUFFD0 U41 ( .I(n7), .Z(n6) );
  BUFFD0 U42 ( .I(n8), .Z(n7) );
  BUFFD0 U43 ( .I(n9), .Z(n8) );
  BUFFD0 U44 ( .I(n10), .Z(n9) );
  BUFFD0 U45 ( .I(n11), .Z(n10) );
  BUFFD0 U46 ( .I(n12), .Z(n11) );
  BUFFD0 U47 ( .I(n13), .Z(n12) );
  BUFFD0 U48 ( .I(n14), .Z(n13) );
  BUFFD0 U49 ( .I(n15), .Z(n14) );
  BUFFD0 U50 ( .I(n16), .Z(n15) );
  BUFFD0 U51 ( .I(n17), .Z(n16) );
  BUFFD0 U52 ( .I(n18), .Z(n17) );
  BUFFD0 U53 ( .I(n19), .Z(n18) );
  BUFFD0 U54 ( .I(n20), .Z(n19) );
  BUFFD0 U55 ( .I(n21), .Z(n20) );
  BUFFD0 U56 ( .I(n22), .Z(n21) );
  BUFFD0 U57 ( .I(n23), .Z(n22) );
  BUFFD0 U58 ( .I(n24), .Z(n23) );
  BUFFD0 U59 ( .I(n25), .Z(n24) );
  BUFFD0 U60 ( .I(n26), .Z(n25) );
  BUFFD0 U61 ( .I(n27), .Z(n26) );
  BUFFD0 U62 ( .I(n28), .Z(n27) );
  BUFFD0 U63 ( .I(n512), .Z(n28) );
  BUFFD0 U64 ( .I(n459), .Z(n29) );
  BUFFD0 U65 ( .I(n29), .Z(n30) );
  INVD5 U66 ( .I(n522), .ZN(n523) );
  BUFFD0 U67 ( .I(n32), .Z(n31) );
  BUFFD0 U68 ( .I(n33), .Z(n32) );
  BUFFD0 U69 ( .I(n34), .Z(n33) );
  BUFFD0 U70 ( .I(n35), .Z(n34) );
  BUFFD0 U71 ( .I(n36), .Z(n35) );
  BUFFD0 U72 ( .I(n37), .Z(n36) );
  BUFFD0 U73 ( .I(n38), .Z(n37) );
  BUFFD0 U74 ( .I(n39), .Z(n38) );
  BUFFD0 U75 ( .I(n40), .Z(n39) );
  BUFFD0 U76 ( .I(n41), .Z(n40) );
  BUFFD0 U77 ( .I(n42), .Z(n41) );
  BUFFD0 U78 ( .I(n43), .Z(n42) );
  BUFFD0 U79 ( .I(n44), .Z(n43) );
  BUFFD0 U80 ( .I(n45), .Z(n44) );
  BUFFD0 U81 ( .I(n521), .Z(n45) );
  BUFFD0 U82 ( .I(n458), .Z(n46) );
  BUFFD0 U83 ( .I(n46), .Z(n47) );
  BUFFD0 U84 ( .I(n47), .Z(n48) );
  BUFFD0 U85 ( .I(n48), .Z(n49) );
  BUFFD0 U86 ( .I(n49), .Z(n50) );
  BUFFD0 U87 ( .I(n50), .Z(n51) );
  BUFFD0 U88 ( .I(n51), .Z(n52) );
  BUFFD0 U89 ( .I(n52), .Z(n53) );
  BUFFD0 U90 ( .I(n53), .Z(n54) );
  BUFFD0 U91 ( .I(n54), .Z(n55) );
  BUFFD0 U92 ( .I(n55), .Z(n56) );
  BUFFD0 U93 ( .I(n56), .Z(n57) );
  INVD5 U94 ( .I(n531), .ZN(n532) );
  BUFFD0 U95 ( .I(n59), .Z(n58) );
  BUFFD0 U96 ( .I(n60), .Z(n59) );
  BUFFD0 U97 ( .I(n61), .Z(n60) );
  BUFFD0 U98 ( .I(n62), .Z(n61) );
  BUFFD0 U99 ( .I(n63), .Z(n62) );
  BUFFD0 U100 ( .I(n64), .Z(n63) );
  BUFFD0 U101 ( .I(n65), .Z(n64) );
  BUFFD0 U102 ( .I(n66), .Z(n65) );
  BUFFD0 U103 ( .I(n67), .Z(n66) );
  BUFFD0 U104 ( .I(n68), .Z(n67) );
  BUFFD0 U105 ( .I(n69), .Z(n68) );
  BUFFD0 U106 ( .I(n70), .Z(n69) );
  BUFFD0 U107 ( .I(n71), .Z(n70) );
  BUFFD0 U108 ( .I(n72), .Z(n71) );
  BUFFD0 U109 ( .I(n530), .Z(n72) );
  BUFFD0 U110 ( .I(n457), .Z(n73) );
  BUFFD0 U111 ( .I(n73), .Z(n74) );
  BUFFD0 U112 ( .I(n74), .Z(n75) );
  BUFFD0 U113 ( .I(n75), .Z(n76) );
  BUFFD0 U114 ( .I(n76), .Z(n77) );
  BUFFD0 U115 ( .I(n77), .Z(n78) );
  BUFFD0 U116 ( .I(n78), .Z(n79) );
  BUFFD0 U117 ( .I(n79), .Z(n80) );
  BUFFD0 U118 ( .I(n80), .Z(n81) );
  BUFFD0 U119 ( .I(n81), .Z(n82) );
  BUFFD0 U120 ( .I(n82), .Z(n83) );
  BUFFD0 U121 ( .I(n83), .Z(n84) );
  INVD5 U122 ( .I(n540), .ZN(n541) );
  BUFFD0 U123 ( .I(n86), .Z(n85) );
  BUFFD0 U124 ( .I(n87), .Z(n86) );
  BUFFD0 U125 ( .I(n88), .Z(n87) );
  BUFFD0 U126 ( .I(n89), .Z(n88) );
  BUFFD0 U127 ( .I(n90), .Z(n89) );
  BUFFD0 U128 ( .I(n91), .Z(n90) );
  BUFFD0 U129 ( .I(n92), .Z(n91) );
  BUFFD0 U130 ( .I(n93), .Z(n92) );
  BUFFD0 U131 ( .I(n94), .Z(n93) );
  BUFFD0 U132 ( .I(n95), .Z(n94) );
  BUFFD0 U133 ( .I(n96), .Z(n95) );
  BUFFD0 U134 ( .I(n97), .Z(n96) );
  BUFFD0 U135 ( .I(n98), .Z(n97) );
  BUFFD0 U136 ( .I(n99), .Z(n98) );
  BUFFD0 U137 ( .I(n539), .Z(n99) );
  BUFFD0 U138 ( .I(n456), .Z(n100) );
  BUFFD0 U139 ( .I(n100), .Z(n101) );
  BUFFD0 U140 ( .I(n101), .Z(n102) );
  BUFFD0 U141 ( .I(n102), .Z(n103) );
  BUFFD0 U142 ( .I(n103), .Z(n104) );
  BUFFD0 U143 ( .I(n104), .Z(n105) );
  BUFFD0 U144 ( .I(n105), .Z(n106) );
  BUFFD0 U145 ( .I(n106), .Z(n107) );
  BUFFD0 U146 ( .I(n107), .Z(n108) );
  BUFFD0 U147 ( .I(n108), .Z(n109) );
  BUFFD0 U148 ( .I(n109), .Z(n110) );
  BUFFD0 U149 ( .I(n110), .Z(n111) );
  INVD5 U150 ( .I(n549), .ZN(n550) );
  BUFFD0 U151 ( .I(n113), .Z(n112) );
  BUFFD0 U152 ( .I(n114), .Z(n113) );
  BUFFD0 U153 ( .I(n115), .Z(n114) );
  BUFFD0 U154 ( .I(n116), .Z(n115) );
  BUFFD0 U155 ( .I(n117), .Z(n116) );
  BUFFD0 U156 ( .I(n118), .Z(n117) );
  BUFFD0 U157 ( .I(n119), .Z(n118) );
  BUFFD0 U158 ( .I(n120), .Z(n119) );
  BUFFD0 U159 ( .I(n121), .Z(n120) );
  BUFFD0 U160 ( .I(n122), .Z(n121) );
  BUFFD0 U161 ( .I(n123), .Z(n122) );
  BUFFD0 U162 ( .I(n124), .Z(n123) );
  BUFFD0 U163 ( .I(n125), .Z(n124) );
  BUFFD0 U164 ( .I(n126), .Z(n125) );
  BUFFD0 U165 ( .I(n127), .Z(n126) );
  BUFFD0 U166 ( .I(n128), .Z(n127) );
  BUFFD0 U167 ( .I(n129), .Z(n128) );
  BUFFD0 U168 ( .I(n130), .Z(n129) );
  BUFFD0 U169 ( .I(n131), .Z(n130) );
  BUFFD0 U170 ( .I(n132), .Z(n131) );
  BUFFD0 U171 ( .I(n133), .Z(n132) );
  BUFFD0 U172 ( .I(n134), .Z(n133) );
  BUFFD0 U173 ( .I(n135), .Z(n134) );
  BUFFD0 U174 ( .I(n136), .Z(n135) );
  BUFFD0 U175 ( .I(n548), .Z(n136) );
  BUFFD0 U176 ( .I(n455), .Z(n137) );
  BUFFD0 U177 ( .I(n137), .Z(n138) );
  INVD5 U178 ( .I(n558), .ZN(n559) );
  BUFFD0 U179 ( .I(n140), .Z(n139) );
  BUFFD0 U180 ( .I(n141), .Z(n140) );
  BUFFD0 U181 ( .I(n142), .Z(n141) );
  BUFFD0 U182 ( .I(n143), .Z(n142) );
  BUFFD0 U183 ( .I(n144), .Z(n143) );
  BUFFD0 U184 ( .I(n145), .Z(n144) );
  BUFFD0 U185 ( .I(n146), .Z(n145) );
  BUFFD0 U186 ( .I(n147), .Z(n146) );
  BUFFD0 U187 ( .I(n148), .Z(n147) );
  BUFFD0 U188 ( .I(n149), .Z(n148) );
  BUFFD0 U189 ( .I(n150), .Z(n149) );
  BUFFD0 U190 ( .I(n151), .Z(n150) );
  BUFFD0 U191 ( .I(n152), .Z(n151) );
  BUFFD0 U192 ( .I(n153), .Z(n152) );
  BUFFD0 U193 ( .I(n557), .Z(n153) );
  BUFFD0 U194 ( .I(n454), .Z(n154) );
  BUFFD0 U195 ( .I(n154), .Z(n155) );
  BUFFD0 U196 ( .I(n155), .Z(n156) );
  BUFFD0 U197 ( .I(n156), .Z(n157) );
  BUFFD0 U198 ( .I(n157), .Z(n158) );
  BUFFD0 U199 ( .I(n158), .Z(n159) );
  BUFFD0 U200 ( .I(n159), .Z(n160) );
  BUFFD0 U201 ( .I(n160), .Z(n161) );
  BUFFD0 U202 ( .I(n161), .Z(n162) );
  BUFFD0 U203 ( .I(n162), .Z(n163) );
  BUFFD0 U204 ( .I(n163), .Z(n164) );
  BUFFD0 U205 ( .I(n164), .Z(n165) );
  INVD5 U206 ( .I(n567), .ZN(n568) );
  BUFFD0 U207 ( .I(n167), .Z(n166) );
  BUFFD0 U208 ( .I(n168), .Z(n167) );
  BUFFD0 U209 ( .I(n169), .Z(n168) );
  BUFFD0 U210 ( .I(n170), .Z(n169) );
  BUFFD0 U211 ( .I(n171), .Z(n170) );
  BUFFD0 U212 ( .I(n172), .Z(n171) );
  BUFFD0 U213 ( .I(n173), .Z(n172) );
  BUFFD0 U214 ( .I(n174), .Z(n173) );
  BUFFD0 U215 ( .I(n175), .Z(n174) );
  BUFFD0 U216 ( .I(n176), .Z(n175) );
  BUFFD0 U217 ( .I(n177), .Z(n176) );
  BUFFD0 U218 ( .I(n178), .Z(n177) );
  BUFFD0 U219 ( .I(n179), .Z(n178) );
  BUFFD0 U220 ( .I(n180), .Z(n179) );
  BUFFD0 U221 ( .I(n181), .Z(n180) );
  BUFFD0 U222 ( .I(n182), .Z(n181) );
  BUFFD0 U223 ( .I(n183), .Z(n182) );
  BUFFD0 U224 ( .I(n184), .Z(n183) );
  BUFFD0 U225 ( .I(n185), .Z(n184) );
  BUFFD0 U226 ( .I(n186), .Z(n185) );
  BUFFD0 U227 ( .I(n187), .Z(n186) );
  BUFFD0 U228 ( .I(n188), .Z(n187) );
  BUFFD0 U229 ( .I(n189), .Z(n188) );
  BUFFD0 U230 ( .I(n190), .Z(n189) );
  BUFFD0 U231 ( .I(n566), .Z(n190) );
  BUFFD0 U232 ( .I(n453), .Z(n191) );
  BUFFD0 U233 ( .I(n191), .Z(n192) );
  INVD5 U234 ( .I(n576), .ZN(n577) );
  BUFFD0 U235 ( .I(n194), .Z(n193) );
  BUFFD0 U236 ( .I(n195), .Z(n194) );
  BUFFD0 U237 ( .I(n196), .Z(n195) );
  BUFFD0 U238 ( .I(n197), .Z(n196) );
  BUFFD0 U239 ( .I(n198), .Z(n197) );
  BUFFD0 U240 ( .I(n199), .Z(n198) );
  BUFFD0 U241 ( .I(n200), .Z(n199) );
  BUFFD0 U242 ( .I(n201), .Z(n200) );
  BUFFD0 U243 ( .I(n202), .Z(n201) );
  BUFFD0 U244 ( .I(n203), .Z(n202) );
  BUFFD0 U245 ( .I(n204), .Z(n203) );
  BUFFD0 U246 ( .I(n205), .Z(n204) );
  BUFFD0 U247 ( .I(n206), .Z(n205) );
  BUFFD0 U248 ( .I(n207), .Z(n206) );
  BUFFD0 U249 ( .I(n575), .Z(n207) );
  BUFFD0 U250 ( .I(n452), .Z(n208) );
  BUFFD0 U251 ( .I(n208), .Z(n209) );
  BUFFD0 U252 ( .I(n209), .Z(n210) );
  BUFFD0 U253 ( .I(n210), .Z(n211) );
  BUFFD0 U254 ( .I(n211), .Z(n212) );
  BUFFD0 U255 ( .I(n212), .Z(n213) );
  BUFFD0 U256 ( .I(n213), .Z(n214) );
  BUFFD0 U257 ( .I(n214), .Z(n215) );
  BUFFD0 U258 ( .I(n215), .Z(n216) );
  BUFFD0 U259 ( .I(n216), .Z(n217) );
  BUFFD0 U260 ( .I(n217), .Z(n218) );
  BUFFD0 U261 ( .I(n218), .Z(n219) );
  CKND8 U262 ( .CLK(n476), .CN(n584) );
  CKND2D0 U263 ( .A1(FIFO_Out[23]), .A2(n871), .ZN(n476) );
  CKND8 U264 ( .CLK(n475), .CN(n593) );
  CKND2D0 U265 ( .A1(FIFO_Out[22]), .A2(n871), .ZN(n475) );
  CKND2D0 U266 ( .A1(FIFO_Out[21]), .A2(n871), .ZN(n474) );
  INVD5 U267 ( .I(n610), .ZN(n611) );
  BUFFD0 U268 ( .I(n221), .Z(n220) );
  BUFFD0 U269 ( .I(n222), .Z(n221) );
  BUFFD0 U270 ( .I(n223), .Z(n222) );
  BUFFD0 U271 ( .I(n224), .Z(n223) );
  BUFFD0 U272 ( .I(n225), .Z(n224) );
  BUFFD0 U273 ( .I(n226), .Z(n225) );
  BUFFD0 U274 ( .I(n227), .Z(n226) );
  BUFFD0 U275 ( .I(n228), .Z(n227) );
  BUFFD0 U276 ( .I(n229), .Z(n228) );
  BUFFD0 U277 ( .I(n230), .Z(n229) );
  BUFFD0 U278 ( .I(n231), .Z(n230) );
  BUFFD0 U279 ( .I(n232), .Z(n231) );
  BUFFD0 U280 ( .I(n233), .Z(n232) );
  BUFFD0 U281 ( .I(n234), .Z(n233) );
  BUFFD0 U282 ( .I(n609), .Z(n234) );
  BUFFD0 U283 ( .I(n451), .Z(n235) );
  BUFFD0 U284 ( .I(n235), .Z(n236) );
  BUFFD0 U285 ( .I(n236), .Z(n237) );
  BUFFD0 U286 ( .I(n237), .Z(n238) );
  BUFFD0 U287 ( .I(n238), .Z(n239) );
  BUFFD0 U288 ( .I(n239), .Z(n240) );
  BUFFD0 U289 ( .I(n240), .Z(n241) );
  BUFFD0 U290 ( .I(n241), .Z(n242) );
  BUFFD0 U291 ( .I(n242), .Z(n243) );
  BUFFD0 U292 ( .I(n243), .Z(n244) );
  BUFFD0 U293 ( .I(n244), .Z(n245) );
  BUFFD0 U294 ( .I(n245), .Z(n246) );
  INVD5 U295 ( .I(n619), .ZN(n620) );
  BUFFD0 U296 ( .I(n248), .Z(n247) );
  BUFFD0 U297 ( .I(n249), .Z(n248) );
  BUFFD0 U298 ( .I(n250), .Z(n249) );
  BUFFD0 U299 ( .I(n251), .Z(n250) );
  BUFFD0 U300 ( .I(n252), .Z(n251) );
  BUFFD0 U301 ( .I(n253), .Z(n252) );
  BUFFD0 U302 ( .I(n254), .Z(n253) );
  BUFFD0 U303 ( .I(n255), .Z(n254) );
  BUFFD0 U304 ( .I(n256), .Z(n255) );
  BUFFD0 U305 ( .I(n257), .Z(n256) );
  BUFFD0 U306 ( .I(n258), .Z(n257) );
  BUFFD0 U307 ( .I(n259), .Z(n258) );
  BUFFD0 U308 ( .I(n260), .Z(n259) );
  BUFFD0 U309 ( .I(n261), .Z(n260) );
  BUFFD0 U310 ( .I(n262), .Z(n261) );
  BUFFD0 U311 ( .I(n263), .Z(n262) );
  BUFFD0 U312 ( .I(n264), .Z(n263) );
  BUFFD0 U313 ( .I(n265), .Z(n264) );
  BUFFD0 U314 ( .I(n266), .Z(n265) );
  BUFFD0 U315 ( .I(n267), .Z(n266) );
  BUFFD0 U316 ( .I(n268), .Z(n267) );
  BUFFD0 U317 ( .I(n269), .Z(n268) );
  BUFFD0 U318 ( .I(n270), .Z(n269) );
  BUFFD0 U319 ( .I(n271), .Z(n270) );
  BUFFD0 U320 ( .I(n618), .Z(n271) );
  BUFFD0 U321 ( .I(n450), .Z(n272) );
  BUFFD0 U322 ( .I(n272), .Z(n273) );
  CKND8 U323 ( .CLK(n473), .CN(n627) );
  CKND2D0 U324 ( .A1(FIFO_Out[18]), .A2(n871), .ZN(n473) );
  CKND8 U325 ( .CLK(n472), .CN(n636) );
  CKND2D0 U326 ( .A1(FIFO_Out[17]), .A2(n871), .ZN(n472) );
  CKBD0 U327 ( .CLK(n480), .C(n479) );
  CKBD0 U328 ( .CLK(n646), .C(n480) );
  CKND2D0 U329 ( .A1(FIFO_Out[16]), .A2(n871), .ZN(n471) );
  INVD5 U330 ( .I(n653), .ZN(n654) );
  BUFFD0 U331 ( .I(n275), .Z(n274) );
  BUFFD0 U332 ( .I(n276), .Z(n275) );
  BUFFD0 U333 ( .I(n277), .Z(n276) );
  BUFFD0 U334 ( .I(n278), .Z(n277) );
  BUFFD0 U335 ( .I(n279), .Z(n278) );
  BUFFD0 U336 ( .I(n280), .Z(n279) );
  BUFFD0 U337 ( .I(n281), .Z(n280) );
  BUFFD0 U338 ( .I(n282), .Z(n281) );
  BUFFD0 U339 ( .I(n283), .Z(n282) );
  BUFFD0 U340 ( .I(n284), .Z(n283) );
  BUFFD0 U341 ( .I(n285), .Z(n284) );
  BUFFD0 U342 ( .I(n286), .Z(n285) );
  BUFFD0 U343 ( .I(n287), .Z(n286) );
  BUFFD0 U344 ( .I(n288), .Z(n287) );
  BUFFD0 U345 ( .I(n289), .Z(n288) );
  BUFFD0 U346 ( .I(n290), .Z(n289) );
  BUFFD0 U347 ( .I(n291), .Z(n290) );
  BUFFD0 U348 ( .I(n292), .Z(n291) );
  BUFFD0 U349 ( .I(n293), .Z(n292) );
  BUFFD0 U350 ( .I(n294), .Z(n293) );
  BUFFD0 U351 ( .I(n295), .Z(n294) );
  BUFFD0 U352 ( .I(n296), .Z(n295) );
  BUFFD0 U353 ( .I(n297), .Z(n296) );
  BUFFD0 U354 ( .I(n298), .Z(n297) );
  BUFFD0 U355 ( .I(n652), .Z(n298) );
  BUFFD0 U356 ( .I(n449), .Z(n299) );
  BUFFD0 U357 ( .I(n299), .Z(n300) );
  INVD5 U358 ( .I(n662), .ZN(n663) );
  BUFFD0 U359 ( .I(n302), .Z(n301) );
  BUFFD0 U360 ( .I(n303), .Z(n302) );
  BUFFD0 U361 ( .I(n304), .Z(n303) );
  BUFFD0 U362 ( .I(n305), .Z(n304) );
  BUFFD0 U363 ( .I(n306), .Z(n305) );
  BUFFD0 U364 ( .I(n307), .Z(n306) );
  BUFFD0 U365 ( .I(n308), .Z(n307) );
  BUFFD0 U366 ( .I(n309), .Z(n308) );
  BUFFD0 U367 ( .I(n310), .Z(n309) );
  BUFFD0 U368 ( .I(n311), .Z(n310) );
  BUFFD0 U369 ( .I(n312), .Z(n311) );
  BUFFD0 U370 ( .I(n313), .Z(n312) );
  BUFFD0 U371 ( .I(n314), .Z(n313) );
  BUFFD0 U372 ( .I(n315), .Z(n314) );
  BUFFD0 U373 ( .I(n661), .Z(n315) );
  BUFFD0 U374 ( .I(n448), .Z(n316) );
  BUFFD0 U375 ( .I(n316), .Z(n317) );
  BUFFD0 U376 ( .I(n317), .Z(n318) );
  BUFFD0 U377 ( .I(n318), .Z(n319) );
  BUFFD0 U378 ( .I(n319), .Z(n320) );
  BUFFD0 U379 ( .I(n320), .Z(n321) );
  BUFFD0 U380 ( .I(n321), .Z(n322) );
  BUFFD0 U381 ( .I(n322), .Z(n323) );
  BUFFD0 U382 ( .I(n323), .Z(n324) );
  BUFFD0 U383 ( .I(n324), .Z(n325) );
  BUFFD0 U384 ( .I(n325), .Z(n326) );
  BUFFD0 U385 ( .I(n326), .Z(n327) );
  CKND8 U386 ( .CLK(n470), .CN(n670) );
  CKND2D0 U387 ( .A1(FIFO_Out[13]), .A2(n871), .ZN(n470) );
  CKND8 U388 ( .CLK(n469), .CN(n679) );
  CKND2D0 U389 ( .A1(FIFO_Out[12]), .A2(n871), .ZN(n469) );
  CKND2D0 U390 ( .A1(FIFO_Out[11]), .A2(n871), .ZN(n468) );
  INVD5 U391 ( .I(n696), .ZN(n697) );
  BUFFD0 U392 ( .I(n329), .Z(n328) );
  BUFFD0 U393 ( .I(n330), .Z(n329) );
  BUFFD0 U394 ( .I(n331), .Z(n330) );
  BUFFD0 U395 ( .I(n332), .Z(n331) );
  BUFFD0 U396 ( .I(n333), .Z(n332) );
  BUFFD0 U397 ( .I(n334), .Z(n333) );
  BUFFD0 U398 ( .I(n335), .Z(n334) );
  BUFFD0 U399 ( .I(n336), .Z(n335) );
  BUFFD0 U400 ( .I(n337), .Z(n336) );
  BUFFD0 U401 ( .I(n338), .Z(n337) );
  BUFFD0 U402 ( .I(n339), .Z(n338) );
  BUFFD0 U403 ( .I(n340), .Z(n339) );
  BUFFD0 U404 ( .I(n341), .Z(n340) );
  BUFFD0 U405 ( .I(n342), .Z(n341) );
  BUFFD0 U406 ( .I(n695), .Z(n342) );
  BUFFD0 U407 ( .I(n447), .Z(n343) );
  BUFFD0 U408 ( .I(n343), .Z(n344) );
  BUFFD0 U409 ( .I(n344), .Z(n345) );
  BUFFD0 U410 ( .I(n345), .Z(n346) );
  BUFFD0 U411 ( .I(n346), .Z(n347) );
  BUFFD0 U412 ( .I(n347), .Z(n348) );
  BUFFD0 U413 ( .I(n348), .Z(n349) );
  BUFFD0 U414 ( .I(n349), .Z(n350) );
  BUFFD0 U415 ( .I(n350), .Z(n351) );
  BUFFD0 U416 ( .I(n351), .Z(n352) );
  BUFFD0 U417 ( .I(n352), .Z(n353) );
  BUFFD0 U418 ( .I(n353), .Z(n354) );
  INVD5 U419 ( .I(n705), .ZN(n706) );
  BUFFD0 U420 ( .I(n356), .Z(n355) );
  BUFFD0 U421 ( .I(n357), .Z(n356) );
  BUFFD0 U422 ( .I(n358), .Z(n357) );
  BUFFD0 U423 ( .I(n359), .Z(n358) );
  BUFFD0 U424 ( .I(n360), .Z(n359) );
  BUFFD0 U425 ( .I(n361), .Z(n360) );
  BUFFD0 U426 ( .I(n362), .Z(n361) );
  BUFFD0 U427 ( .I(n363), .Z(n362) );
  BUFFD0 U428 ( .I(n364), .Z(n363) );
  BUFFD0 U429 ( .I(n365), .Z(n364) );
  BUFFD0 U430 ( .I(n366), .Z(n365) );
  BUFFD0 U431 ( .I(n367), .Z(n366) );
  BUFFD0 U432 ( .I(n368), .Z(n367) );
  BUFFD0 U433 ( .I(n369), .Z(n368) );
  BUFFD0 U434 ( .I(n370), .Z(n369) );
  BUFFD0 U435 ( .I(n371), .Z(n370) );
  BUFFD0 U436 ( .I(n372), .Z(n371) );
  BUFFD0 U437 ( .I(n373), .Z(n372) );
  BUFFD0 U438 ( .I(n374), .Z(n373) );
  BUFFD0 U439 ( .I(n375), .Z(n374) );
  BUFFD0 U440 ( .I(n376), .Z(n375) );
  BUFFD0 U441 ( .I(n377), .Z(n376) );
  BUFFD0 U442 ( .I(n378), .Z(n377) );
  BUFFD0 U443 ( .I(n379), .Z(n378) );
  BUFFD0 U444 ( .I(n704), .Z(n379) );
  BUFFD0 U445 ( .I(n446), .Z(n380) );
  BUFFD0 U446 ( .I(n380), .Z(n381) );
  CKND8 U447 ( .CLK(n467), .CN(n713) );
  CKND2D0 U448 ( .A1(FIFO_Out[8]), .A2(n871), .ZN(n467) );
  CKND8 U449 ( .CLK(n466), .CN(n722) );
  CKND2D0 U450 ( .A1(FIFO_Out[7]), .A2(n871), .ZN(n466) );
  CKND8 U451 ( .CLK(n465), .CN(n731) );
  CKND2D0 U452 ( .A1(FIFO_Out[6]), .A2(n871), .ZN(n465) );
  CKND2D0 U453 ( .A1(FIFO_Out[5]), .A2(n871), .ZN(n464) );
  INVD5 U454 ( .I(n748), .ZN(n749) );
  BUFFD0 U455 ( .I(n383), .Z(n382) );
  BUFFD0 U456 ( .I(n384), .Z(n383) );
  BUFFD0 U457 ( .I(n385), .Z(n384) );
  BUFFD0 U458 ( .I(n386), .Z(n385) );
  BUFFD0 U459 ( .I(n387), .Z(n386) );
  BUFFD0 U460 ( .I(n388), .Z(n387) );
  BUFFD0 U461 ( .I(n389), .Z(n388) );
  BUFFD0 U462 ( .I(n390), .Z(n389) );
  BUFFD0 U463 ( .I(n391), .Z(n390) );
  BUFFD0 U464 ( .I(n392), .Z(n391) );
  BUFFD0 U465 ( .I(n393), .Z(n392) );
  BUFFD0 U466 ( .I(n394), .Z(n393) );
  BUFFD0 U467 ( .I(n395), .Z(n394) );
  BUFFD0 U468 ( .I(n396), .Z(n395) );
  BUFFD0 U469 ( .I(n747), .Z(n396) );
  BUFFD0 U470 ( .I(n445), .Z(n397) );
  BUFFD0 U471 ( .I(n397), .Z(n398) );
  BUFFD0 U472 ( .I(n398), .Z(n399) );
  BUFFD0 U473 ( .I(n399), .Z(n400) );
  BUFFD0 U474 ( .I(n400), .Z(n401) );
  BUFFD0 U475 ( .I(n401), .Z(n402) );
  BUFFD0 U476 ( .I(n402), .Z(n403) );
  BUFFD0 U477 ( .I(n403), .Z(n404) );
  BUFFD0 U478 ( .I(n404), .Z(n405) );
  BUFFD0 U479 ( .I(n405), .Z(n406) );
  BUFFD0 U480 ( .I(n406), .Z(n407) );
  BUFFD0 U481 ( .I(n407), .Z(n408) );
  INVD5 U482 ( .I(n757), .ZN(n758) );
  BUFFD0 U483 ( .I(n410), .Z(n409) );
  BUFFD0 U484 ( .I(n411), .Z(n410) );
  BUFFD0 U485 ( .I(n412), .Z(n411) );
  BUFFD0 U486 ( .I(n413), .Z(n412) );
  BUFFD0 U487 ( .I(n414), .Z(n413) );
  BUFFD0 U488 ( .I(n415), .Z(n414) );
  BUFFD0 U489 ( .I(n416), .Z(n415) );
  BUFFD0 U490 ( .I(n417), .Z(n416) );
  BUFFD0 U491 ( .I(n418), .Z(n417) );
  BUFFD0 U492 ( .I(n419), .Z(n418) );
  BUFFD0 U493 ( .I(n420), .Z(n419) );
  BUFFD0 U494 ( .I(n421), .Z(n420) );
  BUFFD0 U495 ( .I(n422), .Z(n421) );
  BUFFD0 U496 ( .I(n423), .Z(n422) );
  BUFFD0 U497 ( .I(n424), .Z(n423) );
  BUFFD0 U498 ( .I(n425), .Z(n424) );
  BUFFD0 U499 ( .I(n426), .Z(n425) );
  BUFFD0 U500 ( .I(n427), .Z(n426) );
  BUFFD0 U501 ( .I(n428), .Z(n427) );
  BUFFD0 U502 ( .I(n429), .Z(n428) );
  BUFFD0 U503 ( .I(n430), .Z(n429) );
  BUFFD0 U504 ( .I(n431), .Z(n430) );
  BUFFD0 U505 ( .I(n432), .Z(n431) );
  BUFFD0 U506 ( .I(n433), .Z(n432) );
  BUFFD0 U507 ( .I(n756), .Z(n433) );
  BUFFD0 U508 ( .I(n444), .Z(n434) );
  BUFFD0 U509 ( .I(n434), .Z(n435) );
  CKND8 U510 ( .CLK(n463), .CN(n765) );
  CKND2D0 U511 ( .A1(FIFO_Out[2]), .A2(n871), .ZN(n463) );
  CKND8 U512 ( .CLK(n462), .CN(n774) );
  CKND2D0 U513 ( .A1(FIFO_Out[1]), .A2(n871), .ZN(n462) );
  CKND8 U514 ( .CLK(n461), .CN(n783) );
  CKND2D0 U515 ( .A1(FIFO_Out[0]), .A2(n871), .ZN(n461) );
  BUFFD0 U516 ( .I(n437), .Z(n436) );
  BUFFD0 U517 ( .I(n438), .Z(n437) );
  BUFFD0 U518 ( .I(n439), .Z(n438) );
  BUFFD0 U519 ( .I(n440), .Z(n439) );
  BUFFD0 U520 ( .I(n441), .Z(n440) );
  BUFFD0 U521 ( .I(n442), .Z(n441) );
  BUFFD0 U522 ( .I(n443), .Z(n442) );
  BUFFD0 U523 ( .I(n868), .Z(n443) );
  AN2D1 U524 ( .A1(FIFO_Out[3]), .A2(n871), .Z(n444) );
  AN2D1 U525 ( .A1(FIFO_Out[4]), .A2(n871), .Z(n445) );
  AN2D1 U526 ( .A1(FIFO_Out[9]), .A2(n871), .Z(n446) );
  AN2D1 U527 ( .A1(FIFO_Out[10]), .A2(n871), .Z(n447) );
  AN2D1 U528 ( .A1(FIFO_Out[14]), .A2(n871), .Z(n448) );
  AN2D1 U529 ( .A1(FIFO_Out[15]), .A2(n871), .Z(n449) );
  AN2D1 U530 ( .A1(FIFO_Out[19]), .A2(n871), .Z(n450) );
  AN2D1 U531 ( .A1(FIFO_Out[20]), .A2(n871), .Z(n451) );
  AN2D1 U532 ( .A1(FIFO_Out[24]), .A2(n871), .Z(n452) );
  AN2D1 U533 ( .A1(FIFO_Out[25]), .A2(n871), .Z(n453) );
  AN2D1 U534 ( .A1(FIFO_Out[26]), .A2(n871), .Z(n454) );
  AN2D1 U535 ( .A1(FIFO_Out[27]), .A2(n871), .Z(n455) );
  AN2D1 U536 ( .A1(FIFO_Out[28]), .A2(n871), .Z(n456) );
  AN2D1 U537 ( .A1(FIFO_Out[29]), .A2(n871), .Z(n457) );
  AN2D1 U538 ( .A1(FIFO_Out[30]), .A2(n871), .Z(n458) );
  AN2D1 U539 ( .A1(FIFO_Out[31]), .A2(n871), .Z(n459) );
  OR2D1 U540 ( .A1(FIFOEmpty), .A2(n792), .Z(n460) );
  BUFFD0 U541 ( .I(n478), .Z(n477) );
  BUFFD0 U542 ( .I(n603), .Z(n478) );
  BUFFD0 U543 ( .I(n482), .Z(n481) );
  BUFFD0 U544 ( .I(n689), .Z(n482) );
  BUFFD0 U545 ( .I(n484), .Z(n483) );
  BUFFD0 U546 ( .I(n741), .Z(n484) );
  INVD1 U547 ( .I(n460), .ZN(n868) );
  BUFFD0 U548 ( .I(n486), .Z(n485) );
  BUFFD0 U549 ( .I(n487), .Z(n486) );
  BUFFD0 U550 ( .I(n488), .Z(n487) );
  BUFFD0 U551 ( .I(n489), .Z(n488) );
  BUFFD0 U552 ( .I(n490), .Z(n489) );
  BUFFD0 U553 ( .I(n491), .Z(n490) );
  BUFFD0 U554 ( .I(n492), .Z(n491) );
  BUFFD0 U555 ( .I(n493), .Z(n492) );
  BUFFD0 U556 ( .I(n494), .Z(n493) );
  BUFFD0 U557 ( .I(n495), .Z(n494) );
  BUFFD0 U558 ( .I(n496), .Z(n495) );
  BUFFD0 U559 ( .I(n497), .Z(n496) );
  BUFFD0 U560 ( .I(n498), .Z(n497) );
  BUFFD0 U561 ( .I(n499), .Z(n498) );
  BUFFD0 U562 ( .I(n500), .Z(n499) );
  BUFFD0 U563 ( .I(n501), .Z(n500) );
  BUFFD0 U564 ( .I(n502), .Z(n501) );
  BUFFD0 U565 ( .I(n503), .Z(n502) );
  BUFFD0 U566 ( .I(n504), .Z(n503) );
  BUFFD0 U567 ( .I(n505), .Z(n504) );
  BUFFD0 U568 ( .I(n506), .Z(n505) );
  BUFFD0 U569 ( .I(n507), .Z(n506) );
  BUFFD0 U570 ( .I(n508), .Z(n507) );
  BUFFD0 U571 ( .I(n511), .Z(n508) );
  INVD0 U572 ( .I(n509), .ZN(n510) );
  CKNXD16 U573 ( .I(Reset), .ZN(n509) );
  BUFFD0 U574 ( .I(n869), .Z(n511) );
  BUFFD0 U575 ( .I(n514), .Z(n512) );
  INVD0 U576 ( .I(n516), .ZN(n513) );
  CKNXD16 U577 ( .I(n515), .ZN(n516) );
  INVD0 U578 ( .I(n518), .ZN(n515) );
  CKNXD16 U579 ( .I(n517), .ZN(n518) );
  INVD0 U580 ( .I(n520), .ZN(n517) );
  CKNXD16 U581 ( .I(n519), .ZN(n520) );
  INVD0 U582 ( .I(n30), .ZN(n519) );
  BUFFD0 U583 ( .I(n523), .Z(n521) );
  INVD0 U584 ( .I(n525), .ZN(n522) );
  CKNXD16 U585 ( .I(n524), .ZN(n525) );
  INVD0 U586 ( .I(n527), .ZN(n524) );
  CKNXD16 U587 ( .I(n526), .ZN(n527) );
  INVD0 U588 ( .I(n529), .ZN(n526) );
  CKNXD16 U589 ( .I(n528), .ZN(n529) );
  INVD0 U590 ( .I(n57), .ZN(n528) );
  BUFFD0 U591 ( .I(n532), .Z(n530) );
  INVD0 U592 ( .I(n534), .ZN(n531) );
  CKNXD16 U593 ( .I(n533), .ZN(n534) );
  INVD0 U594 ( .I(n536), .ZN(n533) );
  CKNXD16 U595 ( .I(n535), .ZN(n536) );
  INVD0 U596 ( .I(n538), .ZN(n535) );
  CKNXD16 U597 ( .I(n537), .ZN(n538) );
  INVD0 U598 ( .I(n84), .ZN(n537) );
  BUFFD0 U599 ( .I(n541), .Z(n539) );
  INVD0 U600 ( .I(n543), .ZN(n540) );
  CKNXD16 U601 ( .I(n542), .ZN(n543) );
  INVD0 U602 ( .I(n545), .ZN(n542) );
  CKNXD16 U603 ( .I(n544), .ZN(n545) );
  INVD0 U604 ( .I(n547), .ZN(n544) );
  CKNXD16 U605 ( .I(n546), .ZN(n547) );
  INVD0 U606 ( .I(n111), .ZN(n546) );
  BUFFD0 U607 ( .I(n550), .Z(n548) );
  INVD0 U608 ( .I(n552), .ZN(n549) );
  CKNXD16 U609 ( .I(n551), .ZN(n552) );
  INVD0 U610 ( .I(n554), .ZN(n551) );
  CKNXD16 U611 ( .I(n553), .ZN(n554) );
  INVD0 U612 ( .I(n556), .ZN(n553) );
  CKNXD16 U613 ( .I(n555), .ZN(n556) );
  INVD0 U614 ( .I(n138), .ZN(n555) );
  BUFFD0 U615 ( .I(n559), .Z(n557) );
  INVD0 U616 ( .I(n561), .ZN(n558) );
  CKNXD16 U617 ( .I(n560), .ZN(n561) );
  INVD0 U618 ( .I(n563), .ZN(n560) );
  CKNXD16 U619 ( .I(n562), .ZN(n563) );
  INVD0 U620 ( .I(n565), .ZN(n562) );
  CKNXD16 U621 ( .I(n564), .ZN(n565) );
  INVD0 U622 ( .I(n165), .ZN(n564) );
  BUFFD0 U623 ( .I(n568), .Z(n566) );
  INVD0 U624 ( .I(n570), .ZN(n567) );
  CKNXD16 U625 ( .I(n569), .ZN(n570) );
  INVD0 U626 ( .I(n572), .ZN(n569) );
  CKNXD16 U627 ( .I(n571), .ZN(n572) );
  INVD0 U628 ( .I(n574), .ZN(n571) );
  CKNXD16 U629 ( .I(n573), .ZN(n574) );
  INVD0 U630 ( .I(n192), .ZN(n573) );
  BUFFD0 U631 ( .I(n577), .Z(n575) );
  INVD0 U632 ( .I(n579), .ZN(n576) );
  CKNXD16 U633 ( .I(n578), .ZN(n579) );
  INVD0 U634 ( .I(n581), .ZN(n578) );
  CKNXD16 U635 ( .I(n580), .ZN(n581) );
  INVD0 U636 ( .I(n583), .ZN(n580) );
  CKNXD16 U637 ( .I(n582), .ZN(n583) );
  INVD0 U638 ( .I(n219), .ZN(n582) );
  CKNXD16 U639 ( .I(n585), .ZN(n586) );
  INVD0 U640 ( .I(n588), .ZN(n585) );
  CKNXD16 U641 ( .I(n587), .ZN(n588) );
  INVD0 U642 ( .I(n590), .ZN(n587) );
  CKNXD16 U643 ( .I(n589), .ZN(n590) );
  INVD0 U644 ( .I(n592), .ZN(n589) );
  CKNXD16 U645 ( .I(n591), .ZN(n592) );
  INVD0 U646 ( .I(n584), .ZN(n591) );
  CKNXD16 U647 ( .I(n594), .ZN(n595) );
  INVD0 U648 ( .I(n597), .ZN(n594) );
  CKNXD16 U649 ( .I(n596), .ZN(n597) );
  INVD0 U650 ( .I(n599), .ZN(n596) );
  CKNXD16 U651 ( .I(n598), .ZN(n599) );
  INVD0 U652 ( .I(n601), .ZN(n598) );
  CKNXD16 U653 ( .I(n600), .ZN(n601) );
  INVD0 U654 ( .I(n593), .ZN(n600) );
  CKNXD16 U655 ( .I(n602), .ZN(n603) );
  INVD0 U656 ( .I(n605), .ZN(n602) );
  CKNXD16 U657 ( .I(n604), .ZN(n605) );
  INVD0 U658 ( .I(n607), .ZN(n604) );
  CKNXD16 U659 ( .I(n606), .ZN(n607) );
  INVD0 U660 ( .I(n608), .ZN(n606) );
  CKNXD16 U661 ( .I(n474), .ZN(n608) );
  BUFFD0 U662 ( .I(n611), .Z(n609) );
  INVD0 U663 ( .I(n613), .ZN(n610) );
  CKNXD16 U664 ( .I(n612), .ZN(n613) );
  INVD0 U665 ( .I(n615), .ZN(n612) );
  CKNXD16 U666 ( .I(n614), .ZN(n615) );
  INVD0 U667 ( .I(n617), .ZN(n614) );
  CKNXD16 U668 ( .I(n616), .ZN(n617) );
  INVD0 U669 ( .I(n246), .ZN(n616) );
  BUFFD0 U670 ( .I(n620), .Z(n618) );
  INVD0 U671 ( .I(n622), .ZN(n619) );
  CKNXD16 U672 ( .I(n621), .ZN(n622) );
  INVD0 U673 ( .I(n624), .ZN(n621) );
  CKNXD16 U674 ( .I(n623), .ZN(n624) );
  INVD0 U675 ( .I(n626), .ZN(n623) );
  CKNXD16 U676 ( .I(n625), .ZN(n626) );
  INVD0 U677 ( .I(n273), .ZN(n625) );
  CKNXD16 U678 ( .I(n628), .ZN(n629) );
  INVD0 U679 ( .I(n631), .ZN(n628) );
  CKNXD16 U680 ( .I(n630), .ZN(n631) );
  INVD0 U681 ( .I(n633), .ZN(n630) );
  CKNXD16 U682 ( .I(n632), .ZN(n633) );
  INVD0 U683 ( .I(n635), .ZN(n632) );
  CKNXD16 U684 ( .I(n634), .ZN(n635) );
  INVD0 U685 ( .I(n627), .ZN(n634) );
  CKNXD16 U686 ( .I(n637), .ZN(n638) );
  INVD0 U687 ( .I(n640), .ZN(n637) );
  CKNXD16 U688 ( .I(n639), .ZN(n640) );
  INVD0 U689 ( .I(n642), .ZN(n639) );
  CKNXD16 U690 ( .I(n641), .ZN(n642) );
  INVD0 U691 ( .I(n644), .ZN(n641) );
  CKNXD16 U692 ( .I(n643), .ZN(n644) );
  INVD0 U693 ( .I(n636), .ZN(n643) );
  CKNXD16 U694 ( .I(n645), .ZN(n646) );
  INVD0 U695 ( .I(n648), .ZN(n645) );
  CKNXD16 U696 ( .I(n647), .ZN(n648) );
  INVD0 U697 ( .I(n650), .ZN(n647) );
  CKNXD16 U698 ( .I(n649), .ZN(n650) );
  INVD0 U699 ( .I(n651), .ZN(n649) );
  CKNXD16 U700 ( .I(n471), .ZN(n651) );
  BUFFD0 U701 ( .I(n654), .Z(n652) );
  INVD0 U702 ( .I(n656), .ZN(n653) );
  CKNXD16 U703 ( .I(n655), .ZN(n656) );
  INVD0 U704 ( .I(n658), .ZN(n655) );
  CKNXD16 U705 ( .I(n657), .ZN(n658) );
  INVD0 U706 ( .I(n660), .ZN(n657) );
  CKNXD16 U707 ( .I(n659), .ZN(n660) );
  INVD0 U708 ( .I(n300), .ZN(n659) );
  BUFFD0 U709 ( .I(n663), .Z(n661) );
  INVD0 U710 ( .I(n665), .ZN(n662) );
  CKNXD16 U711 ( .I(n664), .ZN(n665) );
  INVD0 U712 ( .I(n667), .ZN(n664) );
  CKNXD16 U713 ( .I(n666), .ZN(n667) );
  INVD0 U714 ( .I(n669), .ZN(n666) );
  CKNXD16 U715 ( .I(n668), .ZN(n669) );
  INVD0 U716 ( .I(n327), .ZN(n668) );
  CKNXD16 U717 ( .I(n671), .ZN(n672) );
  INVD0 U718 ( .I(n674), .ZN(n671) );
  CKNXD16 U719 ( .I(n673), .ZN(n674) );
  INVD0 U720 ( .I(n676), .ZN(n673) );
  CKNXD16 U721 ( .I(n675), .ZN(n676) );
  INVD0 U722 ( .I(n678), .ZN(n675) );
  CKNXD16 U723 ( .I(n677), .ZN(n678) );
  INVD0 U724 ( .I(n670), .ZN(n677) );
  CKNXD16 U725 ( .I(n680), .ZN(n681) );
  INVD0 U726 ( .I(n683), .ZN(n680) );
  CKNXD16 U727 ( .I(n682), .ZN(n683) );
  INVD0 U728 ( .I(n685), .ZN(n682) );
  CKNXD16 U729 ( .I(n684), .ZN(n685) );
  INVD0 U730 ( .I(n687), .ZN(n684) );
  CKNXD16 U731 ( .I(n686), .ZN(n687) );
  INVD0 U732 ( .I(n679), .ZN(n686) );
  CKNXD16 U733 ( .I(n688), .ZN(n689) );
  INVD0 U734 ( .I(n691), .ZN(n688) );
  CKNXD16 U735 ( .I(n690), .ZN(n691) );
  INVD0 U736 ( .I(n693), .ZN(n690) );
  CKNXD16 U737 ( .I(n692), .ZN(n693) );
  INVD0 U738 ( .I(n694), .ZN(n692) );
  CKNXD16 U739 ( .I(n468), .ZN(n694) );
  BUFFD0 U740 ( .I(n697), .Z(n695) );
  INVD0 U741 ( .I(n699), .ZN(n696) );
  CKNXD16 U742 ( .I(n698), .ZN(n699) );
  INVD0 U743 ( .I(n701), .ZN(n698) );
  CKNXD16 U744 ( .I(n700), .ZN(n701) );
  INVD0 U745 ( .I(n703), .ZN(n700) );
  CKNXD16 U746 ( .I(n702), .ZN(n703) );
  INVD0 U747 ( .I(n354), .ZN(n702) );
  BUFFD0 U748 ( .I(n706), .Z(n704) );
  INVD0 U749 ( .I(n708), .ZN(n705) );
  CKNXD16 U750 ( .I(n707), .ZN(n708) );
  INVD0 U751 ( .I(n710), .ZN(n707) );
  CKNXD16 U752 ( .I(n709), .ZN(n710) );
  INVD0 U753 ( .I(n712), .ZN(n709) );
  CKNXD16 U754 ( .I(n711), .ZN(n712) );
  INVD0 U755 ( .I(n381), .ZN(n711) );
  CKNXD16 U756 ( .I(n714), .ZN(n715) );
  INVD0 U757 ( .I(n717), .ZN(n714) );
  CKNXD16 U758 ( .I(n716), .ZN(n717) );
  INVD0 U759 ( .I(n719), .ZN(n716) );
  CKNXD16 U760 ( .I(n718), .ZN(n719) );
  INVD0 U761 ( .I(n721), .ZN(n718) );
  CKNXD16 U762 ( .I(n720), .ZN(n721) );
  INVD0 U763 ( .I(n713), .ZN(n720) );
  CKNXD16 U764 ( .I(n723), .ZN(n724) );
  INVD0 U765 ( .I(n726), .ZN(n723) );
  CKNXD16 U766 ( .I(n725), .ZN(n726) );
  INVD0 U767 ( .I(n728), .ZN(n725) );
  CKNXD16 U768 ( .I(n727), .ZN(n728) );
  INVD0 U769 ( .I(n730), .ZN(n727) );
  CKNXD16 U770 ( .I(n729), .ZN(n730) );
  INVD0 U771 ( .I(n722), .ZN(n729) );
  CKNXD16 U772 ( .I(n732), .ZN(n733) );
  INVD0 U773 ( .I(n735), .ZN(n732) );
  CKNXD16 U774 ( .I(n734), .ZN(n735) );
  INVD0 U775 ( .I(n737), .ZN(n734) );
  CKNXD16 U776 ( .I(n736), .ZN(n737) );
  INVD0 U777 ( .I(n739), .ZN(n736) );
  CKNXD16 U778 ( .I(n738), .ZN(n739) );
  INVD0 U779 ( .I(n731), .ZN(n738) );
  CKNXD16 U780 ( .I(n740), .ZN(n741) );
  INVD0 U781 ( .I(n743), .ZN(n740) );
  CKNXD16 U782 ( .I(n742), .ZN(n743) );
  INVD0 U783 ( .I(n745), .ZN(n742) );
  CKNXD16 U784 ( .I(n744), .ZN(n745) );
  INVD0 U785 ( .I(n746), .ZN(n744) );
  CKNXD16 U786 ( .I(n464), .ZN(n746) );
  BUFFD0 U787 ( .I(n749), .Z(n747) );
  INVD0 U788 ( .I(n751), .ZN(n748) );
  CKNXD16 U789 ( .I(n750), .ZN(n751) );
  INVD0 U790 ( .I(n753), .ZN(n750) );
  CKNXD16 U791 ( .I(n752), .ZN(n753) );
  INVD0 U792 ( .I(n755), .ZN(n752) );
  CKNXD16 U793 ( .I(n754), .ZN(n755) );
  INVD0 U794 ( .I(n408), .ZN(n754) );
  BUFFD0 U795 ( .I(n758), .Z(n756) );
  INVD0 U796 ( .I(n760), .ZN(n757) );
  CKNXD16 U797 ( .I(n759), .ZN(n760) );
  INVD0 U798 ( .I(n762), .ZN(n759) );
  CKNXD16 U799 ( .I(n761), .ZN(n762) );
  INVD0 U800 ( .I(n764), .ZN(n761) );
  CKNXD16 U801 ( .I(n763), .ZN(n764) );
  INVD0 U802 ( .I(n435), .ZN(n763) );
  CKNXD16 U803 ( .I(n766), .ZN(n767) );
  INVD0 U804 ( .I(n769), .ZN(n766) );
  CKNXD16 U805 ( .I(n768), .ZN(n769) );
  INVD0 U806 ( .I(n771), .ZN(n768) );
  CKNXD16 U807 ( .I(n770), .ZN(n771) );
  INVD0 U808 ( .I(n773), .ZN(n770) );
  CKNXD16 U809 ( .I(n772), .ZN(n773) );
  INVD0 U810 ( .I(n765), .ZN(n772) );
  CKNXD16 U811 ( .I(n775), .ZN(n776) );
  INVD0 U812 ( .I(n778), .ZN(n775) );
  CKNXD16 U813 ( .I(n777), .ZN(n778) );
  INVD0 U814 ( .I(n780), .ZN(n777) );
  CKNXD16 U815 ( .I(n779), .ZN(n780) );
  INVD0 U816 ( .I(n782), .ZN(n779) );
  CKNXD16 U817 ( .I(n781), .ZN(n782) );
  INVD0 U818 ( .I(n774), .ZN(n781) );
  CKNXD16 U819 ( .I(n784), .ZN(n785) );
  INVD0 U820 ( .I(n787), .ZN(n784) );
  CKNXD16 U821 ( .I(n786), .ZN(n787) );
  INVD0 U822 ( .I(n789), .ZN(n786) );
  CKNXD16 U823 ( .I(n788), .ZN(n789) );
  INVD0 U824 ( .I(n791), .ZN(n788) );
  CKNXD16 U825 ( .I(n790), .ZN(n791) );
  INVD0 U826 ( .I(n783), .ZN(n790) );
  BUFFD0 U827 ( .I(n793), .Z(n792) );
  BUFFD0 U828 ( .I(n794), .Z(n793) );
  BUFFD0 U829 ( .I(n795), .Z(n794) );
  BUFFD0 U830 ( .I(n796), .Z(n795) );
  BUFFD0 U831 ( .I(n797), .Z(n796) );
  BUFFD0 U832 ( .I(n798), .Z(n797) );
  BUFFD0 U833 ( .I(n799), .Z(n798) );
  BUFFD0 U834 ( .I(n800), .Z(n799) );
  BUFFD0 U835 ( .I(n801), .Z(n800) );
  BUFFD0 U836 ( .I(n802), .Z(n801) );
  BUFFD0 U837 ( .I(n803), .Z(n802) );
  BUFFD0 U838 ( .I(n804), .Z(n803) );
  BUFFD0 U839 ( .I(n805), .Z(n804) );
  BUFFD0 U840 ( .I(n806), .Z(n805) );
  BUFFD0 U841 ( .I(n807), .Z(n806) );
  BUFFD0 U842 ( .I(n808), .Z(n807) );
  BUFFD0 U843 ( .I(n809), .Z(n808) );
  BUFFD0 U844 ( .I(n810), .Z(n809) );
  BUFFD0 U845 ( .I(n811), .Z(n810) );
  BUFFD0 U846 ( .I(n812), .Z(n811) );
  BUFFD0 U847 ( .I(n813), .Z(n812) );
  BUFFD0 U848 ( .I(n814), .Z(n813) );
  BUFFD0 U849 ( .I(n815), .Z(n814) );
  BUFFD0 U850 ( .I(n816), .Z(n815) );
  BUFFD0 U851 ( .I(n817), .Z(n816) );
  BUFFD0 U852 ( .I(n818), .Z(n817) );
  BUFFD0 U853 ( .I(n819), .Z(n818) );
  BUFFD0 U854 ( .I(n820), .Z(n819) );
  BUFFD0 U855 ( .I(n821), .Z(n820) );
  BUFFD0 U856 ( .I(n822), .Z(n821) );
  BUFFD0 U857 ( .I(n823), .Z(n822) );
  BUFFD0 U858 ( .I(n824), .Z(n823) );
  BUFFD0 U859 ( .I(n825), .Z(n824) );
  BUFFD0 U860 ( .I(n826), .Z(n825) );
  BUFFD0 U861 ( .I(n827), .Z(n826) );
  BUFFD0 U862 ( .I(n828), .Z(n827) );
  BUFFD0 U863 ( .I(n829), .Z(n828) );
  BUFFD0 U864 ( .I(n830), .Z(n829) );
  BUFFD0 U865 ( .I(n831), .Z(n830) );
  BUFFD0 U866 ( .I(n832), .Z(n831) );
  BUFFD0 U867 ( .I(n833), .Z(n832) );
  BUFFD0 U868 ( .I(n834), .Z(n833) );
  BUFFD0 U869 ( .I(n835), .Z(n834) );
  BUFFD0 U870 ( .I(n836), .Z(n835) );
  BUFFD0 U871 ( .I(n837), .Z(n836) );
  BUFFD0 U872 ( .I(n838), .Z(n837) );
  BUFFD0 U873 ( .I(n839), .Z(n838) );
  BUFFD0 U874 ( .I(n840), .Z(n839) );
  BUFFD0 U875 ( .I(n841), .Z(n840) );
  BUFFD0 U876 ( .I(n842), .Z(n841) );
  BUFFD0 U877 ( .I(n843), .Z(n842) );
  BUFFD0 U878 ( .I(n844), .Z(n843) );
  BUFFD0 U879 ( .I(n845), .Z(n844) );
  BUFFD0 U880 ( .I(n846), .Z(n845) );
  BUFFD0 U881 ( .I(n847), .Z(n846) );
  BUFFD0 U882 ( .I(n848), .Z(n847) );
  BUFFD0 U883 ( .I(n849), .Z(n848) );
  BUFFD0 U884 ( .I(n850), .Z(n849) );
  BUFFD0 U885 ( .I(n851), .Z(n850) );
  BUFFD0 U886 ( .I(n852), .Z(n851) );
  BUFFD0 U887 ( .I(n853), .Z(n852) );
  BUFFD0 U888 ( .I(n856), .Z(n853) );
  INVD0 U889 ( .I(n854), .ZN(n855) );
  CKNXD16 U890 ( .I(ReadReq), .ZN(n854) );
  BUFFD0 U891 ( .I(n857), .Z(n856) );
  BUFFD0 U892 ( .I(n858), .Z(n857) );
  BUFFD0 U893 ( .I(n859), .Z(n858) );
  BUFFD0 U894 ( .I(n860), .Z(n859) );
  BUFFD0 U895 ( .I(n861), .Z(n860) );
  BUFFD0 U896 ( .I(n862), .Z(n861) );
  BUFFD0 U897 ( .I(n863), .Z(n862) );
  BUFFD0 U898 ( .I(n864), .Z(n863) );
  BUFFD0 U899 ( .I(n865), .Z(n864) );
  BUFFD0 U900 ( .I(n866), .Z(n865) );
  BUFFD0 U901 ( .I(n867), .Z(n866) );
  BUFFD0 U902 ( .I(n872), .Z(n867) );
  INVD4 U903 ( .I(n869), .ZN(n2) );
  CKBXD0 U904 ( .I(n510), .Z(n869) );
  INVD1 U905 ( .I(n792), .ZN(n871) );
  INVD1 U906 ( .I(n855), .ZN(n872) );
  BUFFD1 U907 ( .I(ParOutClk), .Z(n870) );
endmodule


module FIFOTop_AWid5_DWid32 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(n3), .WriteReq(WriteIn), .ClkR(
        ClkR), .ClkW(ClkW), .Reset(Reseter) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({Din[31:2], n2, 
        Din[0]}), .AddrR(SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), 
        .ClkW(ClkW), .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), 
        .Reset(Reseter) );
  CKBD0 U2 ( .CLK(SM_MemReadCmd), .C(n1) );
  BUFFD1 U3 ( .I(ReadIn), .Z(n3) );
  BUFFD1 U4 ( .I(Din[1]), .Z(n2) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   N4, UnLoad, doParSync, N51, N52, N53, N54, N55, N64, N66, N67, N68,
         N69, N70, N71, N72, net420, net419, net418, net417, net416, net415,
         net414, net413, net412, net411, net410, net409, net408, net407,
         net406, net405, net404, net403, net402, net401, net400, net399,
         net398, net397, net396, net395, net394, net393, net392, net391,
         net390, net389, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n1, n4, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196;
  wire   [31:0] DecodeReg;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  LHD1 SerClock_reg ( .E(N71), .D(N66), .QN(N4) );
  LHQD1 \Count32_reg[0]  ( .E(N71), .D(N67), .Q(Count32[0]) );
  LHQD1 \Count32_reg[1]  ( .E(N71), .D(N68), .Q(Count32[1]) );
  LHQD1 \Count32_reg[2]  ( .E(N71), .D(N69), .Q(Count32[2]) );
  LHQD1 \Count32_reg[3]  ( .E(N71), .D(N70), .Q(Count32[3]) );
  LHQD1 \Count32_reg[4]  ( .E(N71), .D(N72), .Q(Count32[4]) );
  MOAI22D1 U6 ( .A1(n192), .A2(net398), .B1(DecodeReg[9]), .B2(n193), .ZN(n47)
         );
  MOAI22D1 U7 ( .A1(n192), .A2(net397), .B1(n193), .B2(DecodeReg[8]), .ZN(n48)
         );
  MOAI22D1 U8 ( .A1(UnLoad), .A2(net396), .B1(n192), .B2(DecodeReg[7]), .ZN(
        n49) );
  MOAI22D1 U9 ( .A1(n192), .A2(net395), .B1(n192), .B2(DecodeReg[6]), .ZN(n50)
         );
  MOAI22D1 U10 ( .A1(n193), .A2(net394), .B1(n192), .B2(DecodeReg[5]), .ZN(n51) );
  MOAI22D1 U11 ( .A1(UnLoad), .A2(net393), .B1(n193), .B2(DecodeReg[4]), .ZN(
        n52) );
  MOAI22D1 U12 ( .A1(UnLoad), .A2(net392), .B1(n193), .B2(DecodeReg[3]), .ZN(
        n53) );
  MOAI22D1 U13 ( .A1(UnLoad), .A2(net420), .B1(n193), .B2(DecodeReg[31]), .ZN(
        n25) );
  MOAI22D1 U14 ( .A1(UnLoad), .A2(net419), .B1(UnLoad), .B2(DecodeReg[30]), 
        .ZN(n26) );
  MOAI22D1 U15 ( .A1(UnLoad), .A2(net391), .B1(n193), .B2(DecodeReg[2]), .ZN(
        n54) );
  MOAI22D1 U16 ( .A1(n192), .A2(net418), .B1(n193), .B2(DecodeReg[29]), .ZN(
        n27) );
  MOAI22D1 U17 ( .A1(n192), .A2(net417), .B1(n193), .B2(DecodeReg[28]), .ZN(
        n28) );
  MOAI22D1 U18 ( .A1(n192), .A2(net416), .B1(n193), .B2(DecodeReg[27]), .ZN(
        n29) );
  MOAI22D1 U19 ( .A1(UnLoad), .A2(net415), .B1(n193), .B2(DecodeReg[26]), .ZN(
        n30) );
  MOAI22D1 U20 ( .A1(n192), .A2(net414), .B1(n193), .B2(DecodeReg[25]), .ZN(
        n31) );
  MOAI22D1 U21 ( .A1(n193), .A2(net413), .B1(n193), .B2(DecodeReg[24]), .ZN(
        n32) );
  MOAI22D1 U22 ( .A1(UnLoad), .A2(net412), .B1(n192), .B2(DecodeReg[23]), .ZN(
        n33) );
  MOAI22D1 U23 ( .A1(n192), .A2(net411), .B1(n193), .B2(DecodeReg[22]), .ZN(
        n34) );
  MOAI22D1 U24 ( .A1(UnLoad), .A2(net410), .B1(n193), .B2(DecodeReg[21]), .ZN(
        n35) );
  MOAI22D1 U25 ( .A1(UnLoad), .A2(net409), .B1(n193), .B2(DecodeReg[20]), .ZN(
        n36) );
  MOAI22D1 U26 ( .A1(n192), .A2(net390), .B1(n193), .B2(DecodeReg[1]), .ZN(n55) );
  MOAI22D1 U27 ( .A1(UnLoad), .A2(net408), .B1(UnLoad), .B2(DecodeReg[19]), 
        .ZN(n37) );
  MOAI22D1 U28 ( .A1(n193), .A2(net407), .B1(UnLoad), .B2(DecodeReg[18]), .ZN(
        n38) );
  MOAI22D1 U29 ( .A1(n192), .A2(net406), .B1(UnLoad), .B2(DecodeReg[17]), .ZN(
        n39) );
  MOAI22D1 U30 ( .A1(UnLoad), .A2(net405), .B1(n192), .B2(DecodeReg[16]), .ZN(
        n40) );
  MOAI22D1 U31 ( .A1(n192), .A2(net404), .B1(n192), .B2(DecodeReg[15]), .ZN(
        n41) );
  MOAI22D1 U32 ( .A1(UnLoad), .A2(net403), .B1(n193), .B2(DecodeReg[14]), .ZN(
        n42) );
  MOAI22D1 U33 ( .A1(n193), .A2(net402), .B1(UnLoad), .B2(DecodeReg[13]), .ZN(
        n43) );
  MOAI22D1 U34 ( .A1(n193), .A2(net401), .B1(UnLoad), .B2(DecodeReg[12]), .ZN(
        n44) );
  MOAI22D1 U35 ( .A1(UnLoad), .A2(net400), .B1(n192), .B2(DecodeReg[11]), .ZN(
        n45) );
  MOAI22D1 U36 ( .A1(n192), .A2(net399), .B1(n192), .B2(DecodeReg[10]), .ZN(
        n46) );
  MOAI22D1 U37 ( .A1(n192), .A2(net389), .B1(UnLoad), .B2(DecodeReg[0]), .ZN(
        n56) );
  OR3D1 U46 ( .A1(doParSync), .A2(Reset), .A3(n6), .Z(n5) );
  OR3D1 U90 ( .A1(FrameSR[55]), .A2(FrameSR[54]), .A3(FrameSR[53]), .Z(n16) );
  OR3D1 U92 ( .A1(FrameSR[39]), .A2(FrameSR[38]), .A3(FrameSR[37]), .Z(n17) );
  OR3D1 U94 ( .A1(FrameSR[32]), .A2(FrameSR[23]), .A3(FrameSR[22]), .Z(n18) );
  DesDecoder_DWid32_DW01_inc_0 \SerClockGen/add_170  ( .A(Count32), .SUM({N55, 
        N54, N53, N52, N51}) );
  DFCND1 \FrameSR_reg[63]  ( .D(FrameSR[62]), .CP(n196), .CDN(n189), .Q(
        FrameSR[63]) );
  DFCND1 \FrameSR_reg[22]  ( .D(FrameSR[21]), .CP(N4), .CDN(n22), .Q(
        FrameSR[22]) );
  DFCND1 \FrameSR_reg[23]  ( .D(FrameSR[22]), .CP(n196), .CDN(n187), .Q(
        FrameSR[23]) );
  DFCND1 \FrameSR_reg[37]  ( .D(FrameSR[36]), .CP(n194), .CDN(n187), .Q(
        FrameSR[37]) );
  DFCND1 \FrameSR_reg[38]  ( .D(FrameSR[37]), .CP(n196), .CDN(n190), .Q(
        FrameSR[38]) );
  DFCND1 \FrameSR_reg[53]  ( .D(FrameSR[52]), .CP(n196), .CDN(n187), .Q(
        FrameSR[53]) );
  DFCND1 \FrameSR_reg[54]  ( .D(FrameSR[53]), .CP(n195), .CDN(n189), .Q(
        FrameSR[54]) );
  DFCND1 \FrameSR_reg[32]  ( .D(FrameSR[31]), .CP(n194), .CDN(n190), .Q(
        FrameSR[32]) );
  DFCND1 \FrameSR_reg[39]  ( .D(FrameSR[38]), .CP(N4), .CDN(n190), .Q(
        FrameSR[39]) );
  DFCND1 \FrameSR_reg[55]  ( .D(FrameSR[54]), .CP(n195), .CDN(n22), .Q(
        FrameSR[55]) );
  DFCND1 \FrameSR_reg[8]  ( .D(FrameSR[7]), .CP(N4), .CDN(n189), .Q(FrameSR[8]) );
  DFCND1 \FrameSR_reg[9]  ( .D(FrameSR[8]), .CP(n196), .CDN(n187), .Q(
        FrameSR[9]) );
  DFCND1 \FrameSR_reg[10]  ( .D(FrameSR[9]), .CP(n195), .CDN(n22), .Q(
        FrameSR[10]) );
  DFCND1 \FrameSR_reg[11]  ( .D(FrameSR[10]), .CP(n195), .CDN(n190), .Q(
        FrameSR[11]) );
  DFCND1 \FrameSR_reg[12]  ( .D(FrameSR[11]), .CP(n195), .CDN(n190), .Q(
        FrameSR[12]) );
  DFCND1 \FrameSR_reg[13]  ( .D(FrameSR[12]), .CP(n195), .CDN(n190), .Q(
        FrameSR[13]) );
  DFCND1 \FrameSR_reg[14]  ( .D(FrameSR[13]), .CP(n195), .CDN(n189), .Q(
        FrameSR[14]) );
  DFCND1 \FrameSR_reg[15]  ( .D(FrameSR[14]), .CP(n195), .CDN(n188), .Q(
        FrameSR[15]) );
  DFCND1 \FrameSR_reg[19]  ( .D(FrameSR[18]), .CP(n195), .CDN(n22), .Q(
        FrameSR[19]) );
  DFCND1 \FrameSR_reg[24]  ( .D(FrameSR[23]), .CP(n196), .CDN(n187), .Q(
        FrameSR[24]) );
  DFCND1 \FrameSR_reg[25]  ( .D(FrameSR[24]), .CP(N4), .CDN(n22), .Q(
        FrameSR[25]) );
  DFCND1 \FrameSR_reg[26]  ( .D(FrameSR[25]), .CP(n194), .CDN(n22), .Q(
        FrameSR[26]) );
  DFCND1 \FrameSR_reg[27]  ( .D(FrameSR[26]), .CP(n195), .CDN(n190), .Q(
        FrameSR[27]) );
  DFCND1 \FrameSR_reg[28]  ( .D(FrameSR[27]), .CP(n196), .CDN(n187), .Q(
        FrameSR[28]) );
  DFCND1 \FrameSR_reg[29]  ( .D(FrameSR[28]), .CP(n196), .CDN(n22), .Q(
        FrameSR[29]) );
  DFCND1 \FrameSR_reg[30]  ( .D(FrameSR[29]), .CP(n195), .CDN(n187), .Q(
        FrameSR[30]) );
  DFCND1 \FrameSR_reg[31]  ( .D(FrameSR[30]), .CP(N4), .CDN(n187), .Q(
        FrameSR[31]) );
  DFCND1 \FrameSR_reg[40]  ( .D(FrameSR[39]), .CP(n196), .CDN(n189), .Q(
        FrameSR[40]) );
  DFCND1 \FrameSR_reg[41]  ( .D(FrameSR[40]), .CP(n194), .CDN(n187), .Q(
        FrameSR[41]) );
  DFCND1 \FrameSR_reg[42]  ( .D(FrameSR[41]), .CP(n196), .CDN(n22), .Q(
        FrameSR[42]) );
  DFCND1 \FrameSR_reg[43]  ( .D(FrameSR[42]), .CP(n195), .CDN(n190), .Q(
        FrameSR[43]) );
  DFCND1 \FrameSR_reg[44]  ( .D(FrameSR[43]), .CP(n195), .CDN(n190), .Q(
        FrameSR[44]) );
  DFCND1 \FrameSR_reg[45]  ( .D(FrameSR[44]), .CP(n195), .CDN(n188), .Q(
        FrameSR[45]) );
  DFCND1 \FrameSR_reg[46]  ( .D(FrameSR[45]), .CP(n195), .CDN(n188), .Q(
        FrameSR[46]) );
  DFCND1 \FrameSR_reg[47]  ( .D(FrameSR[46]), .CP(n196), .CDN(n190), .Q(
        FrameSR[47]) );
  DFCND1 \FrameSR_reg[56]  ( .D(FrameSR[55]), .CP(n194), .CDN(n190), .Q(
        FrameSR[56]) );
  DFCND1 \FrameSR_reg[57]  ( .D(FrameSR[56]), .CP(n196), .CDN(n188), .Q(
        FrameSR[57]) );
  DFCND1 \FrameSR_reg[58]  ( .D(FrameSR[57]), .CP(n195), .CDN(n190), .Q(
        FrameSR[58]) );
  DFCND1 \FrameSR_reg[59]  ( .D(FrameSR[58]), .CP(N4), .CDN(n22), .Q(
        FrameSR[59]) );
  DFCND1 \FrameSR_reg[60]  ( .D(FrameSR[59]), .CP(n195), .CDN(n187), .Q(
        FrameSR[60]) );
  DFCND1 \FrameSR_reg[61]  ( .D(FrameSR[60]), .CP(n194), .CDN(n189), .Q(
        FrameSR[61]) );
  DFCND1 \FrameSR_reg[62]  ( .D(FrameSR[61]), .CP(n194), .CDN(n189), .Q(
        FrameSR[62]) );
  DFCND1 \DecodeReg_reg[9]  ( .D(n68), .CP(n194), .CDN(n187), .Q(DecodeReg[9])
         );
  DFCND1 \DecodeReg_reg[31]  ( .D(n90), .CP(n195), .CDN(n189), .Q(
        DecodeReg[31]) );
  DFCND1 \DecodeReg_reg[30]  ( .D(n89), .CP(N4), .CDN(n189), .Q(DecodeReg[30])
         );
  DFCND1 \DecodeReg_reg[29]  ( .D(n88), .CP(n194), .CDN(n189), .Q(
        DecodeReg[29]) );
  DFCND1 \DecodeReg_reg[28]  ( .D(n87), .CP(n196), .CDN(n189), .Q(
        DecodeReg[28]) );
  DFCND1 \DecodeReg_reg[27]  ( .D(n86), .CP(N4), .CDN(n189), .Q(DecodeReg[27])
         );
  DFCND1 \DecodeReg_reg[26]  ( .D(n85), .CP(n194), .CDN(n189), .Q(
        DecodeReg[26]) );
  DFCND1 \DecodeReg_reg[25]  ( .D(n84), .CP(N4), .CDN(n189), .Q(DecodeReg[25])
         );
  DFCND1 \DecodeReg_reg[24]  ( .D(n83), .CP(n196), .CDN(n189), .Q(
        DecodeReg[24]) );
  DFCND1 \DecodeReg_reg[23]  ( .D(n82), .CP(N4), .CDN(n188), .Q(DecodeReg[23])
         );
  DFCND1 \DecodeReg_reg[22]  ( .D(n81), .CP(n196), .CDN(n188), .Q(
        DecodeReg[22]) );
  DFCND1 \DecodeReg_reg[21]  ( .D(n80), .CP(N4), .CDN(n188), .Q(DecodeReg[21])
         );
  DFCND1 \DecodeReg_reg[20]  ( .D(n79), .CP(n195), .CDN(n188), .Q(
        DecodeReg[20]) );
  DFCND1 \DecodeReg_reg[19]  ( .D(n78), .CP(n195), .CDN(n188), .Q(
        DecodeReg[19]) );
  DFCND1 \DecodeReg_reg[18]  ( .D(n77), .CP(n194), .CDN(n188), .Q(
        DecodeReg[18]) );
  DFCND1 \DecodeReg_reg[17]  ( .D(n76), .CP(N4), .CDN(n188), .Q(DecodeReg[17])
         );
  DFCND1 \DecodeReg_reg[16]  ( .D(n75), .CP(n196), .CDN(n188), .Q(
        DecodeReg[16]) );
  DFCND1 \DecodeReg_reg[15]  ( .D(n74), .CP(n196), .CDN(n188), .Q(
        DecodeReg[15]) );
  DFCND1 \DecodeReg_reg[14]  ( .D(n73), .CP(n196), .CDN(n188), .Q(
        DecodeReg[14]) );
  DFCND1 \DecodeReg_reg[13]  ( .D(n72), .CP(n194), .CDN(n188), .Q(
        DecodeReg[13]) );
  DFCND1 \DecodeReg_reg[12]  ( .D(n71), .CP(n196), .CDN(n188), .Q(
        DecodeReg[12]) );
  DFCND1 \DecodeReg_reg[11]  ( .D(n70), .CP(n194), .CDN(n22), .Q(DecodeReg[11]) );
  DFCND1 \DecodeReg_reg[10]  ( .D(n69), .CP(N4), .CDN(n22), .Q(DecodeReg[10])
         );
  DFCND1 \DecodeReg_reg[8]  ( .D(n67), .CP(n194), .CDN(n190), .Q(DecodeReg[8])
         );
  DFCND1 \DecodeReg_reg[7]  ( .D(n66), .CP(N4), .CDN(n22), .Q(DecodeReg[7]) );
  DFCND1 \DecodeReg_reg[6]  ( .D(n65), .CP(N4), .CDN(n187), .Q(DecodeReg[6])
         );
  DFCND1 \DecodeReg_reg[5]  ( .D(n64), .CP(n196), .CDN(n187), .Q(DecodeReg[5])
         );
  DFCND1 \DecodeReg_reg[4]  ( .D(n63), .CP(n194), .CDN(n22), .Q(DecodeReg[4])
         );
  DFCND1 \DecodeReg_reg[3]  ( .D(n62), .CP(n196), .CDN(n22), .Q(DecodeReg[3])
         );
  DFCND1 \DecodeReg_reg[2]  ( .D(n61), .CP(N4), .CDN(n190), .Q(DecodeReg[2])
         );
  DFCND1 \DecodeReg_reg[1]  ( .D(n60), .CP(n194), .CDN(n187), .Q(DecodeReg[1])
         );
  DFCND1 \DecodeReg_reg[0]  ( .D(n59), .CP(N4), .CDN(n190), .Q(DecodeReg[0])
         );
  DFCND1 \FrameSR_reg[0]  ( .D(SerIn), .CP(n194), .CDN(n188), .Q(FrameSR[0])
         );
  DFCND1 \FrameSR_reg[4]  ( .D(FrameSR[3]), .CP(N4), .CDN(n188), .Q(FrameSR[4]) );
  DFCND1 \FrameSR_reg[20]  ( .D(FrameSR[19]), .CP(n196), .CDN(n190), .Q(
        FrameSR[20]) );
  DFCND1 \FrameSR_reg[34]  ( .D(FrameSR[33]), .CP(n195), .CDN(n189), .Q(
        FrameSR[34]) );
  DFCND1 \FrameSR_reg[49]  ( .D(FrameSR[48]), .CP(N4), .CDN(n189), .Q(
        FrameSR[49]) );
  DFCND1 \FrameSR_reg[2]  ( .D(FrameSR[1]), .CP(n195), .CDN(n187), .Q(
        FrameSR[2]) );
  DFCND1 \FrameSR_reg[6]  ( .D(FrameSR[5]), .CP(n196), .CDN(n189), .Q(
        FrameSR[6]) );
  DFCND1 \FrameSR_reg[18]  ( .D(FrameSR[17]), .CP(n195), .CDN(n189), .Q(
        FrameSR[18]) );
  DFCND1 \FrameSR_reg[33]  ( .D(FrameSR[32]), .CP(n195), .CDN(n189), .Q(
        FrameSR[33]) );
  DFCND1 \FrameSR_reg[48]  ( .D(FrameSR[47]), .CP(N4), .CDN(n188), .Q(
        FrameSR[48]) );
  DFCND1 \FrameSR_reg[1]  ( .D(FrameSR[0]), .CP(n194), .CDN(n188), .Q(
        FrameSR[1]) );
  DFCND1 \FrameSR_reg[3]  ( .D(FrameSR[2]), .CP(N4), .CDN(n187), .Q(FrameSR[3]) );
  DFCND1 \FrameSR_reg[5]  ( .D(FrameSR[4]), .CP(n195), .CDN(n190), .Q(
        FrameSR[5]) );
  DFCND1 \FrameSR_reg[7]  ( .D(FrameSR[6]), .CP(n196), .CDN(n22), .Q(
        FrameSR[7]) );
  DFCND1 \FrameSR_reg[21]  ( .D(FrameSR[20]), .CP(n194), .CDN(n188), .Q(
        FrameSR[21]) );
  DFCND1 \FrameSR_reg[35]  ( .D(FrameSR[34]), .CP(n195), .CDN(n187), .Q(
        FrameSR[35]) );
  DFCND1 \FrameSR_reg[50]  ( .D(FrameSR[49]), .CP(n194), .CDN(n187), .Q(
        FrameSR[50]) );
  DFCND1 doParSync_reg ( .D(n58), .CP(n194), .CDN(n188), .Q(doParSync) );
  DFCND1 \FrameSR_reg[51]  ( .D(FrameSR[50]), .CP(N4), .CDN(n22), .Q(
        FrameSR[51]) );
  DFCND1 \FrameSR_reg[36]  ( .D(FrameSR[35]), .CP(N4), .CDN(n22), .Q(
        FrameSR[36]) );
  DFCND1 \FrameSR_reg[52]  ( .D(FrameSR[51]), .CP(n194), .CDN(n187), .Q(
        FrameSR[52]) );
  DFCND1 \FrameSR_reg[17]  ( .D(FrameSR[16]), .CP(n195), .CDN(n22), .Q(
        FrameSR[17]) );
  DFCND1 \FrameSR_reg[16]  ( .D(FrameSR[15]), .CP(n195), .CDN(n187), .Q(
        FrameSR[16]) );
  DFCND1 \ParOutReg_reg[0]  ( .D(n56), .CP(n194), .CDN(n188), .Q(ParOut[0]), 
        .QN(net389) );
  DFCND1 \ParOutReg_reg[1]  ( .D(n55), .CP(n194), .CDN(n190), .Q(ParOut[1]), 
        .QN(net390) );
  DFCND1 \ParOutReg_reg[2]  ( .D(n54), .CP(n196), .CDN(n189), .Q(ParOut[2]), 
        .QN(net391) );
  DFCND1 \ParOutReg_reg[3]  ( .D(n53), .CP(n194), .CDN(n190), .Q(ParOut[3]), 
        .QN(net392) );
  DFCND1 \ParOutReg_reg[4]  ( .D(n52), .CP(n195), .CDN(n22), .Q(ParOut[4]), 
        .QN(net393) );
  DFCND1 \ParOutReg_reg[5]  ( .D(n51), .CP(n195), .CDN(n190), .Q(ParOut[5]), 
        .QN(net394) );
  DFCND1 \ParOutReg_reg[6]  ( .D(n50), .CP(n194), .CDN(n187), .Q(ParOut[6]), 
        .QN(net395) );
  DFCND1 \ParOutReg_reg[7]  ( .D(n49), .CP(N4), .CDN(n187), .Q(ParOut[7]), 
        .QN(net396) );
  DFCND1 \ParOutReg_reg[8]  ( .D(n48), .CP(n194), .CDN(n187), .Q(ParOut[8]), 
        .QN(net397) );
  DFCND1 \ParOutReg_reg[9]  ( .D(n47), .CP(n196), .CDN(n190), .Q(ParOut[9]), 
        .QN(net398) );
  DFCND1 \ParOutReg_reg[10]  ( .D(n46), .CP(n194), .CDN(n22), .Q(ParOut[10]), 
        .QN(net399) );
  DFCND1 \ParOutReg_reg[11]  ( .D(n45), .CP(n195), .CDN(n22), .Q(ParOut[11]), 
        .QN(net400) );
  DFCND1 \ParOutReg_reg[12]  ( .D(n44), .CP(n196), .CDN(n189), .Q(ParOut[12]), 
        .QN(net401) );
  DFCND1 \ParOutReg_reg[13]  ( .D(n43), .CP(n194), .CDN(n188), .Q(ParOut[13]), 
        .QN(net402) );
  DFCND1 \ParOutReg_reg[14]  ( .D(n42), .CP(n196), .CDN(n190), .Q(ParOut[14]), 
        .QN(net403) );
  DFCND1 \ParOutReg_reg[15]  ( .D(n41), .CP(n196), .CDN(n189), .Q(ParOut[15]), 
        .QN(net404) );
  DFCND1 \ParOutReg_reg[16]  ( .D(n40), .CP(n196), .CDN(n188), .Q(ParOut[16]), 
        .QN(net405) );
  DFCND1 \ParOutReg_reg[17]  ( .D(n39), .CP(n194), .CDN(n22), .Q(ParOut[17]), 
        .QN(net406) );
  DFCND1 \ParOutReg_reg[18]  ( .D(n38), .CP(N4), .CDN(n187), .Q(ParOut[18]), 
        .QN(net407) );
  DFCND1 \ParOutReg_reg[19]  ( .D(n37), .CP(N4), .CDN(n190), .Q(ParOut[19]), 
        .QN(net408) );
  DFCND1 \ParOutReg_reg[20]  ( .D(n36), .CP(n194), .CDN(n22), .Q(ParOut[20]), 
        .QN(net409) );
  DFCND1 \ParOutReg_reg[21]  ( .D(n35), .CP(n194), .CDN(n190), .Q(ParOut[21]), 
        .QN(net410) );
  DFCND1 \ParOutReg_reg[22]  ( .D(n34), .CP(n195), .CDN(n187), .Q(ParOut[22]), 
        .QN(net411) );
  DFCND1 \ParOutReg_reg[23]  ( .D(n33), .CP(n196), .CDN(n189), .Q(ParOut[23]), 
        .QN(net412) );
  DFCND1 \ParOutReg_reg[24]  ( .D(n32), .CP(N4), .CDN(n187), .Q(ParOut[24]), 
        .QN(net413) );
  DFCND1 \ParOutReg_reg[25]  ( .D(n31), .CP(N4), .CDN(n22), .Q(ParOut[25]), 
        .QN(net414) );
  DFCND1 \ParOutReg_reg[26]  ( .D(n30), .CP(N4), .CDN(n190), .Q(ParOut[26]), 
        .QN(net415) );
  DFCND1 \ParOutReg_reg[27]  ( .D(n29), .CP(N4), .CDN(n22), .Q(ParOut[27]), 
        .QN(net416) );
  DFCND1 \ParOutReg_reg[28]  ( .D(n28), .CP(N4), .CDN(n189), .Q(ParOut[28]), 
        .QN(net417) );
  DFCND1 \ParOutReg_reg[29]  ( .D(n27), .CP(N4), .CDN(n188), .Q(ParOut[29]), 
        .QN(net418) );
  DFCND1 \ParOutReg_reg[30]  ( .D(n26), .CP(n195), .CDN(n189), .Q(ParOut[30]), 
        .QN(net419) );
  DFCND1 \ParOutReg_reg[31]  ( .D(n25), .CP(N4), .CDN(n22), .Q(ParOut[31]), 
        .QN(net420) );
  DFCND1 ParValidReg_reg ( .D(n24), .CP(n194), .CDN(n190), .Q(ParValid) );
  DFCND1 UnLoad_reg ( .D(n191), .CP(n196), .CDN(n189), .Q(UnLoad) );
  LHQD4 ParClkReg_reg ( .E(N64), .D(n4), .Q(ParClk) );
  AO21D0 U3 ( .A1(ParClk), .A2(ParValid), .B(n192), .Z(n24) );
  OR2D0 U4 ( .A1(ParClk), .A2(n5), .Z(n1) );
  INVD0 U5 ( .I(n1), .ZN(n4) );
  BUFFD1 U38 ( .I(n190), .Z(n188) );
  BUFFD1 U39 ( .I(n190), .Z(n189) );
  BUFFD1 U40 ( .I(n187), .Z(n190) );
  INVD1 U41 ( .I(n11), .ZN(n191) );
  BUFFD1 U42 ( .I(n22), .Z(n187) );
  IND2D1 U43 ( .A1(n3), .B1(n2), .ZN(n11) );
  INVD1 U44 ( .I(Reset), .ZN(n22) );
  ND2D1 U45 ( .A1(n6), .A2(n188), .ZN(N71) );
  INR2D1 U47 ( .A1(N55), .B1(n5), .ZN(N72) );
  INR2D1 U48 ( .A1(N54), .B1(n5), .ZN(N70) );
  INR2D1 U49 ( .A1(N53), .B1(n5), .ZN(N69) );
  NR2D1 U50 ( .A1(n5), .A2(n7), .ZN(N68) );
  NR2D1 U51 ( .A1(n5), .A2(n8), .ZN(N67) );
  INVD1 U52 ( .I(N52), .ZN(n7) );
  NR2D1 U53 ( .A1(n2), .A2(n3), .ZN(n58) );
  BUFFD1 U54 ( .I(n192), .Z(n193) );
  BUFFD1 U55 ( .I(n196), .Z(n195) );
  NR4D0 U56 ( .A1(n16), .A2(FrameSR[48]), .A3(FrameSR[50]), .A4(FrameSR[49]), 
        .ZN(n15) );
  INVD1 U57 ( .I(SerValid), .ZN(n6) );
  ND2D1 U58 ( .A1(n20), .A2(n21), .ZN(n3) );
  NR4D0 U59 ( .A1(FrameSR[3]), .A2(FrameSR[2]), .A3(FrameSR[1]), .A4(
        FrameSR[0]), .ZN(n20) );
  NR4D0 U60 ( .A1(FrameSR[7]), .A2(FrameSR[6]), .A3(FrameSR[5]), .A4(
        FrameSR[4]), .ZN(n21) );
  INR3D0 U61 ( .A1(SerClk), .B1(Reset), .B2(n6), .ZN(N66) );
  AN4D1 U62 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .Z(n2) );
  INR4D0 U63 ( .A1(FrameSR[19]), .B1(n19), .B2(FrameSR[17]), .B3(FrameSR[16]), 
        .ZN(n12) );
  NR4D0 U64 ( .A1(n18), .A2(FrameSR[18]), .A3(FrameSR[21]), .A4(FrameSR[20]), 
        .ZN(n13) );
  NR4D0 U65 ( .A1(n17), .A2(FrameSR[33]), .A3(FrameSR[35]), .A4(FrameSR[34]), 
        .ZN(n14) );
  OAI21D1 U66 ( .A1(n9), .A2(n6), .B(n187), .ZN(N64) );
  AOI31D0 U67 ( .A1(n8), .A2(n7), .A3(n10), .B(doParSync), .ZN(n9) );
  NR3D0 U68 ( .A1(N53), .A2(N55), .A3(N54), .ZN(n10) );
  INVD1 U69 ( .I(N51), .ZN(n8) );
  ND3D1 U70 ( .A1(FrameSR[51]), .A2(FrameSR[36]), .A3(FrameSR[52]), .ZN(n19)
         );
  AO22D0 U71 ( .A1(FrameSR[8]), .A2(n191), .B1(DecodeReg[0]), .B2(n11), .Z(n59) );
  AO22D0 U72 ( .A1(FrameSR[9]), .A2(n191), .B1(DecodeReg[1]), .B2(n11), .Z(n60) );
  AO22D0 U73 ( .A1(FrameSR[10]), .A2(n191), .B1(DecodeReg[2]), .B2(n11), .Z(
        n61) );
  AO22D0 U74 ( .A1(FrameSR[11]), .A2(n191), .B1(DecodeReg[3]), .B2(n11), .Z(
        n62) );
  AO22D0 U75 ( .A1(FrameSR[12]), .A2(n191), .B1(DecodeReg[4]), .B2(n11), .Z(
        n63) );
  AO22D0 U76 ( .A1(FrameSR[13]), .A2(n191), .B1(DecodeReg[5]), .B2(n11), .Z(
        n64) );
  AO22D0 U77 ( .A1(FrameSR[14]), .A2(n191), .B1(DecodeReg[6]), .B2(n11), .Z(
        n65) );
  AO22D0 U78 ( .A1(FrameSR[15]), .A2(n191), .B1(DecodeReg[7]), .B2(n11), .Z(
        n66) );
  AO22D0 U79 ( .A1(FrameSR[24]), .A2(n191), .B1(DecodeReg[8]), .B2(n11), .Z(
        n67) );
  AO22D0 U80 ( .A1(FrameSR[25]), .A2(n191), .B1(DecodeReg[9]), .B2(n11), .Z(
        n68) );
  AO22D0 U81 ( .A1(FrameSR[26]), .A2(n191), .B1(DecodeReg[10]), .B2(n11), .Z(
        n69) );
  AO22D0 U82 ( .A1(FrameSR[27]), .A2(n191), .B1(DecodeReg[11]), .B2(n11), .Z(
        n70) );
  AO22D0 U83 ( .A1(FrameSR[28]), .A2(n191), .B1(DecodeReg[12]), .B2(n11), .Z(
        n71) );
  AO22D0 U84 ( .A1(FrameSR[29]), .A2(n191), .B1(DecodeReg[13]), .B2(n11), .Z(
        n72) );
  AO22D0 U85 ( .A1(FrameSR[30]), .A2(n191), .B1(DecodeReg[14]), .B2(n11), .Z(
        n73) );
  AO22D0 U86 ( .A1(FrameSR[31]), .A2(n191), .B1(DecodeReg[15]), .B2(n11), .Z(
        n74) );
  AO22D0 U87 ( .A1(FrameSR[40]), .A2(n191), .B1(DecodeReg[16]), .B2(n11), .Z(
        n75) );
  AO22D0 U88 ( .A1(FrameSR[41]), .A2(n191), .B1(DecodeReg[17]), .B2(n11), .Z(
        n76) );
  AO22D0 U89 ( .A1(FrameSR[42]), .A2(n191), .B1(DecodeReg[18]), .B2(n11), .Z(
        n77) );
  AO22D0 U91 ( .A1(FrameSR[43]), .A2(n191), .B1(DecodeReg[19]), .B2(n11), .Z(
        n78) );
  AO22D0 U93 ( .A1(FrameSR[44]), .A2(n191), .B1(DecodeReg[20]), .B2(n11), .Z(
        n79) );
  AO22D0 U95 ( .A1(FrameSR[45]), .A2(n191), .B1(DecodeReg[21]), .B2(n11), .Z(
        n80) );
  AO22D0 U96 ( .A1(FrameSR[46]), .A2(n191), .B1(DecodeReg[22]), .B2(n11), .Z(
        n81) );
  AO22D0 U97 ( .A1(FrameSR[47]), .A2(n191), .B1(DecodeReg[23]), .B2(n11), .Z(
        n82) );
  AO22D0 U98 ( .A1(FrameSR[56]), .A2(n191), .B1(DecodeReg[24]), .B2(n11), .Z(
        n83) );
  AO22D0 U99 ( .A1(FrameSR[57]), .A2(n191), .B1(DecodeReg[25]), .B2(n11), .Z(
        n84) );
  AO22D0 U100 ( .A1(FrameSR[58]), .A2(n191), .B1(DecodeReg[26]), .B2(n11), .Z(
        n85) );
  AO22D0 U101 ( .A1(FrameSR[59]), .A2(n191), .B1(DecodeReg[27]), .B2(n11), .Z(
        n86) );
  AO22D0 U102 ( .A1(FrameSR[60]), .A2(n191), .B1(DecodeReg[28]), .B2(n11), .Z(
        n87) );
  AO22D0 U103 ( .A1(FrameSR[61]), .A2(n191), .B1(DecodeReg[29]), .B2(n11), .Z(
        n88) );
  AO22D0 U104 ( .A1(FrameSR[62]), .A2(n191), .B1(DecodeReg[30]), .B2(n11), .Z(
        n89) );
  AO22D0 U105 ( .A1(FrameSR[63]), .A2(n191), .B1(DecodeReg[31]), .B2(n11), .Z(
        n90) );
  BUFFD1 U106 ( .I(UnLoad), .Z(n192) );
  BUFFD1 U107 ( .I(n194), .Z(n196) );
  BUFFD1 U108 ( .I(N4), .Z(n194) );
endmodule


module SerialRx ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;


  PLLTop PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(Reset) );
  BUFFD1 U1 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n828, n829, n830, n831, n832, StateClockRaw, StateClock, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N68, N69, N70, N71, N72, N73,
         N78, N176, N177, N178, N330, N332, N333, N334, n6, n8, n9, n10, n12,
         n15, n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n86, n87, n88, n89, n90,
         n91, n93, n94, n96, n98, n99, n100, n101, n103, n104, n105, n106,
         n107, n108, n109, n121, n123, n124, n127, n128, n130, n131, n132,
         n133, n134, n136, n143, n144, \add_388/carry[2] , \add_388/carry[3] ,
         \add_388/carry[4] , \add_307/carry[3] , \add_307/carry[4] , n1, n2,
         n3, n4, n5, n7, n11, n13, n14, n21, n69, n70, n71, n84, n85, n92, n95,
         n97, n102, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n122, n125, n126, n129, n135, n137, n138, n139, n140, n141,
         n142, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n798, n799, n800, n801, n802, n803, n804, n820, n822, n823,
         n825, n826, n827;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [4:0] OldReadAr;
  wire   [4:0] OldWriteAr;
  assign WriteAddr[0] = N330;
  assign WriteAddr[1] = \add_388/carry[2] ;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  MOAI22D1 U24 ( .A1(n29), .A2(n30), .B1(n31), .B2(CurState[2]), .ZN(n27) );
  OR3D1 U41 ( .A1(n49), .A2(CurState[2]), .A3(n50), .Z(n47) );
  OA21D1 U111 ( .A1(CurState[2]), .A2(n29), .B(n83), .Z(n35) );
  FIFOStateM_AWid5_DW01_inc_0 r110 ( .A({WriteAddr[4:2], \add_388/carry[2] , 
        n650}), .SUM({N72, N71, N70, N69, N68}) );
  FIFOStateM_AWid5_DW01_inc_1 r109 ( .A({ReadAddr[4], n625, ReadAddr[2], n682, 
        n645}), .SUM({N48, N47, N46, N45, N44}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n388), .CPN(StateClock), .CDN(n820), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n1), .CPN(StateClock), .CDN(n143), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n400), .CPN(StateClock), .CDN(n820), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n11), .CPN(StateClock), .CDN(n820), .Q(
        OldReadAr[1]) );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n13), .CPN(StateClock), .CDN(n820), .Q(
        OldWriteAr[4]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n434), .CPN(StateClock), .CDN(n143), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n449), .CPN(StateClock), .CDN(n820), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n462), .CPN(StateClock), .CDN(n820), .Q(
        OldReadAr[4]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n92), .CPN(StateClock), .CDN(n820), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n111), .CPN(StateClock), .CDN(n820), .Q(
        OldReadAr[3]) );
  DFNCND1 \NextState_reg[1]  ( .D(n116), .CPN(StateClock), .CDN(n820), .Q(
        NextState[1]), .QN(n124) );
  DFNCND1 \NextState_reg[0]  ( .D(n514), .CPN(StateClock), .CDN(n143), .Q(
        NextState[0]), .QN(n123) );
  DFNCND1 \NextState_reg[2]  ( .D(n129), .CPN(StateClock), .CDN(n143), .Q(
        NextState[2]), .QN(n121) );
  DFNCND1 ReadCmdr_reg ( .D(n541), .CPN(StateClock), .CDN(n143), .Q(n831) );
  DFNCND1 WriteCmdr_reg ( .D(n152), .CPN(StateClock), .CDN(n820), .Q(n832) );
  EDFCNQD1 \WriteAr_reg[4]  ( .D(n157), .E(n651), .CP(StateClock), .CDN(n820), 
        .Q(WriteAddr[4]) );
  EDFCNQD1 \WriteAr_reg[3]  ( .D(n159), .E(n651), .CP(StateClock), .CDN(n820), 
        .Q(WriteAddr[3]) );
  EDFCNQD1 \ReadAr_reg[2]  ( .D(n593), .E(N53), .CP(StateClock), .CDN(n820), 
        .Q(n829) );
  EDFCNQD1 \ReadAr_reg[4]  ( .D(n162), .E(N53), .CP(StateClock), .CDN(n143), 
        .Q(n828) );
  EDFCNQD1 \WriteAr_reg[2]  ( .D(n168), .E(n651), .CP(StateClock), .CDN(n820), 
        .Q(n830) );
  EDFCNQD1 \ReadAr_reg[3]  ( .D(n175), .E(N53), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[3]) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(n627), .E(n651), .CP(StateClock), .CDN(n143), 
        .Q(\add_388/carry[2] ) );
  EDFCNQD1 \WriteAr_reg[0]  ( .D(n176), .E(n651), .CP(StateClock), .CDN(n143), 
        .Q(N330) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[2]), .QN(n96) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[1]), .QN(n29) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[0]), .QN(n55) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n185), .E(N53), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[1]), .QN(n825) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n687), .E(N53), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[0]), .QN(n822) );
  DFND1 FullFIFOr_reg ( .D(n132), .CPN(StateClock), .QN(n206) );
  DFND4 EmptyFIFOr_reg ( .D(n127), .CPN(StateClock), .Q(EmptyFIFO) );
  BUFFD0 U3 ( .I(n3), .Z(n1) );
  XOR2D0 U4 ( .A1(WriteAddr[3]), .A2(n562), .Z(n39) );
  XOR2D0 U5 ( .A1(WriteAddr[2]), .A2(n560), .Z(n40) );
  BUFFD0 U6 ( .I(n5), .Z(n428) );
  BUFFD0 U7 ( .I(n195), .Z(n2) );
  BUFFD0 U8 ( .I(n208), .Z(n3) );
  BUFFD0 U9 ( .I(OldWriteAr[0]), .Z(n4) );
  BUFFD0 U10 ( .I(n4), .Z(n5) );
  CKNXD0 U11 ( .I(n418), .ZN(n419) );
  INVD8 U12 ( .I(n202), .ZN(n7) );
  INVD1 U13 ( .I(n7), .ZN(n11) );
  INVD0 U14 ( .I(OldReadAr[1]), .ZN(n413) );
  BUFFD0 U15 ( .I(n14), .Z(n13) );
  BUFFD0 U16 ( .I(n21), .Z(n14) );
  BUFFD0 U17 ( .I(n69), .Z(n21) );
  BUFFD0 U18 ( .I(n70), .Z(n69) );
  BUFFD0 U19 ( .I(n71), .Z(n70) );
  BUFFD0 U20 ( .I(n84), .Z(n71) );
  BUFFD0 U21 ( .I(n85), .Z(n84) );
  BUFFD0 U22 ( .I(n216), .Z(n85) );
  INVD3 U23 ( .I(n464), .ZN(n461) );
  INVD0 U25 ( .I(n131), .ZN(n463) );
  CKNXD16 U26 ( .I(n201), .ZN(n131) );
  CKND12 U27 ( .CLK(n475), .CN(n476) );
  BUFFD0 U28 ( .I(n476), .Z(n92) );
  BUFFD0 U29 ( .I(n97), .Z(n95) );
  BUFFD0 U30 ( .I(n102), .Z(n97) );
  BUFFD0 U31 ( .I(n482), .Z(n102) );
  CKBD0 U32 ( .CLK(n484), .C(n110) );
  BUFFD16 U33 ( .I(n110), .Z(n479) );
  CKND12 U34 ( .CLK(n488), .CN(n489) );
  BUFFD0 U35 ( .I(n112), .Z(n111) );
  MOAI22D0 U36 ( .A1(n199), .A2(n113), .B1(n625), .B2(n8), .ZN(n128) );
  BUFFD0 U37 ( .I(n489), .Z(n112) );
  BUFFD0 U38 ( .I(n114), .Z(n113) );
  BUFFD0 U39 ( .I(n495), .Z(n114) );
  CKBD0 U40 ( .CLK(n497), .C(n115) );
  BUFFD16 U42 ( .I(n115), .Z(n492) );
  BUFFD0 U43 ( .I(n501), .Z(n116) );
  BUFFD0 U44 ( .I(n124), .Z(n117) );
  BUFFD0 U45 ( .I(n117), .Z(n118) );
  BUFFD0 U46 ( .I(n118), .Z(n119) );
  BUFFD0 U47 ( .I(n119), .Z(n120) );
  BUFFD0 U48 ( .I(n120), .Z(n122) );
  BUFFD0 U49 ( .I(n122), .Z(n125) );
  BUFFD0 U50 ( .I(n125), .Z(n126) );
  OA21D0 U51 ( .A1(n24), .A2(n518), .B(n42), .Z(n197) );
  BUFFD0 U52 ( .I(n528), .Z(n129) );
  BUFFD0 U53 ( .I(n121), .Z(n135) );
  BUFFD0 U54 ( .I(n135), .Z(n137) );
  BUFFD0 U55 ( .I(n137), .Z(n138) );
  BUFFD0 U56 ( .I(n138), .Z(n139) );
  BUFFD0 U57 ( .I(n139), .Z(n140) );
  BUFFD0 U58 ( .I(n140), .Z(n141) );
  BUFFD0 U59 ( .I(n141), .Z(n142) );
  INVD4 U60 ( .I(n542), .ZN(n145) );
  CKBXD0 U61 ( .I(n544), .Z(n542) );
  CKNXD0 U62 ( .I(n543), .ZN(n544) );
  CKNXD16 U63 ( .I(n546), .ZN(n543) );
  INVD1 U64 ( .I(n145), .ZN(n146) );
  BUFFD0 U65 ( .I(n204), .Z(n147) );
  BUFFD0 U66 ( .I(n147), .Z(n148) );
  BUFFD0 U67 ( .I(OldReadAr[4]), .Z(n149) );
  BUFFD0 U68 ( .I(OldReadAr[0]), .Z(n150) );
  CKXOR2D0 U69 ( .A1(ReadAddr[4]), .A2(n474), .Z(n108) );
  CKBXD0 U70 ( .I(n150), .Z(n397) );
  ND3D0 U71 ( .A1(n103), .A2(n104), .A3(n105), .ZN(n194) );
  CKBD0 U72 ( .CLK(n34), .C(n151) );
  BUFFD0 U73 ( .I(n154), .Z(n152) );
  BUFFD0 U74 ( .I(n566), .Z(n153) );
  BUFFD0 U75 ( .I(n552), .Z(n154) );
  BUFFD0 U76 ( .I(n186), .Z(n155) );
  BUFFD0 U77 ( .I(n153), .Z(n156) );
  CKND2D0 U78 ( .A1(n156), .A2(n653), .ZN(n34) );
  INVD2P5 U79 ( .I(n190), .ZN(n567) );
  BUFFD0 U80 ( .I(n158), .Z(n157) );
  BUFFD0 U81 ( .I(n569), .Z(n158) );
  BUFFD0 U82 ( .I(n160), .Z(n159) );
  CKBD0 U83 ( .CLK(n581), .C(n160) );
  INVD0 U84 ( .I(n189), .ZN(n590) );
  OAI22D4 U85 ( .A1(n826), .A2(n653), .B1(n161), .B2(n34), .ZN(n189) );
  BUFFD0 U86 ( .I(n74), .Z(n161) );
  INVD10 U87 ( .I(n599), .ZN(n600) );
  CKND2D0 U88 ( .A1(N48), .A2(n193), .ZN(n192) );
  BUFFD0 U89 ( .I(n163), .Z(n162) );
  BUFFD0 U90 ( .I(n164), .Z(n163) );
  BUFFD0 U91 ( .I(n598), .Z(n164) );
  BUFFD0 U92 ( .I(n828), .Z(n165) );
  BUFFD0 U93 ( .I(n188), .Z(n166) );
  BUFFD0 U94 ( .I(n166), .Z(n167) );
  BUFFD0 U95 ( .I(n609), .Z(n168) );
  INVD16 U96 ( .I(N52), .ZN(n169) );
  INVD1 U97 ( .I(n169), .ZN(n170) );
  BUFFD0 U98 ( .I(n172), .Z(n171) );
  BUFFD0 U99 ( .I(n173), .Z(n172) );
  BUFFD0 U100 ( .I(n174), .Z(n173) );
  BUFFD0 U101 ( .I(n622), .Z(n174) );
  BUFFD0 U102 ( .I(n621), .Z(n175) );
  INR2D0 U103 ( .A1(n171), .B1(n99), .ZN(N52) );
  CKBXD0 U104 ( .I(n649), .Z(n650) );
  CKND1 U105 ( .CLK(n648), .CN(n649) );
  BUFFD0 U106 ( .I(n177), .Z(n176) );
  BUFFD0 U107 ( .I(n178), .Z(n177) );
  CKBD0 U108 ( .CLK(n640), .C(n178) );
  CKNXD16 U109 ( .I(n639), .ZN(n640) );
  CKNXD0 U110 ( .I(n644), .ZN(n639) );
  INVD0 U112 ( .I(n647), .ZN(n643) );
  INVD0 U113 ( .I(n641), .ZN(n642) );
  CKNXD16 U114 ( .I(N73), .ZN(n641) );
  CKBD0 U115 ( .CLK(n674), .C(n672) );
  INVD16 U116 ( .I(N50), .ZN(n179) );
  INVD1 U117 ( .I(n179), .ZN(n180) );
  BUFFD0 U118 ( .I(n182), .Z(n181) );
  BUFFD0 U119 ( .I(n183), .Z(n182) );
  BUFFD0 U120 ( .I(n184), .Z(n183) );
  BUFFD0 U121 ( .I(n678), .Z(n184) );
  BUFFD0 U122 ( .I(n677), .Z(n185) );
  INR2D0 U123 ( .A1(n181), .B1(n99), .ZN(N50) );
  INVD0 U124 ( .I(n686), .ZN(n687) );
  INVD5 U125 ( .I(N49), .ZN(n686) );
  INR2D0 U126 ( .A1(n683), .B1(n99), .ZN(N49) );
  CKBXD0 U127 ( .I(n688), .Z(n645) );
  CKBXD0 U128 ( .I(n685), .Z(n689) );
  INVD3 U129 ( .I(n99), .ZN(n193) );
  OAI32D1 U130 ( .A1(n23), .A2(n32), .A3(n33), .B1(n151), .B2(n22), .ZN(n186)
         );
  CKNXD12 U131 ( .I(n9), .ZN(n200) );
  AOI22D0 U132 ( .A1(n682), .A2(n28), .B1(N69), .B2(n109), .ZN(n187) );
  AO22D0 U133 ( .A1(N70), .A2(n109), .B1(ReadAddr[2]), .B2(n28), .Z(n188) );
  AOI22D0 U134 ( .A1(N72), .A2(n109), .B1(ReadAddr[4]), .B2(n28), .ZN(n190) );
  AOI22D0 U135 ( .A1(WriteAddr[4]), .A2(n16), .B1(n17), .B2(n218), .ZN(n191)
         );
  OA22D0 U136 ( .A1(n16), .A2(n212), .B1(n648), .B2(n17), .Z(n195) );
  CKNXD12 U137 ( .I(n596), .ZN(n597) );
  OAI22D0 U138 ( .A1(n24), .A2(n538), .B1(n25), .B2(n26), .ZN(n196) );
  OAI22D0 U139 ( .A1(n24), .A2(n511), .B1(n25), .B2(n57), .ZN(n198) );
  CKND16 U140 ( .CLK(n9), .CN(n199) );
  MOAI22D1 U141 ( .A1(n200), .A2(n95), .B1(ReadAddr[2]), .B2(n8), .ZN(n130) );
  AOI22D0 U142 ( .A1(ReadAddr[4]), .A2(n8), .B1(n9), .B2(n469), .ZN(n201) );
  OAI22D0 U143 ( .A1(n8), .A2(n419), .B1(n825), .B2(n9), .ZN(n202) );
  AO22D0 U144 ( .A1(WriteAddr[2]), .A2(n16), .B1(n17), .B2(n560), .Z(n136) );
  AO22D0 U145 ( .A1(n645), .A2(n28), .B1(N68), .B2(n109), .Z(N73) );
  CKND2D0 U146 ( .A1(n798), .A2(FullFIFO), .ZN(n203) );
  OA32D0 U147 ( .A1(n146), .A2(n98), .A3(n827), .B1(n99), .B2(n100), .Z(n204)
         );
  AO21D1 U148 ( .A1(CurState[2]), .A2(CurState[0]), .B(n15), .Z(n205) );
  INVD0 U149 ( .I(n2), .ZN(n207) );
  BUFFD0 U150 ( .I(n399), .Z(n214) );
  BUFFD0 U151 ( .I(n209), .Z(n208) );
  BUFFD0 U152 ( .I(n211), .Z(n209) );
  CKNXD16 U153 ( .I(n210), .ZN(n211) );
  INVD0 U154 ( .I(n214), .ZN(n210) );
  INVD0 U155 ( .I(n398), .ZN(n399) );
  BUFFD0 U156 ( .I(n213), .Z(n212) );
  BUFFD0 U157 ( .I(n215), .Z(n213) );
  BUFFD0 U158 ( .I(n424), .Z(n215) );
  BUFFD0 U159 ( .I(n219), .Z(n216) );
  BUFFD0 U160 ( .I(OldWriteAr[4]), .Z(n217) );
  BUFFD0 U161 ( .I(n426), .Z(n218) );
  ND3D0 U162 ( .A1(n22), .A2(n23), .A3(WriteReq), .ZN(n17) );
  BUFFD0 U163 ( .I(n220), .Z(n219) );
  BUFFD0 U164 ( .I(n221), .Z(n220) );
  BUFFD0 U165 ( .I(n222), .Z(n221) );
  BUFFD0 U166 ( .I(n223), .Z(n222) );
  BUFFD0 U167 ( .I(n224), .Z(n223) );
  BUFFD0 U168 ( .I(n225), .Z(n224) );
  BUFFD0 U169 ( .I(n226), .Z(n225) );
  BUFFD0 U170 ( .I(n227), .Z(n226) );
  BUFFD0 U171 ( .I(n228), .Z(n227) );
  BUFFD0 U172 ( .I(n229), .Z(n228) );
  BUFFD0 U173 ( .I(n427), .Z(n229) );
  ND3D0 U174 ( .A1(n657), .A2(CurState[0]), .A3(CurState[2]), .ZN(n230) );
  CKBD0 U175 ( .CLK(n144), .C(n231) );
  CKBD0 U176 ( .CLK(n206), .C(n232) );
  CKNXD16 U177 ( .I(n232), .ZN(FullFIFO) );
  BUFFD0 U178 ( .I(n566), .Z(n235) );
  BUFFD0 U179 ( .I(n235), .Z(n236) );
  BUFFD0 U180 ( .I(n236), .Z(n237) );
  BUFFD0 U181 ( .I(n237), .Z(n238) );
  BUFFD0 U182 ( .I(n238), .Z(n239) );
  BUFFD0 U183 ( .I(n239), .Z(n240) );
  BUFFD0 U184 ( .I(n240), .Z(n241) );
  BUFFD0 U185 ( .I(n241), .Z(n242) );
  BUFFD0 U186 ( .I(n242), .Z(n243) );
  BUFFD0 U187 ( .I(n243), .Z(n244) );
  BUFFD0 U188 ( .I(n244), .Z(n245) );
  BUFFD0 U189 ( .I(n245), .Z(n246) );
  BUFFD0 U190 ( .I(n246), .Z(n247) );
  BUFFD0 U191 ( .I(n247), .Z(n248) );
  BUFFD0 U192 ( .I(n248), .Z(n249) );
  BUFFD0 U193 ( .I(n249), .Z(n250) );
  BUFFD0 U194 ( .I(n250), .Z(n251) );
  BUFFD0 U195 ( .I(n251), .Z(n252) );
  BUFFD0 U196 ( .I(n252), .Z(n253) );
  BUFFD0 U197 ( .I(n253), .Z(n254) );
  BUFFD0 U198 ( .I(n254), .Z(n255) );
  BUFFD0 U199 ( .I(n255), .Z(n256) );
  BUFFD0 U200 ( .I(n256), .Z(n257) );
  BUFFD0 U201 ( .I(n257), .Z(n258) );
  BUFFD0 U202 ( .I(n258), .Z(n259) );
  BUFFD0 U203 ( .I(n259), .Z(n260) );
  BUFFD0 U204 ( .I(n260), .Z(n261) );
  BUFFD0 U205 ( .I(n261), .Z(n262) );
  BUFFD0 U206 ( .I(n262), .Z(n263) );
  BUFFD0 U207 ( .I(n263), .Z(n264) );
  BUFFD0 U208 ( .I(n264), .Z(n265) );
  BUFFD0 U209 ( .I(n265), .Z(n266) );
  BUFFD0 U210 ( .I(n266), .Z(n267) );
  BUFFD0 U211 ( .I(n267), .Z(n268) );
  BUFFD0 U212 ( .I(n268), .Z(n269) );
  BUFFD0 U213 ( .I(n269), .Z(n270) );
  BUFFD0 U214 ( .I(n270), .Z(n271) );
  BUFFD0 U215 ( .I(n271), .Z(n272) );
  BUFFD0 U216 ( .I(n272), .Z(n273) );
  BUFFD0 U217 ( .I(n273), .Z(n274) );
  BUFFD0 U218 ( .I(n274), .Z(n275) );
  BUFFD0 U219 ( .I(n275), .Z(n276) );
  BUFFD0 U220 ( .I(n276), .Z(n277) );
  BUFFD0 U221 ( .I(n277), .Z(n278) );
  BUFFD0 U222 ( .I(n278), .Z(n279) );
  BUFFD0 U223 ( .I(n279), .Z(n280) );
  BUFFD0 U224 ( .I(n280), .Z(n281) );
  BUFFD0 U225 ( .I(n281), .Z(n282) );
  BUFFD0 U226 ( .I(n282), .Z(n283) );
  BUFFD0 U227 ( .I(n283), .Z(n284) );
  BUFFD0 U228 ( .I(n284), .Z(n285) );
  BUFFD0 U229 ( .I(n285), .Z(n286) );
  BUFFD0 U230 ( .I(n286), .Z(n287) );
  BUFFD0 U231 ( .I(n287), .Z(n288) );
  BUFFD0 U232 ( .I(n288), .Z(n289) );
  BUFFD0 U233 ( .I(n289), .Z(n290) );
  BUFFD0 U234 ( .I(n290), .Z(n291) );
  BUFFD0 U235 ( .I(n291), .Z(n292) );
  BUFFD0 U236 ( .I(n292), .Z(n293) );
  BUFFD0 U237 ( .I(n293), .Z(n294) );
  BUFFD0 U238 ( .I(n294), .Z(n295) );
  BUFFD0 U239 ( .I(n295), .Z(n296) );
  BUFFD0 U240 ( .I(n296), .Z(n297) );
  BUFFD0 U241 ( .I(n297), .Z(n298) );
  BUFFD0 U242 ( .I(n298), .Z(n299) );
  BUFFD0 U243 ( .I(n299), .Z(n300) );
  BUFFD0 U244 ( .I(n300), .Z(n301) );
  BUFFD0 U245 ( .I(n301), .Z(n302) );
  BUFFD0 U246 ( .I(n302), .Z(n303) );
  BUFFD0 U247 ( .I(n303), .Z(n304) );
  BUFFD0 U248 ( .I(n304), .Z(n305) );
  BUFFD0 U249 ( .I(n305), .Z(n306) );
  BUFFD0 U250 ( .I(n306), .Z(n307) );
  BUFFD0 U251 ( .I(n307), .Z(n308) );
  BUFFD0 U252 ( .I(n308), .Z(n309) );
  BUFFD0 U253 ( .I(n309), .Z(n310) );
  BUFFD0 U254 ( .I(n310), .Z(n311) );
  BUFFD0 U255 ( .I(n311), .Z(n312) );
  BUFFD0 U256 ( .I(n312), .Z(n313) );
  BUFFD0 U257 ( .I(n313), .Z(n314) );
  BUFFD0 U258 ( .I(n314), .Z(n315) );
  BUFFD0 U259 ( .I(n315), .Z(n316) );
  BUFFD0 U260 ( .I(n316), .Z(n317) );
  BUFFD0 U261 ( .I(n317), .Z(n318) );
  BUFFD0 U262 ( .I(n318), .Z(n319) );
  BUFFD0 U263 ( .I(n319), .Z(n320) );
  BUFFD0 U264 ( .I(n320), .Z(n321) );
  BUFFD0 U265 ( .I(n321), .Z(n322) );
  BUFFD0 U266 ( .I(n322), .Z(n323) );
  BUFFD0 U267 ( .I(n323), .Z(n324) );
  BUFFD0 U268 ( .I(n324), .Z(n325) );
  BUFFD0 U269 ( .I(n325), .Z(n326) );
  BUFFD0 U270 ( .I(n326), .Z(n327) );
  BUFFD0 U271 ( .I(n327), .Z(n328) );
  BUFFD0 U272 ( .I(n328), .Z(n329) );
  BUFFD0 U273 ( .I(n329), .Z(n330) );
  BUFFD0 U274 ( .I(n330), .Z(n331) );
  BUFFD0 U275 ( .I(n331), .Z(n332) );
  BUFFD0 U276 ( .I(n332), .Z(n333) );
  BUFFD0 U277 ( .I(n333), .Z(n334) );
  BUFFD0 U278 ( .I(n334), .Z(n335) );
  BUFFD0 U279 ( .I(n335), .Z(n336) );
  BUFFD0 U280 ( .I(n336), .Z(n337) );
  BUFFD0 U281 ( .I(n337), .Z(n338) );
  BUFFD0 U282 ( .I(n338), .Z(n339) );
  BUFFD0 U283 ( .I(n339), .Z(n340) );
  BUFFD0 U284 ( .I(n340), .Z(n341) );
  BUFFD0 U285 ( .I(n341), .Z(n342) );
  BUFFD0 U286 ( .I(n342), .Z(n343) );
  BUFFD0 U287 ( .I(n343), .Z(n344) );
  BUFFD0 U288 ( .I(n344), .Z(n345) );
  BUFFD0 U289 ( .I(n345), .Z(n346) );
  BUFFD0 U290 ( .I(n346), .Z(n347) );
  BUFFD0 U291 ( .I(n347), .Z(n348) );
  BUFFD0 U292 ( .I(n348), .Z(n349) );
  BUFFD0 U293 ( .I(n349), .Z(n350) );
  BUFFD0 U294 ( .I(n350), .Z(n351) );
  BUFFD0 U295 ( .I(n351), .Z(n352) );
  BUFFD0 U296 ( .I(n352), .Z(n353) );
  BUFFD0 U297 ( .I(n353), .Z(n354) );
  BUFFD0 U298 ( .I(n354), .Z(n355) );
  BUFFD0 U299 ( .I(n355), .Z(n356) );
  BUFFD0 U300 ( .I(n356), .Z(n357) );
  BUFFD0 U301 ( .I(n357), .Z(n358) );
  BUFFD0 U302 ( .I(n358), .Z(n359) );
  BUFFD0 U303 ( .I(n359), .Z(n360) );
  BUFFD0 U304 ( .I(n360), .Z(n361) );
  BUFFD0 U305 ( .I(n361), .Z(n362) );
  BUFFD0 U306 ( .I(n362), .Z(n363) );
  BUFFD0 U307 ( .I(n363), .Z(n364) );
  BUFFD0 U308 ( .I(n364), .Z(n365) );
  BUFFD0 U309 ( .I(n365), .Z(n366) );
  BUFFD0 U310 ( .I(n366), .Z(n367) );
  BUFFD0 U311 ( .I(n367), .Z(n368) );
  BUFFD0 U312 ( .I(n368), .Z(n369) );
  BUFFD0 U313 ( .I(n369), .Z(n370) );
  BUFFD0 U314 ( .I(n370), .Z(n371) );
  BUFFD0 U315 ( .I(n371), .Z(n372) );
  BUFFD0 U316 ( .I(n372), .Z(n373) );
  BUFFD0 U317 ( .I(n373), .Z(n374) );
  BUFFD0 U318 ( .I(n374), .Z(n375) );
  BUFFD0 U319 ( .I(n375), .Z(n376) );
  BUFFD0 U320 ( .I(n376), .Z(n377) );
  BUFFD0 U321 ( .I(n377), .Z(n378) );
  BUFFD0 U322 ( .I(n378), .Z(n379) );
  BUFFD0 U323 ( .I(n379), .Z(n380) );
  BUFFD0 U324 ( .I(n380), .Z(n381) );
  BUFFD0 U325 ( .I(n381), .Z(n382) );
  BUFFD0 U326 ( .I(n382), .Z(n383) );
  BUFFD0 U327 ( .I(n832), .Z(n384) );
  BUFFD0 U328 ( .I(n384), .Z(n385) );
  CKBD0 U329 ( .CLK(n383), .C(WriteCmd) );
  INVD16 U330 ( .I(n231), .ZN(n387) );
  INVD1 U331 ( .I(n387), .ZN(n388) );
  CKNXD16 U332 ( .I(n389), .ZN(n390) );
  INVD0 U333 ( .I(n394), .ZN(n389) );
  CKBXD0 U334 ( .I(n101), .Z(n548) );
  INVD0 U335 ( .I(n391), .ZN(n392) );
  CKNXD16 U336 ( .I(n548), .ZN(n391) );
  INVD0 U337 ( .I(n393), .ZN(n394) );
  CKNXD16 U338 ( .I(n396), .ZN(n393) );
  INVD0 U339 ( .I(n395), .ZN(n396) );
  CKNXD16 U340 ( .I(n392), .ZN(n395) );
  BUFFD0 U341 ( .I(n20), .Z(n564) );
  CKNXD16 U342 ( .I(n207), .ZN(n398) );
  INVD16 U343 ( .I(n402), .ZN(n403) );
  CKND12 U344 ( .CLK(n410), .CN(n411) );
  BUFFD0 U345 ( .I(n401), .Z(n400) );
  BUFFD0 U346 ( .I(n403), .Z(n401) );
  CKNXD0 U347 ( .I(n405), .ZN(n402) );
  CKNXD16 U348 ( .I(n404), .ZN(n405) );
  CKNXD0 U349 ( .I(n407), .ZN(n404) );
  CKNXD16 U350 ( .I(n406), .ZN(n407) );
  CKNXD0 U351 ( .I(n409), .ZN(n406) );
  CKNXD16 U352 ( .I(n408), .ZN(n409) );
  CKNXD0 U353 ( .I(n411), .ZN(n408) );
  INVD0 U354 ( .I(n134), .ZN(n410) );
  OAI22D4 U355 ( .A1(n16), .A2(n550), .B1(n19), .B2(n17), .ZN(n134) );
  BUFFD0 U356 ( .I(OldWriteAr[1]), .Z(n412) );
  CKNXD0 U357 ( .I(n421), .ZN(n422) );
  CKNXD16 U358 ( .I(n413), .ZN(n414) );
  CKBXD0 U359 ( .I(n422), .Z(n415) );
  INVD0 U360 ( .I(n416), .ZN(n417) );
  CKNXD16 U361 ( .I(n415), .ZN(n416) );
  CKBD0 U362 ( .CLK(n10), .C(n547) );
  CKNXD16 U363 ( .I(n417), .ZN(n418) );
  BUFFD0 U364 ( .I(n414), .Z(n420) );
  CKNXD16 U365 ( .I(n547), .ZN(n421) );
  CKNXD16 U366 ( .I(n420), .ZN(n10) );
  INVD0 U367 ( .I(n423), .ZN(n424) );
  CKNXD16 U368 ( .I(n564), .ZN(n423) );
  CKNXD16 U369 ( .I(n425), .ZN(n426) );
  INVD0 U370 ( .I(n432), .ZN(n425) );
  INVD0 U371 ( .I(n191), .ZN(n427) );
  CKNXD16 U372 ( .I(n429), .ZN(n430) );
  INVD0 U373 ( .I(n217), .ZN(n429) );
  CKNXD16 U374 ( .I(n431), .ZN(n432) );
  CKNXD0 U375 ( .I(n430), .ZN(n431) );
  INVD12 U376 ( .I(n433), .ZN(n434) );
  INVD0 U377 ( .I(n436), .ZN(n433) );
  CKNXD16 U378 ( .I(n435), .ZN(n436) );
  CKNXD0 U379 ( .I(n438), .ZN(n435) );
  CKNXD16 U380 ( .I(n437), .ZN(n438) );
  CKNXD0 U381 ( .I(n440), .ZN(n437) );
  CKNXD16 U382 ( .I(n439), .ZN(n440) );
  CKNXD0 U383 ( .I(n442), .ZN(n439) );
  CKNXD16 U384 ( .I(n441), .ZN(n442) );
  INVD0 U385 ( .I(n444), .ZN(n441) );
  INVD0 U386 ( .I(n443), .ZN(n444) );
  CKNXD16 U387 ( .I(n445), .ZN(n443) );
  BUFFD0 U388 ( .I(n136), .Z(n445) );
  CKBXD0 U389 ( .I(OldWriteAr[2]), .Z(n446) );
  INVD0 U390 ( .I(n458), .ZN(n459) );
  CKND12 U391 ( .CLK(n447), .CN(n458) );
  BUFFD0 U392 ( .I(n133), .Z(n447) );
  INVD0 U393 ( .I(n561), .ZN(n562) );
  CKNXD16 U394 ( .I(n448), .ZN(n449) );
  CKNXD0 U395 ( .I(n451), .ZN(n448) );
  CKNXD16 U396 ( .I(n450), .ZN(n451) );
  INVD0 U397 ( .I(n453), .ZN(n450) );
  CKNXD16 U398 ( .I(n452), .ZN(n453) );
  CKNXD0 U399 ( .I(n455), .ZN(n452) );
  CKNXD16 U400 ( .I(n454), .ZN(n455) );
  CKNXD0 U401 ( .I(n457), .ZN(n454) );
  CKNXD16 U402 ( .I(n456), .ZN(n457) );
  CKNXD0 U403 ( .I(n459), .ZN(n456) );
  AO22D4 U404 ( .A1(WriteAddr[3]), .A2(n16), .B1(n17), .B2(n562), .Z(n133) );
  CKBXD0 U405 ( .I(OldWriteAr[3]), .Z(n460) );
  INVD1 U406 ( .I(n461), .ZN(n462) );
  INVD0 U407 ( .I(n463), .ZN(n464) );
  CKBXD0 U408 ( .I(n474), .Z(n465) );
  CKBXD0 U409 ( .I(n471), .Z(n472) );
  INVD0 U410 ( .I(n466), .ZN(n467) );
  CKNXD16 U411 ( .I(n465), .ZN(n466) );
  INVD0 U412 ( .I(n468), .ZN(n469) );
  CKNXD16 U413 ( .I(n467), .ZN(n468) );
  INVD0 U414 ( .I(n473), .ZN(n474) );
  INVD0 U415 ( .I(n149), .ZN(n470) );
  CKNXD16 U416 ( .I(n470), .ZN(n471) );
  CKNXD16 U417 ( .I(n472), .ZN(n473) );
  CKNXD0 U418 ( .I(n478), .ZN(n475) );
  CKNXD16 U419 ( .I(n477), .ZN(n478) );
  INVD0 U420 ( .I(n130), .ZN(n477) );
  BUFFD0 U421 ( .I(n481), .Z(n485) );
  INVD0 U422 ( .I(OldReadAr[2]), .ZN(n480) );
  CKNXD16 U423 ( .I(n480), .ZN(n481) );
  INVD0 U424 ( .I(n479), .ZN(n482) );
  INVD0 U425 ( .I(n483), .ZN(n484) );
  CKNXD16 U426 ( .I(n487), .ZN(n483) );
  INVD0 U427 ( .I(n486), .ZN(n487) );
  CKNXD16 U428 ( .I(n485), .ZN(n486) );
  CKNXD0 U429 ( .I(n491), .ZN(n488) );
  CKNXD16 U430 ( .I(n490), .ZN(n491) );
  INVD0 U431 ( .I(n128), .ZN(n490) );
  BUFFD0 U432 ( .I(n494), .Z(n498) );
  INVD0 U433 ( .I(OldReadAr[3]), .ZN(n493) );
  CKNXD16 U434 ( .I(n493), .ZN(n494) );
  INVD0 U435 ( .I(n492), .ZN(n495) );
  INVD0 U436 ( .I(n496), .ZN(n497) );
  CKNXD16 U437 ( .I(n500), .ZN(n496) );
  INVD0 U438 ( .I(n499), .ZN(n500) );
  CKNXD16 U439 ( .I(n498), .ZN(n499) );
  BUFFD0 U440 ( .I(n503), .Z(n501) );
  BUFFD0 U441 ( .I(n126), .Z(n502) );
  BUFFD0 U442 ( .I(n507), .Z(n503) );
  CKNXD16 U443 ( .I(n504), .ZN(n505) );
  INVD0 U444 ( .I(n502), .ZN(n504) );
  CKNXD16 U445 ( .I(n506), .ZN(n507) );
  INVD0 U446 ( .I(n198), .ZN(n506) );
  CKNXD16 U447 ( .I(n508), .ZN(n509) );
  INVD0 U448 ( .I(n505), .ZN(n508) );
  CKNXD16 U449 ( .I(n510), .ZN(n511) );
  INVD0 U450 ( .I(n513), .ZN(n510) );
  CKNXD16 U451 ( .I(n512), .ZN(n513) );
  CKNXD0 U452 ( .I(n509), .ZN(n512) );
  BUFFD0 U453 ( .I(n515), .Z(n514) );
  BUFFD0 U454 ( .I(n520), .Z(n515) );
  BUFFD0 U455 ( .I(n123), .Z(n516) );
  CKNXD16 U456 ( .I(n517), .ZN(n518) );
  INVD0 U457 ( .I(n522), .ZN(n517) );
  CKNXD16 U458 ( .I(n519), .ZN(n520) );
  INVD0 U459 ( .I(n525), .ZN(n519) );
  CKNXD16 U460 ( .I(n521), .ZN(n522) );
  INVD0 U461 ( .I(n527), .ZN(n521) );
  CKNXD16 U462 ( .I(n523), .ZN(n524) );
  CKNXD0 U463 ( .I(n516), .ZN(n523) );
  CKNXD16 U464 ( .I(n197), .ZN(n525) );
  CKNXD16 U465 ( .I(n526), .ZN(n527) );
  INVD0 U466 ( .I(n524), .ZN(n526) );
  BUFFD0 U467 ( .I(n530), .Z(n528) );
  BUFFD0 U468 ( .I(n142), .Z(n529) );
  BUFFD0 U469 ( .I(n534), .Z(n530) );
  CKNXD16 U470 ( .I(n531), .ZN(n532) );
  INVD0 U471 ( .I(n529), .ZN(n531) );
  CKNXD16 U472 ( .I(n533), .ZN(n534) );
  INVD0 U473 ( .I(n196), .ZN(n533) );
  CKNXD16 U474 ( .I(n535), .ZN(n536) );
  INVD0 U475 ( .I(n532), .ZN(n535) );
  CKNXD16 U476 ( .I(n537), .ZN(n538) );
  INVD0 U477 ( .I(n540), .ZN(n537) );
  CKNXD16 U478 ( .I(n539), .ZN(n540) );
  CKNXD0 U479 ( .I(n536), .ZN(n539) );
  INVD1 U480 ( .I(n148), .ZN(n541) );
  INVD0 U481 ( .I(n545), .ZN(n546) );
  CKNXD16 U482 ( .I(n194), .ZN(n545) );
  CKNXD16 U483 ( .I(n397), .ZN(n101) );
  ND3D0 U484 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n23) );
  CKNXD0 U485 ( .I(n549), .ZN(n550) );
  CKNXD16 U486 ( .I(n563), .ZN(n549) );
  CKNXD16 U487 ( .I(n412), .ZN(n18) );
  INVD0 U488 ( .I(n551), .ZN(n552) );
  CKNXD16 U489 ( .I(n554), .ZN(n551) );
  CKBXD0 U490 ( .I(n556), .Z(n565) );
  INVD0 U491 ( .I(n553), .ZN(n554) );
  CKNXD16 U492 ( .I(n558), .ZN(n553) );
  CKNXD16 U493 ( .I(n555), .ZN(n556) );
  INVD0 U494 ( .I(n155), .ZN(n555) );
  INVD0 U495 ( .I(n557), .ZN(n558) );
  CKNXD16 U496 ( .I(n565), .ZN(n557) );
  CKNXD0 U497 ( .I(n559), .ZN(n560) );
  CKNXD16 U498 ( .I(n446), .ZN(n559) );
  CKNXD16 U499 ( .I(n460), .ZN(n561) );
  BUFFD0 U500 ( .I(n18), .Z(n563) );
  CKNXD16 U501 ( .I(n428), .ZN(n20) );
  CKBXD0 U502 ( .I(n385), .Z(n566) );
  CKNXD16 U503 ( .I(n568), .ZN(n569) );
  CKNXD0 U504 ( .I(n571), .ZN(n568) );
  CKNXD16 U505 ( .I(n570), .ZN(n571) );
  CKNXD0 U506 ( .I(n573), .ZN(n570) );
  CKNXD16 U507 ( .I(n572), .ZN(n573) );
  CKNXD0 U508 ( .I(n575), .ZN(n572) );
  CKNXD16 U509 ( .I(n574), .ZN(n575) );
  CKNXD0 U510 ( .I(n577), .ZN(n574) );
  CKNXD16 U511 ( .I(n576), .ZN(n577) );
  CKNXD0 U512 ( .I(n579), .ZN(n576) );
  CKNXD16 U513 ( .I(n578), .ZN(n579) );
  INVD0 U514 ( .I(n567), .ZN(n578) );
  CKNXD16 U515 ( .I(n580), .ZN(n581) );
  CKNXD0 U516 ( .I(n583), .ZN(n580) );
  CKNXD16 U517 ( .I(n582), .ZN(n583) );
  CKNXD0 U518 ( .I(n585), .ZN(n582) );
  CKNXD16 U519 ( .I(n584), .ZN(n585) );
  CKNXD0 U520 ( .I(n587), .ZN(n584) );
  CKNXD16 U521 ( .I(n586), .ZN(n587) );
  CKNXD0 U522 ( .I(n589), .ZN(n586) );
  CKNXD16 U523 ( .I(n588), .ZN(n589) );
  CKNXD0 U524 ( .I(n591), .ZN(n588) );
  CKNXD16 U525 ( .I(n590), .ZN(n591) );
  CKND8 U526 ( .CLK(n592), .CN(n593) );
  INVD0 U527 ( .I(n595), .ZN(n592) );
  CKNXD16 U528 ( .I(n594), .ZN(n595) );
  INVD0 U529 ( .I(n597), .ZN(n594) );
  INVD0 U530 ( .I(N51), .ZN(n596) );
  INR2D0 U531 ( .A1(N46), .B1(n99), .ZN(N51) );
  CKBD0 U532 ( .CLK(n600), .C(n598) );
  INVD0 U533 ( .I(n602), .ZN(n599) );
  INVD0 U534 ( .I(n604), .ZN(n601) );
  INVD0 U535 ( .I(n605), .ZN(n606) );
  CKNXD16 U536 ( .I(n607), .ZN(n605) );
  INVD0 U537 ( .I(n606), .ZN(n603) );
  INVD0 U538 ( .I(n192), .ZN(n607) );
  CKNXD16 U539 ( .I(n601), .ZN(n602) );
  CKNXD16 U540 ( .I(n603), .ZN(n604) );
  CKBD0 U541 ( .CLK(n165), .C(ReadAddr[4]) );
  CKNXD16 U542 ( .I(n608), .ZN(n609) );
  CKNXD0 U543 ( .I(n611), .ZN(n608) );
  CKNXD16 U544 ( .I(n610), .ZN(n611) );
  CKNXD0 U545 ( .I(n613), .ZN(n610) );
  CKNXD16 U546 ( .I(n612), .ZN(n613) );
  CKNXD0 U547 ( .I(n615), .ZN(n612) );
  CKNXD16 U548 ( .I(n614), .ZN(n615) );
  CKNXD0 U549 ( .I(n617), .ZN(n614) );
  CKNXD16 U550 ( .I(n616), .ZN(n617) );
  CKNXD0 U551 ( .I(n619), .ZN(n616) );
  CKNXD16 U552 ( .I(n618), .ZN(n619) );
  INVD0 U553 ( .I(n167), .ZN(n618) );
  CKNXD16 U554 ( .I(n620), .ZN(n621) );
  INVD0 U555 ( .I(n624), .ZN(n620) );
  INVD0 U556 ( .I(n73), .ZN(n622) );
  INVD0 U557 ( .I(N47), .ZN(n73) );
  CKNXD16 U558 ( .I(n623), .ZN(n624) );
  INVD0 U559 ( .I(n170), .ZN(n623) );
  BUFFD0 U560 ( .I(ReadAddr[3]), .Z(n625) );
  CKBD0 U561 ( .CLK(n829), .C(ReadAddr[2]) );
  INVD12 U562 ( .I(n626), .ZN(n627) );
  INVD0 U563 ( .I(n629), .ZN(n626) );
  CKNXD16 U564 ( .I(n628), .ZN(n629) );
  CKNXD0 U565 ( .I(n631), .ZN(n628) );
  CKNXD16 U566 ( .I(n630), .ZN(n631) );
  CKNXD0 U567 ( .I(n633), .ZN(n630) );
  CKNXD16 U568 ( .I(n632), .ZN(n633) );
  CKNXD0 U569 ( .I(n635), .ZN(n632) );
  CKNXD16 U570 ( .I(n634), .ZN(n635) );
  CKNXD0 U571 ( .I(n637), .ZN(n634) );
  CKNXD16 U572 ( .I(n636), .ZN(n637) );
  CKNXD0 U573 ( .I(n638), .ZN(n636) );
  CKNXD16 U574 ( .I(n187), .ZN(n638) );
  CKNXD16 U575 ( .I(n643), .ZN(n644) );
  CKBD16 U576 ( .CLK(n689), .C(n688) );
  CKNXD16 U577 ( .I(n646), .ZN(n647) );
  INVD0 U578 ( .I(n642), .ZN(n646) );
  INVD0 U579 ( .I(N330), .ZN(n648) );
  BUFFD0 U580 ( .I(n652), .Z(n651) );
  BUFFD0 U581 ( .I(N78), .Z(n652) );
  BUFFD0 U582 ( .I(n654), .Z(n653) );
  BUFFD0 U583 ( .I(n655), .Z(n654) );
  BUFFD0 U584 ( .I(n656), .Z(n655) );
  BUFFD0 U585 ( .I(n658), .Z(n656) );
  BUFFD0 U586 ( .I(n675), .Z(n657) );
  BUFFD0 U587 ( .I(n659), .Z(n658) );
  BUFFD0 U588 ( .I(n660), .Z(n659) );
  BUFFD0 U589 ( .I(n661), .Z(n660) );
  BUFFD0 U590 ( .I(n662), .Z(n661) );
  BUFFD0 U591 ( .I(n663), .Z(n662) );
  BUFFD0 U592 ( .I(n664), .Z(n663) );
  BUFFD0 U593 ( .I(n665), .Z(n664) );
  BUFFD0 U594 ( .I(n666), .Z(n665) );
  BUFFD0 U595 ( .I(n667), .Z(n666) );
  BUFFD0 U596 ( .I(n668), .Z(n667) );
  BUFFD0 U597 ( .I(n669), .Z(n668) );
  BUFFD0 U598 ( .I(n670), .Z(n669) );
  BUFFD0 U599 ( .I(n671), .Z(n670) );
  BUFFD0 U600 ( .I(n672), .Z(n671) );
  INVD0 U601 ( .I(n673), .ZN(n674) );
  CKNXD16 U602 ( .I(n12), .ZN(n673) );
  BUFFD0 U603 ( .I(CurState[1]), .Z(n675) );
  ND3D0 U604 ( .A1(n657), .A2(CurState[0]), .A3(CurState[2]), .ZN(n12) );
  CKNXD16 U605 ( .I(n676), .ZN(n677) );
  INVD0 U606 ( .I(n680), .ZN(n676) );
  INVD0 U607 ( .I(n72), .ZN(n678) );
  INVD0 U608 ( .I(N45), .ZN(n72) );
  CKNXD16 U609 ( .I(n679), .ZN(n680) );
  INVD0 U610 ( .I(n180), .ZN(n679) );
  BUFFD0 U611 ( .I(ReadAddr[1]), .Z(n681) );
  CKBD0 U612 ( .CLK(n681), .C(n682) );
  INVD0 U613 ( .I(n823), .ZN(n683) );
  CKNXD0 U614 ( .I(N44), .ZN(n823) );
  CKNXD16 U615 ( .I(n684), .ZN(n685) );
  INVD0 U616 ( .I(ReadAddr[0]), .ZN(n684) );
  BUFFD0 U617 ( .I(n691), .Z(n690) );
  BUFFD0 U618 ( .I(n692), .Z(n691) );
  BUFFD0 U619 ( .I(n693), .Z(n692) );
  BUFFD0 U620 ( .I(n694), .Z(n693) );
  BUFFD0 U621 ( .I(n695), .Z(n694) );
  BUFFD0 U622 ( .I(n696), .Z(n695) );
  BUFFD0 U623 ( .I(n697), .Z(n696) );
  BUFFD0 U624 ( .I(n698), .Z(n697) );
  BUFFD0 U625 ( .I(n699), .Z(n698) );
  BUFFD0 U626 ( .I(n700), .Z(n699) );
  BUFFD0 U627 ( .I(n701), .Z(n700) );
  BUFFD0 U628 ( .I(n702), .Z(n701) );
  BUFFD0 U629 ( .I(n703), .Z(n702) );
  BUFFD0 U630 ( .I(n704), .Z(n703) );
  BUFFD0 U631 ( .I(n705), .Z(n704) );
  BUFFD0 U632 ( .I(n706), .Z(n705) );
  BUFFD0 U633 ( .I(n707), .Z(n706) );
  BUFFD0 U634 ( .I(n708), .Z(n707) );
  BUFFD0 U635 ( .I(n709), .Z(n708) );
  BUFFD0 U636 ( .I(n711), .Z(n709) );
  INVD0 U637 ( .I(n710), .ZN(n711) );
  CKNXD16 U638 ( .I(n6), .ZN(n710) );
  ND2D0 U639 ( .A1(n690), .A2(n99), .ZN(N53) );
  ND3D0 U640 ( .A1(n29), .A2(n96), .A3(n55), .ZN(n6) );
  BUFFD0 U641 ( .I(n831), .Z(n712) );
  BUFFD0 U642 ( .I(n712), .Z(n713) );
  BUFFD0 U643 ( .I(n713), .Z(n714) );
  BUFFD0 U644 ( .I(n714), .Z(n715) );
  BUFFD0 U645 ( .I(n715), .Z(n716) );
  BUFFD0 U646 ( .I(n716), .Z(n717) );
  BUFFD0 U647 ( .I(n717), .Z(n718) );
  BUFFD0 U648 ( .I(n718), .Z(n719) );
  BUFFD0 U649 ( .I(n719), .Z(n720) );
  BUFFD0 U650 ( .I(n720), .Z(n721) );
  BUFFD0 U651 ( .I(n721), .Z(n722) );
  BUFFD0 U652 ( .I(n722), .Z(n723) );
  BUFFD0 U653 ( .I(n723), .Z(n724) );
  BUFFD0 U654 ( .I(n724), .Z(n725) );
  BUFFD0 U655 ( .I(n725), .Z(n726) );
  BUFFD0 U656 ( .I(n726), .Z(n727) );
  BUFFD0 U657 ( .I(n727), .Z(n728) );
  BUFFD0 U658 ( .I(n728), .Z(n729) );
  BUFFD0 U659 ( .I(n729), .Z(n730) );
  BUFFD0 U660 ( .I(n730), .Z(n731) );
  BUFFD0 U661 ( .I(n731), .Z(n732) );
  BUFFD0 U662 ( .I(n732), .Z(n733) );
  BUFFD0 U663 ( .I(n733), .Z(n734) );
  BUFFD0 U664 ( .I(n734), .Z(n735) );
  BUFFD0 U665 ( .I(n735), .Z(n736) );
  BUFFD0 U666 ( .I(n736), .Z(n737) );
  BUFFD0 U667 ( .I(n737), .Z(n738) );
  BUFFD0 U668 ( .I(n738), .Z(n739) );
  BUFFD0 U669 ( .I(n739), .Z(n740) );
  BUFFD0 U670 ( .I(n740), .Z(n741) );
  BUFFD0 U671 ( .I(n741), .Z(n742) );
  BUFFD0 U672 ( .I(n742), .Z(n743) );
  BUFFD0 U673 ( .I(n743), .Z(n744) );
  BUFFD0 U674 ( .I(n744), .Z(n745) );
  BUFFD0 U675 ( .I(n745), .Z(n746) );
  BUFFD0 U676 ( .I(n746), .Z(n747) );
  BUFFD0 U677 ( .I(n747), .Z(n748) );
  BUFFD0 U678 ( .I(n748), .Z(n749) );
  BUFFD0 U679 ( .I(n749), .Z(n750) );
  BUFFD0 U680 ( .I(n750), .Z(n751) );
  BUFFD0 U681 ( .I(n751), .Z(n752) );
  BUFFD0 U682 ( .I(n752), .Z(n753) );
  BUFFD0 U683 ( .I(n753), .Z(n754) );
  BUFFD0 U684 ( .I(n754), .Z(n755) );
  BUFFD0 U685 ( .I(n755), .Z(n756) );
  BUFFD0 U686 ( .I(n756), .Z(n757) );
  BUFFD0 U687 ( .I(n757), .Z(n758) );
  BUFFD0 U688 ( .I(n758), .Z(n759) );
  BUFFD0 U689 ( .I(n759), .Z(n760) );
  BUFFD0 U690 ( .I(n760), .Z(n761) );
  BUFFD0 U691 ( .I(n761), .Z(n762) );
  BUFFD0 U692 ( .I(n762), .Z(n763) );
  BUFFD0 U693 ( .I(n763), .Z(n764) );
  BUFFD0 U694 ( .I(n764), .Z(n765) );
  BUFFD0 U695 ( .I(n765), .Z(n766) );
  BUFFD0 U696 ( .I(n766), .Z(n767) );
  BUFFD0 U697 ( .I(n767), .Z(n768) );
  BUFFD0 U698 ( .I(n768), .Z(n769) );
  BUFFD0 U699 ( .I(n769), .Z(n770) );
  BUFFD0 U700 ( .I(n770), .Z(n771) );
  BUFFD0 U701 ( .I(n771), .Z(n772) );
  BUFFD0 U702 ( .I(n772), .Z(n773) );
  BUFFD0 U703 ( .I(n773), .Z(n774) );
  BUFFD0 U704 ( .I(n774), .Z(n775) );
  BUFFD0 U705 ( .I(n775), .Z(n776) );
  BUFFD0 U706 ( .I(n776), .Z(n777) );
  BUFFD0 U707 ( .I(n777), .Z(n778) );
  BUFFD0 U708 ( .I(n778), .Z(n779) );
  BUFFD0 U709 ( .I(n779), .Z(n780) );
  BUFFD0 U710 ( .I(n780), .Z(n781) );
  BUFFD0 U711 ( .I(n781), .Z(n782) );
  BUFFD0 U712 ( .I(n782), .Z(n783) );
  BUFFD0 U713 ( .I(n783), .Z(n784) );
  BUFFD0 U714 ( .I(n784), .Z(n785) );
  BUFFD0 U715 ( .I(n785), .Z(n786) );
  BUFFD0 U716 ( .I(n786), .Z(n787) );
  BUFFD0 U717 ( .I(n787), .Z(n788) );
  BUFFD0 U718 ( .I(n788), .Z(n789) );
  BUFFD0 U719 ( .I(n789), .Z(n790) );
  BUFFD0 U720 ( .I(n790), .Z(n791) );
  BUFFD0 U721 ( .I(n791), .Z(n792) );
  BUFFD0 U722 ( .I(n792), .Z(n793) );
  BUFFD0 U723 ( .I(n793), .Z(n794) );
  BUFFD0 U724 ( .I(n794), .Z(n795) );
  BUFFD0 U725 ( .I(n795), .Z(n796) );
  CKBD0 U726 ( .CLK(n796), .C(ReadCmd) );
  CKND2D0 U727 ( .A1(ClkR), .A2(ClkW), .ZN(StateClockRaw) );
  OAI31D0 U728 ( .A1(n12), .A2(Reset), .A3(ReadReq), .B(n203), .ZN(n132) );
  CKND2D0 U729 ( .A1(n143), .A2(n205), .ZN(n798) );
  OA31D0 U730 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(EmptyFIFO), 
        .Z(n799) );
  INVD1 U731 ( .I(n799), .ZN(n800) );
  OAI31D0 U732 ( .A1(n711), .A2(WriteReq), .A3(Reset), .B(n800), .ZN(n127) );
  INVD1 U733 ( .I(n9), .ZN(n8) );
  INVD1 U734 ( .I(n6), .ZN(n15) );
  ND3D1 U735 ( .A1(n100), .A2(n542), .A3(ReadReq), .ZN(n9) );
  INVD1 U736 ( .I(ReadReq), .ZN(n827) );
  INVD1 U737 ( .I(Reset), .ZN(n820) );
  NR3D0 U738 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n53) );
  ND4D1 U739 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(n30) );
  XOR2D1 U740 ( .A1(n625), .A2(n74), .Z(n62) );
  NR3D0 U741 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n65) );
  XNR2D1 U742 ( .A1(ReadAddr[4]), .A2(N72), .ZN(n64) );
  XNR2D1 U743 ( .A1(N177), .A2(n81), .ZN(n49) );
  XOR2D1 U744 ( .A1(WriteAddr[2]), .A2(N46), .Z(n54) );
  ND3D1 U745 ( .A1(n86), .A2(n87), .A3(n88), .ZN(n31) );
  XOR2D1 U746 ( .A1(n19), .A2(n825), .Z(n87) );
  XOR2D1 U747 ( .A1(N333), .A2(n826), .Z(n86) );
  NR3D0 U748 ( .A1(n89), .A2(n90), .A3(n91), .ZN(n88) );
  IIND4D1 U749 ( .A1(n54), .A2(n56), .B1(n51), .B2(n52), .ZN(n63) );
  XOR2D1 U750 ( .A1(ReadAddr[1]), .A2(N69), .Z(n66) );
  XOR2D1 U751 ( .A1(ReadAddr[2]), .A2(N70), .Z(n68) );
  INVD1 U752 ( .I(N71), .ZN(n74) );
  ND3D1 U753 ( .A1(n653), .A2(n690), .A3(n34), .ZN(N78) );
  INVD1 U754 ( .I(n100), .ZN(n98) );
  ND2D1 U755 ( .A1(n35), .A2(n230), .ZN(n100) );
  ND2D1 U756 ( .A1(n35), .A2(n6), .ZN(n22) );
  INVD1 U757 ( .I(n653), .ZN(n28) );
  OAI22D0 U758 ( .A1(n8), .A2(n390), .B1(n822), .B2(n9), .ZN(n144) );
  INVD1 U759 ( .I(n17), .ZN(n16) );
  INVD1 U760 ( .I(n24), .ZN(n25) );
  XOR2D1 U761 ( .A1(ReadAddr[1]), .A2(n19), .Z(n78) );
  NR2D1 U762 ( .A1(n801), .A2(n802), .ZN(n76) );
  XNR2D1 U763 ( .A1(n625), .A2(n81), .ZN(n801) );
  XOR2D1 U764 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .Z(n802) );
  INVD1 U765 ( .I(n34), .ZN(n109) );
  XOR2D1 U766 ( .A1(ReadAddr[0]), .A2(n548), .Z(n103) );
  XOR2D1 U767 ( .A1(ReadAddr[1]), .A2(n422), .Z(n104) );
  NR3D0 U768 ( .A1(n106), .A2(n107), .A3(n108), .ZN(n105) );
  XOR2D1 U769 ( .A1(N176), .A2(WriteAddr[2]), .Z(n50) );
  XOR2D1 U770 ( .A1(n825), .A2(n19), .Z(n45) );
  IND4D1 U771 ( .A1(n80), .B1(n75), .B2(n76), .B3(n78), .ZN(n82) );
  XOR2D1 U772 ( .A1(ReadAddr[0]), .A2(N68), .Z(n67) );
  INVD1 U773 ( .I(Reset), .ZN(n143) );
  AOI22D0 U774 ( .A1(n61), .A2(n55), .B1(CurState[0]), .B2(n30), .ZN(n60) );
  ND4D1 U775 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(n61) );
  AOI31D0 U776 ( .A1(n46), .A2(n45), .A3(n79), .B(n80), .ZN(n77) );
  NR3D0 U777 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n79) );
  AOI21D1 U778 ( .A1(CurState[0]), .A2(n27), .B(n28), .ZN(n26) );
  NR3D0 U779 ( .A1(n58), .A2(n15), .A3(n59), .ZN(n57) );
  AOI21D1 U780 ( .A1(n31), .A2(n82), .B(n83), .ZN(n58) );
  NR3D0 U781 ( .A1(n29), .A2(CurState[2]), .A3(n60), .ZN(n59) );
  OAI221D0 U782 ( .A1(CurState[2]), .A2(n43), .B1(CurState[0]), .B2(n44), .C(
        n24), .ZN(n42) );
  IINR4D0 U783 ( .A1(n45), .A2(n46), .B1(n47), .B2(n48), .ZN(n44) );
  AOI31D0 U784 ( .A1(n51), .A2(n52), .A3(n53), .B(n29), .ZN(n43) );
  XOR2D1 U785 ( .A1(WriteAddr[3]), .A2(n73), .Z(n51) );
  XOR2D1 U786 ( .A1(WriteAddr[4]), .A2(N48), .Z(n56) );
  XOR2D1 U787 ( .A1(ReadAddr[4]), .A2(N334), .Z(n90) );
  XNR2D1 U788 ( .A1(N178), .A2(WriteAddr[4]), .ZN(n46) );
  INVD1 U789 ( .I(n625), .ZN(n826) );
  BUFFD1 U790 ( .I(n830), .Z(WriteAddr[2]) );
  NR2D1 U791 ( .A1(n803), .A2(n804), .ZN(n52) );
  XNR2D1 U792 ( .A1(\add_388/carry[2] ), .A2(n72), .ZN(n803) );
  XNR2D1 U793 ( .A1(N330), .A2(n823), .ZN(n804) );
  OAI211D1 U794 ( .A1(CurState[1]), .A2(n55), .B(n35), .C(n93), .ZN(n24) );
  AOI21D1 U795 ( .A1(WriteReq), .A2(n15), .B(n94), .ZN(n93) );
  AOI21D1 U796 ( .A1(CurState[0]), .A2(n827), .B(n96), .ZN(n94) );
  ND2D1 U797 ( .A1(ReadCmd), .A2(n690), .ZN(n99) );
  INVD1 U798 ( .I(WriteReq), .ZN(n33) );
  INVD1 U799 ( .I(n22), .ZN(n32) );
  INVD1 U800 ( .I(\add_388/carry[2] ), .ZN(n19) );
  XOR2D1 U801 ( .A1(ReadAddr[0]), .A2(N330), .Z(n48) );
  XOR2D1 U802 ( .A1(N330), .A2(n212), .Z(n36) );
  XOR2D1 U803 ( .A1(\add_388/carry[2] ), .A2(n550), .Z(n37) );
  NR3D0 U804 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n38) );
  XNR2D1 U805 ( .A1(ReadAddr[4]), .A2(WriteAddr[4]), .ZN(n75) );
  ND3D1 U806 ( .A1(CurState[0]), .A2(n29), .A3(CurState[2]), .ZN(n83) );
  INVD1 U807 ( .I(WriteAddr[3]), .ZN(n81) );
  XOR2D1 U808 ( .A1(ReadAddr[2]), .A2(N332), .Z(n89) );
  XOR2D1 U809 ( .A1(ReadAddr[0]), .A2(N330), .Z(n80) );
  XOR2D1 U810 ( .A1(ReadAddr[0]), .A2(N330), .Z(n91) );
  XOR2D1 U811 ( .A1(n625), .A2(n497), .Z(n106) );
  XOR2D1 U812 ( .A1(WriteAddr[4]), .A2(n218), .Z(n41) );
  XOR2D1 U813 ( .A1(ReadAddr[2]), .A2(n484), .Z(n107) );
  CKXOR2D0 U814 ( .A1(ReadAddr[4]), .A2(\add_307/carry[4] ), .Z(N178) );
  AN2D0 U815 ( .A1(n625), .A2(\add_307/carry[3] ), .Z(\add_307/carry[4] ) );
  CKXOR2D0 U816 ( .A1(\add_307/carry[3] ), .A2(n625), .Z(N177) );
  AN2D0 U817 ( .A1(ReadAddr[2]), .A2(ReadAddr[1]), .Z(\add_307/carry[3] ) );
  CKXOR2D0 U818 ( .A1(ReadAddr[1]), .A2(ReadAddr[2]), .Z(N176) );
  CKXOR2D0 U819 ( .A1(WriteAddr[4]), .A2(\add_388/carry[4] ), .Z(N334) );
  AN2D0 U820 ( .A1(WriteAddr[3]), .A2(\add_388/carry[3] ), .Z(
        \add_388/carry[4] ) );
  CKXOR2D0 U821 ( .A1(\add_388/carry[3] ), .A2(WriteAddr[3]), .Z(N333) );
  AN2D0 U822 ( .A1(WriteAddr[2]), .A2(\add_388/carry[2] ), .Z(
        \add_388/carry[3] ) );
  CKXOR2D0 U823 ( .A1(\add_388/carry[2] ), .A2(WriteAddr[2]), .Z(N332) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, ClockR, ClockW, Dreadyr,
         \Storage[31][32] , \Storage[31][31] , \Storage[31][30] ,
         \Storage[31][29] , \Storage[31][28] , \Storage[31][27] ,
         \Storage[31][26] , \Storage[31][25] , \Storage[31][24] ,
         \Storage[31][23] , \Storage[31][22] , \Storage[31][21] ,
         \Storage[31][20] , \Storage[31][19] , \Storage[31][18] ,
         \Storage[31][17] , \Storage[31][16] , \Storage[31][15] ,
         \Storage[31][14] , \Storage[31][13] , \Storage[31][12] ,
         \Storage[31][11] , \Storage[31][10] , \Storage[31][9] ,
         \Storage[31][8] , \Storage[31][7] , \Storage[31][6] ,
         \Storage[31][5] , \Storage[31][4] , \Storage[31][3] ,
         \Storage[31][2] , \Storage[31][1] , \Storage[31][0] ,
         \Storage[30][32] , \Storage[30][31] , \Storage[30][30] ,
         \Storage[30][29] , \Storage[30][28] , \Storage[30][27] ,
         \Storage[30][26] , \Storage[30][25] , \Storage[30][24] ,
         \Storage[30][23] , \Storage[30][22] , \Storage[30][21] ,
         \Storage[30][20] , \Storage[30][19] , \Storage[30][18] ,
         \Storage[30][17] , \Storage[30][16] , \Storage[30][15] ,
         \Storage[30][14] , \Storage[30][13] , \Storage[30][12] ,
         \Storage[30][11] , \Storage[30][10] , \Storage[30][9] ,
         \Storage[30][8] , \Storage[30][7] , \Storage[30][6] ,
         \Storage[30][5] , \Storage[30][4] , \Storage[30][3] ,
         \Storage[30][2] , \Storage[30][1] , \Storage[30][0] ,
         \Storage[29][32] , \Storage[29][31] , \Storage[29][30] ,
         \Storage[29][29] , \Storage[29][28] , \Storage[29][27] ,
         \Storage[29][26] , \Storage[29][25] , \Storage[29][24] ,
         \Storage[29][23] , \Storage[29][22] , \Storage[29][21] ,
         \Storage[29][20] , \Storage[29][19] , \Storage[29][18] ,
         \Storage[29][17] , \Storage[29][16] , \Storage[29][15] ,
         \Storage[29][14] , \Storage[29][13] , \Storage[29][12] ,
         \Storage[29][11] , \Storage[29][10] , \Storage[29][9] ,
         \Storage[29][8] , \Storage[29][7] , \Storage[29][6] ,
         \Storage[29][5] , \Storage[29][4] , \Storage[29][3] ,
         \Storage[29][2] , \Storage[29][1] , \Storage[29][0] ,
         \Storage[28][32] , \Storage[28][31] , \Storage[28][30] ,
         \Storage[28][29] , \Storage[28][28] , \Storage[28][27] ,
         \Storage[28][26] , \Storage[28][25] , \Storage[28][24] ,
         \Storage[28][23] , \Storage[28][22] , \Storage[28][21] ,
         \Storage[28][20] , \Storage[28][19] , \Storage[28][18] ,
         \Storage[28][17] , \Storage[28][16] , \Storage[28][15] ,
         \Storage[28][14] , \Storage[28][13] , \Storage[28][12] ,
         \Storage[28][11] , \Storage[28][10] , \Storage[28][9] ,
         \Storage[28][8] , \Storage[28][7] , \Storage[28][6] ,
         \Storage[28][5] , \Storage[28][4] , \Storage[28][3] ,
         \Storage[28][2] , \Storage[28][1] , \Storage[28][0] ,
         \Storage[27][32] , \Storage[27][31] , \Storage[27][30] ,
         \Storage[27][29] , \Storage[27][28] , \Storage[27][27] ,
         \Storage[27][26] , \Storage[27][25] , \Storage[27][24] ,
         \Storage[27][23] , \Storage[27][22] , \Storage[27][21] ,
         \Storage[27][20] , \Storage[27][19] , \Storage[27][18] ,
         \Storage[27][17] , \Storage[27][16] , \Storage[27][15] ,
         \Storage[27][14] , \Storage[27][13] , \Storage[27][12] ,
         \Storage[27][11] , \Storage[27][10] , \Storage[27][9] ,
         \Storage[27][8] , \Storage[27][7] , \Storage[27][6] ,
         \Storage[27][5] , \Storage[27][4] , \Storage[27][3] ,
         \Storage[27][2] , \Storage[27][1] , \Storage[27][0] ,
         \Storage[26][32] , \Storage[26][31] , \Storage[26][30] ,
         \Storage[26][29] , \Storage[26][28] , \Storage[26][27] ,
         \Storage[26][26] , \Storage[26][25] , \Storage[26][24] ,
         \Storage[26][23] , \Storage[26][22] , \Storage[26][21] ,
         \Storage[26][20] , \Storage[26][19] , \Storage[26][18] ,
         \Storage[26][17] , \Storage[26][16] , \Storage[26][15] ,
         \Storage[26][14] , \Storage[26][13] , \Storage[26][12] ,
         \Storage[26][11] , \Storage[26][10] , \Storage[26][9] ,
         \Storage[26][8] , \Storage[26][7] , \Storage[26][6] ,
         \Storage[26][5] , \Storage[26][4] , \Storage[26][3] ,
         \Storage[26][2] , \Storage[26][1] , \Storage[26][0] ,
         \Storage[25][32] , \Storage[25][31] , \Storage[25][30] ,
         \Storage[25][29] , \Storage[25][28] , \Storage[25][27] ,
         \Storage[25][26] , \Storage[25][25] , \Storage[25][24] ,
         \Storage[25][23] , \Storage[25][22] , \Storage[25][21] ,
         \Storage[25][20] , \Storage[25][19] , \Storage[25][18] ,
         \Storage[25][17] , \Storage[25][16] , \Storage[25][15] ,
         \Storage[25][14] , \Storage[25][13] , \Storage[25][12] ,
         \Storage[25][11] , \Storage[25][10] , \Storage[25][9] ,
         \Storage[25][8] , \Storage[25][7] , \Storage[25][6] ,
         \Storage[25][5] , \Storage[25][4] , \Storage[25][3] ,
         \Storage[25][2] , \Storage[25][1] , \Storage[25][0] ,
         \Storage[24][32] , \Storage[24][31] , \Storage[24][30] ,
         \Storage[24][29] , \Storage[24][28] , \Storage[24][27] ,
         \Storage[24][26] , \Storage[24][25] , \Storage[24][24] ,
         \Storage[24][23] , \Storage[24][22] , \Storage[24][21] ,
         \Storage[24][20] , \Storage[24][19] , \Storage[24][18] ,
         \Storage[24][17] , \Storage[24][16] , \Storage[24][15] ,
         \Storage[24][14] , \Storage[24][13] , \Storage[24][12] ,
         \Storage[24][11] , \Storage[24][10] , \Storage[24][9] ,
         \Storage[24][8] , \Storage[24][7] , \Storage[24][6] ,
         \Storage[24][5] , \Storage[24][4] , \Storage[24][3] ,
         \Storage[24][2] , \Storage[24][1] , \Storage[24][0] ,
         \Storage[23][32] , \Storage[23][31] , \Storage[23][30] ,
         \Storage[23][29] , \Storage[23][28] , \Storage[23][27] ,
         \Storage[23][26] , \Storage[23][25] , \Storage[23][24] ,
         \Storage[23][23] , \Storage[23][22] , \Storage[23][21] ,
         \Storage[23][20] , \Storage[23][19] , \Storage[23][18] ,
         \Storage[23][17] , \Storage[23][16] , \Storage[23][15] ,
         \Storage[23][14] , \Storage[23][13] , \Storage[23][12] ,
         \Storage[23][11] , \Storage[23][10] , \Storage[23][9] ,
         \Storage[23][8] , \Storage[23][7] , \Storage[23][6] ,
         \Storage[23][5] , \Storage[23][4] , \Storage[23][3] ,
         \Storage[23][2] , \Storage[23][1] , \Storage[23][0] ,
         \Storage[22][32] , \Storage[22][31] , \Storage[22][30] ,
         \Storage[22][29] , \Storage[22][28] , \Storage[22][27] ,
         \Storage[22][26] , \Storage[22][25] , \Storage[22][24] ,
         \Storage[22][23] , \Storage[22][22] , \Storage[22][21] ,
         \Storage[22][20] , \Storage[22][19] , \Storage[22][18] ,
         \Storage[22][17] , \Storage[22][16] , \Storage[22][15] ,
         \Storage[22][14] , \Storage[22][13] , \Storage[22][12] ,
         \Storage[22][11] , \Storage[22][10] , \Storage[22][9] ,
         \Storage[22][8] , \Storage[22][7] , \Storage[22][6] ,
         \Storage[22][5] , \Storage[22][4] , \Storage[22][3] ,
         \Storage[22][2] , \Storage[22][1] , \Storage[22][0] ,
         \Storage[21][32] , \Storage[21][31] , \Storage[21][30] ,
         \Storage[21][29] , \Storage[21][28] , \Storage[21][27] ,
         \Storage[21][26] , \Storage[21][25] , \Storage[21][24] ,
         \Storage[21][23] , \Storage[21][22] , \Storage[21][21] ,
         \Storage[21][20] , \Storage[21][19] , \Storage[21][18] ,
         \Storage[21][17] , \Storage[21][16] , \Storage[21][15] ,
         \Storage[21][14] , \Storage[21][13] , \Storage[21][12] ,
         \Storage[21][11] , \Storage[21][10] , \Storage[21][9] ,
         \Storage[21][8] , \Storage[21][7] , \Storage[21][6] ,
         \Storage[21][5] , \Storage[21][4] , \Storage[21][3] ,
         \Storage[21][2] , \Storage[21][1] , \Storage[21][0] ,
         \Storage[20][32] , \Storage[20][31] , \Storage[20][30] ,
         \Storage[20][29] , \Storage[20][28] , \Storage[20][27] ,
         \Storage[20][26] , \Storage[20][25] , \Storage[20][24] ,
         \Storage[20][23] , \Storage[20][22] , \Storage[20][21] ,
         \Storage[20][20] , \Storage[20][19] , \Storage[20][18] ,
         \Storage[20][17] , \Storage[20][16] , \Storage[20][15] ,
         \Storage[20][14] , \Storage[20][13] , \Storage[20][12] ,
         \Storage[20][11] , \Storage[20][10] , \Storage[20][9] ,
         \Storage[20][8] , \Storage[20][7] , \Storage[20][6] ,
         \Storage[20][5] , \Storage[20][4] , \Storage[20][3] ,
         \Storage[20][2] , \Storage[20][1] , \Storage[20][0] ,
         \Storage[19][32] , \Storage[19][31] , \Storage[19][30] ,
         \Storage[19][29] , \Storage[19][28] , \Storage[19][27] ,
         \Storage[19][26] , \Storage[19][25] , \Storage[19][24] ,
         \Storage[19][23] , \Storage[19][22] , \Storage[19][21] ,
         \Storage[19][20] , \Storage[19][19] , \Storage[19][18] ,
         \Storage[19][17] , \Storage[19][16] , \Storage[19][15] ,
         \Storage[19][14] , \Storage[19][13] , \Storage[19][12] ,
         \Storage[19][11] , \Storage[19][10] , \Storage[19][9] ,
         \Storage[19][8] , \Storage[19][7] , \Storage[19][6] ,
         \Storage[19][5] , \Storage[19][4] , \Storage[19][3] ,
         \Storage[19][2] , \Storage[19][1] , \Storage[19][0] ,
         \Storage[18][32] , \Storage[18][31] , \Storage[18][30] ,
         \Storage[18][29] , \Storage[18][28] , \Storage[18][27] ,
         \Storage[18][26] , \Storage[18][25] , \Storage[18][24] ,
         \Storage[18][23] , \Storage[18][22] , \Storage[18][21] ,
         \Storage[18][20] , \Storage[18][19] , \Storage[18][18] ,
         \Storage[18][17] , \Storage[18][16] , \Storage[18][15] ,
         \Storage[18][14] , \Storage[18][13] , \Storage[18][12] ,
         \Storage[18][11] , \Storage[18][10] , \Storage[18][9] ,
         \Storage[18][8] , \Storage[18][7] , \Storage[18][6] ,
         \Storage[18][5] , \Storage[18][4] , \Storage[18][3] ,
         \Storage[18][2] , \Storage[18][1] , \Storage[18][0] ,
         \Storage[17][32] , \Storage[17][31] , \Storage[17][30] ,
         \Storage[17][29] , \Storage[17][28] , \Storage[17][27] ,
         \Storage[17][26] , \Storage[17][25] , \Storage[17][24] ,
         \Storage[17][23] , \Storage[17][22] , \Storage[17][21] ,
         \Storage[17][20] , \Storage[17][19] , \Storage[17][18] ,
         \Storage[17][17] , \Storage[17][16] , \Storage[17][15] ,
         \Storage[17][14] , \Storage[17][13] , \Storage[17][12] ,
         \Storage[17][11] , \Storage[17][10] , \Storage[17][9] ,
         \Storage[17][8] , \Storage[17][7] , \Storage[17][6] ,
         \Storage[17][5] , \Storage[17][4] , \Storage[17][3] ,
         \Storage[17][2] , \Storage[17][1] , \Storage[17][0] ,
         \Storage[16][32] , \Storage[16][31] , \Storage[16][30] ,
         \Storage[16][29] , \Storage[16][28] , \Storage[16][27] ,
         \Storage[16][26] , \Storage[16][25] , \Storage[16][24] ,
         \Storage[16][23] , \Storage[16][22] , \Storage[16][21] ,
         \Storage[16][20] , \Storage[16][19] , \Storage[16][18] ,
         \Storage[16][17] , \Storage[16][16] , \Storage[16][15] ,
         \Storage[16][14] , \Storage[16][13] , \Storage[16][12] ,
         \Storage[16][11] , \Storage[16][10] , \Storage[16][9] ,
         \Storage[16][8] , \Storage[16][7] , \Storage[16][6] ,
         \Storage[16][5] , \Storage[16][4] , \Storage[16][3] ,
         \Storage[16][2] , \Storage[16][1] , \Storage[16][0] ,
         \Storage[15][32] , \Storage[15][31] , \Storage[15][30] ,
         \Storage[15][29] , \Storage[15][28] , \Storage[15][27] ,
         \Storage[15][26] , \Storage[15][25] , \Storage[15][24] ,
         \Storage[15][23] , \Storage[15][22] , \Storage[15][21] ,
         \Storage[15][20] , \Storage[15][19] , \Storage[15][18] ,
         \Storage[15][17] , \Storage[15][16] , \Storage[15][15] ,
         \Storage[15][14] , \Storage[15][13] , \Storage[15][12] ,
         \Storage[15][11] , \Storage[15][10] , \Storage[15][9] ,
         \Storage[15][8] , \Storage[15][7] , \Storage[15][6] ,
         \Storage[15][5] , \Storage[15][4] , \Storage[15][3] ,
         \Storage[15][2] , \Storage[15][1] , \Storage[15][0] ,
         \Storage[14][32] , \Storage[14][31] , \Storage[14][30] ,
         \Storage[14][29] , \Storage[14][28] , \Storage[14][27] ,
         \Storage[14][26] , \Storage[14][25] , \Storage[14][24] ,
         \Storage[14][23] , \Storage[14][22] , \Storage[14][21] ,
         \Storage[14][20] , \Storage[14][19] , \Storage[14][18] ,
         \Storage[14][17] , \Storage[14][16] , \Storage[14][15] ,
         \Storage[14][14] , \Storage[14][13] , \Storage[14][12] ,
         \Storage[14][11] , \Storage[14][10] , \Storage[14][9] ,
         \Storage[14][8] , \Storage[14][7] , \Storage[14][6] ,
         \Storage[14][5] , \Storage[14][4] , \Storage[14][3] ,
         \Storage[14][2] , \Storage[14][1] , \Storage[14][0] ,
         \Storage[13][32] , \Storage[13][31] , \Storage[13][30] ,
         \Storage[13][29] , \Storage[13][28] , \Storage[13][27] ,
         \Storage[13][26] , \Storage[13][25] , \Storage[13][24] ,
         \Storage[13][23] , \Storage[13][22] , \Storage[13][21] ,
         \Storage[13][20] , \Storage[13][19] , \Storage[13][18] ,
         \Storage[13][17] , \Storage[13][16] , \Storage[13][15] ,
         \Storage[13][14] , \Storage[13][13] , \Storage[13][12] ,
         \Storage[13][11] , \Storage[13][10] , \Storage[13][9] ,
         \Storage[13][8] , \Storage[13][7] , \Storage[13][6] ,
         \Storage[13][5] , \Storage[13][4] , \Storage[13][3] ,
         \Storage[13][2] , \Storage[13][1] , \Storage[13][0] ,
         \Storage[12][32] , \Storage[12][31] , \Storage[12][30] ,
         \Storage[12][29] , \Storage[12][28] , \Storage[12][27] ,
         \Storage[12][26] , \Storage[12][25] , \Storage[12][24] ,
         \Storage[12][23] , \Storage[12][22] , \Storage[12][21] ,
         \Storage[12][20] , \Storage[12][19] , \Storage[12][18] ,
         \Storage[12][17] , \Storage[12][16] , \Storage[12][15] ,
         \Storage[12][14] , \Storage[12][13] , \Storage[12][12] ,
         \Storage[12][11] , \Storage[12][10] , \Storage[12][9] ,
         \Storage[12][8] , \Storage[12][7] , \Storage[12][6] ,
         \Storage[12][5] , \Storage[12][4] , \Storage[12][3] ,
         \Storage[12][2] , \Storage[12][1] , \Storage[12][0] ,
         \Storage[11][32] , \Storage[11][31] , \Storage[11][30] ,
         \Storage[11][29] , \Storage[11][28] , \Storage[11][27] ,
         \Storage[11][26] , \Storage[11][25] , \Storage[11][24] ,
         \Storage[11][23] , \Storage[11][22] , \Storage[11][21] ,
         \Storage[11][20] , \Storage[11][19] , \Storage[11][18] ,
         \Storage[11][17] , \Storage[11][16] , \Storage[11][15] ,
         \Storage[11][14] , \Storage[11][13] , \Storage[11][12] ,
         \Storage[11][11] , \Storage[11][10] , \Storage[11][9] ,
         \Storage[11][8] , \Storage[11][7] , \Storage[11][6] ,
         \Storage[11][5] , \Storage[11][4] , \Storage[11][3] ,
         \Storage[11][2] , \Storage[11][1] , \Storage[11][0] ,
         \Storage[10][32] , \Storage[10][31] , \Storage[10][30] ,
         \Storage[10][29] , \Storage[10][28] , \Storage[10][27] ,
         \Storage[10][26] , \Storage[10][25] , \Storage[10][24] ,
         \Storage[10][23] , \Storage[10][22] , \Storage[10][21] ,
         \Storage[10][20] , \Storage[10][19] , \Storage[10][18] ,
         \Storage[10][17] , \Storage[10][16] , \Storage[10][15] ,
         \Storage[10][14] , \Storage[10][13] , \Storage[10][12] ,
         \Storage[10][11] , \Storage[10][10] , \Storage[10][9] ,
         \Storage[10][8] , \Storage[10][7] , \Storage[10][6] ,
         \Storage[10][5] , \Storage[10][4] , \Storage[10][3] ,
         \Storage[10][2] , \Storage[10][1] , \Storage[10][0] ,
         \Storage[9][32] , \Storage[9][31] , \Storage[9][30] ,
         \Storage[9][29] , \Storage[9][28] , \Storage[9][27] ,
         \Storage[9][26] , \Storage[9][25] , \Storage[9][24] ,
         \Storage[9][23] , \Storage[9][22] , \Storage[9][21] ,
         \Storage[9][20] , \Storage[9][19] , \Storage[9][18] ,
         \Storage[9][17] , \Storage[9][16] , \Storage[9][15] ,
         \Storage[9][14] , \Storage[9][13] , \Storage[9][12] ,
         \Storage[9][11] , \Storage[9][10] , \Storage[9][9] , \Storage[9][8] ,
         \Storage[9][7] , \Storage[9][6] , \Storage[9][5] , \Storage[9][4] ,
         \Storage[9][3] , \Storage[9][2] , \Storage[9][1] , \Storage[9][0] ,
         \Storage[8][32] , \Storage[8][31] , \Storage[8][30] ,
         \Storage[8][29] , \Storage[8][28] , \Storage[8][27] ,
         \Storage[8][26] , \Storage[8][25] , \Storage[8][24] ,
         \Storage[8][23] , \Storage[8][22] , \Storage[8][21] ,
         \Storage[8][20] , \Storage[8][19] , \Storage[8][18] ,
         \Storage[8][17] , \Storage[8][16] , \Storage[8][15] ,
         \Storage[8][14] , \Storage[8][13] , \Storage[8][12] ,
         \Storage[8][11] , \Storage[8][10] , \Storage[8][9] , \Storage[8][8] ,
         \Storage[8][7] , \Storage[8][6] , \Storage[8][5] , \Storage[8][4] ,
         \Storage[8][3] , \Storage[8][2] , \Storage[8][1] , \Storage[8][0] ,
         \Storage[7][32] , \Storage[7][31] , \Storage[7][30] ,
         \Storage[7][29] , \Storage[7][28] , \Storage[7][27] ,
         \Storage[7][26] , \Storage[7][25] , \Storage[7][24] ,
         \Storage[7][23] , \Storage[7][22] , \Storage[7][21] ,
         \Storage[7][20] , \Storage[7][19] , \Storage[7][18] ,
         \Storage[7][17] , \Storage[7][16] , \Storage[7][15] ,
         \Storage[7][14] , \Storage[7][13] , \Storage[7][12] ,
         \Storage[7][11] , \Storage[7][10] , \Storage[7][9] , \Storage[7][8] ,
         \Storage[7][7] , \Storage[7][6] , \Storage[7][5] , \Storage[7][4] ,
         \Storage[7][3] , \Storage[7][2] , \Storage[7][1] , \Storage[7][0] ,
         \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N50, N67, N68, N71, N72, N73, N77, N78, N79, N81, N82, N83, N85, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n90, n92, n107, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n122, n123, n124,
         n126, n127, n128, n130, n131, n132, n134, n135, n136, n138, n139,
         n140, n142, n143, n144, n146, n147, n148, n150, n151, n152, n154,
         n155, n156, n158, n159, n160, n162, n163, n164, n166, n167, n168,
         n170, n171, n172, n174, n175, n176, n178, n179, n180, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n241, n243, n245, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  XNR4D1 U18 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n84) );
  XOR4D1 U19 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n83) );
  XOR4D1 U20 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n80) );
  XOR4D1 U21 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n77) );
  XNR4D1 U22 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n74) );
  XNR4D1 U28 ( .A1(n951), .A2(n885), .A3(n994), .A4(n986), .ZN(n91) );
  XOR4D1 U34 ( .A1(n453), .A2(n389), .A3(n494), .A4(n488), .Z(n96) );
  XNR4D1 U35 ( .A1(n699), .A2(n634), .A3(n740), .A4(n734), .ZN(n93) );
  XNR4D1 U36 ( .A1(n1354), .A2(n1251), .A3(n1397), .A4(n1361), .ZN(n87) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(DataI[9]), .E(n239), .CP(n2206), .CDN(
        n2171), .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(DataI[8]), .E(n239), .CP(n2206), .CDN(
        n2160), .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(DataI[3]), .E(n239), .CP(n2207), .CDN(
        n2148), .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(DataI[9]), .E(n238), .CP(n2213), .CDN(
        n2176), .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(DataI[8]), .E(n238), .CP(n2213), .CDN(
        n2156), .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(DataI[3]), .E(n238), .CP(n2214), .CDN(
        n2157), .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(DataI[9]), .E(n237), .CP(n2193), .CDN(
        n2160), .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n237), .CP(n2193), .CDN(
        n2161), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(n237), .CP(n2194), .CDN(
        n2162), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(n236), .CP(n2196), .CDN(
        n2153), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(n236), .CP(n2197), .CDN(
        n2155), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(n236), .CP(n2197), .CDN(
        n2156), .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(DataI[9]), .E(n235), .CP(n2200), .CDN(
        n2148), .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(DataI[8]), .E(n235), .CP(n2200), .CDN(
        n2180), .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(DataI[3]), .E(n235), .CP(n2200), .CDN(
        n2148), .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(n234), .CP(n2203), .CDN(
        n2178), .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(n234), .CP(n2203), .CDN(
        n2155), .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(DataI[3]), .E(n234), .CP(n2204), .CDN(
        n2157), .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(DataI[9]), .E(n233), .CP(n2210), .CDN(
        n2157), .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(DataI[8]), .E(n233), .CP(n2210), .CDN(
        n2153), .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(n233), .CP(n2210), .CDN(
        n2157), .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(DataI[9]), .E(n232), .CP(n2220), .CDN(
        n2167), .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(DataI[8]), .E(n232), .CP(n2220), .CDN(
        n2168), .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(DataI[3]), .E(n232), .CP(n2220), .CDN(
        n2169), .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(DataI[9]), .E(n231), .CP(n2223), .CDN(
        n2180), .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(DataI[8]), .E(n231), .CP(n2223), .CDN(
        n2181), .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(DataI[3]), .E(n231), .CP(n2223), .CDN(
        n2171), .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(DataI[9]), .E(n230), .CP(n2229), .CDN(
        n108), .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(DataI[8]), .E(n230), .CP(n2229), .CDN(
        n2148), .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(n230), .CP(n2229), .CDN(
        n2175), .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(DataI[9]), .E(n229), .CP(n2228), .CDN(
        n2183), .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(DataI[8]), .E(n229), .CP(n2227), .CDN(
        n2178), .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(DataI[3]), .E(n229), .CP(n2187), .CDN(
        n2183), .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(n228), .CP(n2224), .CDN(
        n2155), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n228), .CP(n2211), .CDN(
        n2156), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(n228), .CP(n2202), .CDN(
        n2182), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(n227), .CP(n2255), .CDN(
        n108), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(n227), .CP(n2188), .CDN(
        n2162), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(n227), .CP(n2241), .CDN(
        n2162), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(n226), .CP(n2240), .CDN(
        n2152), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(n226), .CP(n2241), .CDN(
        n2164), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(n226), .CP(n2204), .CDN(
        n2149), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(n225), .CP(n2230), .CDN(
        n2166), .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(n225), .CP(n2247), .CDN(
        n2179), .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(n225), .CP(n2245), .CDN(
        n2164), .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n224), .CP(n2248), .CDN(
        n2169), .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n224), .CP(n2232), .CDN(
        n2169), .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n224), .CP(n2243), .CDN(
        n2169), .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n223), .CP(n2242), .CDN(
        n2166), .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n223), .CP(n2255), .CDN(
        n2166), .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n223), .CP(n2235), .CDN(
        n2166), .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n222), .CP(n2186), .CDN(
        n2157), .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n222), .CP(n2241), .CDN(
        n2157), .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n222), .CP(n2233), .CDN(
        n2157), .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n221), .CP(n2186), .CDN(
        n2154), .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n221), .CP(n2227), .CDN(
        n2154), .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n221), .CP(n2196), .CDN(
        n2154), .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(DataI[9]), .E(n220), .CP(n2216), .CDN(
        n108), .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(DataI[8]), .E(n220), .CP(n2216), .CDN(
        n108), .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(DataI[3]), .E(n220), .CP(n2217), .CDN(
        n2178), .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(DataI[9]), .E(n219), .CP(n2255), .CDN(
        n2164), .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(n219), .CP(n2221), .CDN(
        n2152), .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(DataI[3]), .E(n219), .CP(n2219), .CDN(
        n2181), .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(DataI[9]), .E(n218), .CP(n2225), .CDN(
        n2156), .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(DataI[8]), .E(n218), .CP(n2226), .CDN(
        n2185), .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(n218), .CP(n2226), .CDN(
        n2178), .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(DataI[9]), .E(n217), .CP(n2251), .CDN(
        n2173), .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(DataI[8]), .E(n217), .CP(n2190), .CDN(
        n2157), .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(DataI[3]), .E(n217), .CP(n2245), .CDN(
        n2185), .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(n216), .CP(n2194), .CDN(
        n2174), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(n216), .CP(n2225), .CDN(
        n2150), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(n216), .CP(n2215), .CDN(
        n2158), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(n215), .CP(n2240), .CDN(
        n2171), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(n215), .CP(n2197), .CDN(
        n2169), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(n215), .CP(n2247), .CDN(
        n2172), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(n214), .CP(n2223), .CDN(
        n2180), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(n214), .CP(n2250), .CDN(
        n2174), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(n214), .CP(n2245), .CDN(
        n2170), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(n213), .CP(n2234), .CDN(
        n2158), .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(n213), .CP(n2207), .CDN(
        n2177), .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(n213), .CP(n2249), .CDN(
        n2155), .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n212), .CP(n2205), .CDN(
        n2172), .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n212), .CP(n2241), .CDN(
        n2172), .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n212), .CP(n2232), .CDN(
        n2172), .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n211), .CP(n2210), .CDN(
        n2163), .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n211), .CP(n2187), .CDN(
        n2163), .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n211), .CP(n2247), .CDN(
        n2163), .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n210), .CP(n2250), .CDN(
        n2160), .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n210), .CP(n2192), .CDN(
        n2160), .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n210), .CP(n2252), .CDN(
        n2160), .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n209), .CP(n2235), .CDN(
        n2151), .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n209), .CP(n2238), .CDN(
        n2151), .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n209), .CP(n2253), .CDN(
        n2151), .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(n208), .CP(n2190), .CDN(
        n2148), .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(n208), .CP(n2190), .CDN(
        n2179), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(n208), .CP(n2190), .CDN(
        n2181), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(N85), .E(n239), .CP(n2204), .CDN(n2151), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(n239), .CP(n2204), .CDN(
        n2174), .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(DataI[30]), .E(n239), .CP(n2204), .CDN(
        n2148), .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(DataI[29]), .E(n239), .CP(n2204), .CDN(
        n2177), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(n239), .CP(n2204), .CDN(
        n2185), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(n239), .CP(n2205), .CDN(
        n2148), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(DataI[26]), .E(n239), .CP(n2205), .CDN(
        n2177), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(DataI[25]), .E(n239), .CP(n2205), .CDN(
        n2175), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(n239), .CP(n2205), .CDN(
        n2169), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(n239), .CP(n2205), .CDN(
        n2154), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(DataI[22]), .E(n239), .CP(n2205), .CDN(
        n2177), .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(DataI[21]), .E(n239), .CP(n2205), .CDN(
        n2176), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(n239), .CP(n2205), .CDN(
        n2150), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(n239), .CP(n2205), .CDN(
        n2182), .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(DataI[18]), .E(n239), .CP(n2205), .CDN(
        n2152), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(DataI[17]), .E(n239), .CP(n2206), .CDN(
        n2185), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(n239), .CP(n2206), .CDN(
        n2182), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(DataI[15]), .E(n239), .CP(n2206), .CDN(
        n2151), .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(DataI[14]), .E(n239), .CP(n2206), .CDN(
        n2184), .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(n239), .CP(n2206), .CDN(
        n2181), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(DataI[12]), .E(n239), .CP(n2206), .CDN(
        n2167), .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(DataI[11]), .E(n239), .CP(n2206), .CDN(
        n2159), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(DataI[10]), .E(n239), .CP(n2206), .CDN(
        n2148), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(DataI[7]), .E(n239), .CP(n2207), .CDN(
        n2180), .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(DataI[6]), .E(n239), .CP(n2207), .CDN(
        n2156), .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(DataI[5]), .E(n239), .CP(n2207), .CDN(
        n2161), .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(DataI[4]), .E(n239), .CP(n2207), .CDN(
        n2182), .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(DataI[2]), .E(n239), .CP(n2207), .CDN(
        n2180), .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(n239), .CP(n2207), .CDN(
        n2158), .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(DataI[0]), .E(n239), .CP(n2207), .CDN(
        n2163), .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(N85), .E(n238), .CP(n2211), .CDN(n2158), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(DataI[31]), .E(n238), .CP(n2211), .CDN(
        n2166), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(DataI[30]), .E(n238), .CP(n2211), .CDN(
        n2162), .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(DataI[29]), .E(n238), .CP(n2211), .CDN(
        n2163), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(DataI[28]), .E(n238), .CP(n2211), .CDN(
        n2164), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(DataI[27]), .E(n238), .CP(n2211), .CDN(
        n2159), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(DataI[26]), .E(n238), .CP(n2211), .CDN(
        n2160), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(DataI[25]), .E(n238), .CP(n2211), .CDN(
        n2161), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(DataI[24]), .E(n238), .CP(n2211), .CDN(
        n2184), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(DataI[23]), .E(n238), .CP(n2212), .CDN(
        n2184), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(DataI[22]), .E(n238), .CP(n2212), .CDN(
        n2184), .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(DataI[21]), .E(n238), .CP(n2212), .CDN(
        n2178), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(DataI[20]), .E(n238), .CP(n2212), .CDN(
        n2153), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(DataI[19]), .E(n238), .CP(n2212), .CDN(
        n2182), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(DataI[18]), .E(n238), .CP(n2212), .CDN(
        n2167), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(DataI[17]), .E(n238), .CP(n2212), .CDN(
        n2169), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(DataI[16]), .E(n238), .CP(n2212), .CDN(
        n2166), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(DataI[15]), .E(n238), .CP(n2212), .CDN(
        n2148), .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(DataI[14]), .E(n238), .CP(n2212), .CDN(
        n2174), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(DataI[13]), .E(n238), .CP(n2213), .CDN(
        n2180), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(DataI[12]), .E(n238), .CP(n2213), .CDN(
        n2179), .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(DataI[11]), .E(n238), .CP(n2213), .CDN(
        n2182), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(DataI[10]), .E(n238), .CP(n2213), .CDN(
        n2181), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(DataI[7]), .E(n238), .CP(n2213), .CDN(
        n2150), .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(DataI[6]), .E(n238), .CP(n2213), .CDN(
        n2153), .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(DataI[5]), .E(n238), .CP(n2213), .CDN(
        n2158), .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(DataI[4]), .E(n238), .CP(n2213), .CDN(
        n2150), .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(DataI[2]), .E(n238), .CP(n2214), .CDN(
        n2184), .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(DataI[1]), .E(n238), .CP(n2214), .CDN(
        n2161), .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(DataI[0]), .E(n238), .CP(n2214), .CDN(
        n2160), .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(N85), .E(n237), .CP(n2191), .CDN(n2182), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(n237), .CP(n2191), .CDN(
        n2179), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n237), .CP(n2191), .CDN(
        n2170), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(n237), .CP(n2191), .CDN(
        n2167), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(n237), .CP(n2191), .CDN(
        n2168), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(n237), .CP(n2191), .CDN(
        n2169), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n237), .CP(n2191), .CDN(
        n2178), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n237), .CP(n2192), .CDN(
        n2181), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(n237), .CP(n2192), .CDN(
        n2182), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(n237), .CP(n2192), .CDN(
        n2179), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(n237), .CP(n2192), .CDN(
        n2180), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n237), .CP(n2192), .CDN(
        n2178), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(n237), .CP(n2192), .CDN(
        n2181), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(n237), .CP(n2192), .CDN(
        n2182), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n237), .CP(n2192), .CDN(
        n2181), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(n237), .CP(n2192), .CDN(
        n2170), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(n237), .CP(n2192), .CDN(
        n2160), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(n237), .CP(n2193), .CDN(
        n2161), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n237), .CP(n2193), .CDN(
        n2162), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(n237), .CP(n2193), .CDN(
        n2163), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(DataI[12]), .E(n237), .CP(n2193), .CDN(
        n2164), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n237), .CP(n2193), .CDN(
        n2165), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(n237), .CP(n2193), .CDN(
        n2159), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(n237), .CP(n2193), .CDN(
        n2163), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(DataI[6]), .E(n237), .CP(n2193), .CDN(
        n2164), .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(DataI[5]), .E(n237), .CP(n2194), .CDN(
        n2165), .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(n237), .CP(n2194), .CDN(
        n2159), .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(DataI[2]), .E(n237), .CP(n2194), .CDN(
        n2167), .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(n237), .CP(n2194), .CDN(
        n2168), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(DataI[0]), .E(n237), .CP(n2194), .CDN(
        n2169), .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n2147), .E(n236), .CP(n2194), .CDN(n2166), .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(n236), .CP(n2194), .CDN(
        n2159), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(n236), .CP(n2194), .CDN(
        n2151), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(n236), .CP(n2194), .CDN(
        n2167), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(n236), .CP(n2195), .CDN(
        n2168), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(DataI[27]), .E(n236), .CP(n2195), .CDN(
        n2169), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(n236), .CP(n2195), .CDN(
        n2158), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(n236), .CP(n2195), .CDN(
        n2166), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(n236), .CP(n2195), .CDN(
        n2170), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(DataI[23]), .E(n236), .CP(n2195), .CDN(
        n2157), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(n236), .CP(n2195), .CDN(
        n2156), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(n236), .CP(n2195), .CDN(
        n2160), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(n236), .CP(n2195), .CDN(
        n2175), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(n236), .CP(n2195), .CDN(
        n2175), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(DataI[13]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(n236), .CP(n2196), .CDN(
        n2175), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(n236), .CP(n2197), .CDN(
        n2154), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(DataI[6]), .E(n236), .CP(n2197), .CDN(
        n2183), .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(DataI[5]), .E(n236), .CP(n2197), .CDN(
        n2159), .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(n236), .CP(n2197), .CDN(
        n2161), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(n236), .CP(n2197), .CDN(
        n2162), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(n236), .CP(n2197), .CDN(
        n2163), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(DataI[0]), .E(n236), .CP(n2197), .CDN(
        n2160), .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(N85), .E(n235), .CP(n2197), .CDN(n2164), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(n235), .CP(n2198), .CDN(
        n2153), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(DataI[30]), .E(n235), .CP(n2198), .CDN(
        n2155), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(DataI[29]), .E(n235), .CP(n2198), .CDN(
        n2152), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(n235), .CP(n2198), .CDN(
        n2157), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(n235), .CP(n2198), .CDN(
        n2158), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(DataI[26]), .E(n235), .CP(n2198), .CDN(
        n2151), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(DataI[25]), .E(n235), .CP(n2198), .CDN(
        n2156), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(n235), .CP(n2198), .CDN(
        n2185), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(n235), .CP(n2198), .CDN(
        n2148), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(DataI[22]), .E(n235), .CP(n2198), .CDN(
        n2176), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(DataI[21]), .E(n235), .CP(n2199), .CDN(
        n2175), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(n235), .CP(n2199), .CDN(
        n2174), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(n235), .CP(n2199), .CDN(
        n2173), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(DataI[18]), .E(n235), .CP(n2199), .CDN(
        n2183), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(DataI[17]), .E(n235), .CP(n2199), .CDN(
        n2180), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(n235), .CP(n2199), .CDN(
        n2179), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(DataI[15]), .E(n235), .CP(n2199), .CDN(
        n2171), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(DataI[14]), .E(n235), .CP(n2199), .CDN(
        n2185), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(n235), .CP(n2199), .CDN(
        n2148), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(DataI[12]), .E(n235), .CP(n2199), .CDN(
        n2179), .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(DataI[11]), .E(n235), .CP(n2200), .CDN(
        n2172), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(DataI[10]), .E(n235), .CP(n2200), .CDN(
        n2183), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(DataI[7]), .E(n235), .CP(n2200), .CDN(
        n2171), .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(DataI[6]), .E(n235), .CP(n2200), .CDN(
        n2176), .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(DataI[5]), .E(n235), .CP(n2200), .CDN(
        n2150), .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(DataI[4]), .E(n235), .CP(n2200), .CDN(
        n2185), .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(DataI[2]), .E(n235), .CP(n2200), .CDN(
        n2180), .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(DataI[1]), .E(n235), .CP(n2201), .CDN(
        n2179), .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(DataI[0]), .E(n235), .CP(n2201), .CDN(
        n2176), .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n2147), .E(n234), .CP(n2201), .CDN(n2175), .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(n234), .CP(n2201), .CDN(
        n2159), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(n234), .CP(n2201), .CDN(
        n2183), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(DataI[29]), .E(n234), .CP(n2201), .CDN(
        n2183), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(n234), .CP(n2201), .CDN(
        n2176), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(n234), .CP(n2201), .CDN(
        n2171), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(n234), .CP(n2201), .CDN(
        n2174), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(n234), .CP(n2201), .CDN(
        n2167), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(n234), .CP(n2202), .CDN(
        n2168), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(n234), .CP(n2202), .CDN(
        n2169), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(DataI[22]), .E(n234), .CP(n2202), .CDN(
        n2170), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(n234), .CP(n2202), .CDN(
        n2173), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(n234), .CP(n2202), .CDN(
        n2160), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(n234), .CP(n2202), .CDN(
        n2181), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(n234), .CP(n2202), .CDN(
        n2148), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(DataI[17]), .E(n234), .CP(n2202), .CDN(
        n2177), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(n234), .CP(n2202), .CDN(
        n2180), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(DataI[15]), .E(n234), .CP(n2202), .CDN(
        n2179), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(DataI[14]), .E(n234), .CP(n2203), .CDN(
        n2182), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(n234), .CP(n2203), .CDN(
        n2181), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(n234), .CP(n2203), .CDN(
        n2171), .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(n234), .CP(n2203), .CDN(
        n2159), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(DataI[10]), .E(n234), .CP(n2203), .CDN(
        n2170), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(DataI[7]), .E(n234), .CP(n2203), .CDN(
        n2148), .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(DataI[6]), .E(n234), .CP(n2203), .CDN(
        n2161), .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(n234), .CP(n2203), .CDN(
        n2154), .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(DataI[4]), .E(n234), .CP(n2204), .CDN(
        n2179), .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(DataI[2]), .E(n234), .CP(n2204), .CDN(
        n2158), .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(DataI[1]), .E(n234), .CP(n2204), .CDN(
        n2157), .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(n234), .CP(n2204), .CDN(
        n2156), .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n2147), .E(n233), .CP(n2207), .CDN(n2164), .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(n233), .CP(n2207), .CDN(
        n2170), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(DataI[30]), .E(n233), .CP(n2208), .CDN(
        n2148), .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(n233), .CP(n2208), .CDN(
        n2174), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(n233), .CP(n2208), .CDN(
        n2165), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(n233), .CP(n2208), .CDN(
        n2184), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(DataI[26]), .E(n233), .CP(n2208), .CDN(
        n2166), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(DataI[25]), .E(n233), .CP(n2208), .CDN(
        n2159), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(n233), .CP(n2208), .CDN(
        n2160), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(n233), .CP(n2208), .CDN(
        n2165), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(DataI[22]), .E(n233), .CP(n2208), .CDN(
        n2164), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(DataI[21]), .E(n233), .CP(n2208), .CDN(
        n2161), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(n233), .CP(n2209), .CDN(
        n2168), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(n233), .CP(n2209), .CDN(
        n2150), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(DataI[18]), .E(n233), .CP(n2209), .CDN(
        n2184), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(n233), .CP(n2209), .CDN(
        n2166), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(n233), .CP(n2209), .CDN(
        n2159), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(n233), .CP(n2209), .CDN(
        n2160), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(DataI[14]), .E(n233), .CP(n2209), .CDN(
        n2165), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(n233), .CP(n2209), .CDN(
        n2164), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(DataI[12]), .E(n233), .CP(n2209), .CDN(
        n2163), .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(DataI[11]), .E(n233), .CP(n2209), .CDN(
        n2162), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(n233), .CP(n2210), .CDN(
        n2161), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(n233), .CP(n2210), .CDN(
        n2153), .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(DataI[6]), .E(n233), .CP(n2210), .CDN(
        n2167), .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(DataI[5]), .E(n233), .CP(n2210), .CDN(
        n2176), .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(DataI[4]), .E(n233), .CP(n2210), .CDN(
        n2160), .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(n233), .CP(n2210), .CDN(
        n2156), .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(n233), .CP(n2210), .CDN(
        n2173), .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(DataI[0]), .E(n233), .CP(n2211), .CDN(
        n2176), .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(N85), .E(n232), .CP(n2217), .CDN(n2183), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(DataI[31]), .E(n232), .CP(n2217), .CDN(
        n2176), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(DataI[30]), .E(n232), .CP(n2217), .CDN(
        n2174), .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(DataI[29]), .E(n232), .CP(n2218), .CDN(
        n2148), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(DataI[28]), .E(n232), .CP(n2218), .CDN(
        n108), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(DataI[27]), .E(n232), .CP(n2218), .CDN(
        n2183), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(DataI[26]), .E(n232), .CP(n2218), .CDN(
        n2148), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(DataI[25]), .E(n232), .CP(n2218), .CDN(
        n2184), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(DataI[24]), .E(n232), .CP(n2218), .CDN(
        n2173), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(DataI[23]), .E(n232), .CP(n2218), .CDN(
        n108), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(DataI[22]), .E(n232), .CP(n2218), .CDN(
        n2167), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(DataI[21]), .E(n232), .CP(n2218), .CDN(
        n2184), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(DataI[20]), .E(n232), .CP(n2218), .CDN(
        n2175), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(DataI[19]), .E(n232), .CP(n2219), .CDN(
        n2148), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(DataI[18]), .E(n232), .CP(n2219), .CDN(
        n2156), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(DataI[17]), .E(n232), .CP(n2219), .CDN(
        n2176), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(DataI[16]), .E(n232), .CP(n2219), .CDN(
        n2172), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(DataI[15]), .E(n232), .CP(n2219), .CDN(
        n2169), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(DataI[14]), .E(n232), .CP(n2219), .CDN(
        n2161), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(DataI[13]), .E(n232), .CP(n2219), .CDN(
        n2181), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(DataI[12]), .E(n232), .CP(n2219), .CDN(
        n2173), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(DataI[11]), .E(n232), .CP(n2219), .CDN(
        n2181), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(DataI[10]), .E(n232), .CP(n2219), .CDN(
        n2161), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(DataI[7]), .E(n232), .CP(n2220), .CDN(
        n2170), .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(DataI[6]), .E(n232), .CP(n2220), .CDN(
        n2178), .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(DataI[5]), .E(n232), .CP(n2220), .CDN(
        n2177), .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(DataI[4]), .E(n232), .CP(n2220), .CDN(
        n2153), .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(DataI[2]), .E(n232), .CP(n2220), .CDN(
        n2176), .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(DataI[1]), .E(n232), .CP(n2220), .CDN(
        n2156), .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(DataI[0]), .E(n232), .CP(n2220), .CDN(
        n2158), .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(n2147), .E(n231), .CP(n2221), .CDN(n2151), .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(DataI[31]), .E(n231), .CP(n2221), .CDN(
        n108), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(DataI[30]), .E(n231), .CP(n2221), .CDN(
        n108), .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(DataI[29]), .E(n231), .CP(n2221), .CDN(
        n108), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(DataI[28]), .E(n231), .CP(n2221), .CDN(
        n2150), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(n231), .CP(n2221), .CDN(
        n2178), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(DataI[26]), .E(n231), .CP(n2221), .CDN(
        n2177), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(DataI[25]), .E(n231), .CP(n2221), .CDN(
        n2166), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(DataI[24]), .E(n231), .CP(n2221), .CDN(
        n2182), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(n231), .CP(n2221), .CDN(
        n2152), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(DataI[22]), .E(n231), .CP(n2222), .CDN(
        n2170), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(DataI[21]), .E(n231), .CP(n2222), .CDN(
        n2184), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(DataI[20]), .E(n231), .CP(n2222), .CDN(
        n2176), .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(DataI[19]), .E(n231), .CP(n2222), .CDN(
        n2185), .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(n231), .CP(n2222), .CDN(
        n2149), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(DataI[17]), .E(n231), .CP(n2222), .CDN(
        n2166), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(DataI[16]), .E(n231), .CP(n2222), .CDN(
        n2167), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(DataI[15]), .E(n231), .CP(n2222), .CDN(
        n2168), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(DataI[14]), .E(n231), .CP(n2222), .CDN(
        n2169), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(DataI[13]), .E(n231), .CP(n2222), .CDN(
        n2170), .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(DataI[12]), .E(n231), .CP(n2223), .CDN(
        n2178), .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(DataI[11]), .E(n231), .CP(n2223), .CDN(
        n2177), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(DataI[10]), .E(n231), .CP(n2223), .CDN(
        n2170), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(DataI[7]), .E(n231), .CP(n2223), .CDN(
        n2179), .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(DataI[6]), .E(n231), .CP(n2223), .CDN(
        n2185), .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(DataI[5]), .E(n231), .CP(n2223), .CDN(
        n2177), .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(DataI[4]), .E(n231), .CP(n2223), .CDN(
        n2182), .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(DataI[2]), .E(n231), .CP(n2246), .CDN(
        n2181), .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(DataI[1]), .E(n231), .CP(n2231), .CDN(
        n2180), .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(DataI[0]), .E(n231), .CP(n2255), .CDN(
        n2171), .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N85), .E(n230), .CP(n2226), .CDN(n2168), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(DataI[31]), .E(n230), .CP(n2227), .CDN(
        n2172), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(DataI[30]), .E(n230), .CP(n2227), .CDN(
        n2183), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(n230), .CP(n2227), .CDN(
        n2176), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(DataI[28]), .E(n230), .CP(n2227), .CDN(
        n2183), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(DataI[27]), .E(n230), .CP(n2227), .CDN(
        n2154), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(DataI[26]), .E(n230), .CP(n2227), .CDN(
        n2153), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(DataI[25]), .E(n230), .CP(n2227), .CDN(
        n2152), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(DataI[24]), .E(n230), .CP(n2227), .CDN(
        n2151), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(DataI[23]), .E(n230), .CP(n2227), .CDN(
        n2181), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(DataI[22]), .E(n230), .CP(n2227), .CDN(
        n2185), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(DataI[21]), .E(n230), .CP(n2228), .CDN(
        n2154), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(n230), .CP(n2228), .CDN(
        n108), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(DataI[19]), .E(n230), .CP(n2228), .CDN(
        n2150), .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(DataI[18]), .E(n230), .CP(n2228), .CDN(
        n2168), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(n230), .CP(n2228), .CDN(
        n2167), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(DataI[16]), .E(n230), .CP(n2228), .CDN(
        n2161), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(n230), .CP(n2228), .CDN(
        n2180), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(DataI[14]), .E(n230), .CP(n2228), .CDN(
        n108), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(DataI[13]), .E(n230), .CP(n2228), .CDN(
        n2149), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(DataI[12]), .E(n230), .CP(n2228), .CDN(
        n2162), .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(DataI[11]), .E(n230), .CP(n2229), .CDN(
        n2148), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(n230), .CP(n2229), .CDN(
        n2185), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(n230), .CP(n2229), .CDN(
        n2185), .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(DataI[6]), .E(n230), .CP(n2229), .CDN(
        n2175), .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(DataI[5]), .E(n230), .CP(n2229), .CDN(
        n108), .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(DataI[4]), .E(n230), .CP(n2229), .CDN(
        n2150), .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(DataI[2]), .E(n230), .CP(n2229), .CDN(
        n2183), .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(n230), .CP(n2195), .CDN(
        n2151), .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(DataI[0]), .E(n230), .CP(n2194), .CDN(
        n2162), .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n2147), .E(n229), .CP(n2188), .CDN(n108), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(DataI[31]), .E(n229), .CP(n2189), .CDN(
        n2162), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(DataI[30]), .E(n229), .CP(n2193), .CDN(
        n2161), .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(DataI[29]), .E(n229), .CP(n2192), .CDN(
        n2150), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(DataI[28]), .E(n229), .CP(n2196), .CDN(
        n2150), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(DataI[27]), .E(n229), .CP(n2228), .CDN(
        n2177), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(DataI[26]), .E(n229), .CP(n2226), .CDN(
        n108), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(DataI[25]), .E(n229), .CP(n2191), .CDN(
        n2169), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(DataI[24]), .E(n229), .CP(n2222), .CDN(
        n2181), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(DataI[23]), .E(n229), .CP(n2205), .CDN(
        n2149), .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(DataI[22]), .E(n229), .CP(n2212), .CDN(
        n2150), .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(DataI[21]), .E(n229), .CP(n2213), .CDN(
        n2150), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(DataI[20]), .E(n229), .CP(n2214), .CDN(
        n2185), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(DataI[19]), .E(n229), .CP(n2215), .CDN(
        n2164), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(DataI[18]), .E(n229), .CP(n2216), .CDN(
        n2183), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(DataI[17]), .E(n229), .CP(n2217), .CDN(
        n2177), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(DataI[16]), .E(n229), .CP(n2218), .CDN(
        n2150), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(DataI[15]), .E(n229), .CP(n2219), .CDN(
        n2170), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(DataI[14]), .E(n229), .CP(n2226), .CDN(
        n2183), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(DataI[13]), .E(n229), .CP(n2225), .CDN(
        n2176), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(DataI[12]), .E(n229), .CP(n2224), .CDN(
        n2165), .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(DataI[11]), .E(n229), .CP(n2189), .CDN(
        n2159), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(DataI[10]), .E(n229), .CP(n2246), .CDN(
        n2153), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(DataI[7]), .E(n229), .CP(n2238), .CDN(
        n2173), .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(DataI[6]), .E(n229), .CP(n2248), .CDN(
        n2184), .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(DataI[5]), .E(n229), .CP(n2199), .CDN(
        n2158), .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(DataI[4]), .E(n229), .CP(n2243), .CDN(
        n2148), .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(DataI[2]), .E(n229), .CP(n2251), .CDN(
        n2177), .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(DataI[1]), .E(n229), .CP(n2250), .CDN(
        n2149), .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(DataI[0]), .E(n229), .CP(n2187), .CDN(
        n2154), .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N85), .E(n228), .CP(n2210), .CDN(n2149), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(n228), .CP(n2200), .CDN(
        n2160), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(n228), .CP(n2201), .CDN(
        n2183), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(n228), .CP(n2202), .CDN(
        n2172), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n228), .CP(n2203), .CDN(
        n2150), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n228), .CP(n2204), .CDN(
        n2152), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n228), .CP(n2205), .CDN(
        n2150), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(n228), .CP(n2206), .CDN(
        n2182), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n228), .CP(n2207), .CDN(
        n2166), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n228), .CP(n2211), .CDN(
        n2158), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(n228), .CP(n2207), .CDN(
        n2171), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n228), .CP(n2206), .CDN(
        n2184), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(n228), .CP(n2209), .CDN(
        n2173), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n228), .CP(n2208), .CDN(
        n2177), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(n228), .CP(n2202), .CDN(
        n2185), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(n228), .CP(n2203), .CDN(
        n2176), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(n228), .CP(n2200), .CDN(
        n2180), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(n228), .CP(n2201), .CDN(
        n2178), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(n228), .CP(n2205), .CDN(
        n2152), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(n228), .CP(n2204), .CDN(
        n2181), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(n228), .CP(n2209), .CDN(
        n2172), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n228), .CP(n2198), .CDN(
        n2184), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(n228), .CP(n2199), .CDN(
        n2150), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(n228), .CP(n2228), .CDN(
        n2181), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(n228), .CP(n2240), .CDN(
        n2162), .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(n228), .CP(n2187), .CDN(
        n2176), .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(n228), .CP(ClockW), .CDN(
        n2149), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(n228), .CP(n2225), .CDN(
        n2185), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(n228), .CP(n2226), .CDN(
        n2163), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(n228), .CP(n2227), .CDN(
        n2177), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n2147), .E(n227), .CP(n2228), .CDN(n108), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(n227), .CP(n2229), .CDN(
        n2154), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(n227), .CP(n2221), .CDN(
        n2171), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n227), .CP(n2220), .CDN(
        n2166), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(n227), .CP(n2200), .CDN(
        n2176), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(n227), .CP(n2201), .CDN(
        n2148), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(n227), .CP(n2211), .CDN(
        n2165), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(n227), .CP(ClockW), .CDN(
        n2151), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(n227), .CP(n2212), .CDN(
        n2176), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(n227), .CP(n2213), .CDN(
        n2182), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(n227), .CP(n2214), .CDN(
        n2155), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(n227), .CP(n2215), .CDN(
        n2172), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n227), .CP(n2216), .CDN(
        n2157), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(n227), .CP(n2217), .CDN(
        n2168), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(n227), .CP(n2198), .CDN(
        n2154), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n227), .CP(n2214), .CDN(
        n2169), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(n227), .CP(n2237), .CDN(
        n2155), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n227), .CP(n2213), .CDN(
        n108), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(n227), .CP(n2223), .CDN(
        n2169), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(n227), .CP(n2197), .CDN(
        n2181), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(n227), .CP(ClockW), .CDN(
        n2154), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(n227), .CP(n2251), .CDN(
        n2166), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n227), .CP(n2254), .CDN(
        n2176), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(n227), .CP(n2187), .CDN(
        n108), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(DataI[6]), .E(n227), .CP(n2225), .CDN(
        n2151), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(n227), .CP(n2236), .CDN(
        n2175), .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(n227), .CP(n2237), .CDN(
        n2174), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(n227), .CP(n2244), .CDN(
        n2185), .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n227), .CP(n2231), .CDN(
        n2174), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(n227), .CP(n2224), .CDN(
        n2171), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N85), .E(n226), .CP(n2252), .CDN(n2168), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(n226), .CP(n2231), .CDN(
        n2183), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(n226), .CP(n2220), .CDN(
        n2184), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(n226), .CP(n2186), .CDN(
        n2180), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(n226), .CP(n2208), .CDN(
        n2179), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(n226), .CP(n2232), .CDN(
        n2181), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(n226), .CP(n2252), .CDN(
        n2182), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(n226), .CP(n2246), .CDN(
        n2162), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(n226), .CP(n2240), .CDN(
        n2161), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(n226), .CP(n2247), .CDN(
        n2160), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(n226), .CP(n2231), .CDN(
        n2159), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(n226), .CP(n2248), .CDN(
        n2166), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(n226), .CP(ClockW), .CDN(
        n2176), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(n226), .CP(n2226), .CDN(
        n2151), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(n226), .CP(n2249), .CDN(
        n2177), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(n226), .CP(n2248), .CDN(
        n2185), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(n226), .CP(n2247), .CDN(
        n2184), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(DataI[15]), .E(n226), .CP(n2245), .CDN(
        n2155), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(DataI[14]), .E(n226), .CP(n2244), .CDN(
        n2183), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(DataI[13]), .E(n226), .CP(n2186), .CDN(
        n2178), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(n226), .CP(n2243), .CDN(
        n2185), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(n226), .CP(n2242), .CDN(
        n2165), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(n226), .CP(n2241), .CDN(
        n2173), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(DataI[7]), .E(n226), .CP(n2238), .CDN(
        n2164), .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(DataI[6]), .E(n226), .CP(n2239), .CDN(
        n2170), .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(DataI[5]), .E(n226), .CP(n2204), .CDN(
        n2152), .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(n226), .CP(n2255), .CDN(
        n2172), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(n226), .CP(n2210), .CDN(
        n2181), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(n226), .CP(n2247), .CDN(
        n2183), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(n226), .CP(n2255), .CDN(
        n2163), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n2147), .E(n225), .CP(n2234), .CDN(n2171), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(n225), .CP(n2201), .CDN(
        n2183), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(n225), .CP(n2199), .CDN(
        n2153), .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(n225), .CP(n2230), .CDN(
        n2173), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(n225), .CP(n2246), .CDN(
        n2155), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(n225), .CP(n2255), .CDN(
        n2177), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(n225), .CP(n2196), .CDN(
        n2184), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(n225), .CP(n2186), .CDN(
        n2165), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(n225), .CP(n2213), .CDN(
        n2154), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(n225), .CP(ClockW), .CDN(
        n2182), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n225), .CP(n2246), .CDN(
        n2168), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(n225), .CP(n2232), .CDN(
        n2178), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(n225), .CP(n2190), .CDN(
        n2163), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(n225), .CP(n2252), .CDN(
        n2167), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(n225), .CP(n2247), .CDN(
        n2183), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(n225), .CP(n2186), .CDN(
        n2172), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(n225), .CP(n2243), .CDN(
        n2179), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(DataI[15]), .E(n225), .CP(n2235), .CDN(
        n2155), .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(n225), .CP(n2188), .CDN(
        n2161), .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(n225), .CP(n2241), .CDN(
        n2172), .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n225), .CP(n2199), .CDN(
        n2166), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(n225), .CP(n2192), .CDN(
        n2175), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(n225), .CP(n2206), .CDN(
        n2175), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(DataI[7]), .E(n225), .CP(n2224), .CDN(
        n2184), .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(n225), .CP(n2191), .CDN(
        n2177), .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(n225), .CP(n2187), .CDN(
        n2151), .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n225), .CP(n2201), .CDN(
        n2157), .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(n225), .CP(n2248), .CDN(
        n2172), .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(n225), .CP(n2186), .CDN(
        n2148), .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n225), .CP(n2198), .CDN(
        n2165), .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N85), .E(n224), .CP(n2255), .CDN(n2172), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n224), .CP(n2240), .CDN(
        n2171), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n224), .CP(n2239), .CDN(
        n2171), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n224), .CP(n2238), .CDN(
        n2171), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n224), .CP(n2234), .CDN(
        n2171), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n224), .CP(n2216), .CDN(
        n2171), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n224), .CP(n2253), .CDN(
        n2171), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n224), .CP(n2235), .CDN(
        n2171), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n224), .CP(n2199), .CDN(
        n2171), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n224), .CP(n2244), .CDN(
        n2171), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n224), .CP(n2253), .CDN(
        n2171), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n224), .CP(n2232), .CDN(
        n2171), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n224), .CP(n2237), .CDN(
        n2170), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n224), .CP(n2254), .CDN(
        n2170), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n224), .CP(n2187), .CDN(
        n2170), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n224), .CP(n2241), .CDN(
        n2170), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n224), .CP(n2240), .CDN(
        n2170), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n224), .CP(n2239), .CDN(
        n2170), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n224), .CP(n2238), .CDN(
        n2170), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n224), .CP(n2242), .CDN(
        n2170), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n224), .CP(n2243), .CDN(
        n2170), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n224), .CP(n2241), .CDN(
        n2170), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n224), .CP(n2247), .CDN(
        n2170), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n224), .CP(n2254), .CDN(
        n2169), .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n224), .CP(n2209), .CDN(
        n2169), .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n224), .CP(n2249), .CDN(
        n2169), .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n224), .CP(n2248), .CDN(
        n2169), .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n224), .CP(n2247), .CDN(
        n2169), .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n224), .CP(n2246), .CDN(
        n2169), .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n224), .CP(n2245), .CDN(
        n2169), .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n2147), .E(n223), .CP(n2244), .CDN(n2169), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n223), .CP(n2186), .CDN(
        n2168), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n223), .CP(n2233), .CDN(
        n2168), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n223), .CP(n2238), .CDN(
        n2168), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n223), .CP(n2241), .CDN(
        n2168), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n223), .CP(n2231), .CDN(
        n2168), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n223), .CP(n2192), .CDN(
        n2168), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n223), .CP(n2232), .CDN(
        n2168), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n223), .CP(n2231), .CDN(
        n2168), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n223), .CP(n2230), .CDN(
        n2168), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n223), .CP(n2245), .CDN(
        n2168), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n223), .CP(n2231), .CDN(
        n2168), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n223), .CP(n2239), .CDN(
        n2167), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n223), .CP(n2205), .CDN(
        n2167), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n223), .CP(n2193), .CDN(
        n2167), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n223), .CP(n2243), .CDN(
        n2167), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n223), .CP(n2197), .CDN(
        n2167), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n223), .CP(n2190), .CDN(
        n2167), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n223), .CP(n2204), .CDN(
        n2167), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n223), .CP(n2242), .CDN(
        n2167), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n223), .CP(n2241), .CDN(
        n2167), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n223), .CP(n2240), .CDN(
        n2167), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n223), .CP(n2236), .CDN(
        n2167), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n223), .CP(ClockW), .CDN(
        n2166), .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n223), .CP(n2242), .CDN(
        n2166), .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n223), .CP(n2234), .CDN(
        n2166), .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n223), .CP(n2225), .CDN(
        n2166), .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n223), .CP(n2253), .CDN(
        n2166), .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n223), .CP(n2244), .CDN(
        n2166), .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n223), .CP(n2236), .CDN(
        n2166), .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(n222), .CP(n2250), .CDN(n2160), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n222), .CP(n2253), .CDN(
        n2159), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n222), .CP(n2254), .CDN(
        n2159), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(n222), .CP(n2241), .CDN(
        n2159), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n222), .CP(n2253), .CDN(
        n2159), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n222), .CP(n2251), .CDN(
        n2159), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n222), .CP(n2186), .CDN(
        n2159), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n222), .CP(n2210), .CDN(
        n2159), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n222), .CP(n2239), .CDN(
        n2159), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n222), .CP(n2242), .CDN(
        n2159), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n222), .CP(n2240), .CDN(
        n2159), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n222), .CP(n2239), .CDN(
        n2159), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n222), .CP(n2238), .CDN(
        n2158), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n222), .CP(n2233), .CDN(
        n2158), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n222), .CP(n2236), .CDN(
        n2158), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n222), .CP(n2237), .CDN(
        n2158), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n222), .CP(n2227), .CDN(
        n2158), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n222), .CP(n2238), .CDN(
        n2158), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n222), .CP(n2203), .CDN(
        n2158), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n222), .CP(n2187), .CDN(
        n2158), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n222), .CP(n2233), .CDN(
        n2158), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n222), .CP(n2250), .CDN(
        n2158), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n222), .CP(n2202), .CDN(
        n2158), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n222), .CP(n2211), .CDN(
        n2157), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n222), .CP(n2249), .CDN(
        n2157), .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n222), .CP(n2248), .CDN(
        n2157), .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n222), .CP(n2247), .CDN(
        n2157), .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n222), .CP(n2246), .CDN(
        n2157), .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n222), .CP(n2245), .CDN(
        n2157), .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n222), .CP(n2244), .CDN(
        n2157), .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n2147), .E(n221), .CP(n2242), .CDN(n2157), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n221), .CP(n2240), .CDN(
        n2156), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n221), .CP(n2218), .CDN(
        n2156), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n221), .CP(n2237), .CDN(
        n2156), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n221), .CP(n2236), .CDN(
        n2156), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n221), .CP(n2235), .CDN(
        n2156), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n221), .CP(n2234), .CDN(
        n2156), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n221), .CP(n2233), .CDN(
        n2156), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n221), .CP(n2203), .CDN(
        n2156), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n221), .CP(n2243), .CDN(
        n2156), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n221), .CP(n2202), .CDN(
        n2156), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n221), .CP(n2233), .CDN(
        n2156), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n221), .CP(n2238), .CDN(
        n2155), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n221), .CP(n2239), .CDN(
        n2155), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n221), .CP(n2251), .CDN(
        n2155), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n221), .CP(n2255), .CDN(
        n2155), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n221), .CP(n2190), .CDN(
        n2155), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n221), .CP(n2232), .CDN(
        n2155), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n221), .CP(n2231), .CDN(
        n2155), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n221), .CP(n2230), .CDN(
        n2155), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n221), .CP(n2222), .CDN(
        n2155), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n221), .CP(n2250), .CDN(
        n2155), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n221), .CP(n2235), .CDN(
        n2155), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n221), .CP(n2234), .CDN(
        n2154), .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n221), .CP(n2253), .CDN(
        n2154), .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n221), .CP(n2233), .CDN(
        n2154), .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n221), .CP(n2242), .CDN(
        n2154), .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n221), .CP(n2193), .CDN(
        n2154), .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n221), .CP(n2206), .CDN(
        n2154), .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n221), .CP(ClockW), .CDN(
        n2154), .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n2147), .E(n220), .CP(n2214), .CDN(n2159), .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(DataI[31]), .E(n220), .CP(n2214), .CDN(
        n2172), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(DataI[30]), .E(n220), .CP(n2214), .CDN(
        n2177), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(DataI[29]), .E(n220), .CP(n2214), .CDN(
        n2149), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(DataI[28]), .E(n220), .CP(n2214), .CDN(
        n2184), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(DataI[27]), .E(n220), .CP(n2214), .CDN(
        n2153), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(DataI[26]), .E(n220), .CP(n2215), .CDN(
        n2158), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(DataI[25]), .E(n220), .CP(n2215), .CDN(
        n108), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(DataI[24]), .E(n220), .CP(n2215), .CDN(
        n2163), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(DataI[23]), .E(n220), .CP(n2215), .CDN(
        n2180), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(DataI[22]), .E(n220), .CP(n2215), .CDN(
        n2181), .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(DataI[21]), .E(n220), .CP(n2215), .CDN(
        n108), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(DataI[20]), .E(n220), .CP(n2215), .CDN(
        n2177), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(DataI[19]), .E(n220), .CP(n2215), .CDN(
        n108), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(DataI[18]), .E(n220), .CP(n2215), .CDN(
        n2152), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(DataI[17]), .E(n220), .CP(n2215), .CDN(
        n2168), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(DataI[16]), .E(n220), .CP(n2216), .CDN(
        n2185), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(DataI[15]), .E(n220), .CP(n2216), .CDN(
        n2170), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(DataI[14]), .E(n220), .CP(n2216), .CDN(
        n2148), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(DataI[13]), .E(n220), .CP(n2216), .CDN(
        n2175), .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(DataI[12]), .E(n220), .CP(n2216), .CDN(
        n108), .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(DataI[11]), .E(n220), .CP(n2216), .CDN(
        n2160), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(DataI[10]), .E(n220), .CP(n2216), .CDN(
        n2179), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(DataI[7]), .E(n220), .CP(n2216), .CDN(
        n2178), .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(DataI[6]), .E(n220), .CP(n2217), .CDN(
        n2184), .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(DataI[5]), .E(n220), .CP(n2217), .CDN(
        n108), .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(DataI[4]), .E(n220), .CP(n2217), .CDN(
        n108), .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(DataI[2]), .E(n220), .CP(n2217), .CDN(
        n2150), .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(DataI[1]), .E(n220), .CP(n2217), .CDN(
        n2171), .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(DataI[0]), .E(n220), .CP(n2217), .CDN(
        n2182), .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N85), .E(n219), .CP(n2252), .CDN(n2155), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(n219), .CP(n2250), .CDN(
        n2181), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(n219), .CP(n2254), .CDN(
        n2158), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(DataI[29]), .E(n219), .CP(n2229), .CDN(
        n2155), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(n219), .CP(n2253), .CDN(
        n2183), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(n219), .CP(n2243), .CDN(
        n2179), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(n219), .CP(n2186), .CDN(
        n2175), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(n219), .CP(n2242), .CDN(
        n2157), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(n219), .CP(n2196), .CDN(
        n2163), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(n219), .CP(n2245), .CDN(
        n2149), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(DataI[22]), .E(n219), .CP(n2244), .CDN(
        n2149), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(n219), .CP(n2234), .CDN(
        n2170), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(DataI[20]), .E(n219), .CP(n2233), .CDN(
        n2157), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(n219), .CP(n2200), .CDN(
        n2153), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(n219), .CP(n2235), .CDN(
        n2185), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(DataI[17]), .E(n219), .CP(n2236), .CDN(
        n2173), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(n219), .CP(n2237), .CDN(
        n2163), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(DataI[15]), .E(n219), .CP(n2220), .CDN(
        n2182), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(n219), .CP(n2217), .CDN(
        n2165), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(n219), .CP(n2214), .CDN(
        n2178), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(DataI[12]), .E(n219), .CP(n2215), .CDN(
        n2174), .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(n219), .CP(n2212), .CDN(
        n2178), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(DataI[10]), .E(n219), .CP(n2213), .CDN(
        n2155), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(DataI[7]), .E(n219), .CP(n2254), .CDN(
        n2157), .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(DataI[6]), .E(n219), .CP(n2234), .CDN(
        n2151), .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(DataI[5]), .E(n219), .CP(n2233), .CDN(
        n2173), .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(DataI[4]), .E(n219), .CP(n2247), .CDN(
        n2159), .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(DataI[2]), .E(n219), .CP(n2248), .CDN(
        n2173), .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(DataI[1]), .E(n219), .CP(n2249), .CDN(
        n2175), .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(DataI[0]), .E(n219), .CP(n2235), .CDN(
        n2150), .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(n2147), .E(n218), .CP(n2236), .CDN(n2160), .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(DataI[31]), .E(n218), .CP(n2237), .CDN(
        n2164), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(DataI[30]), .E(n218), .CP(n2232), .CDN(
        n2156), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(n218), .CP(n2230), .CDN(
        n2165), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(DataI[28]), .E(n218), .CP(n2224), .CDN(
        n2166), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(DataI[27]), .E(n218), .CP(n2224), .CDN(
        n2158), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(DataI[26]), .E(n218), .CP(n2224), .CDN(
        n2153), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(DataI[25]), .E(n218), .CP(n2224), .CDN(
        n2182), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(DataI[24]), .E(n218), .CP(n2224), .CDN(
        n2180), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(DataI[23]), .E(n218), .CP(n2224), .CDN(
        n2179), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(DataI[22]), .E(n218), .CP(n2224), .CDN(
        n2184), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(DataI[21]), .E(n218), .CP(n2224), .CDN(
        n2154), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(n218), .CP(n2224), .CDN(
        n2183), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(DataI[19]), .E(n218), .CP(n2224), .CDN(
        n2148), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(DataI[18]), .E(n218), .CP(n2225), .CDN(
        n2156), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(n218), .CP(n2225), .CDN(
        n2168), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(DataI[16]), .E(n218), .CP(n2225), .CDN(
        n2151), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(n218), .CP(n2225), .CDN(
        n2176), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(DataI[14]), .E(n218), .CP(n2225), .CDN(
        n2171), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(DataI[13]), .E(n218), .CP(n2225), .CDN(
        n2148), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(DataI[12]), .E(n218), .CP(n2225), .CDN(
        n2177), .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(DataI[11]), .E(n218), .CP(n2225), .CDN(
        n2179), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(n218), .CP(n2225), .CDN(
        n2150), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(n218), .CP(n2226), .CDN(
        n2170), .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(DataI[6]), .E(n218), .CP(n2226), .CDN(
        n2169), .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(DataI[5]), .E(n218), .CP(n2226), .CDN(
        n2167), .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(DataI[4]), .E(n218), .CP(n2226), .CDN(
        n2178), .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(DataI[2]), .E(n218), .CP(n2226), .CDN(
        n2185), .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(n218), .CP(n2226), .CDN(
        n2184), .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(DataI[0]), .E(n218), .CP(n2226), .CDN(
        n2157), .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(n217), .CP(n2252), .CDN(n2152), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(DataI[31]), .E(n217), .CP(n2253), .CDN(
        n2177), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(DataI[30]), .E(n217), .CP(n2254), .CDN(
        n2164), .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(DataI[29]), .E(n217), .CP(n2228), .CDN(
        n2175), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(DataI[28]), .E(n217), .CP(n2255), .CDN(
        n2151), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(DataI[27]), .E(n217), .CP(n2197), .CDN(
        n2185), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(DataI[26]), .E(n217), .CP(n2223), .CDN(
        n2153), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(DataI[25]), .E(n217), .CP(n2188), .CDN(
        n2148), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(DataI[24]), .E(n217), .CP(n2189), .CDN(
        n2162), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(DataI[23]), .E(n217), .CP(n2229), .CDN(
        n2157), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(DataI[22]), .E(n217), .CP(n2236), .CDN(
        n2154), .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(DataI[21]), .E(n217), .CP(n2191), .CDN(
        n2162), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(DataI[20]), .E(n217), .CP(n2192), .CDN(
        n2172), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(DataI[19]), .E(n217), .CP(n2193), .CDN(
        n2184), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(DataI[18]), .E(n217), .CP(n2194), .CDN(
        n2172), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(DataI[17]), .E(n217), .CP(n2229), .CDN(
        n2172), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(DataI[16]), .E(n217), .CP(n2197), .CDN(
        n108), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(DataI[15]), .E(n217), .CP(n2198), .CDN(
        n2159), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(DataI[14]), .E(n217), .CP(n2199), .CDN(
        n2179), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(DataI[13]), .E(n217), .CP(n2208), .CDN(
        n2178), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(DataI[12]), .E(n217), .CP(n2209), .CDN(
        n2152), .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(DataI[11]), .E(n217), .CP(n2206), .CDN(
        n2169), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(DataI[10]), .E(n217), .CP(n2207), .CDN(
        n2180), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(DataI[7]), .E(n217), .CP(n2221), .CDN(
        n2166), .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(DataI[6]), .E(n217), .CP(n2251), .CDN(
        n2176), .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(DataI[5]), .E(n217), .CP(n2238), .CDN(
        n2180), .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(DataI[4]), .E(n217), .CP(n2253), .CDN(
        n2174), .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(DataI[2]), .E(n217), .CP(n2187), .CDN(
        n2181), .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(DataI[1]), .E(n217), .CP(n2250), .CDN(
        n2163), .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(DataI[0]), .E(n217), .CP(n2255), .CDN(
        n2174), .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n2147), .E(n216), .CP(n2232), .CDN(n2154), .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n216), .CP(n2254), .CDN(
        n2179), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(n216), .CP(n2246), .CDN(
        n2182), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(n216), .CP(n2249), .CDN(
        n2180), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(n216), .CP(n2247), .CDN(
        n2185), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(n216), .CP(n2200), .CDN(
        n2154), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(n216), .CP(n2195), .CDN(
        n2165), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(n216), .CP(n2223), .CDN(
        n2165), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(n216), .CP(n2232), .CDN(
        n108), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(n216), .CP(n2230), .CDN(
        n108), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(n216), .CP(n2231), .CDN(
        n108), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n216), .CP(n2242), .CDN(
        n2180), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(n216), .CP(n2214), .CDN(
        n2182), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n216), .CP(n2248), .CDN(
        n2158), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n216), .CP(n2211), .CDN(
        n2156), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(n216), .CP(n2190), .CDN(
        n2174), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n216), .CP(n2237), .CDN(
        n2173), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(n216), .CP(n2196), .CDN(
        n2177), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n216), .CP(n2210), .CDN(
        n2154), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n216), .CP(n2252), .CDN(
        n2176), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(n216), .CP(n2235), .CDN(
        n2184), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n216), .CP(n2212), .CDN(
        n2163), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(n216), .CP(n2216), .CDN(
        n2175), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(n216), .CP(n2217), .CDN(
        n2184), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(n216), .CP(n2218), .CDN(
        n2179), .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(n216), .CP(n2219), .CDN(
        n2175), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(n216), .CP(n2220), .CDN(
        n2178), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(n216), .CP(n2221), .CDN(
        n2171), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(n216), .CP(n2222), .CDN(
        n2181), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(n216), .CP(n2208), .CDN(
        n2182), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(n215), .CP(n2249), .CDN(n2177), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(n215), .CP(ClockW), .CDN(
        n2153), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(n215), .CP(n2196), .CDN(
        n2153), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(n215), .CP(n2251), .CDN(
        n2172), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(n215), .CP(n2244), .CDN(
        n2166), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(n215), .CP(n2222), .CDN(
        n2171), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(n215), .CP(n2197), .CDN(
        n2172), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(n215), .CP(n2231), .CDN(
        n2164), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(n215), .CP(n2230), .CDN(
        n2184), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(n215), .CP(n2241), .CDN(
        n2156), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(n215), .CP(ClockW), .CDN(
        n2162), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(n215), .CP(n2193), .CDN(
        n2178), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(n215), .CP(n2190), .CDN(
        n2151), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(n215), .CP(n2244), .CDN(
        n2183), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(n215), .CP(n2234), .CDN(
        n2151), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(n215), .CP(n2245), .CDN(
        n2155), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(n215), .CP(n2232), .CDN(
        n2182), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(DataI[15]), .E(n215), .CP(n2195), .CDN(
        n2175), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(DataI[14]), .E(n215), .CP(n2225), .CDN(
        n2155), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(n215), .CP(n2230), .CDN(
        n2174), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(n215), .CP(n2231), .CDN(
        n2179), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(n215), .CP(n2245), .CDN(
        n2171), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(n215), .CP(n2246), .CDN(
        n2165), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(DataI[7]), .E(n215), .CP(n2248), .CDN(
        n2185), .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(DataI[6]), .E(n215), .CP(n2249), .CDN(
        n2164), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(DataI[5]), .E(n215), .CP(n2241), .CDN(
        n2177), .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(n215), .CP(n2243), .CDN(
        n2150), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(n215), .CP(n2242), .CDN(
        n2148), .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(n215), .CP(n2238), .CDN(
        n2185), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(n215), .CP(n2239), .CDN(
        n2183), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n2147), .E(n214), .CP(n2239), .CDN(n2184), .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(n214), .CP(n2209), .CDN(
        n2177), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(n214), .CP(n2187), .CDN(
        n2148), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(n214), .CP(n2186), .CDN(
        n2150), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(n214), .CP(n2243), .CDN(
        n2173), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(n214), .CP(n2242), .CDN(
        n2157), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(n214), .CP(n2241), .CDN(
        n2168), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(n214), .CP(n2240), .CDN(
        n2163), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(n214), .CP(n2239), .CDN(
        n2150), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(n214), .CP(n2238), .CDN(
        n2167), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(n214), .CP(n2195), .CDN(
        n2169), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(n214), .CP(n2245), .CDN(
        n2171), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(n214), .CP(n2237), .CDN(
        n2157), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(n214), .CP(n2236), .CDN(
        n2155), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(n214), .CP(n2235), .CDN(
        n2152), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(n214), .CP(n2254), .CDN(
        n2165), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(n214), .CP(n2249), .CDN(
        n2158), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(DataI[15]), .E(n214), .CP(n2191), .CDN(
        n2156), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(DataI[14]), .E(n214), .CP(n2229), .CDN(
        n2176), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(n214), .CP(n2227), .CDN(
        n2167), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(n214), .CP(n2195), .CDN(
        n2151), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(n214), .CP(n2250), .CDN(
        n2154), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(n214), .CP(n2218), .CDN(
        n108), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(DataI[7]), .E(n214), .CP(n2219), .CDN(
        n2174), .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(DataI[6]), .E(n214), .CP(n2220), .CDN(
        n2169), .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(DataI[5]), .E(n214), .CP(n2221), .CDN(
        n2172), .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(n214), .CP(n2222), .CDN(
        n2168), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(n214), .CP(n2187), .CDN(
        n2167), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(n214), .CP(n2250), .CDN(
        n2160), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(n214), .CP(n2251), .CDN(
        n2174), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(n213), .CP(n2239), .CDN(n2185), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(n213), .CP(n2255), .CDN(
        n2165), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(n213), .CP(n2239), .CDN(
        n2153), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(n213), .CP(n2240), .CDN(
        n2152), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(n213), .CP(n2231), .CDN(
        n2185), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(n213), .CP(n2205), .CDN(
        n2165), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(n213), .CP(n2187), .CDN(
        n2150), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(n213), .CP(n2198), .CDN(
        n2151), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(n213), .CP(n2250), .CDN(
        n2154), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(n213), .CP(n2251), .CDN(
        n2168), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(n213), .CP(n2248), .CDN(
        n2149), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(n213), .CP(n2246), .CDN(
        n2154), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(n213), .CP(n2236), .CDN(
        n2150), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(n213), .CP(n2215), .CDN(
        n2184), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(n213), .CP(n2187), .CDN(
        n2164), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(n213), .CP(ClockW), .CDN(
        n2152), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(n213), .CP(n2206), .CDN(
        n2163), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(DataI[15]), .E(n213), .CP(n2247), .CDN(
        n2156), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(n213), .CP(n2248), .CDN(
        n2178), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(n213), .CP(n2249), .CDN(
        n2166), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n213), .CP(n2244), .CDN(
        n2149), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(n213), .CP(n2246), .CDN(
        n2158), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(n213), .CP(n2245), .CDN(
        n2162), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(DataI[7]), .E(n213), .CP(n2244), .CDN(
        n2162), .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(n213), .CP(n2186), .CDN(
        n2152), .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(n213), .CP(n2237), .CDN(
        n2150), .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(n213), .CP(n2236), .CDN(
        n2159), .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(n213), .CP(n2235), .CDN(
        n2155), .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(n213), .CP(n2249), .CDN(
        n2158), .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n213), .CP(n2238), .CDN(
        n2151), .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n2147), .E(n212), .CP(n2237), .CDN(n2163), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n212), .CP(n2240), .CDN(
        n2174), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n212), .CP(n2194), .CDN(
        n2174), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n212), .CP(n2239), .CDN(
        n2174), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n212), .CP(n2243), .CDN(
        n2174), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n212), .CP(n2228), .CDN(
        n2174), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n212), .CP(n2207), .CDN(
        n2174), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n212), .CP(n2193), .CDN(
        n2174), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n212), .CP(n2232), .CDN(
        n2174), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(n212), .CP(n2249), .CDN(
        n2174), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n212), .CP(n2252), .CDN(
        n2174), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n212), .CP(n2212), .CDN(
        n2174), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n212), .CP(n2227), .CDN(
        n2173), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n212), .CP(n2229), .CDN(
        n2173), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n212), .CP(n2235), .CDN(
        n2173), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n212), .CP(n2249), .CDN(
        n2173), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n212), .CP(ClockW), .CDN(
        n2173), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n212), .CP(n2236), .CDN(
        n2173), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n212), .CP(n2231), .CDN(
        n2173), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n212), .CP(n2230), .CDN(
        n2173), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n212), .CP(n2216), .CDN(
        n2173), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n212), .CP(n2234), .CDN(
        n2173), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n212), .CP(n2192), .CDN(
        n2173), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n212), .CP(n2242), .CDN(
        n2172), .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n212), .CP(n2198), .CDN(
        n2172), .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n212), .CP(n2191), .CDN(
        n2172), .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n212), .CP(n2233), .CDN(
        n2172), .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n212), .CP(n2204), .CDN(
        n2172), .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n212), .CP(n2236), .CDN(
        n2172), .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n212), .CP(n2235), .CDN(
        n2172), .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(n211), .CP(n2250), .CDN(n2166), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n211), .CP(n2230), .CDN(
        n2165), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n211), .CP(n2223), .CDN(
        n2165), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n211), .CP(n2189), .CDN(
        n2165), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n211), .CP(n2217), .CDN(
        n2165), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n211), .CP(n2251), .CDN(
        n2165), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n211), .CP(n2252), .CDN(
        n2165), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n211), .CP(ClockW), .CDN(
        n2165), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n211), .CP(n2186), .CDN(
        n2165), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n211), .CP(n2244), .CDN(
        n2165), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n211), .CP(n2232), .CDN(
        n2165), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n211), .CP(n2253), .CDN(
        n2165), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n211), .CP(n2251), .CDN(
        n2164), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n211), .CP(n2237), .CDN(
        n2164), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n211), .CP(n2186), .CDN(
        n2164), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n211), .CP(n2243), .CDN(
        n2164), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n211), .CP(n2208), .CDN(
        n2164), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n211), .CP(n2246), .CDN(
        n2164), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n211), .CP(n2245), .CDN(
        n2164), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n211), .CP(n2191), .CDN(
        n2164), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n211), .CP(n2232), .CDN(
        n2164), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n211), .CP(n2231), .CDN(
        n2164), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n211), .CP(n2230), .CDN(
        n2164), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n211), .CP(n2203), .CDN(
        n2163), .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n211), .CP(n2210), .CDN(
        n2163), .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n211), .CP(n2226), .CDN(
        n2163), .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n211), .CP(n2219), .CDN(
        n2163), .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n211), .CP(n2233), .CDN(
        n2163), .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n211), .CP(n2208), .CDN(
        n2163), .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n211), .CP(n2254), .CDN(
        n2163), .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n2147), .E(n210), .CP(n2209), .CDN(n2163), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n210), .CP(n2252), .CDN(
        n2162), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n210), .CP(n2254), .CDN(
        n2162), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n210), .CP(n2236), .CDN(
        n2162), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n210), .CP(n2249), .CDN(
        n2162), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n210), .CP(n2248), .CDN(
        n2162), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n210), .CP(n2230), .CDN(
        n2162), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n210), .CP(n2234), .CDN(
        n2162), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n210), .CP(n2246), .CDN(
        n2162), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(n210), .CP(n2245), .CDN(
        n2162), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n210), .CP(n2244), .CDN(
        n2162), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n210), .CP(n2243), .CDN(
        n2162), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n210), .CP(n2242), .CDN(
        n2161), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n210), .CP(n2211), .CDN(
        n2161), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n210), .CP(n2252), .CDN(
        n2161), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n210), .CP(n2233), .CDN(
        n2161), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n210), .CP(n2235), .CDN(
        n2161), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n210), .CP(n2253), .CDN(
        n2161), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n210), .CP(n2187), .CDN(
        n2161), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n210), .CP(n2230), .CDN(
        n2161), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n210), .CP(n2255), .CDN(
        n2161), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n210), .CP(n2218), .CDN(
        n2161), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n210), .CP(n2246), .CDN(
        n2161), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n210), .CP(n2207), .CDN(
        n2160), .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n210), .CP(n2237), .CDN(
        n2160), .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n210), .CP(n2243), .CDN(
        n2160), .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n210), .CP(n2237), .CDN(
        n2160), .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n210), .CP(ClockW), .CDN(
        n2160), .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n210), .CP(n2234), .CDN(
        n2160), .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n210), .CP(n2240), .CDN(
        n2160), .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(n209), .CP(ClockW), .CDN(n2154), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n209), .CP(n2233), .CDN(
        n2153), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n209), .CP(n2254), .CDN(
        n2153), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n209), .CP(n2234), .CDN(
        n2153), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(n209), .CP(n2240), .CDN(
        n2153), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n209), .CP(n2248), .CDN(
        n2153), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(n209), .CP(n2194), .CDN(
        n2153), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n209), .CP(n2230), .CDN(
        n2153), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n209), .CP(n2188), .CDN(
        n2153), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n209), .CP(n2253), .CDN(
        n2153), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n209), .CP(n2252), .CDN(
        n2153), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n209), .CP(n2234), .CDN(
        n2153), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n209), .CP(n2238), .CDN(
        n2152), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n209), .CP(n2189), .CDN(
        n2152), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n209), .CP(n2247), .CDN(
        n2152), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n209), .CP(n2251), .CDN(
        n2152), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n209), .CP(n2194), .CDN(
        n2152), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n209), .CP(n2254), .CDN(
        n2152), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n209), .CP(n2226), .CDN(
        n2152), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n209), .CP(n2255), .CDN(
        n2152), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n209), .CP(n2219), .CDN(
        n2152), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n209), .CP(n2233), .CDN(
        n2152), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n209), .CP(n2239), .CDN(
        n2152), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n209), .CP(n2244), .CDN(
        n2151), .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n209), .CP(n2195), .CDN(
        n2151), .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n209), .CP(ClockW), .CDN(
        n2151), .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n209), .CP(n2187), .CDN(
        n2151), .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n209), .CP(n2250), .CDN(
        n2151), .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n209), .CP(n2251), .CDN(
        n2151), .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n209), .CP(n2252), .CDN(
        n2151), .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n2147), .E(n208), .CP(n2188), .CDN(n2150), .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(n208), .CP(n2188), .CDN(
        n2179), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(n208), .CP(n2188), .CDN(
        n2175), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(n208), .CP(n2188), .CDN(
        n2152), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(n208), .CP(n2188), .CDN(
        n2170), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(n208), .CP(n2188), .CDN(
        n2182), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(n208), .CP(n2188), .CDN(
        n2175), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(n208), .CP(n2188), .CDN(
        n2153), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(n208), .CP(n2188), .CDN(
        n2176), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(n208), .CP(n2188), .CDN(
        n2176), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(n208), .CP(n2189), .CDN(
        n2179), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(n208), .CP(n2189), .CDN(
        n2180), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(n208), .CP(n2189), .CDN(
        n2149), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(n208), .CP(n2189), .CDN(
        n2180), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(n208), .CP(n2189), .CDN(
        n2168), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(n208), .CP(n2189), .CDN(
        n2169), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(n208), .CP(n2189), .CDN(
        n2170), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(n208), .CP(n2189), .CDN(
        n2167), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(n208), .CP(n2189), .CDN(
        n2178), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(n208), .CP(n2189), .CDN(
        n2181), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(n208), .CP(n2190), .CDN(
        n2182), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(n208), .CP(n2190), .CDN(
        n2180), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(n208), .CP(n2190), .CDN(
        n2179), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(n208), .CP(n2190), .CDN(
        n2179), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(DataI[6]), .E(n208), .CP(n2190), .CDN(
        n2180), .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(n208), .CP(n2190), .CDN(
        n2181), .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(n208), .CP(n2190), .CDN(
        n2182), .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(n208), .CP(n2191), .CDN(
        n2179), .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(n208), .CP(n2191), .CDN(
        n2180), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(n208), .CP(n2191), .CDN(
        n2173), .Q(\Storage[31][0] ) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(n2290) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(n2289) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(n2288) );
  BUFTD0 \DataO_tri[3]  ( .I(n180), .OE(ChipEna), .Z(n2287) );
  BUFTD0 \DataO_tri[4]  ( .I(n176), .OE(ChipEna), .Z(n2286) );
  BUFTD0 \DataO_tri[5]  ( .I(n247), .OE(ChipEna), .Z(n2285) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(n2284) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(n2283) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(n2282) );
  BUFTD0 \DataO_tri[9]  ( .I(n172), .OE(ChipEna), .Z(n2281) );
  BUFTD0 \DataO_tri[10]  ( .I(n168), .OE(ChipEna), .Z(n2280) );
  BUFTD0 \DataO_tri[11]  ( .I(n245), .OE(ChipEna), .Z(n2279) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(n2278) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(n2277) );
  BUFTD0 \DataO_tri[14]  ( .I(n164), .OE(ChipEna), .Z(n2276) );
  BUFTD0 \DataO_tri[15]  ( .I(n160), .OE(ChipEna), .Z(n2275) );
  BUFTD0 \DataO_tri[16]  ( .I(n243), .OE(ChipEna), .Z(n2274) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(n2273) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(n2272) );
  BUFTD0 \DataO_tri[19]  ( .I(n156), .OE(ChipEna), .Z(n2271) );
  BUFTD0 \DataO_tri[20]  ( .I(n152), .OE(ChipEna), .Z(n2270) );
  BUFTD0 \DataO_tri[21]  ( .I(n241), .OE(ChipEna), .Z(n2269) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(n2268) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(n2267) );
  BUFTD0 \DataO_tri[24]  ( .I(n148), .OE(ChipEna), .Z(n2266) );
  BUFTD0 \DataO_tri[25]  ( .I(n144), .OE(ChipEna), .Z(n2265) );
  BUFTD0 \DataO_tri[26]  ( .I(n140), .OE(ChipEna), .Z(n2264) );
  BUFTD0 \DataO_tri[27]  ( .I(n136), .OE(ChipEna), .Z(n2263) );
  BUFTD0 \DataO_tri[28]  ( .I(n132), .OE(ChipEna), .Z(n2262) );
  BUFTD0 \DataO_tri[29]  ( .I(n128), .OE(ChipEna), .Z(n2261) );
  BUFTD0 \DataO_tri[30]  ( .I(n124), .OE(ChipEna), .Z(n2260) );
  BUFTD0 \DataO_tri[31]  ( .I(n120), .OE(ChipEna), .Z(n2259) );
  EDFCNQD1 Parityr_reg ( .D(n274), .E(n1427), .CP(ClockR), .CDN(n2161), .Q(
        ParityErr) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n7), .E(Read), .CP(ClockR), .CDN(n2156), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n12), .E(n1427), .CP(ClockR), .CDN(n2150), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n351), .E(Read), .CP(ClockR), .CDN(n2183), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n386), .E(n2256), .CP(ClockR), .CDN(n2173), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n17), .E(n1427), .CP(ClockR), .CDN(n2178), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n22), .E(n2256), .CP(ClockR), .CDN(n2149), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n491), .E(n2256), .CP(ClockR), .CDN(n2173), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n27), .E(Read), .CP(ClockR), .CDN(n2174), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n30), .E(Read), .CP(ClockR), .CDN(n2176), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n595), .E(Read), .CP(ClockR), .CDN(n2180), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n631), .E(Read), .CP(ClockR), .CDN(n2178), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n37), .E(n1427), .CP(ClockR), .CDN(n2183), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n42), .E(n2256), .CP(ClockR), .CDN(n2160), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n737), .E(Read), .CP(ClockR), .CDN(n2176), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n46), .E(Read), .CP(ClockR), .CDN(n2185), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n49), .E(Read), .CP(ClockR), .CDN(n2184), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n840), .E(Read), .CP(ClockR), .CDN(n2177), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n879), .E(Read), .CP(ClockR), .CDN(n2159), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n55), .E(Read), .CP(ClockR), .CDN(n2160), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n60), .E(n2256), .CP(ClockR), .CDN(n2167), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n988), .E(n1427), .CP(ClockR), .CDN(n2183), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n1028), .E(n2256), .CP(ClockR), .CDN(n2159), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n1064), .E(n1427), .CP(ClockR), .CDN(n2163), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n1105), .E(n1427), .CP(ClockR), .CDN(n2152), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n90), .E(n2256), .CP(ClockR), .CDN(n2157), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n111), .E(n2256), .CP(ClockR), .CDN(n2178), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n1211), .E(n2256), .CP(ClockR), .CDN(n2161), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n1248), .E(n2256), .CP(ClockR), .CDN(n2178), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n1285), .E(n2256), .CP(ClockR), .CDN(n2155), 
        .Q(DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n117), .E(n2256), .CP(ClockR), .CDN(n2164), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n1357), .E(n2256), .CP(ClockR), .CDN(n2162), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n1391), .E(n1427), .CP(ClockR), .CDN(n2161), 
        .Q(DataOr[0]) );
  EDFCNQD1 Dreadyr_reg ( .D(n1684), .E(n1427), .CP(ClockR), .CDN(n2183), .Q(
        Dreadyr) );
  TIEH U3 ( .Z(n1684) );
  INVD12 U4 ( .I(n263), .ZN(n1) );
  CKNXD0 U5 ( .I(n262), .ZN(n263) );
  CKBD0 U6 ( .CLK(n268), .C(n266) );
  CKNXD0 U7 ( .I(n275), .ZN(n276) );
  INVD0 U8 ( .I(n254), .ZN(n255) );
  CKNXD0 U9 ( .I(n253), .ZN(n254) );
  CKNXD16 U10 ( .I(n206), .ZN(n253) );
  INVD1 U11 ( .I(n1), .ZN(n2) );
  XNR3D0 U12 ( .A1(n775), .A2(n93), .A3(n94), .ZN(n207) );
  BUFFD0 U13 ( .I(n207), .Z(n3) );
  BUFFD0 U14 ( .I(n95), .Z(n4) );
  XOR3D0 U15 ( .A1(n846), .A2(n809), .A3(n3), .Z(n206) );
  XOR3D0 U16 ( .A1(n1070), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D0 U17 ( .A1(n598), .A2(n563), .A3(n4), .Z(n94) );
  INVD0 U23 ( .I(n269), .ZN(n270) );
  CKBXD0 U24 ( .I(n272), .Z(n279) );
  MUX3ND1 U25 ( .I0(n2098), .I1(n2099), .I2(n2100), .S0(N47), .S1(n2115), .ZN(
        n195) );
  BUFFD0 U26 ( .I(n313), .Z(n5) );
  CKBD0 U27 ( .CLK(n195), .C(n8) );
  BUFFD0 U29 ( .I(n5), .Z(n6) );
  BUFFD0 U30 ( .I(n281), .Z(n7) );
  INVD0 U31 ( .I(n312), .ZN(n313) );
  CKBXD0 U32 ( .I(n286), .Z(n287) );
  CKBXD0 U33 ( .I(n8), .Z(n282) );
  BUFFD0 U37 ( .I(n6), .Z(n9) );
  MUX3ND1 U38 ( .I0(n2085), .I1(n2086), .I2(n2087), .S0(n2257), .S1(n2115), 
        .ZN(n194) );
  BUFFD0 U39 ( .I(n348), .Z(n10) );
  BUFFD0 U40 ( .I(n10), .Z(n11) );
  BUFFD0 U41 ( .I(n316), .Z(n12) );
  BUFFD0 U42 ( .I(n194), .Z(n13) );
  INVD0 U43 ( .I(n347), .ZN(n348) );
  CKBXD0 U44 ( .I(n321), .Z(n322) );
  CKBXD0 U45 ( .I(n13), .Z(n317) );
  BUFFD0 U46 ( .I(n11), .Z(n14) );
  INVD16 U47 ( .I(n354), .ZN(n350) );
  INVD0 U48 ( .I(n353), .ZN(n354) );
  CKBXD0 U49 ( .I(n356), .Z(n357) );
  MUX3D0 U50 ( .I0(n2072), .I1(n2073), .I2(n2074), .S0(n2117), .S1(n2115), .Z(
        n205) );
  INVD16 U51 ( .I(n389), .ZN(n385) );
  INVD0 U52 ( .I(n388), .ZN(n389) );
  CKBXD0 U53 ( .I(n391), .Z(n392) );
  MUX3D0 U54 ( .I0(n2059), .I1(n2060), .I2(n2061), .S0(n2117), .S1(n2115), .Z(
        n204) );
  INVD0 U55 ( .I(n15), .ZN(n16) );
  INVD10 U56 ( .I(n193), .ZN(n15) );
  MUX3ND0 U57 ( .I0(n2046), .I1(n2047), .I2(n2048), .S0(n2116), .S1(n2115), 
        .ZN(n193) );
  BUFFD0 U58 ( .I(n421), .Z(n17) );
  BUFFD0 U59 ( .I(n16), .Z(n18) );
  INVD0 U60 ( .I(n452), .ZN(n453) );
  CKBXD0 U61 ( .I(n426), .Z(n427) );
  CKBXD0 U62 ( .I(n18), .Z(n422) );
  BUFFD0 U63 ( .I(n453), .Z(n19) );
  MUX3ND1 U64 ( .I0(n2033), .I1(n2034), .I2(n2035), .S0(N47), .S1(n2115), .ZN(
        n192) );
  BUFFD0 U65 ( .I(n488), .Z(n20) );
  CKBD0 U66 ( .CLK(n192), .C(n23) );
  BUFFD0 U67 ( .I(n20), .Z(n21) );
  BUFFD0 U68 ( .I(n456), .Z(n22) );
  INVD0 U69 ( .I(n487), .ZN(n488) );
  CKBXD0 U70 ( .I(n461), .Z(n462) );
  CKBXD0 U71 ( .I(n23), .Z(n457) );
  BUFFD0 U72 ( .I(n21), .Z(n24) );
  INVD16 U73 ( .I(n494), .ZN(n490) );
  INVD0 U74 ( .I(n493), .ZN(n494) );
  CKBXD0 U75 ( .I(n496), .Z(n497) );
  MUX3D0 U76 ( .I0(n2020), .I1(n2021), .I2(n2022), .S0(n2116), .S1(n2115), .Z(
        n203) );
  MUX3ND1 U77 ( .I0(n2007), .I1(n2008), .I2(n2009), .S0(N47), .S1(n2115), .ZN(
        n191) );
  BUFFD0 U78 ( .I(n558), .Z(n25) );
  CKBD0 U79 ( .CLK(n191), .C(n28) );
  BUFFD0 U80 ( .I(n25), .Z(n26) );
  BUFFD0 U81 ( .I(n526), .Z(n27) );
  INVD0 U82 ( .I(n557), .ZN(n558) );
  CKBXD0 U83 ( .I(n531), .Z(n532) );
  CKBXD0 U84 ( .I(n28), .Z(n527) );
  BUFFD0 U85 ( .I(n26), .Z(n29) );
  BUFFD12 U86 ( .I(n583), .Z(n584) );
  BUFFD0 U87 ( .I(n31), .Z(n30) );
  BUFFD0 U88 ( .I(n33), .Z(n31) );
  BUFFD0 U89 ( .I(n198), .Z(n32) );
  BUFFD0 U90 ( .I(n563), .Z(n33) );
  MUX3D0 U91 ( .I0(n1981), .I1(n1982), .I2(n1983), .S0(n2257), .S1(n2115), .Z(
        n202) );
  BUFFD0 U92 ( .I(n201), .Z(n34) );
  MUX3ND1 U93 ( .I0(n1955), .I1(n1956), .I2(n1957), .S0(N47), .S1(n2115), .ZN(
        n190) );
  BUFFD0 U94 ( .I(n699), .Z(n35) );
  CKBD0 U95 ( .CLK(n190), .C(n38) );
  BUFFD0 U96 ( .I(n35), .Z(n36) );
  BUFFD0 U97 ( .I(n667), .Z(n37) );
  INVD0 U98 ( .I(n698), .ZN(n699) );
  CKBXD0 U99 ( .I(n672), .Z(n673) );
  CKBXD0 U100 ( .I(n38), .Z(n668) );
  BUFFD0 U101 ( .I(n36), .Z(n39) );
  MUX3ND1 U102 ( .I0(n1942), .I1(n1943), .I2(n1944), .S0(N47), .S1(n2258), 
        .ZN(n189) );
  BUFFD0 U103 ( .I(n734), .Z(n40) );
  CKBD0 U104 ( .CLK(n189), .C(n43) );
  BUFFD0 U105 ( .I(n40), .Z(n41) );
  BUFFD0 U106 ( .I(n702), .Z(n42) );
  INVD0 U107 ( .I(n733), .ZN(n734) );
  CKBXD0 U108 ( .I(n707), .Z(n708) );
  CKBXD0 U109 ( .I(n43), .Z(n703) );
  BUFFD0 U110 ( .I(n41), .Z(n44) );
  BUFFD0 U111 ( .I(n200), .Z(n45) );
  BUFFD16 U112 ( .I(n796), .Z(n797) );
  MUX3ND1 U113 ( .I0(n1916), .I1(n1917), .I2(n805), .S0(n2117), .S1(N48), .ZN(
        n197) );
  BUFFD0 U114 ( .I(n48), .Z(n46) );
  BUFFD0 U115 ( .I(n197), .Z(n47) );
  BUFFD0 U116 ( .I(n775), .Z(n48) );
  BUFFD12 U117 ( .I(n829), .Z(n830) );
  BUFFD0 U118 ( .I(n50), .Z(n49) );
  BUFFD0 U119 ( .I(n52), .Z(n50) );
  BUFFD0 U120 ( .I(n196), .Z(n51) );
  BUFFD0 U121 ( .I(n809), .Z(n52) );
  MUX3ND1 U122 ( .I0(n1864), .I1(n1865), .I2(n1866), .S0(n2257), .S1(N48), 
        .ZN(n188) );
  BUFFD0 U123 ( .I(n951), .Z(n53) );
  CKBD0 U124 ( .CLK(n188), .C(n56) );
  BUFFD0 U125 ( .I(n53), .Z(n54) );
  BUFFD0 U126 ( .I(n919), .Z(n55) );
  INVD0 U127 ( .I(n950), .ZN(n951) );
  CKBXD0 U128 ( .I(n924), .Z(n925) );
  CKBXD0 U129 ( .I(n56), .Z(n920) );
  BUFFD0 U130 ( .I(n54), .Z(n57) );
  INVD0 U131 ( .I(n58), .ZN(n59) );
  INVD10 U132 ( .I(n187), .ZN(n58) );
  MUX3ND0 U133 ( .I0(n1851), .I1(n1852), .I2(n1853), .S0(n2116), .S1(n2258), 
        .ZN(n187) );
  BUFFD0 U134 ( .I(n954), .Z(n60) );
  BUFFD0 U135 ( .I(n59), .Z(n61) );
  INVD0 U136 ( .I(n985), .ZN(n986) );
  CKBXD0 U137 ( .I(n959), .Z(n960) );
  CKBXD0 U138 ( .I(n61), .Z(n955) );
  BUFFD0 U139 ( .I(n986), .Z(n62) );
  MUX3ND1 U140 ( .I0(n1825), .I1(n1826), .I2(n63), .S0(n2116), .S1(n2258), 
        .ZN(N72) );
  BUFFD0 U141 ( .I(n1827), .Z(n63) );
  BUFFD10 U142 ( .I(n1129), .Z(n1130) );
  INVD10 U143 ( .I(n199), .ZN(n1103) );
  MUX3D0 U144 ( .I0(n1799), .I1(n1800), .I2(n1139), .S0(n2117), .S1(n2258), 
        .Z(n199) );
  INVD0 U145 ( .I(n64), .ZN(n65) );
  INVD10 U146 ( .I(n186), .ZN(n64) );
  MUX3ND0 U147 ( .I0(n1786), .I1(n1787), .I2(n1788), .S0(n2116), .S1(n2258), 
        .ZN(n186) );
  BUFFD0 U148 ( .I(n1141), .Z(n90) );
  BUFFD0 U149 ( .I(n65), .Z(n92) );
  INVD0 U150 ( .I(n1172), .ZN(n1173) );
  CKBXD0 U151 ( .I(n1146), .Z(n1147) );
  CKBXD0 U152 ( .I(n92), .Z(n1142) );
  BUFFD0 U153 ( .I(n1173), .Z(n107) );
  CKNXD0 U154 ( .I(n109), .ZN(n110) );
  INVD10 U155 ( .I(n185), .ZN(n109) );
  MUX3ND0 U156 ( .I0(n1773), .I1(n1774), .I2(n1775), .S0(n2116), .S1(n2258), 
        .ZN(n185) );
  BUFFD0 U157 ( .I(n1176), .Z(n111) );
  BUFFD0 U158 ( .I(n110), .Z(n112) );
  INVD0 U159 ( .I(n1207), .ZN(n1208) );
  CKBXD0 U160 ( .I(n1181), .Z(n1182) );
  CKBXD0 U161 ( .I(n112), .Z(n1177) );
  BUFFD0 U162 ( .I(n1208), .Z(n113) );
  MUX3ND1 U163 ( .I0(n1747), .I1(n1748), .I2(n114), .S0(n2116), .S1(n2258), 
        .ZN(N78) );
  BUFFD0 U164 ( .I(n1749), .Z(n114) );
  INVD0 U165 ( .I(n115), .ZN(n116) );
  INVD10 U166 ( .I(n184), .ZN(n115) );
  MUX3ND0 U167 ( .I0(n1721), .I1(n1722), .I2(n1723), .S0(n2117), .S1(n2258), 
        .ZN(n184) );
  BUFFD0 U168 ( .I(n1322), .Z(n117) );
  BUFFD0 U169 ( .I(n116), .Z(n118) );
  INVD0 U170 ( .I(n1353), .ZN(n1354) );
  CKBXD0 U171 ( .I(n1327), .Z(n1328) );
  CKBXD0 U172 ( .I(n118), .Z(n1323) );
  BUFFD0 U173 ( .I(n1354), .Z(n119) );
  BUFFD0 U174 ( .I(n122), .Z(n120) );
  BUFFD0 U175 ( .I(n123), .Z(DataO[31]) );
  BUFFD0 U176 ( .I(DataOr[31]), .Z(n122) );
  BUFFD0 U177 ( .I(n1429), .Z(n123) );
  BUFFD0 U178 ( .I(n126), .Z(n124) );
  BUFFD0 U179 ( .I(n127), .Z(DataO[30]) );
  BUFFD0 U180 ( .I(DataOr[30]), .Z(n126) );
  BUFFD0 U181 ( .I(n1437), .Z(n127) );
  BUFFD0 U182 ( .I(n130), .Z(n128) );
  BUFFD0 U183 ( .I(n131), .Z(DataO[29]) );
  BUFFD0 U184 ( .I(DataOr[29]), .Z(n130) );
  BUFFD0 U185 ( .I(n1445), .Z(n131) );
  BUFFD0 U186 ( .I(n134), .Z(n132) );
  BUFFD0 U187 ( .I(n135), .Z(DataO[28]) );
  BUFFD0 U188 ( .I(DataOr[28]), .Z(n134) );
  BUFFD0 U189 ( .I(n1453), .Z(n135) );
  BUFFD0 U190 ( .I(n138), .Z(n136) );
  BUFFD0 U191 ( .I(n139), .Z(DataO[27]) );
  BUFFD0 U192 ( .I(DataOr[27]), .Z(n138) );
  BUFFD0 U193 ( .I(n1461), .Z(n139) );
  BUFFD0 U194 ( .I(n142), .Z(n140) );
  BUFFD0 U195 ( .I(n143), .Z(DataO[26]) );
  BUFFD0 U196 ( .I(DataOr[26]), .Z(n142) );
  BUFFD0 U197 ( .I(n1469), .Z(n143) );
  BUFFD0 U198 ( .I(n146), .Z(n144) );
  BUFFD0 U199 ( .I(n147), .Z(DataO[25]) );
  BUFFD0 U200 ( .I(DataOr[25]), .Z(n146) );
  BUFFD0 U201 ( .I(n1477), .Z(n147) );
  BUFFD0 U202 ( .I(n150), .Z(n148) );
  BUFFD0 U203 ( .I(n151), .Z(DataO[24]) );
  BUFFD0 U204 ( .I(DataOr[24]), .Z(n150) );
  BUFFD0 U205 ( .I(n1485), .Z(n151) );
  BUFFD0 U206 ( .I(n154), .Z(n152) );
  BUFFD0 U207 ( .I(n155), .Z(DataO[20]) );
  BUFFD0 U208 ( .I(DataOr[20]), .Z(n154) );
  BUFFD0 U209 ( .I(n1517), .Z(n155) );
  BUFFD0 U210 ( .I(n158), .Z(n156) );
  BUFFD0 U211 ( .I(n159), .Z(DataO[19]) );
  BUFFD0 U212 ( .I(DataOr[19]), .Z(n158) );
  BUFFD0 U213 ( .I(n1525), .Z(n159) );
  BUFFD0 U214 ( .I(n162), .Z(n160) );
  BUFFD0 U215 ( .I(n163), .Z(DataO[15]) );
  BUFFD0 U216 ( .I(DataOr[15]), .Z(n162) );
  BUFFD0 U217 ( .I(n1557), .Z(n163) );
  BUFFD0 U218 ( .I(n166), .Z(n164) );
  BUFFD0 U219 ( .I(n167), .Z(DataO[14]) );
  BUFFD0 U220 ( .I(DataOr[14]), .Z(n166) );
  BUFFD0 U221 ( .I(n1565), .Z(n167) );
  BUFFD0 U222 ( .I(n170), .Z(n168) );
  BUFFD0 U223 ( .I(n171), .Z(DataO[10]) );
  BUFFD0 U224 ( .I(DataOr[10]), .Z(n170) );
  BUFFD0 U225 ( .I(n1597), .Z(n171) );
  BUFFD0 U226 ( .I(n174), .Z(n172) );
  BUFFD0 U227 ( .I(n175), .Z(DataO[9]) );
  BUFFD0 U228 ( .I(DataOr[9]), .Z(n174) );
  BUFFD0 U229 ( .I(n1605), .Z(n175) );
  BUFFD0 U230 ( .I(n178), .Z(n176) );
  BUFFD0 U231 ( .I(n179), .Z(DataO[4]) );
  BUFFD0 U232 ( .I(DataOr[4]), .Z(n178) );
  BUFFD0 U233 ( .I(n1645), .Z(n179) );
  BUFFD0 U234 ( .I(n182), .Z(n180) );
  BUFFD0 U235 ( .I(n183), .Z(DataO[3]) );
  BUFFD0 U236 ( .I(DataOr[3]), .Z(n182) );
  BUFFD0 U237 ( .I(n1653), .Z(n183) );
  MUX3ND0 U238 ( .I0(n1903), .I1(n1904), .I2(n839), .S0(n2257), .S1(N48), .ZN(
        n196) );
  MUX3ND0 U239 ( .I0(n1994), .I1(n1995), .I2(n593), .S0(N47), .S1(n2115), .ZN(
        n198) );
  MUX3D1 U240 ( .I0(n1929), .I1(n1930), .I2(n1931), .S0(N47), .S1(n2258), .Z(
        n200) );
  MUX3D1 U241 ( .I0(n1968), .I1(n1969), .I2(n1970), .S0(N47), .S1(n2115), .Z(
        n201) );
  INVD1 U242 ( .I(n1659), .ZN(n1656) );
  INVD1 U243 ( .I(n2287), .ZN(n1658) );
  INVD1 U244 ( .I(n1651), .ZN(n1648) );
  INVD1 U245 ( .I(n2286), .ZN(n1650) );
  INVD1 U246 ( .I(n1611), .ZN(n1608) );
  INVD1 U247 ( .I(n2281), .ZN(n1610) );
  INVD1 U248 ( .I(n1603), .ZN(n1600) );
  INVD1 U249 ( .I(n2280), .ZN(n1602) );
  INVD1 U250 ( .I(n1571), .ZN(n1568) );
  INVD1 U251 ( .I(n2276), .ZN(n1570) );
  INVD1 U252 ( .I(n1563), .ZN(n1560) );
  INVD1 U253 ( .I(n2275), .ZN(n1562) );
  INVD1 U254 ( .I(n1531), .ZN(n1528) );
  INVD1 U255 ( .I(n2271), .ZN(n1530) );
  INVD1 U256 ( .I(n1523), .ZN(n1520) );
  INVD1 U257 ( .I(n2270), .ZN(n1522) );
  INVD1 U258 ( .I(n1491), .ZN(n1488) );
  INVD1 U259 ( .I(n2266), .ZN(n1490) );
  INVD1 U260 ( .I(n1483), .ZN(n1480) );
  INVD1 U261 ( .I(n2265), .ZN(n1482) );
  INVD1 U262 ( .I(n1475), .ZN(n1472) );
  INVD1 U263 ( .I(n2264), .ZN(n1474) );
  INVD1 U264 ( .I(n1467), .ZN(n1464) );
  INVD1 U265 ( .I(n2263), .ZN(n1466) );
  INVD1 U266 ( .I(n1459), .ZN(n1456) );
  INVD1 U267 ( .I(n2262), .ZN(n1458) );
  INVD1 U268 ( .I(n1451), .ZN(n1448) );
  INVD1 U269 ( .I(n2261), .ZN(n1450) );
  INVD1 U270 ( .I(n1443), .ZN(n1440) );
  INVD1 U271 ( .I(n2260), .ZN(n1442) );
  INVD1 U272 ( .I(n1435), .ZN(n1432) );
  INVD1 U273 ( .I(n2259), .ZN(n1434) );
  INVD1 U274 ( .I(n1655), .ZN(n1652) );
  INVD1 U275 ( .I(n1657), .ZN(n1654) );
  INVD1 U276 ( .I(n1647), .ZN(n1644) );
  INVD1 U277 ( .I(n1649), .ZN(n1646) );
  INVD1 U278 ( .I(n1607), .ZN(n1604) );
  INVD1 U279 ( .I(n1609), .ZN(n1606) );
  INVD1 U280 ( .I(n1599), .ZN(n1596) );
  INVD1 U281 ( .I(n1601), .ZN(n1598) );
  INVD1 U282 ( .I(n1567), .ZN(n1564) );
  INVD1 U283 ( .I(n1569), .ZN(n1566) );
  INVD1 U284 ( .I(n1559), .ZN(n1556) );
  INVD1 U285 ( .I(n1561), .ZN(n1558) );
  INVD1 U286 ( .I(n1527), .ZN(n1524) );
  INVD1 U287 ( .I(n1529), .ZN(n1526) );
  INVD1 U288 ( .I(n1519), .ZN(n1516) );
  INVD1 U289 ( .I(n1521), .ZN(n1518) );
  INVD1 U290 ( .I(n1487), .ZN(n1484) );
  INVD1 U291 ( .I(n1489), .ZN(n1486) );
  INVD1 U292 ( .I(n1479), .ZN(n1476) );
  INVD1 U293 ( .I(n1481), .ZN(n1478) );
  INVD1 U294 ( .I(n1471), .ZN(n1468) );
  INVD1 U295 ( .I(n1473), .ZN(n1470) );
  INVD1 U296 ( .I(n1463), .ZN(n1460) );
  INVD1 U297 ( .I(n1465), .ZN(n1462) );
  INVD1 U298 ( .I(n1455), .ZN(n1452) );
  INVD1 U299 ( .I(n1457), .ZN(n1454) );
  INVD1 U300 ( .I(n1447), .ZN(n1444) );
  INVD1 U301 ( .I(n1449), .ZN(n1446) );
  INVD1 U302 ( .I(n1439), .ZN(n1436) );
  INVD1 U303 ( .I(n1441), .ZN(n1438) );
  INVD1 U304 ( .I(n1431), .ZN(n1428) );
  INVD1 U305 ( .I(n1433), .ZN(n1430) );
  XNR3D1 U306 ( .A1(n1214), .A2(n1208), .A3(n264), .ZN(n88) );
  INVD1 U307 ( .I(n265), .ZN(n264) );
  NR2D1 U308 ( .A1(n66), .A2(n71), .ZN(n208) );
  NR2D1 U309 ( .A1(n69), .A2(n103), .ZN(n209) );
  NR2D1 U310 ( .A1(n99), .A2(n103), .ZN(n210) );
  NR2D1 U311 ( .A1(n98), .A2(n103), .ZN(n211) );
  NR2D1 U312 ( .A1(n71), .A2(n103), .ZN(n212) );
  NR2D1 U313 ( .A1(n69), .A2(n101), .ZN(n213) );
  NR2D1 U314 ( .A1(n99), .A2(n101), .ZN(n214) );
  NR2D1 U315 ( .A1(n98), .A2(n101), .ZN(n215) );
  NR2D1 U316 ( .A1(n71), .A2(n101), .ZN(n216) );
  NR2D1 U317 ( .A1(n69), .A2(n70), .ZN(n217) );
  NR2D1 U318 ( .A1(n70), .A2(n99), .ZN(n218) );
  NR2D1 U319 ( .A1(n70), .A2(n98), .ZN(n219) );
  NR2D1 U320 ( .A1(n70), .A2(n71), .ZN(n220) );
  NR2D1 U321 ( .A1(n68), .A2(n103), .ZN(n221) );
  NR2D1 U322 ( .A1(n67), .A2(n103), .ZN(n222) );
  NR2D1 U323 ( .A1(n85), .A2(n103), .ZN(n223) );
  NR2D1 U324 ( .A1(n72), .A2(n103), .ZN(n224) );
  NR2D1 U325 ( .A1(n68), .A2(n101), .ZN(n225) );
  NR2D1 U326 ( .A1(n67), .A2(n101), .ZN(n226) );
  NR2D1 U327 ( .A1(n85), .A2(n101), .ZN(n227) );
  NR2D1 U328 ( .A1(n72), .A2(n101), .ZN(n228) );
  NR2D1 U329 ( .A1(n68), .A2(n70), .ZN(n229) );
  NR2D1 U330 ( .A1(n67), .A2(n70), .ZN(n230) );
  NR2D1 U331 ( .A1(n70), .A2(n85), .ZN(n231) );
  NR2D1 U332 ( .A1(n70), .A2(n72), .ZN(n232) );
  NR2D1 U333 ( .A1(n66), .A2(n68), .ZN(n233) );
  NR2D1 U334 ( .A1(n66), .A2(n99), .ZN(n234) );
  NR2D1 U335 ( .A1(n66), .A2(n98), .ZN(n235) );
  NR2D1 U336 ( .A1(n66), .A2(n85), .ZN(n236) );
  NR2D1 U337 ( .A1(n66), .A2(n72), .ZN(n237) );
  NR2D1 U338 ( .A1(n66), .A2(n69), .ZN(n238) );
  NR2D1 U339 ( .A1(n66), .A2(n67), .ZN(n239) );
  CKBD0 U340 ( .CLK(n2256), .C(n1427) );
  CKBD0 U341 ( .CLK(Read), .C(n2256) );
  BUFFD1 U342 ( .I(n2150), .Z(n2148) );
  BUFFD0 U343 ( .I(n108), .Z(n2149) );
  BUFFD0 U344 ( .I(N46), .Z(n2118) );
  BUFFD0 U345 ( .I(N47), .Z(n2257) );
  BUFFD1 U346 ( .I(n2133), .Z(n2136) );
  CKBD0 U347 ( .CLK(n2134), .C(n2135) );
  CKNXD12 U348 ( .I(n1259), .ZN(n1260) );
  CKNXD12 U349 ( .I(n1039), .ZN(n1040) );
  CKNXD12 U350 ( .I(n1247), .ZN(n1248) );
  CKND8 U351 ( .CLK(n1210), .CN(n1211) );
  CKNXD12 U352 ( .I(n1027), .ZN(n1028) );
  BUFFD0 U353 ( .I(n1509), .Z(DataO[21]) );
  BUFFD0 U354 ( .I(DataOr[21]), .Z(n241) );
  BUFFD0 U355 ( .I(n1549), .Z(DataO[16]) );
  BUFFD0 U356 ( .I(DataOr[16]), .Z(n243) );
  BUFFD0 U357 ( .I(n1589), .Z(DataO[11]) );
  BUFFD0 U358 ( .I(DataOr[11]), .Z(n245) );
  BUFFD0 U359 ( .I(n1637), .Z(DataO[5]) );
  BUFFD0 U360 ( .I(DataOr[5]), .Z(n247) );
  BUFFD0 U361 ( .I(N72), .Z(n248) );
  BUFFD0 U362 ( .I(N78), .Z(n249) );
  BUFFD0 U363 ( .I(N77), .Z(n250) );
  CKND12 U364 ( .CLK(N83), .CN(n251) );
  INVD1 U365 ( .I(n251), .ZN(n252) );
  INVD0 U366 ( .I(n256), .ZN(n257) );
  CKNXD16 U367 ( .I(n270), .ZN(n256) );
  CKNXD16 U368 ( .I(n258), .ZN(n259) );
  INVD0 U369 ( .I(n97), .ZN(n258) );
  XOR4D0 U370 ( .A1(n2), .A2(n1031), .A3(n91), .A4(n1173), .Z(n89) );
  INVD0 U371 ( .I(n260), .ZN(n261) );
  CKNXD16 U372 ( .I(n255), .ZN(n260) );
  CKNXD16 U373 ( .I(n266), .ZN(n262) );
  CKBXD0 U374 ( .I(n89), .Z(n265) );
  INVD0 U375 ( .I(n277), .ZN(n278) );
  CKNXD16 U376 ( .I(n267), .ZN(n268) );
  INVD0 U377 ( .I(n276), .ZN(n267) );
  CKNXD16 U378 ( .I(n278), .ZN(n269) );
  CKNXD16 U379 ( .I(n271), .ZN(n272) );
  INVD0 U380 ( .I(n259), .ZN(n271) );
  CKNXD16 U381 ( .I(n273), .ZN(n274) );
  INVD0 U382 ( .I(n252), .ZN(n273) );
  XOR3D0 U383 ( .A1(n1285), .A2(n1105), .A3(n86), .Z(N83) );
  CKNXD16 U384 ( .I(n261), .ZN(n275) );
  CKNXD16 U385 ( .I(n279), .ZN(n277) );
  XNR4D4 U386 ( .A1(n313), .A2(N50), .A3(n354), .A4(n348), .ZN(n97) );
  INVD12 U387 ( .I(n9), .ZN(n280) );
  BUFFD0 U388 ( .I(n311), .Z(n314) );
  INVD0 U389 ( .I(n298), .ZN(n299) );
  INVD0 U390 ( .I(n288), .ZN(n289) );
  INVD1 U391 ( .I(n280), .ZN(n281) );
  INVD0 U392 ( .I(n283), .ZN(n284) );
  CKNXD16 U393 ( .I(n282), .ZN(n283) );
  CKNXD16 U394 ( .I(n285), .ZN(n286) );
  INVD0 U395 ( .I(n284), .ZN(n285) );
  CKNXD16 U396 ( .I(n287), .ZN(n288) );
  CKNXD16 U397 ( .I(n290), .ZN(n291) );
  INVD0 U398 ( .I(n289), .ZN(n290) );
  BUFFD0 U399 ( .I(n291), .Z(n292) );
  INVD0 U400 ( .I(n293), .ZN(n294) );
  CKNXD16 U401 ( .I(n292), .ZN(n293) );
  CKNXD16 U402 ( .I(n295), .ZN(n296) );
  INVD0 U403 ( .I(n294), .ZN(n295) );
  BUFFD0 U404 ( .I(n296), .Z(n297) );
  CKNXD16 U405 ( .I(n297), .ZN(n298) );
  CKNXD16 U406 ( .I(n300), .ZN(n301) );
  INVD0 U407 ( .I(n299), .ZN(n300) );
  BUFFD0 U408 ( .I(n301), .Z(n302) );
  INVD0 U409 ( .I(n303), .ZN(n304) );
  CKNXD16 U410 ( .I(n302), .ZN(n303) );
  CKNXD16 U411 ( .I(n305), .ZN(n306) );
  INVD0 U412 ( .I(n304), .ZN(n305) );
  BUFFD0 U413 ( .I(n306), .Z(n307) );
  INVD0 U414 ( .I(n308), .ZN(n309) );
  CKNXD16 U415 ( .I(n307), .ZN(n308) );
  CKNXD16 U416 ( .I(n310), .ZN(n311) );
  INVD0 U417 ( .I(n309), .ZN(n310) );
  CKNXD16 U418 ( .I(n314), .ZN(n312) );
  INVD12 U419 ( .I(n14), .ZN(n315) );
  BUFFD0 U420 ( .I(n346), .Z(n349) );
  INVD0 U421 ( .I(n333), .ZN(n334) );
  INVD0 U422 ( .I(n323), .ZN(n324) );
  INVD1 U423 ( .I(n315), .ZN(n316) );
  INVD0 U424 ( .I(n318), .ZN(n319) );
  CKNXD16 U425 ( .I(n317), .ZN(n318) );
  CKNXD16 U426 ( .I(n320), .ZN(n321) );
  INVD0 U427 ( .I(n319), .ZN(n320) );
  CKNXD16 U428 ( .I(n322), .ZN(n323) );
  CKNXD16 U429 ( .I(n325), .ZN(n326) );
  INVD0 U430 ( .I(n324), .ZN(n325) );
  BUFFD0 U431 ( .I(n326), .Z(n327) );
  INVD0 U432 ( .I(n328), .ZN(n329) );
  CKNXD16 U433 ( .I(n327), .ZN(n328) );
  CKNXD16 U434 ( .I(n330), .ZN(n331) );
  INVD0 U435 ( .I(n329), .ZN(n330) );
  BUFFD0 U436 ( .I(n331), .Z(n332) );
  CKNXD16 U437 ( .I(n332), .ZN(n333) );
  CKNXD16 U438 ( .I(n335), .ZN(n336) );
  INVD0 U439 ( .I(n334), .ZN(n335) );
  BUFFD0 U440 ( .I(n336), .Z(n337) );
  INVD0 U441 ( .I(n338), .ZN(n339) );
  CKNXD16 U442 ( .I(n337), .ZN(n338) );
  CKNXD16 U443 ( .I(n340), .ZN(n341) );
  INVD0 U444 ( .I(n339), .ZN(n340) );
  BUFFD0 U445 ( .I(n341), .Z(n342) );
  INVD0 U446 ( .I(n343), .ZN(n344) );
  CKNXD16 U447 ( .I(n342), .ZN(n343) );
  CKNXD16 U448 ( .I(n345), .ZN(n346) );
  INVD0 U449 ( .I(n344), .ZN(n345) );
  CKNXD16 U450 ( .I(n349), .ZN(n347) );
  INVD0 U451 ( .I(n382), .ZN(n383) );
  INVD0 U452 ( .I(n363), .ZN(n364) );
  INVD0 U453 ( .I(n358), .ZN(n359) );
  INVD1 U454 ( .I(n350), .ZN(n351) );
  CKNXD16 U455 ( .I(n205), .ZN(n352) );
  CKNXD16 U456 ( .I(n383), .ZN(n353) );
  BUFFD0 U457 ( .I(n381), .Z(n384) );
  INVD0 U458 ( .I(n368), .ZN(n369) );
  CKNXD16 U459 ( .I(n355), .ZN(n356) );
  INVD0 U460 ( .I(n352), .ZN(n355) );
  CKNXD16 U461 ( .I(n357), .ZN(n358) );
  CKNXD16 U462 ( .I(n360), .ZN(n361) );
  INVD0 U463 ( .I(n359), .ZN(n360) );
  BUFFD0 U464 ( .I(n361), .Z(n362) );
  CKNXD16 U465 ( .I(n362), .ZN(n363) );
  CKNXD16 U466 ( .I(n365), .ZN(n366) );
  INVD0 U467 ( .I(n364), .ZN(n365) );
  BUFFD0 U468 ( .I(n366), .Z(n367) );
  CKNXD16 U469 ( .I(n367), .ZN(n368) );
  CKNXD16 U470 ( .I(n370), .ZN(n371) );
  INVD0 U471 ( .I(n369), .ZN(n370) );
  BUFFD0 U472 ( .I(n371), .Z(n372) );
  INVD0 U473 ( .I(n373), .ZN(n374) );
  CKNXD16 U474 ( .I(n372), .ZN(n373) );
  CKNXD16 U475 ( .I(n375), .ZN(n376) );
  INVD0 U476 ( .I(n374), .ZN(n375) );
  BUFFD0 U477 ( .I(n376), .Z(n377) );
  INVD0 U478 ( .I(n378), .ZN(n379) );
  CKNXD16 U479 ( .I(n377), .ZN(n378) );
  CKNXD16 U480 ( .I(n380), .ZN(n381) );
  INVD0 U481 ( .I(n379), .ZN(n380) );
  CKNXD16 U482 ( .I(n384), .ZN(n382) );
  INVD0 U483 ( .I(n417), .ZN(n418) );
  INVD0 U484 ( .I(n398), .ZN(n399) );
  INVD0 U485 ( .I(n393), .ZN(n394) );
  INVD1 U486 ( .I(n385), .ZN(n386) );
  CKNXD16 U487 ( .I(n204), .ZN(n387) );
  CKNXD16 U488 ( .I(n418), .ZN(n388) );
  BUFFD0 U489 ( .I(n416), .Z(n419) );
  INVD0 U490 ( .I(n403), .ZN(n404) );
  CKNXD16 U491 ( .I(n390), .ZN(n391) );
  INVD0 U492 ( .I(n387), .ZN(n390) );
  CKNXD16 U493 ( .I(n392), .ZN(n393) );
  CKNXD16 U494 ( .I(n395), .ZN(n396) );
  INVD0 U495 ( .I(n394), .ZN(n395) );
  BUFFD0 U496 ( .I(n396), .Z(n397) );
  CKNXD16 U497 ( .I(n397), .ZN(n398) );
  CKNXD16 U498 ( .I(n400), .ZN(n401) );
  INVD0 U499 ( .I(n399), .ZN(n400) );
  BUFFD0 U500 ( .I(n401), .Z(n402) );
  CKNXD16 U501 ( .I(n402), .ZN(n403) );
  CKNXD16 U502 ( .I(n405), .ZN(n406) );
  INVD0 U503 ( .I(n404), .ZN(n405) );
  BUFFD0 U504 ( .I(n406), .Z(n407) );
  INVD0 U505 ( .I(n408), .ZN(n409) );
  CKNXD16 U506 ( .I(n407), .ZN(n408) );
  CKNXD16 U507 ( .I(n410), .ZN(n411) );
  INVD0 U508 ( .I(n409), .ZN(n410) );
  BUFFD0 U509 ( .I(n411), .Z(n412) );
  INVD0 U510 ( .I(n413), .ZN(n414) );
  CKNXD16 U511 ( .I(n412), .ZN(n413) );
  CKNXD16 U512 ( .I(n415), .ZN(n416) );
  INVD0 U513 ( .I(n414), .ZN(n415) );
  CKNXD16 U514 ( .I(n419), .ZN(n417) );
  INVD12 U515 ( .I(n19), .ZN(n420) );
  BUFFD0 U516 ( .I(n451), .Z(n454) );
  INVD0 U517 ( .I(n438), .ZN(n439) );
  INVD0 U518 ( .I(n428), .ZN(n429) );
  INVD1 U519 ( .I(n420), .ZN(n421) );
  INVD0 U520 ( .I(n423), .ZN(n424) );
  CKNXD16 U521 ( .I(n422), .ZN(n423) );
  CKNXD16 U522 ( .I(n425), .ZN(n426) );
  INVD0 U523 ( .I(n424), .ZN(n425) );
  CKNXD16 U524 ( .I(n427), .ZN(n428) );
  CKNXD16 U525 ( .I(n430), .ZN(n431) );
  INVD0 U526 ( .I(n429), .ZN(n430) );
  BUFFD0 U527 ( .I(n431), .Z(n432) );
  INVD0 U528 ( .I(n433), .ZN(n434) );
  CKNXD16 U529 ( .I(n432), .ZN(n433) );
  CKNXD16 U530 ( .I(n435), .ZN(n436) );
  INVD0 U531 ( .I(n434), .ZN(n435) );
  BUFFD0 U532 ( .I(n436), .Z(n437) );
  CKNXD16 U533 ( .I(n437), .ZN(n438) );
  CKNXD16 U534 ( .I(n440), .ZN(n441) );
  INVD0 U535 ( .I(n439), .ZN(n440) );
  BUFFD0 U536 ( .I(n441), .Z(n442) );
  INVD0 U537 ( .I(n443), .ZN(n444) );
  CKNXD16 U538 ( .I(n442), .ZN(n443) );
  CKNXD16 U539 ( .I(n445), .ZN(n446) );
  INVD0 U540 ( .I(n444), .ZN(n445) );
  BUFFD0 U541 ( .I(n446), .Z(n447) );
  INVD0 U542 ( .I(n448), .ZN(n449) );
  CKNXD16 U543 ( .I(n447), .ZN(n448) );
  CKNXD16 U544 ( .I(n450), .ZN(n451) );
  INVD0 U545 ( .I(n449), .ZN(n450) );
  CKNXD16 U546 ( .I(n454), .ZN(n452) );
  INVD12 U547 ( .I(n24), .ZN(n455) );
  BUFFD0 U548 ( .I(n486), .Z(n489) );
  INVD0 U549 ( .I(n473), .ZN(n474) );
  INVD0 U550 ( .I(n463), .ZN(n464) );
  INVD1 U551 ( .I(n455), .ZN(n456) );
  INVD0 U552 ( .I(n458), .ZN(n459) );
  CKNXD16 U553 ( .I(n457), .ZN(n458) );
  CKNXD16 U554 ( .I(n460), .ZN(n461) );
  INVD0 U555 ( .I(n459), .ZN(n460) );
  CKNXD16 U556 ( .I(n462), .ZN(n463) );
  CKNXD16 U557 ( .I(n465), .ZN(n466) );
  INVD0 U558 ( .I(n464), .ZN(n465) );
  BUFFD0 U559 ( .I(n466), .Z(n467) );
  INVD0 U560 ( .I(n468), .ZN(n469) );
  CKNXD16 U561 ( .I(n467), .ZN(n468) );
  CKNXD16 U562 ( .I(n470), .ZN(n471) );
  INVD0 U563 ( .I(n469), .ZN(n470) );
  BUFFD0 U564 ( .I(n471), .Z(n472) );
  CKNXD16 U565 ( .I(n472), .ZN(n473) );
  CKNXD16 U566 ( .I(n475), .ZN(n476) );
  INVD0 U567 ( .I(n474), .ZN(n475) );
  BUFFD0 U568 ( .I(n476), .Z(n477) );
  INVD0 U569 ( .I(n478), .ZN(n479) );
  CKNXD16 U570 ( .I(n477), .ZN(n478) );
  CKNXD16 U571 ( .I(n480), .ZN(n481) );
  INVD0 U572 ( .I(n479), .ZN(n480) );
  BUFFD0 U573 ( .I(n481), .Z(n482) );
  INVD0 U574 ( .I(n483), .ZN(n484) );
  CKNXD16 U575 ( .I(n482), .ZN(n483) );
  CKNXD16 U576 ( .I(n485), .ZN(n486) );
  INVD0 U577 ( .I(n484), .ZN(n485) );
  CKNXD16 U578 ( .I(n489), .ZN(n487) );
  INVD0 U579 ( .I(n522), .ZN(n523) );
  INVD0 U580 ( .I(n503), .ZN(n504) );
  INVD0 U581 ( .I(n498), .ZN(n499) );
  INVD1 U582 ( .I(n490), .ZN(n491) );
  CKNXD16 U583 ( .I(n203), .ZN(n492) );
  CKNXD16 U584 ( .I(n523), .ZN(n493) );
  BUFFD0 U585 ( .I(n521), .Z(n524) );
  INVD0 U586 ( .I(n508), .ZN(n509) );
  CKNXD16 U587 ( .I(n495), .ZN(n496) );
  INVD0 U588 ( .I(n492), .ZN(n495) );
  CKNXD16 U589 ( .I(n497), .ZN(n498) );
  CKNXD16 U590 ( .I(n500), .ZN(n501) );
  INVD0 U591 ( .I(n499), .ZN(n500) );
  BUFFD0 U592 ( .I(n501), .Z(n502) );
  CKNXD16 U593 ( .I(n502), .ZN(n503) );
  CKNXD16 U594 ( .I(n505), .ZN(n506) );
  INVD0 U595 ( .I(n504), .ZN(n505) );
  BUFFD0 U596 ( .I(n506), .Z(n507) );
  CKNXD16 U597 ( .I(n507), .ZN(n508) );
  CKNXD16 U598 ( .I(n510), .ZN(n511) );
  INVD0 U599 ( .I(n509), .ZN(n510) );
  BUFFD0 U600 ( .I(n511), .Z(n512) );
  INVD0 U601 ( .I(n513), .ZN(n514) );
  CKNXD16 U602 ( .I(n512), .ZN(n513) );
  CKNXD16 U603 ( .I(n515), .ZN(n516) );
  INVD0 U604 ( .I(n514), .ZN(n515) );
  BUFFD0 U605 ( .I(n516), .Z(n517) );
  INVD0 U606 ( .I(n518), .ZN(n519) );
  CKNXD16 U607 ( .I(n517), .ZN(n518) );
  CKNXD16 U608 ( .I(n520), .ZN(n521) );
  INVD0 U609 ( .I(n519), .ZN(n520) );
  CKNXD16 U610 ( .I(n524), .ZN(n522) );
  INVD12 U611 ( .I(n29), .ZN(n525) );
  BUFFD0 U612 ( .I(n556), .Z(n559) );
  INVD0 U613 ( .I(n543), .ZN(n544) );
  INVD0 U614 ( .I(n533), .ZN(n534) );
  INVD1 U615 ( .I(n525), .ZN(n526) );
  INVD0 U616 ( .I(n528), .ZN(n529) );
  CKNXD16 U617 ( .I(n527), .ZN(n528) );
  CKNXD16 U618 ( .I(n530), .ZN(n531) );
  INVD0 U619 ( .I(n529), .ZN(n530) );
  CKNXD16 U620 ( .I(n532), .ZN(n533) );
  CKNXD16 U621 ( .I(n535), .ZN(n536) );
  INVD0 U622 ( .I(n534), .ZN(n535) );
  BUFFD0 U623 ( .I(n536), .Z(n537) );
  INVD0 U624 ( .I(n538), .ZN(n539) );
  CKNXD16 U625 ( .I(n537), .ZN(n538) );
  CKNXD16 U626 ( .I(n540), .ZN(n541) );
  INVD0 U627 ( .I(n539), .ZN(n540) );
  BUFFD0 U628 ( .I(n541), .Z(n542) );
  CKNXD16 U629 ( .I(n542), .ZN(n543) );
  CKNXD16 U630 ( .I(n545), .ZN(n546) );
  INVD0 U631 ( .I(n544), .ZN(n545) );
  BUFFD0 U632 ( .I(n546), .Z(n547) );
  INVD0 U633 ( .I(n548), .ZN(n549) );
  CKNXD16 U634 ( .I(n547), .ZN(n548) );
  CKNXD16 U635 ( .I(n550), .ZN(n551) );
  INVD0 U636 ( .I(n549), .ZN(n550) );
  BUFFD0 U637 ( .I(n551), .Z(n552) );
  INVD0 U638 ( .I(n553), .ZN(n554) );
  CKNXD16 U639 ( .I(n552), .ZN(n553) );
  CKNXD16 U640 ( .I(n555), .ZN(n556) );
  INVD0 U641 ( .I(n554), .ZN(n555) );
  CKNXD16 U642 ( .I(n559), .ZN(n557) );
  CKNXD0 U643 ( .I(n562), .ZN(n563) );
  INVD0 U644 ( .I(n566), .ZN(n567) );
  CKNXD16 U645 ( .I(n560), .ZN(n561) );
  INVD0 U646 ( .I(n32), .ZN(n560) );
  CKNXD16 U647 ( .I(n567), .ZN(n562) );
  INVD0 U648 ( .I(n570), .ZN(n571) );
  CKNXD16 U649 ( .I(n564), .ZN(n565) );
  INVD0 U650 ( .I(n561), .ZN(n564) );
  CKNXD16 U651 ( .I(n571), .ZN(n566) );
  INVD0 U652 ( .I(n572), .ZN(n573) );
  CKNXD16 U653 ( .I(n568), .ZN(n569) );
  INVD0 U654 ( .I(n565), .ZN(n568) );
  CKNXD16 U655 ( .I(n573), .ZN(n570) );
  CKNXD16 U656 ( .I(n574), .ZN(n572) );
  CKNXD0 U657 ( .I(n582), .ZN(n583) );
  CKNXD16 U658 ( .I(n575), .ZN(n576) );
  INVD0 U659 ( .I(n578), .ZN(n575) );
  INVD0 U660 ( .I(n577), .ZN(n578) );
  INVD0 U661 ( .I(n590), .ZN(n591) );
  BUFFD0 U662 ( .I(n576), .Z(n574) );
  CKNXD16 U663 ( .I(n585), .ZN(n577) );
  CKNXD16 U664 ( .I(n579), .ZN(n580) );
  INVD0 U665 ( .I(n569), .ZN(n579) );
  BUFFD0 U666 ( .I(n580), .Z(n581) );
  CKNXD16 U667 ( .I(n581), .ZN(n582) );
  CKNXD16 U668 ( .I(n586), .ZN(n587) );
  INVD0 U669 ( .I(n591), .ZN(n586) );
  BUFFD0 U670 ( .I(n587), .Z(n585) );
  BUFFD0 U671 ( .I(n589), .Z(n592) );
  CKNXD16 U672 ( .I(n588), .ZN(n589) );
  INVD0 U673 ( .I(n584), .ZN(n588) );
  CKNXD16 U674 ( .I(n592), .ZN(n590) );
  BUFFD0 U675 ( .I(n1996), .Z(n593) );
  INVD8 U676 ( .I(n597), .ZN(n594) );
  INVD1 U677 ( .I(n594), .ZN(n595) );
  INVD0 U678 ( .I(n596), .ZN(n597) );
  CKNXD16 U679 ( .I(n598), .ZN(n596) );
  CKBXD0 U680 ( .I(n601), .Z(n602) );
  CKNXD16 U681 ( .I(n599), .ZN(n600) );
  INVD0 U682 ( .I(n628), .ZN(n599) );
  INVD0 U683 ( .I(n627), .ZN(n628) );
  INVD0 U684 ( .I(n608), .ZN(n609) );
  INVD0 U685 ( .I(n603), .ZN(n604) );
  BUFFD0 U686 ( .I(n600), .Z(n598) );
  BUFFD0 U687 ( .I(n626), .Z(n629) );
  INVD0 U688 ( .I(n613), .ZN(n614) );
  CKNXD16 U689 ( .I(n202), .ZN(n601) );
  CKNXD16 U690 ( .I(n602), .ZN(n603) );
  CKNXD16 U691 ( .I(n605), .ZN(n606) );
  INVD0 U692 ( .I(n604), .ZN(n605) );
  BUFFD0 U693 ( .I(n606), .Z(n607) );
  CKNXD16 U694 ( .I(n607), .ZN(n608) );
  CKNXD16 U695 ( .I(n610), .ZN(n611) );
  INVD0 U696 ( .I(n609), .ZN(n610) );
  BUFFD0 U697 ( .I(n611), .Z(n612) );
  CKNXD16 U698 ( .I(n612), .ZN(n613) );
  CKNXD16 U699 ( .I(n615), .ZN(n616) );
  INVD0 U700 ( .I(n614), .ZN(n615) );
  BUFFD0 U701 ( .I(n616), .Z(n617) );
  INVD0 U702 ( .I(n618), .ZN(n619) );
  CKNXD16 U703 ( .I(n617), .ZN(n618) );
  CKNXD16 U704 ( .I(n620), .ZN(n621) );
  INVD0 U705 ( .I(n619), .ZN(n620) );
  BUFFD0 U706 ( .I(n621), .Z(n622) );
  INVD0 U707 ( .I(n623), .ZN(n624) );
  CKNXD16 U708 ( .I(n622), .ZN(n623) );
  CKNXD16 U709 ( .I(n625), .ZN(n626) );
  INVD0 U710 ( .I(n624), .ZN(n625) );
  CKNXD16 U711 ( .I(n629), .ZN(n627) );
  INVD8 U712 ( .I(n633), .ZN(n630) );
  INVD1 U713 ( .I(n630), .ZN(n631) );
  INVD0 U714 ( .I(n632), .ZN(n633) );
  CKNXD16 U715 ( .I(n634), .ZN(n632) );
  CKBXD0 U716 ( .I(n637), .Z(n638) );
  CKNXD16 U717 ( .I(n635), .ZN(n636) );
  INVD0 U718 ( .I(n664), .ZN(n635) );
  INVD0 U719 ( .I(n663), .ZN(n664) );
  INVD0 U720 ( .I(n644), .ZN(n645) );
  INVD0 U721 ( .I(n639), .ZN(n640) );
  BUFFD0 U722 ( .I(n636), .Z(n634) );
  BUFFD0 U723 ( .I(n662), .Z(n665) );
  INVD0 U724 ( .I(n649), .ZN(n650) );
  CKNXD16 U725 ( .I(n34), .ZN(n637) );
  CKNXD16 U726 ( .I(n638), .ZN(n639) );
  CKNXD16 U727 ( .I(n641), .ZN(n642) );
  INVD0 U728 ( .I(n640), .ZN(n641) );
  BUFFD0 U729 ( .I(n642), .Z(n643) );
  CKNXD16 U730 ( .I(n643), .ZN(n644) );
  CKNXD16 U731 ( .I(n646), .ZN(n647) );
  INVD0 U732 ( .I(n645), .ZN(n646) );
  BUFFD0 U733 ( .I(n647), .Z(n648) );
  CKNXD16 U734 ( .I(n648), .ZN(n649) );
  CKNXD16 U735 ( .I(n651), .ZN(n652) );
  INVD0 U736 ( .I(n650), .ZN(n651) );
  BUFFD0 U737 ( .I(n652), .Z(n653) );
  INVD0 U738 ( .I(n654), .ZN(n655) );
  CKNXD16 U739 ( .I(n653), .ZN(n654) );
  CKNXD16 U740 ( .I(n656), .ZN(n657) );
  INVD0 U741 ( .I(n655), .ZN(n656) );
  BUFFD0 U742 ( .I(n657), .Z(n658) );
  INVD0 U743 ( .I(n659), .ZN(n660) );
  CKNXD16 U744 ( .I(n658), .ZN(n659) );
  CKNXD16 U745 ( .I(n661), .ZN(n662) );
  INVD0 U746 ( .I(n660), .ZN(n661) );
  CKNXD16 U747 ( .I(n665), .ZN(n663) );
  INVD12 U748 ( .I(n39), .ZN(n666) );
  BUFFD0 U749 ( .I(n697), .Z(n700) );
  INVD0 U750 ( .I(n684), .ZN(n685) );
  INVD0 U751 ( .I(n674), .ZN(n675) );
  INVD1 U752 ( .I(n666), .ZN(n667) );
  INVD0 U753 ( .I(n669), .ZN(n670) );
  CKNXD16 U754 ( .I(n668), .ZN(n669) );
  CKNXD16 U755 ( .I(n671), .ZN(n672) );
  INVD0 U756 ( .I(n670), .ZN(n671) );
  CKNXD16 U757 ( .I(n673), .ZN(n674) );
  CKNXD16 U758 ( .I(n676), .ZN(n677) );
  INVD0 U759 ( .I(n675), .ZN(n676) );
  BUFFD0 U760 ( .I(n677), .Z(n678) );
  INVD0 U761 ( .I(n679), .ZN(n680) );
  CKNXD16 U762 ( .I(n678), .ZN(n679) );
  CKNXD16 U763 ( .I(n681), .ZN(n682) );
  INVD0 U764 ( .I(n680), .ZN(n681) );
  BUFFD0 U765 ( .I(n682), .Z(n683) );
  CKNXD16 U766 ( .I(n683), .ZN(n684) );
  CKNXD16 U767 ( .I(n686), .ZN(n687) );
  INVD0 U768 ( .I(n685), .ZN(n686) );
  BUFFD0 U769 ( .I(n687), .Z(n688) );
  INVD0 U770 ( .I(n689), .ZN(n690) );
  CKNXD16 U771 ( .I(n688), .ZN(n689) );
  CKNXD16 U772 ( .I(n691), .ZN(n692) );
  INVD0 U773 ( .I(n690), .ZN(n691) );
  BUFFD0 U774 ( .I(n692), .Z(n693) );
  INVD0 U775 ( .I(n694), .ZN(n695) );
  CKNXD16 U776 ( .I(n693), .ZN(n694) );
  CKNXD16 U777 ( .I(n696), .ZN(n697) );
  INVD0 U778 ( .I(n695), .ZN(n696) );
  CKNXD16 U779 ( .I(n700), .ZN(n698) );
  INVD12 U780 ( .I(n44), .ZN(n701) );
  BUFFD0 U781 ( .I(n732), .Z(n735) );
  INVD0 U782 ( .I(n719), .ZN(n720) );
  INVD0 U783 ( .I(n709), .ZN(n710) );
  INVD1 U784 ( .I(n701), .ZN(n702) );
  INVD0 U785 ( .I(n704), .ZN(n705) );
  CKNXD16 U786 ( .I(n703), .ZN(n704) );
  CKNXD16 U787 ( .I(n706), .ZN(n707) );
  INVD0 U788 ( .I(n705), .ZN(n706) );
  CKNXD16 U789 ( .I(n708), .ZN(n709) );
  CKNXD16 U790 ( .I(n711), .ZN(n712) );
  INVD0 U791 ( .I(n710), .ZN(n711) );
  BUFFD0 U792 ( .I(n712), .Z(n713) );
  INVD0 U793 ( .I(n714), .ZN(n715) );
  CKNXD16 U794 ( .I(n713), .ZN(n714) );
  CKNXD16 U795 ( .I(n716), .ZN(n717) );
  INVD0 U796 ( .I(n715), .ZN(n716) );
  BUFFD0 U797 ( .I(n717), .Z(n718) );
  CKNXD16 U798 ( .I(n718), .ZN(n719) );
  CKNXD16 U799 ( .I(n721), .ZN(n722) );
  INVD0 U800 ( .I(n720), .ZN(n721) );
  BUFFD0 U801 ( .I(n722), .Z(n723) );
  INVD0 U802 ( .I(n724), .ZN(n725) );
  CKNXD16 U803 ( .I(n723), .ZN(n724) );
  CKNXD16 U804 ( .I(n726), .ZN(n727) );
  INVD0 U805 ( .I(n725), .ZN(n726) );
  BUFFD0 U806 ( .I(n727), .Z(n728) );
  INVD0 U807 ( .I(n729), .ZN(n730) );
  CKNXD16 U808 ( .I(n728), .ZN(n729) );
  CKNXD16 U809 ( .I(n731), .ZN(n732) );
  INVD0 U810 ( .I(n730), .ZN(n731) );
  CKNXD16 U811 ( .I(n735), .ZN(n733) );
  INVD8 U812 ( .I(n739), .ZN(n736) );
  INVD1 U813 ( .I(n736), .ZN(n737) );
  INVD0 U814 ( .I(n738), .ZN(n739) );
  CKNXD16 U815 ( .I(n740), .ZN(n738) );
  CKBXD0 U816 ( .I(n743), .Z(n744) );
  CKNXD16 U817 ( .I(n741), .ZN(n742) );
  INVD0 U818 ( .I(n770), .ZN(n741) );
  INVD0 U819 ( .I(n769), .ZN(n770) );
  INVD0 U820 ( .I(n750), .ZN(n751) );
  INVD0 U821 ( .I(n745), .ZN(n746) );
  BUFFD0 U822 ( .I(n742), .Z(n740) );
  BUFFD0 U823 ( .I(n768), .Z(n771) );
  INVD0 U824 ( .I(n755), .ZN(n756) );
  CKNXD16 U825 ( .I(n45), .ZN(n743) );
  CKNXD16 U826 ( .I(n744), .ZN(n745) );
  CKNXD16 U827 ( .I(n747), .ZN(n748) );
  INVD0 U828 ( .I(n746), .ZN(n747) );
  BUFFD0 U829 ( .I(n748), .Z(n749) );
  CKNXD16 U830 ( .I(n749), .ZN(n750) );
  CKNXD16 U831 ( .I(n752), .ZN(n753) );
  INVD0 U832 ( .I(n751), .ZN(n752) );
  BUFFD0 U833 ( .I(n753), .Z(n754) );
  CKNXD16 U834 ( .I(n754), .ZN(n755) );
  CKNXD16 U835 ( .I(n757), .ZN(n758) );
  INVD0 U836 ( .I(n756), .ZN(n757) );
  BUFFD0 U837 ( .I(n758), .Z(n759) );
  INVD0 U838 ( .I(n760), .ZN(n761) );
  CKNXD16 U839 ( .I(n759), .ZN(n760) );
  CKNXD16 U840 ( .I(n762), .ZN(n763) );
  INVD0 U841 ( .I(n761), .ZN(n762) );
  BUFFD0 U842 ( .I(n763), .Z(n764) );
  INVD0 U843 ( .I(n765), .ZN(n766) );
  CKNXD16 U844 ( .I(n764), .ZN(n765) );
  CKNXD16 U845 ( .I(n767), .ZN(n768) );
  INVD0 U846 ( .I(n766), .ZN(n767) );
  CKNXD16 U847 ( .I(n771), .ZN(n769) );
  CKNXD0 U848 ( .I(n774), .ZN(n775) );
  INVD0 U849 ( .I(n778), .ZN(n779) );
  CKNXD16 U850 ( .I(n772), .ZN(n773) );
  INVD0 U851 ( .I(n47), .ZN(n772) );
  CKNXD16 U852 ( .I(n779), .ZN(n774) );
  INVD0 U853 ( .I(n782), .ZN(n783) );
  CKNXD16 U854 ( .I(n776), .ZN(n777) );
  INVD0 U855 ( .I(n773), .ZN(n776) );
  CKNXD16 U856 ( .I(n783), .ZN(n778) );
  INVD0 U857 ( .I(n784), .ZN(n785) );
  CKNXD16 U858 ( .I(n780), .ZN(n781) );
  INVD0 U859 ( .I(n777), .ZN(n780) );
  CKNXD16 U860 ( .I(n785), .ZN(n782) );
  CKNXD16 U861 ( .I(n786), .ZN(n784) );
  CKNXD0 U862 ( .I(n795), .ZN(n796) );
  CKNXD16 U863 ( .I(n787), .ZN(n788) );
  INVD0 U864 ( .I(n790), .ZN(n787) );
  INVD0 U865 ( .I(n789), .ZN(n790) );
  INVD0 U866 ( .I(n802), .ZN(n803) );
  BUFFD0 U867 ( .I(n788), .Z(n786) );
  CKNXD16 U868 ( .I(n791), .ZN(n789) );
  BUFFD0 U869 ( .I(n793), .Z(n791) );
  CKNXD16 U870 ( .I(n792), .ZN(n793) );
  INVD0 U871 ( .I(n799), .ZN(n792) );
  BUFFD0 U872 ( .I(n781), .Z(n794) );
  CKNXD16 U873 ( .I(n794), .ZN(n795) );
  CKNXD16 U874 ( .I(n798), .ZN(n799) );
  INVD0 U875 ( .I(n803), .ZN(n798) );
  BUFFD0 U876 ( .I(n801), .Z(n804) );
  CKNXD16 U877 ( .I(n800), .ZN(n801) );
  INVD0 U878 ( .I(n797), .ZN(n800) );
  CKNXD16 U879 ( .I(n804), .ZN(n802) );
  BUFFD0 U880 ( .I(n1918), .Z(n805) );
  CKNXD0 U881 ( .I(n808), .ZN(n809) );
  INVD0 U882 ( .I(n812), .ZN(n813) );
  CKNXD16 U883 ( .I(n806), .ZN(n807) );
  INVD0 U884 ( .I(n51), .ZN(n806) );
  CKNXD16 U885 ( .I(n813), .ZN(n808) );
  INVD0 U886 ( .I(n816), .ZN(n817) );
  CKNXD16 U887 ( .I(n810), .ZN(n811) );
  INVD0 U888 ( .I(n807), .ZN(n810) );
  CKNXD16 U889 ( .I(n817), .ZN(n812) );
  INVD0 U890 ( .I(n818), .ZN(n819) );
  CKNXD16 U891 ( .I(n814), .ZN(n815) );
  INVD0 U892 ( .I(n811), .ZN(n814) );
  CKNXD16 U893 ( .I(n819), .ZN(n816) );
  CKNXD16 U894 ( .I(n820), .ZN(n818) );
  CKNXD0 U895 ( .I(n828), .ZN(n829) );
  CKNXD16 U896 ( .I(n821), .ZN(n822) );
  INVD0 U897 ( .I(n824), .ZN(n821) );
  INVD0 U898 ( .I(n823), .ZN(n824) );
  INVD0 U899 ( .I(n836), .ZN(n837) );
  BUFFD0 U900 ( .I(n822), .Z(n820) );
  CKNXD16 U901 ( .I(n831), .ZN(n823) );
  CKNXD16 U902 ( .I(n825), .ZN(n826) );
  INVD0 U903 ( .I(n815), .ZN(n825) );
  BUFFD0 U904 ( .I(n826), .Z(n827) );
  CKNXD16 U905 ( .I(n827), .ZN(n828) );
  CKNXD16 U906 ( .I(n832), .ZN(n833) );
  INVD0 U907 ( .I(n837), .ZN(n832) );
  BUFFD0 U908 ( .I(n833), .Z(n831) );
  BUFFD0 U909 ( .I(n835), .Z(n838) );
  CKNXD16 U910 ( .I(n834), .ZN(n835) );
  INVD0 U911 ( .I(n830), .ZN(n834) );
  CKNXD16 U912 ( .I(n838), .ZN(n836) );
  BUFFD0 U913 ( .I(n1905), .Z(n839) );
  MUX3ND0 U914 ( .I0(n1890), .I1(n1891), .I2(n1892), .S0(n2257), .S1(N48), 
        .ZN(N67) );
  BUFFD0 U915 ( .I(n842), .Z(n840) );
  INVD10 U916 ( .I(n841), .ZN(n842) );
  INVD0 U917 ( .I(n848), .ZN(n841) );
  INVD0 U918 ( .I(n844), .ZN(n845) );
  BUFFD0 U919 ( .I(N67), .Z(n843) );
  CKNXD16 U920 ( .I(n843), .ZN(n844) );
  CKNXD16 U921 ( .I(n847), .ZN(n848) );
  INVD0 U922 ( .I(n877), .ZN(n847) );
  INVD0 U923 ( .I(n876), .ZN(n877) );
  INVD0 U924 ( .I(n857), .ZN(n858) );
  INVD0 U925 ( .I(n852), .ZN(n853) );
  BUFFD0 U926 ( .I(n848), .Z(n846) );
  BUFFD0 U927 ( .I(n875), .Z(n878) );
  INVD0 U928 ( .I(n862), .ZN(n863) );
  CKNXD16 U929 ( .I(n849), .ZN(n850) );
  INVD0 U930 ( .I(n845), .ZN(n849) );
  BUFFD0 U931 ( .I(n850), .Z(n851) );
  CKNXD16 U932 ( .I(n851), .ZN(n852) );
  CKNXD16 U933 ( .I(n854), .ZN(n855) );
  INVD0 U934 ( .I(n853), .ZN(n854) );
  BUFFD0 U935 ( .I(n855), .Z(n856) );
  CKNXD16 U936 ( .I(n856), .ZN(n857) );
  CKNXD16 U937 ( .I(n859), .ZN(n860) );
  INVD0 U938 ( .I(n858), .ZN(n859) );
  BUFFD0 U939 ( .I(n860), .Z(n861) );
  CKNXD16 U940 ( .I(n861), .ZN(n862) );
  CKNXD16 U941 ( .I(n864), .ZN(n865) );
  INVD0 U942 ( .I(n863), .ZN(n864) );
  BUFFD0 U943 ( .I(n865), .Z(n866) );
  INVD0 U944 ( .I(n867), .ZN(n868) );
  CKNXD16 U945 ( .I(n866), .ZN(n867) );
  CKNXD16 U946 ( .I(n869), .ZN(n870) );
  INVD0 U947 ( .I(n868), .ZN(n869) );
  BUFFD0 U948 ( .I(n870), .Z(n871) );
  INVD0 U949 ( .I(n872), .ZN(n873) );
  CKNXD16 U950 ( .I(n871), .ZN(n872) );
  CKNXD16 U951 ( .I(n874), .ZN(n875) );
  INVD0 U952 ( .I(n873), .ZN(n874) );
  CKNXD16 U953 ( .I(n878), .ZN(n876) );
  MUX3ND0 U954 ( .I0(n1877), .I1(n1878), .I2(n1879), .S0(n2257), .S1(n2258), 
        .ZN(N68) );
  BUFFD0 U955 ( .I(n881), .Z(n879) );
  INVD10 U956 ( .I(n880), .ZN(n881) );
  INVD0 U957 ( .I(n887), .ZN(n880) );
  INVD0 U958 ( .I(n883), .ZN(n884) );
  BUFFD0 U959 ( .I(N68), .Z(n882) );
  CKNXD16 U960 ( .I(n882), .ZN(n883) );
  CKNXD16 U961 ( .I(n886), .ZN(n887) );
  INVD0 U962 ( .I(n916), .ZN(n886) );
  INVD0 U963 ( .I(n915), .ZN(n916) );
  INVD0 U964 ( .I(n896), .ZN(n897) );
  INVD0 U965 ( .I(n891), .ZN(n892) );
  BUFFD0 U966 ( .I(n887), .Z(n885) );
  BUFFD0 U967 ( .I(n914), .Z(n917) );
  INVD0 U968 ( .I(n901), .ZN(n902) );
  CKNXD16 U969 ( .I(n888), .ZN(n889) );
  INVD0 U970 ( .I(n884), .ZN(n888) );
  BUFFD0 U971 ( .I(n889), .Z(n890) );
  CKNXD16 U972 ( .I(n890), .ZN(n891) );
  CKNXD16 U973 ( .I(n893), .ZN(n894) );
  INVD0 U974 ( .I(n892), .ZN(n893) );
  BUFFD0 U975 ( .I(n894), .Z(n895) );
  CKNXD16 U976 ( .I(n895), .ZN(n896) );
  CKNXD16 U977 ( .I(n898), .ZN(n899) );
  INVD0 U978 ( .I(n897), .ZN(n898) );
  BUFFD0 U979 ( .I(n899), .Z(n900) );
  CKNXD16 U980 ( .I(n900), .ZN(n901) );
  CKNXD16 U981 ( .I(n903), .ZN(n904) );
  INVD0 U982 ( .I(n902), .ZN(n903) );
  BUFFD0 U983 ( .I(n904), .Z(n905) );
  INVD0 U984 ( .I(n906), .ZN(n907) );
  CKNXD16 U985 ( .I(n905), .ZN(n906) );
  CKNXD16 U986 ( .I(n908), .ZN(n909) );
  INVD0 U987 ( .I(n907), .ZN(n908) );
  BUFFD0 U988 ( .I(n909), .Z(n910) );
  INVD0 U989 ( .I(n911), .ZN(n912) );
  CKNXD16 U990 ( .I(n910), .ZN(n911) );
  CKNXD16 U991 ( .I(n913), .ZN(n914) );
  INVD0 U992 ( .I(n912), .ZN(n913) );
  CKNXD16 U993 ( .I(n917), .ZN(n915) );
  INVD12 U994 ( .I(n57), .ZN(n918) );
  BUFFD0 U995 ( .I(n949), .Z(n952) );
  INVD0 U996 ( .I(n936), .ZN(n937) );
  INVD0 U997 ( .I(n926), .ZN(n927) );
  INVD1 U998 ( .I(n918), .ZN(n919) );
  INVD0 U999 ( .I(n921), .ZN(n922) );
  CKNXD16 U1000 ( .I(n920), .ZN(n921) );
  CKNXD16 U1001 ( .I(n923), .ZN(n924) );
  INVD0 U1002 ( .I(n922), .ZN(n923) );
  CKNXD16 U1003 ( .I(n925), .ZN(n926) );
  CKNXD16 U1004 ( .I(n928), .ZN(n929) );
  INVD0 U1005 ( .I(n927), .ZN(n928) );
  BUFFD0 U1006 ( .I(n929), .Z(n930) );
  INVD0 U1007 ( .I(n931), .ZN(n932) );
  CKNXD16 U1008 ( .I(n930), .ZN(n931) );
  CKNXD16 U1009 ( .I(n933), .ZN(n934) );
  INVD0 U1010 ( .I(n932), .ZN(n933) );
  BUFFD0 U1011 ( .I(n934), .Z(n935) );
  CKNXD16 U1012 ( .I(n935), .ZN(n936) );
  CKNXD16 U1013 ( .I(n938), .ZN(n939) );
  INVD0 U1014 ( .I(n937), .ZN(n938) );
  BUFFD0 U1015 ( .I(n939), .Z(n940) );
  INVD0 U1016 ( .I(n941), .ZN(n942) );
  CKNXD16 U1017 ( .I(n940), .ZN(n941) );
  CKNXD16 U1018 ( .I(n943), .ZN(n944) );
  INVD0 U1019 ( .I(n942), .ZN(n943) );
  BUFFD0 U1020 ( .I(n944), .Z(n945) );
  INVD0 U1021 ( .I(n946), .ZN(n947) );
  CKNXD16 U1022 ( .I(n945), .ZN(n946) );
  CKNXD16 U1023 ( .I(n948), .ZN(n949) );
  INVD0 U1024 ( .I(n947), .ZN(n948) );
  CKNXD16 U1025 ( .I(n952), .ZN(n950) );
  INVD12 U1026 ( .I(n62), .ZN(n953) );
  BUFFD0 U1027 ( .I(n984), .Z(n987) );
  INVD0 U1028 ( .I(n971), .ZN(n972) );
  INVD0 U1029 ( .I(n961), .ZN(n962) );
  INVD1 U1030 ( .I(n953), .ZN(n954) );
  INVD0 U1031 ( .I(n956), .ZN(n957) );
  CKNXD16 U1032 ( .I(n955), .ZN(n956) );
  CKNXD16 U1033 ( .I(n958), .ZN(n959) );
  INVD0 U1034 ( .I(n957), .ZN(n958) );
  CKNXD16 U1035 ( .I(n960), .ZN(n961) );
  CKNXD16 U1036 ( .I(n963), .ZN(n964) );
  INVD0 U1037 ( .I(n962), .ZN(n963) );
  BUFFD0 U1038 ( .I(n964), .Z(n965) );
  INVD0 U1039 ( .I(n966), .ZN(n967) );
  CKNXD16 U1040 ( .I(n965), .ZN(n966) );
  CKNXD16 U1041 ( .I(n968), .ZN(n969) );
  INVD0 U1042 ( .I(n967), .ZN(n968) );
  BUFFD0 U1043 ( .I(n969), .Z(n970) );
  CKNXD16 U1044 ( .I(n970), .ZN(n971) );
  CKNXD16 U1045 ( .I(n973), .ZN(n974) );
  INVD0 U1046 ( .I(n972), .ZN(n973) );
  BUFFD0 U1047 ( .I(n974), .Z(n975) );
  INVD0 U1048 ( .I(n976), .ZN(n977) );
  CKNXD16 U1049 ( .I(n975), .ZN(n976) );
  CKNXD16 U1050 ( .I(n978), .ZN(n979) );
  INVD0 U1051 ( .I(n977), .ZN(n978) );
  BUFFD0 U1052 ( .I(n979), .Z(n980) );
  INVD0 U1053 ( .I(n981), .ZN(n982) );
  CKNXD16 U1054 ( .I(n980), .ZN(n981) );
  CKNXD16 U1055 ( .I(n983), .ZN(n984) );
  INVD0 U1056 ( .I(n982), .ZN(n983) );
  CKNXD16 U1057 ( .I(n987), .ZN(n985) );
  MUX3ND0 U1058 ( .I0(n1838), .I1(n1839), .I2(n1840), .S0(n2116), .S1(n2258), 
        .ZN(N71) );
  BUFFD0 U1059 ( .I(n990), .Z(n988) );
  INVD10 U1060 ( .I(n989), .ZN(n990) );
  INVD0 U1061 ( .I(n996), .ZN(n989) );
  INVD0 U1062 ( .I(n992), .ZN(n993) );
  BUFFD0 U1063 ( .I(N71), .Z(n991) );
  CKNXD16 U1064 ( .I(n991), .ZN(n992) );
  CKNXD16 U1065 ( .I(n995), .ZN(n996) );
  INVD0 U1066 ( .I(n1025), .ZN(n995) );
  INVD0 U1067 ( .I(n1024), .ZN(n1025) );
  INVD0 U1068 ( .I(n1005), .ZN(n1006) );
  INVD0 U1069 ( .I(n1000), .ZN(n1001) );
  BUFFD0 U1070 ( .I(n996), .Z(n994) );
  BUFFD0 U1071 ( .I(n1023), .Z(n1026) );
  INVD0 U1072 ( .I(n1010), .ZN(n1011) );
  CKNXD16 U1073 ( .I(n997), .ZN(n998) );
  INVD0 U1074 ( .I(n993), .ZN(n997) );
  BUFFD0 U1075 ( .I(n998), .Z(n999) );
  CKNXD16 U1076 ( .I(n999), .ZN(n1000) );
  CKNXD16 U1077 ( .I(n1002), .ZN(n1003) );
  INVD0 U1078 ( .I(n1001), .ZN(n1002) );
  BUFFD0 U1079 ( .I(n1003), .Z(n1004) );
  CKNXD16 U1080 ( .I(n1004), .ZN(n1005) );
  CKNXD16 U1081 ( .I(n1007), .ZN(n1008) );
  INVD0 U1082 ( .I(n1006), .ZN(n1007) );
  BUFFD0 U1083 ( .I(n1008), .Z(n1009) );
  CKNXD16 U1084 ( .I(n1009), .ZN(n1010) );
  CKNXD16 U1085 ( .I(n1012), .ZN(n1013) );
  INVD0 U1086 ( .I(n1011), .ZN(n1012) );
  BUFFD0 U1087 ( .I(n1013), .Z(n1014) );
  INVD0 U1088 ( .I(n1015), .ZN(n1016) );
  CKNXD16 U1089 ( .I(n1014), .ZN(n1015) );
  CKNXD16 U1090 ( .I(n1017), .ZN(n1018) );
  INVD0 U1091 ( .I(n1016), .ZN(n1017) );
  BUFFD0 U1092 ( .I(n1018), .Z(n1019) );
  INVD0 U1093 ( .I(n1020), .ZN(n1021) );
  CKNXD16 U1094 ( .I(n1019), .ZN(n1020) );
  CKNXD16 U1095 ( .I(n1022), .ZN(n1023) );
  INVD0 U1096 ( .I(n1021), .ZN(n1022) );
  CKNXD16 U1097 ( .I(n1026), .ZN(n1024) );
  INVD0 U1098 ( .I(n1033), .ZN(n1027) );
  CKND12 U1099 ( .CLK(n1044), .CN(n1045) );
  INVD0 U1100 ( .I(n1029), .ZN(n1030) );
  CKNXD16 U1101 ( .I(n248), .ZN(n1029) );
  CKNXD16 U1102 ( .I(n1032), .ZN(n1033) );
  INVD0 U1103 ( .I(n1062), .ZN(n1032) );
  INVD0 U1104 ( .I(n1061), .ZN(n1062) );
  INVD0 U1105 ( .I(n1042), .ZN(n1043) );
  INVD0 U1106 ( .I(n1037), .ZN(n1038) );
  BUFFD0 U1107 ( .I(n1033), .Z(n1031) );
  BUFFD0 U1108 ( .I(n1060), .Z(n1063) );
  INVD0 U1109 ( .I(n1047), .ZN(n1048) );
  CKNXD16 U1110 ( .I(n1034), .ZN(n1035) );
  INVD0 U1111 ( .I(n1030), .ZN(n1034) );
  BUFFD0 U1112 ( .I(n1035), .Z(n1036) );
  CKNXD16 U1113 ( .I(n1036), .ZN(n1037) );
  INVD0 U1114 ( .I(n1038), .ZN(n1039) );
  BUFFD0 U1115 ( .I(n1040), .Z(n1041) );
  CKNXD16 U1116 ( .I(n1041), .ZN(n1042) );
  INVD0 U1117 ( .I(n1043), .ZN(n1044) );
  BUFFD0 U1118 ( .I(n1045), .Z(n1046) );
  CKNXD16 U1119 ( .I(n1046), .ZN(n1047) );
  CKNXD16 U1120 ( .I(n1049), .ZN(n1050) );
  INVD0 U1121 ( .I(n1048), .ZN(n1049) );
  BUFFD0 U1122 ( .I(n1050), .Z(n1051) );
  INVD0 U1123 ( .I(n1052), .ZN(n1053) );
  CKNXD16 U1124 ( .I(n1051), .ZN(n1052) );
  CKNXD16 U1125 ( .I(n1054), .ZN(n1055) );
  INVD0 U1126 ( .I(n1053), .ZN(n1054) );
  BUFFD0 U1127 ( .I(n1055), .Z(n1056) );
  INVD0 U1128 ( .I(n1057), .ZN(n1058) );
  CKNXD16 U1129 ( .I(n1056), .ZN(n1057) );
  CKNXD16 U1130 ( .I(n1059), .ZN(n1060) );
  INVD0 U1131 ( .I(n1058), .ZN(n1059) );
  CKNXD16 U1132 ( .I(n1063), .ZN(n1061) );
  MUX3ND0 U1133 ( .I0(n1812), .I1(n1813), .I2(n1814), .S0(n2116), .S1(n2258), 
        .ZN(N73) );
  BUFFD0 U1134 ( .I(n1066), .Z(n1064) );
  INVD10 U1135 ( .I(n1065), .ZN(n1066) );
  INVD0 U1136 ( .I(n1072), .ZN(n1065) );
  INVD0 U1137 ( .I(n1068), .ZN(n1069) );
  BUFFD0 U1138 ( .I(N73), .Z(n1067) );
  CKNXD16 U1139 ( .I(n1067), .ZN(n1068) );
  CKNXD16 U1140 ( .I(n1071), .ZN(n1072) );
  INVD0 U1141 ( .I(n1101), .ZN(n1071) );
  INVD0 U1142 ( .I(n1100), .ZN(n1101) );
  INVD0 U1143 ( .I(n1081), .ZN(n1082) );
  INVD0 U1144 ( .I(n1076), .ZN(n1077) );
  BUFFD0 U1145 ( .I(n1072), .Z(n1070) );
  BUFFD0 U1146 ( .I(n1099), .Z(n1102) );
  INVD0 U1147 ( .I(n1086), .ZN(n1087) );
  CKNXD16 U1148 ( .I(n1073), .ZN(n1074) );
  INVD0 U1149 ( .I(n1069), .ZN(n1073) );
  BUFFD0 U1150 ( .I(n1074), .Z(n1075) );
  CKNXD16 U1151 ( .I(n1075), .ZN(n1076) );
  CKNXD16 U1152 ( .I(n1078), .ZN(n1079) );
  INVD0 U1153 ( .I(n1077), .ZN(n1078) );
  BUFFD0 U1154 ( .I(n1079), .Z(n1080) );
  CKNXD16 U1155 ( .I(n1080), .ZN(n1081) );
  CKNXD16 U1156 ( .I(n1083), .ZN(n1084) );
  INVD0 U1157 ( .I(n1082), .ZN(n1083) );
  BUFFD0 U1158 ( .I(n1084), .Z(n1085) );
  CKNXD16 U1159 ( .I(n1085), .ZN(n1086) );
  CKNXD16 U1160 ( .I(n1088), .ZN(n1089) );
  INVD0 U1161 ( .I(n1087), .ZN(n1088) );
  BUFFD0 U1162 ( .I(n1089), .Z(n1090) );
  INVD0 U1163 ( .I(n1091), .ZN(n1092) );
  CKNXD16 U1164 ( .I(n1090), .ZN(n1091) );
  CKNXD16 U1165 ( .I(n1093), .ZN(n1094) );
  INVD0 U1166 ( .I(n1092), .ZN(n1093) );
  BUFFD0 U1167 ( .I(n1094), .Z(n1095) );
  INVD0 U1168 ( .I(n1096), .ZN(n1097) );
  CKNXD16 U1169 ( .I(n1095), .ZN(n1096) );
  CKNXD16 U1170 ( .I(n1098), .ZN(n1099) );
  INVD0 U1171 ( .I(n1097), .ZN(n1098) );
  CKNXD16 U1172 ( .I(n1102), .ZN(n1100) );
  INVD0 U1173 ( .I(n1104), .ZN(n1105) );
  CKNXD16 U1174 ( .I(n1107), .ZN(n1104) );
  CKNXD0 U1175 ( .I(n1106), .ZN(n1107) );
  CKNXD16 U1176 ( .I(n1109), .ZN(n1106) );
  CKNXD0 U1177 ( .I(n1128), .ZN(n1129) );
  CKBD0 U1178 ( .CLK(n1103), .C(n1110) );
  INVD0 U1179 ( .I(n1108), .ZN(n1109) );
  CKNXD16 U1180 ( .I(n1111), .ZN(n1108) );
  CKBD0 U1181 ( .CLK(n1113), .C(n1111) );
  CKNXD16 U1182 ( .I(n1112), .ZN(n1113) );
  INVD0 U1183 ( .I(n1117), .ZN(n1112) );
  INVD0 U1184 ( .I(n1116), .ZN(n1117) );
  INVD0 U1185 ( .I(n1123), .ZN(n1124) );
  INVD0 U1186 ( .I(n1136), .ZN(n1137) );
  BUFFD0 U1187 ( .I(n1126), .Z(n1127) );
  CKNXD16 U1188 ( .I(n1114), .ZN(n1115) );
  INVD0 U1189 ( .I(n1110), .ZN(n1114) );
  CKNXD16 U1190 ( .I(n1119), .ZN(n1116) );
  INVD0 U1191 ( .I(n1118), .ZN(n1119) );
  CKNXD16 U1192 ( .I(n1120), .ZN(n1118) );
  CKNXD16 U1193 ( .I(n1121), .ZN(n1122) );
  INVD0 U1194 ( .I(n1124), .ZN(n1121) );
  BUFFD0 U1195 ( .I(n1122), .Z(n1120) );
  CKNXD16 U1196 ( .I(n1131), .ZN(n1123) );
  CKNXD16 U1197 ( .I(n1125), .ZN(n1126) );
  INVD0 U1198 ( .I(n1115), .ZN(n1125) );
  CKNXD16 U1199 ( .I(n1127), .ZN(n1128) );
  CKNXD16 U1200 ( .I(n1132), .ZN(n1133) );
  INVD0 U1201 ( .I(n1137), .ZN(n1132) );
  BUFFD0 U1202 ( .I(n1133), .Z(n1131) );
  BUFFD0 U1203 ( .I(n1135), .Z(n1138) );
  CKNXD16 U1204 ( .I(n1134), .ZN(n1135) );
  INVD0 U1205 ( .I(n1130), .ZN(n1134) );
  CKNXD16 U1206 ( .I(n1138), .ZN(n1136) );
  BUFFD0 U1207 ( .I(n1801), .Z(n1139) );
  INVD12 U1208 ( .I(n107), .ZN(n1140) );
  BUFFD0 U1209 ( .I(n1171), .Z(n1174) );
  INVD0 U1210 ( .I(n1158), .ZN(n1159) );
  INVD0 U1211 ( .I(n1148), .ZN(n1149) );
  INVD1 U1212 ( .I(n1140), .ZN(n1141) );
  INVD0 U1213 ( .I(n1143), .ZN(n1144) );
  CKNXD16 U1214 ( .I(n1142), .ZN(n1143) );
  CKNXD16 U1215 ( .I(n1145), .ZN(n1146) );
  INVD0 U1216 ( .I(n1144), .ZN(n1145) );
  CKNXD16 U1217 ( .I(n1147), .ZN(n1148) );
  CKNXD16 U1218 ( .I(n1150), .ZN(n1151) );
  INVD0 U1219 ( .I(n1149), .ZN(n1150) );
  BUFFD0 U1220 ( .I(n1151), .Z(n1152) );
  INVD0 U1221 ( .I(n1153), .ZN(n1154) );
  CKNXD16 U1222 ( .I(n1152), .ZN(n1153) );
  CKNXD16 U1223 ( .I(n1155), .ZN(n1156) );
  INVD0 U1224 ( .I(n1154), .ZN(n1155) );
  BUFFD0 U1225 ( .I(n1156), .Z(n1157) );
  CKNXD16 U1226 ( .I(n1157), .ZN(n1158) );
  CKNXD16 U1227 ( .I(n1160), .ZN(n1161) );
  INVD0 U1228 ( .I(n1159), .ZN(n1160) );
  BUFFD0 U1229 ( .I(n1161), .Z(n1162) );
  INVD0 U1230 ( .I(n1163), .ZN(n1164) );
  CKNXD16 U1231 ( .I(n1162), .ZN(n1163) );
  CKNXD16 U1232 ( .I(n1165), .ZN(n1166) );
  INVD0 U1233 ( .I(n1164), .ZN(n1165) );
  BUFFD0 U1234 ( .I(n1166), .Z(n1167) );
  INVD0 U1235 ( .I(n1168), .ZN(n1169) );
  CKNXD16 U1236 ( .I(n1167), .ZN(n1168) );
  CKNXD16 U1237 ( .I(n1170), .ZN(n1171) );
  INVD0 U1238 ( .I(n1169), .ZN(n1170) );
  CKNXD16 U1239 ( .I(n1174), .ZN(n1172) );
  INVD12 U1240 ( .I(n113), .ZN(n1175) );
  BUFFD0 U1241 ( .I(n1206), .Z(n1209) );
  INVD0 U1242 ( .I(n1193), .ZN(n1194) );
  INVD0 U1243 ( .I(n1183), .ZN(n1184) );
  INVD1 U1244 ( .I(n1175), .ZN(n1176) );
  INVD0 U1245 ( .I(n1178), .ZN(n1179) );
  CKNXD16 U1246 ( .I(n1177), .ZN(n1178) );
  CKNXD16 U1247 ( .I(n1180), .ZN(n1181) );
  INVD0 U1248 ( .I(n1179), .ZN(n1180) );
  CKNXD16 U1249 ( .I(n1182), .ZN(n1183) );
  CKNXD16 U1250 ( .I(n1185), .ZN(n1186) );
  INVD0 U1251 ( .I(n1184), .ZN(n1185) );
  BUFFD0 U1252 ( .I(n1186), .Z(n1187) );
  INVD0 U1253 ( .I(n1188), .ZN(n1189) );
  CKNXD16 U1254 ( .I(n1187), .ZN(n1188) );
  CKNXD16 U1255 ( .I(n1190), .ZN(n1191) );
  INVD0 U1256 ( .I(n1189), .ZN(n1190) );
  BUFFD0 U1257 ( .I(n1191), .Z(n1192) );
  CKNXD16 U1258 ( .I(n1192), .ZN(n1193) );
  CKNXD16 U1259 ( .I(n1195), .ZN(n1196) );
  INVD0 U1260 ( .I(n1194), .ZN(n1195) );
  BUFFD0 U1261 ( .I(n1196), .Z(n1197) );
  INVD0 U1262 ( .I(n1198), .ZN(n1199) );
  CKNXD16 U1263 ( .I(n1197), .ZN(n1198) );
  CKNXD16 U1264 ( .I(n1200), .ZN(n1201) );
  INVD0 U1265 ( .I(n1199), .ZN(n1200) );
  BUFFD0 U1266 ( .I(n1201), .Z(n1202) );
  INVD0 U1267 ( .I(n1203), .ZN(n1204) );
  CKNXD16 U1268 ( .I(n1202), .ZN(n1203) );
  CKNXD16 U1269 ( .I(n1205), .ZN(n1206) );
  INVD0 U1270 ( .I(n1204), .ZN(n1205) );
  CKNXD16 U1271 ( .I(n1209), .ZN(n1207) );
  INVD0 U1272 ( .I(n1216), .ZN(n1210) );
  INVD0 U1273 ( .I(n1212), .ZN(n1213) );
  CKNXD16 U1274 ( .I(n250), .ZN(n1212) );
  MUX3ND0 U1275 ( .I0(n1760), .I1(n1761), .I2(n1762), .S0(n2117), .S1(n2258), 
        .ZN(N77) );
  CKNXD16 U1276 ( .I(n1215), .ZN(n1216) );
  INVD0 U1277 ( .I(n1245), .ZN(n1215) );
  INVD0 U1278 ( .I(n1244), .ZN(n1245) );
  INVD0 U1279 ( .I(n1225), .ZN(n1226) );
  INVD0 U1280 ( .I(n1220), .ZN(n1221) );
  BUFFD0 U1281 ( .I(n1216), .Z(n1214) );
  BUFFD0 U1282 ( .I(n1243), .Z(n1246) );
  INVD0 U1283 ( .I(n1230), .ZN(n1231) );
  CKNXD16 U1284 ( .I(n1217), .ZN(n1218) );
  INVD0 U1285 ( .I(n1213), .ZN(n1217) );
  BUFFD0 U1286 ( .I(n1218), .Z(n1219) );
  CKNXD16 U1287 ( .I(n1219), .ZN(n1220) );
  CKNXD16 U1288 ( .I(n1222), .ZN(n1223) );
  INVD0 U1289 ( .I(n1221), .ZN(n1222) );
  BUFFD0 U1290 ( .I(n1223), .Z(n1224) );
  CKNXD16 U1291 ( .I(n1224), .ZN(n1225) );
  CKNXD16 U1292 ( .I(n1227), .ZN(n1228) );
  INVD0 U1293 ( .I(n1226), .ZN(n1227) );
  BUFFD0 U1294 ( .I(n1228), .Z(n1229) );
  CKNXD16 U1295 ( .I(n1229), .ZN(n1230) );
  CKNXD16 U1296 ( .I(n1232), .ZN(n1233) );
  INVD0 U1297 ( .I(n1231), .ZN(n1232) );
  BUFFD0 U1298 ( .I(n1233), .Z(n1234) );
  INVD0 U1299 ( .I(n1235), .ZN(n1236) );
  CKNXD16 U1300 ( .I(n1234), .ZN(n1235) );
  CKNXD16 U1301 ( .I(n1237), .ZN(n1238) );
  INVD0 U1302 ( .I(n1236), .ZN(n1237) );
  BUFFD0 U1303 ( .I(n1238), .Z(n1239) );
  INVD0 U1304 ( .I(n1240), .ZN(n1241) );
  CKNXD16 U1305 ( .I(n1239), .ZN(n1240) );
  CKNXD16 U1306 ( .I(n1242), .ZN(n1243) );
  INVD0 U1307 ( .I(n1241), .ZN(n1242) );
  CKNXD16 U1308 ( .I(n1246), .ZN(n1244) );
  INVD0 U1309 ( .I(n1253), .ZN(n1247) );
  CKND12 U1310 ( .CLK(n1264), .CN(n1265) );
  INVD0 U1311 ( .I(n1249), .ZN(n1250) );
  CKNXD16 U1312 ( .I(n249), .ZN(n1249) );
  CKNXD16 U1313 ( .I(n1252), .ZN(n1253) );
  INVD0 U1314 ( .I(n1282), .ZN(n1252) );
  INVD0 U1315 ( .I(n1281), .ZN(n1282) );
  INVD0 U1316 ( .I(n1262), .ZN(n1263) );
  INVD0 U1317 ( .I(n1257), .ZN(n1258) );
  BUFFD0 U1318 ( .I(n1253), .Z(n1251) );
  BUFFD0 U1319 ( .I(n1280), .Z(n1283) );
  INVD0 U1320 ( .I(n1267), .ZN(n1268) );
  CKNXD16 U1321 ( .I(n1254), .ZN(n1255) );
  INVD0 U1322 ( .I(n1250), .ZN(n1254) );
  BUFFD0 U1323 ( .I(n1255), .Z(n1256) );
  CKNXD16 U1324 ( .I(n1256), .ZN(n1257) );
  INVD0 U1325 ( .I(n1258), .ZN(n1259) );
  BUFFD0 U1326 ( .I(n1260), .Z(n1261) );
  CKNXD16 U1327 ( .I(n1261), .ZN(n1262) );
  INVD0 U1328 ( .I(n1263), .ZN(n1264) );
  BUFFD0 U1329 ( .I(n1265), .Z(n1266) );
  CKNXD16 U1330 ( .I(n1266), .ZN(n1267) );
  CKNXD16 U1331 ( .I(n1269), .ZN(n1270) );
  INVD0 U1332 ( .I(n1268), .ZN(n1269) );
  BUFFD0 U1333 ( .I(n1270), .Z(n1271) );
  INVD0 U1334 ( .I(n1272), .ZN(n1273) );
  CKNXD16 U1335 ( .I(n1271), .ZN(n1272) );
  CKNXD16 U1336 ( .I(n1274), .ZN(n1275) );
  INVD0 U1337 ( .I(n1273), .ZN(n1274) );
  BUFFD0 U1338 ( .I(n1275), .Z(n1276) );
  INVD0 U1339 ( .I(n1277), .ZN(n1278) );
  CKNXD16 U1340 ( .I(n1276), .ZN(n1277) );
  CKNXD16 U1341 ( .I(n1279), .ZN(n1280) );
  INVD0 U1342 ( .I(n1278), .ZN(n1279) );
  CKNXD16 U1343 ( .I(n1283), .ZN(n1281) );
  CKNXD0 U1344 ( .I(n1287), .ZN(n1288) );
  INVD8 U1345 ( .I(n1284), .ZN(n1285) );
  INVD0 U1346 ( .I(n1290), .ZN(n1284) );
  MUX3ND4 U1347 ( .I0(n1734), .I1(n1735), .I2(n1736), .S0(n2116), .S1(n2258), 
        .ZN(N79) );
  BUFFD0 U1348 ( .I(N79), .Z(n1286) );
  CKNXD16 U1349 ( .I(n1286), .ZN(n1287) );
  CKNXD16 U1350 ( .I(n1289), .ZN(n1290) );
  INVD0 U1351 ( .I(n1319), .ZN(n1289) );
  INVD0 U1352 ( .I(n1318), .ZN(n1319) );
  INVD0 U1353 ( .I(n1299), .ZN(n1300) );
  INVD0 U1354 ( .I(n1294), .ZN(n1295) );
  BUFFD0 U1355 ( .I(n1317), .Z(n1320) );
  INVD0 U1356 ( .I(n1304), .ZN(n1305) );
  CKNXD16 U1357 ( .I(n1291), .ZN(n1292) );
  INVD0 U1358 ( .I(n1288), .ZN(n1291) );
  BUFFD0 U1359 ( .I(n1292), .Z(n1293) );
  CKNXD16 U1360 ( .I(n1293), .ZN(n1294) );
  CKNXD16 U1361 ( .I(n1296), .ZN(n1297) );
  INVD0 U1362 ( .I(n1295), .ZN(n1296) );
  BUFFD0 U1363 ( .I(n1297), .Z(n1298) );
  CKNXD16 U1364 ( .I(n1298), .ZN(n1299) );
  CKNXD16 U1365 ( .I(n1301), .ZN(n1302) );
  INVD0 U1366 ( .I(n1300), .ZN(n1301) );
  BUFFD0 U1367 ( .I(n1302), .Z(n1303) );
  CKNXD16 U1368 ( .I(n1303), .ZN(n1304) );
  CKNXD16 U1369 ( .I(n1306), .ZN(n1307) );
  INVD0 U1370 ( .I(n1305), .ZN(n1306) );
  BUFFD0 U1371 ( .I(n1307), .Z(n1308) );
  INVD0 U1372 ( .I(n1309), .ZN(n1310) );
  CKNXD16 U1373 ( .I(n1308), .ZN(n1309) );
  CKNXD16 U1374 ( .I(n1311), .ZN(n1312) );
  INVD0 U1375 ( .I(n1310), .ZN(n1311) );
  BUFFD0 U1376 ( .I(n1312), .Z(n1313) );
  INVD0 U1377 ( .I(n1314), .ZN(n1315) );
  CKNXD16 U1378 ( .I(n1313), .ZN(n1314) );
  CKNXD16 U1379 ( .I(n1316), .ZN(n1317) );
  INVD0 U1380 ( .I(n1315), .ZN(n1316) );
  CKNXD16 U1381 ( .I(n1320), .ZN(n1318) );
  INVD12 U1382 ( .I(n119), .ZN(n1321) );
  BUFFD0 U1383 ( .I(n1352), .Z(n1355) );
  INVD0 U1384 ( .I(n1339), .ZN(n1340) );
  INVD0 U1385 ( .I(n1329), .ZN(n1330) );
  INVD1 U1386 ( .I(n1321), .ZN(n1322) );
  INVD0 U1387 ( .I(n1324), .ZN(n1325) );
  CKNXD16 U1388 ( .I(n1323), .ZN(n1324) );
  CKNXD16 U1389 ( .I(n1326), .ZN(n1327) );
  INVD0 U1390 ( .I(n1325), .ZN(n1326) );
  CKNXD16 U1391 ( .I(n1328), .ZN(n1329) );
  CKNXD16 U1392 ( .I(n1331), .ZN(n1332) );
  INVD0 U1393 ( .I(n1330), .ZN(n1331) );
  BUFFD0 U1394 ( .I(n1332), .Z(n1333) );
  INVD0 U1395 ( .I(n1334), .ZN(n1335) );
  CKNXD16 U1396 ( .I(n1333), .ZN(n1334) );
  CKNXD16 U1397 ( .I(n1336), .ZN(n1337) );
  INVD0 U1398 ( .I(n1335), .ZN(n1336) );
  BUFFD0 U1399 ( .I(n1337), .Z(n1338) );
  CKNXD16 U1400 ( .I(n1338), .ZN(n1339) );
  CKNXD16 U1401 ( .I(n1341), .ZN(n1342) );
  INVD0 U1402 ( .I(n1340), .ZN(n1341) );
  BUFFD0 U1403 ( .I(n1342), .Z(n1343) );
  INVD0 U1404 ( .I(n1344), .ZN(n1345) );
  CKNXD16 U1405 ( .I(n1343), .ZN(n1344) );
  CKNXD16 U1406 ( .I(n1346), .ZN(n1347) );
  INVD0 U1407 ( .I(n1345), .ZN(n1346) );
  BUFFD0 U1408 ( .I(n1347), .Z(n1348) );
  INVD0 U1409 ( .I(n1349), .ZN(n1350) );
  CKNXD16 U1410 ( .I(n1348), .ZN(n1349) );
  CKNXD16 U1411 ( .I(n1351), .ZN(n1352) );
  INVD0 U1412 ( .I(n1350), .ZN(n1351) );
  CKNXD16 U1413 ( .I(n1355), .ZN(n1353) );
  INVD0 U1414 ( .I(n1356), .ZN(n1357) );
  CKNXD16 U1415 ( .I(n1361), .ZN(n1356) );
  CKND12 U1416 ( .CLK(n1379), .CN(n1380) );
  INVD0 U1417 ( .I(N81), .ZN(n1358) );
  CKNXD16 U1418 ( .I(n1358), .ZN(n1359) );
  MUX3ND0 U1419 ( .I0(n1708), .I1(n1709), .I2(n1710), .S0(n2116), .S1(n2258), 
        .ZN(N81) );
  INVD0 U1420 ( .I(n1360), .ZN(n1361) );
  CKNXD16 U1421 ( .I(n1365), .ZN(n1360) );
  INVD0 U1422 ( .I(n1359), .ZN(n1362) );
  CKNXD16 U1423 ( .I(n1362), .ZN(n1363) );
  INVD0 U1424 ( .I(n1364), .ZN(n1365) );
  CKNXD16 U1425 ( .I(n1369), .ZN(n1364) );
  INVD0 U1426 ( .I(n1363), .ZN(n1366) );
  CKNXD16 U1427 ( .I(n1366), .ZN(n1367) );
  INVD0 U1428 ( .I(n1368), .ZN(n1369) );
  CKNXD16 U1429 ( .I(n1374), .ZN(n1368) );
  INVD0 U1430 ( .I(n1367), .ZN(n1370) );
  CKNXD16 U1431 ( .I(n1370), .ZN(n1371) );
  CKBD0 U1432 ( .CLK(n1371), .C(n1372) );
  BUFFD0 U1433 ( .I(n1372), .Z(n1373) );
  BUFFD0 U1434 ( .I(n1376), .Z(n1374) );
  CKNXD16 U1435 ( .I(n1375), .ZN(n1376) );
  INVD0 U1436 ( .I(n1380), .ZN(n1375) );
  INVD0 U1437 ( .I(n1377), .ZN(n1378) );
  CKNXD16 U1438 ( .I(n1373), .ZN(n1377) );
  INVD0 U1439 ( .I(n1389), .ZN(n1379) );
  INVD0 U1440 ( .I(n1388), .ZN(n1389) );
  BUFFD0 U1441 ( .I(n1387), .Z(n1390) );
  CKNXD16 U1442 ( .I(n1381), .ZN(n1382) );
  INVD0 U1443 ( .I(n1378), .ZN(n1381) );
  BUFFD0 U1444 ( .I(n1382), .Z(n1383) );
  INVD0 U1445 ( .I(n1384), .ZN(n1385) );
  CKNXD16 U1446 ( .I(n1383), .ZN(n1384) );
  CKNXD16 U1447 ( .I(n1386), .ZN(n1387) );
  INVD0 U1448 ( .I(n1385), .ZN(n1386) );
  CKNXD16 U1449 ( .I(n1390), .ZN(n1388) );
  INVD16 U1450 ( .I(n1394), .ZN(n1395) );
  BUFFD0 U1451 ( .I(n1393), .Z(n1391) );
  INVD0 U1452 ( .I(n1392), .ZN(n1393) );
  CKNXD16 U1453 ( .I(n1397), .ZN(n1392) );
  INVD0 U1454 ( .I(N82), .ZN(n1394) );
  MUX3ND0 U1455 ( .I0(n1695), .I1(n1696), .I2(n1697), .S0(n2116), .S1(n2258), 
        .ZN(N82) );
  INVD0 U1456 ( .I(n1396), .ZN(n1397) );
  CKNXD16 U1457 ( .I(n1401), .ZN(n1396) );
  INVD0 U1458 ( .I(n1395), .ZN(n1398) );
  CKNXD16 U1459 ( .I(n1398), .ZN(n1399) );
  INVD0 U1460 ( .I(n1400), .ZN(n1401) );
  CKNXD16 U1461 ( .I(n1405), .ZN(n1400) );
  INVD0 U1462 ( .I(n1399), .ZN(n1402) );
  CKNXD16 U1463 ( .I(n1402), .ZN(n1403) );
  INVD0 U1464 ( .I(n1404), .ZN(n1405) );
  CKNXD16 U1465 ( .I(n1410), .ZN(n1404) );
  INVD0 U1466 ( .I(n1403), .ZN(n1406) );
  CKNXD16 U1467 ( .I(n1406), .ZN(n1407) );
  CKBD0 U1468 ( .CLK(n1407), .C(n1408) );
  BUFFD0 U1469 ( .I(n1408), .Z(n1409) );
  BUFFD0 U1470 ( .I(n1412), .Z(n1410) );
  CKNXD16 U1471 ( .I(n1411), .ZN(n1412) );
  INVD0 U1472 ( .I(n1416), .ZN(n1411) );
  INVD0 U1473 ( .I(n1413), .ZN(n1414) );
  CKNXD16 U1474 ( .I(n1409), .ZN(n1413) );
  CKNXD16 U1475 ( .I(n1415), .ZN(n1416) );
  INVD0 U1476 ( .I(n1425), .ZN(n1415) );
  INVD0 U1477 ( .I(n1424), .ZN(n1425) );
  BUFFD0 U1478 ( .I(n1423), .Z(n1426) );
  CKNXD16 U1479 ( .I(n1417), .ZN(n1418) );
  INVD0 U1480 ( .I(n1414), .ZN(n1417) );
  BUFFD0 U1481 ( .I(n1418), .Z(n1419) );
  INVD0 U1482 ( .I(n1420), .ZN(n1421) );
  CKNXD16 U1483 ( .I(n1419), .ZN(n1420) );
  CKNXD16 U1484 ( .I(n1422), .ZN(n1423) );
  INVD0 U1485 ( .I(n1421), .ZN(n1422) );
  CKNXD16 U1486 ( .I(n1426), .ZN(n1424) );
  CKNXD0 U1487 ( .I(n1428), .ZN(n1429) );
  INVD0 U1488 ( .I(n1430), .ZN(n1431) );
  INVD0 U1489 ( .I(n1432), .ZN(n1433) );
  INVD0 U1490 ( .I(n1434), .ZN(n1435) );
  CKNXD0 U1491 ( .I(n1436), .ZN(n1437) );
  INVD0 U1492 ( .I(n1438), .ZN(n1439) );
  INVD0 U1493 ( .I(n1440), .ZN(n1441) );
  INVD0 U1494 ( .I(n1442), .ZN(n1443) );
  CKNXD0 U1495 ( .I(n1444), .ZN(n1445) );
  INVD0 U1496 ( .I(n1446), .ZN(n1447) );
  INVD0 U1497 ( .I(n1448), .ZN(n1449) );
  INVD0 U1498 ( .I(n1450), .ZN(n1451) );
  CKNXD0 U1499 ( .I(n1452), .ZN(n1453) );
  INVD0 U1500 ( .I(n1454), .ZN(n1455) );
  INVD0 U1501 ( .I(n1456), .ZN(n1457) );
  INVD0 U1502 ( .I(n1458), .ZN(n1459) );
  CKNXD0 U1503 ( .I(n1460), .ZN(n1461) );
  INVD0 U1504 ( .I(n1462), .ZN(n1463) );
  INVD0 U1505 ( .I(n1464), .ZN(n1465) );
  INVD0 U1506 ( .I(n1466), .ZN(n1467) );
  CKNXD0 U1507 ( .I(n1468), .ZN(n1469) );
  INVD0 U1508 ( .I(n1470), .ZN(n1471) );
  INVD0 U1509 ( .I(n1472), .ZN(n1473) );
  INVD0 U1510 ( .I(n1474), .ZN(n1475) );
  CKNXD0 U1511 ( .I(n1476), .ZN(n1477) );
  INVD0 U1512 ( .I(n1478), .ZN(n1479) );
  INVD0 U1513 ( .I(n1480), .ZN(n1481) );
  INVD0 U1514 ( .I(n1482), .ZN(n1483) );
  CKNXD0 U1515 ( .I(n1484), .ZN(n1485) );
  INVD0 U1516 ( .I(n1486), .ZN(n1487) );
  INVD0 U1517 ( .I(n1488), .ZN(n1489) );
  INVD0 U1518 ( .I(n1490), .ZN(n1491) );
  CKNXD0 U1519 ( .I(n1492), .ZN(DataO[23]) );
  CKNXD16 U1520 ( .I(n1495), .ZN(n1492) );
  INVD0 U1521 ( .I(n1494), .ZN(n1495) );
  CKNXD16 U1522 ( .I(n1497), .ZN(n1494) );
  INVD0 U1523 ( .I(n1496), .ZN(n1497) );
  CKNXD16 U1524 ( .I(n1499), .ZN(n1496) );
  INVD0 U1525 ( .I(n1498), .ZN(n1499) );
  CKNXD16 U1526 ( .I(n2267), .ZN(n1498) );
  CKNXD0 U1527 ( .I(n1500), .ZN(DataO[22]) );
  CKNXD16 U1528 ( .I(n1503), .ZN(n1500) );
  INVD0 U1529 ( .I(n1502), .ZN(n1503) );
  CKNXD16 U1530 ( .I(n1505), .ZN(n1502) );
  INVD0 U1531 ( .I(n1504), .ZN(n1505) );
  CKNXD16 U1532 ( .I(n1507), .ZN(n1504) );
  INVD0 U1533 ( .I(n1506), .ZN(n1507) );
  CKNXD16 U1534 ( .I(n2268), .ZN(n1506) );
  CKNXD0 U1535 ( .I(n1508), .ZN(n1509) );
  CKNXD16 U1536 ( .I(n1511), .ZN(n1508) );
  INVD0 U1537 ( .I(n1510), .ZN(n1511) );
  CKNXD16 U1538 ( .I(n1513), .ZN(n1510) );
  INVD0 U1539 ( .I(n1512), .ZN(n1513) );
  CKNXD16 U1540 ( .I(n1515), .ZN(n1512) );
  INVD0 U1541 ( .I(n1514), .ZN(n1515) );
  CKNXD16 U1542 ( .I(n2269), .ZN(n1514) );
  CKNXD0 U1543 ( .I(n1516), .ZN(n1517) );
  INVD0 U1544 ( .I(n1518), .ZN(n1519) );
  INVD0 U1545 ( .I(n1520), .ZN(n1521) );
  INVD0 U1546 ( .I(n1522), .ZN(n1523) );
  CKNXD0 U1547 ( .I(n1524), .ZN(n1525) );
  INVD0 U1548 ( .I(n1526), .ZN(n1527) );
  INVD0 U1549 ( .I(n1528), .ZN(n1529) );
  INVD0 U1550 ( .I(n1530), .ZN(n1531) );
  CKNXD0 U1551 ( .I(n1532), .ZN(DataO[18]) );
  CKNXD16 U1552 ( .I(n1535), .ZN(n1532) );
  INVD0 U1553 ( .I(n1534), .ZN(n1535) );
  CKNXD16 U1554 ( .I(n1537), .ZN(n1534) );
  INVD0 U1555 ( .I(n1536), .ZN(n1537) );
  CKNXD16 U1556 ( .I(n1539), .ZN(n1536) );
  INVD0 U1557 ( .I(n1538), .ZN(n1539) );
  CKNXD16 U1558 ( .I(n2272), .ZN(n1538) );
  CKNXD0 U1559 ( .I(n1540), .ZN(DataO[17]) );
  CKNXD16 U1560 ( .I(n1543), .ZN(n1540) );
  INVD0 U1561 ( .I(n1542), .ZN(n1543) );
  CKNXD16 U1562 ( .I(n1545), .ZN(n1542) );
  INVD0 U1563 ( .I(n1544), .ZN(n1545) );
  CKNXD16 U1564 ( .I(n1547), .ZN(n1544) );
  INVD0 U1565 ( .I(n1546), .ZN(n1547) );
  CKNXD16 U1566 ( .I(n2273), .ZN(n1546) );
  CKNXD0 U1567 ( .I(n1548), .ZN(n1549) );
  CKNXD16 U1568 ( .I(n1551), .ZN(n1548) );
  INVD0 U1569 ( .I(n1550), .ZN(n1551) );
  CKNXD16 U1570 ( .I(n1553), .ZN(n1550) );
  INVD0 U1571 ( .I(n1552), .ZN(n1553) );
  CKNXD16 U1572 ( .I(n1555), .ZN(n1552) );
  INVD0 U1573 ( .I(n1554), .ZN(n1555) );
  CKNXD16 U1574 ( .I(n2274), .ZN(n1554) );
  CKNXD0 U1575 ( .I(n1556), .ZN(n1557) );
  INVD0 U1576 ( .I(n1558), .ZN(n1559) );
  INVD0 U1577 ( .I(n1560), .ZN(n1561) );
  INVD0 U1578 ( .I(n1562), .ZN(n1563) );
  CKNXD0 U1579 ( .I(n1564), .ZN(n1565) );
  INVD0 U1580 ( .I(n1566), .ZN(n1567) );
  INVD0 U1581 ( .I(n1568), .ZN(n1569) );
  INVD0 U1582 ( .I(n1570), .ZN(n1571) );
  CKNXD0 U1583 ( .I(n1572), .ZN(DataO[13]) );
  CKNXD16 U1584 ( .I(n1575), .ZN(n1572) );
  INVD0 U1585 ( .I(n1574), .ZN(n1575) );
  CKNXD16 U1586 ( .I(n1577), .ZN(n1574) );
  INVD0 U1587 ( .I(n1576), .ZN(n1577) );
  CKNXD16 U1588 ( .I(n1579), .ZN(n1576) );
  INVD0 U1589 ( .I(n1578), .ZN(n1579) );
  CKNXD16 U1590 ( .I(n2277), .ZN(n1578) );
  CKNXD0 U1591 ( .I(n1580), .ZN(DataO[12]) );
  CKNXD16 U1592 ( .I(n1583), .ZN(n1580) );
  INVD0 U1593 ( .I(n1582), .ZN(n1583) );
  CKNXD16 U1594 ( .I(n1585), .ZN(n1582) );
  INVD0 U1595 ( .I(n1584), .ZN(n1585) );
  CKNXD16 U1596 ( .I(n1587), .ZN(n1584) );
  INVD0 U1597 ( .I(n1586), .ZN(n1587) );
  CKNXD16 U1598 ( .I(n2278), .ZN(n1586) );
  CKNXD0 U1599 ( .I(n1588), .ZN(n1589) );
  CKNXD16 U1600 ( .I(n1591), .ZN(n1588) );
  INVD0 U1601 ( .I(n1590), .ZN(n1591) );
  CKNXD16 U1602 ( .I(n1593), .ZN(n1590) );
  INVD0 U1603 ( .I(n1592), .ZN(n1593) );
  CKNXD16 U1604 ( .I(n1595), .ZN(n1592) );
  INVD0 U1605 ( .I(n1594), .ZN(n1595) );
  CKNXD16 U1606 ( .I(n2279), .ZN(n1594) );
  CKNXD0 U1607 ( .I(n1596), .ZN(n1597) );
  INVD0 U1608 ( .I(n1598), .ZN(n1599) );
  INVD0 U1609 ( .I(n1600), .ZN(n1601) );
  INVD0 U1610 ( .I(n1602), .ZN(n1603) );
  CKNXD0 U1611 ( .I(n1604), .ZN(n1605) );
  INVD0 U1612 ( .I(n1606), .ZN(n1607) );
  INVD0 U1613 ( .I(n1608), .ZN(n1609) );
  INVD0 U1614 ( .I(n1610), .ZN(n1611) );
  CKNXD0 U1615 ( .I(n1612), .ZN(DataO[8]) );
  CKNXD16 U1616 ( .I(n1615), .ZN(n1612) );
  INVD0 U1617 ( .I(n1614), .ZN(n1615) );
  CKNXD16 U1618 ( .I(n1617), .ZN(n1614) );
  INVD0 U1619 ( .I(n1616), .ZN(n1617) );
  CKNXD16 U1620 ( .I(n1619), .ZN(n1616) );
  INVD0 U1621 ( .I(n1618), .ZN(n1619) );
  CKNXD16 U1622 ( .I(n2282), .ZN(n1618) );
  CKNXD0 U1623 ( .I(n1620), .ZN(DataO[7]) );
  CKNXD16 U1624 ( .I(n1623), .ZN(n1620) );
  INVD0 U1625 ( .I(n1622), .ZN(n1623) );
  CKNXD16 U1626 ( .I(n1625), .ZN(n1622) );
  INVD0 U1627 ( .I(n1624), .ZN(n1625) );
  CKNXD16 U1628 ( .I(n1627), .ZN(n1624) );
  INVD0 U1629 ( .I(n1626), .ZN(n1627) );
  CKNXD16 U1630 ( .I(n2283), .ZN(n1626) );
  CKNXD0 U1631 ( .I(n1628), .ZN(DataO[6]) );
  CKNXD16 U1632 ( .I(n1631), .ZN(n1628) );
  INVD0 U1633 ( .I(n1630), .ZN(n1631) );
  CKNXD16 U1634 ( .I(n1633), .ZN(n1630) );
  INVD0 U1635 ( .I(n1632), .ZN(n1633) );
  CKNXD16 U1636 ( .I(n1635), .ZN(n1632) );
  INVD0 U1637 ( .I(n1634), .ZN(n1635) );
  CKNXD16 U1638 ( .I(n2284), .ZN(n1634) );
  CKNXD0 U1639 ( .I(n1636), .ZN(n1637) );
  CKNXD16 U1640 ( .I(n1639), .ZN(n1636) );
  INVD0 U1641 ( .I(n1638), .ZN(n1639) );
  CKNXD16 U1642 ( .I(n1641), .ZN(n1638) );
  INVD0 U1643 ( .I(n1640), .ZN(n1641) );
  CKNXD16 U1644 ( .I(n1643), .ZN(n1640) );
  INVD0 U1645 ( .I(n1642), .ZN(n1643) );
  CKNXD16 U1646 ( .I(n2285), .ZN(n1642) );
  CKNXD0 U1647 ( .I(n1644), .ZN(n1645) );
  INVD0 U1648 ( .I(n1646), .ZN(n1647) );
  INVD0 U1649 ( .I(n1648), .ZN(n1649) );
  INVD0 U1650 ( .I(n1650), .ZN(n1651) );
  CKNXD0 U1651 ( .I(n1652), .ZN(n1653) );
  INVD0 U1652 ( .I(n1654), .ZN(n1655) );
  INVD0 U1653 ( .I(n1656), .ZN(n1657) );
  INVD0 U1654 ( .I(n1658), .ZN(n1659) );
  CKNXD0 U1655 ( .I(n1660), .ZN(DataO[2]) );
  CKNXD16 U1656 ( .I(n1663), .ZN(n1660) );
  INVD0 U1657 ( .I(n1662), .ZN(n1663) );
  CKNXD16 U1658 ( .I(n1665), .ZN(n1662) );
  INVD0 U1659 ( .I(n1664), .ZN(n1665) );
  CKNXD16 U1660 ( .I(n1667), .ZN(n1664) );
  INVD0 U1661 ( .I(n1666), .ZN(n1667) );
  CKNXD16 U1662 ( .I(n2288), .ZN(n1666) );
  CKNXD0 U1663 ( .I(n1668), .ZN(DataO[1]) );
  CKNXD16 U1664 ( .I(n1671), .ZN(n1668) );
  INVD0 U1665 ( .I(n1670), .ZN(n1671) );
  CKNXD16 U1666 ( .I(n1673), .ZN(n1670) );
  INVD0 U1667 ( .I(n1672), .ZN(n1673) );
  CKNXD16 U1668 ( .I(n1675), .ZN(n1672) );
  INVD0 U1669 ( .I(n1674), .ZN(n1675) );
  CKNXD16 U1670 ( .I(n2289), .ZN(n1674) );
  CKNXD0 U1671 ( .I(n1676), .ZN(DataO[0]) );
  CKNXD16 U1672 ( .I(n1679), .ZN(n1676) );
  INVD0 U1673 ( .I(n1678), .ZN(n1679) );
  CKNXD16 U1674 ( .I(n1681), .ZN(n1678) );
  INVD0 U1675 ( .I(n1680), .ZN(n1681) );
  CKNXD16 U1676 ( .I(n1683), .ZN(n1680) );
  INVD0 U1677 ( .I(n1682), .ZN(n1683) );
  CKNXD16 U1678 ( .I(n2290), .ZN(n1682) );
  CKAN2D0 U1679 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U1680 ( .I(n2258), .ZN(n2114) );
  BUFFD1 U1681 ( .I(n2176), .Z(n2175) );
  BUFFD1 U1682 ( .I(n2182), .Z(n2151) );
  BUFFD1 U1683 ( .I(n2182), .Z(n2152) );
  BUFFD1 U1684 ( .I(n2182), .Z(n2153) );
  BUFFD1 U1685 ( .I(n2182), .Z(n2154) );
  BUFFD1 U1686 ( .I(n2181), .Z(n2155) );
  BUFFD1 U1687 ( .I(n2181), .Z(n2156) );
  BUFFD1 U1688 ( .I(n2181), .Z(n2157) );
  BUFFD1 U1689 ( .I(n2181), .Z(n2158) );
  BUFFD1 U1690 ( .I(n2180), .Z(n2159) );
  BUFFD1 U1691 ( .I(n2180), .Z(n2160) );
  BUFFD1 U1692 ( .I(n2180), .Z(n2161) );
  BUFFD1 U1693 ( .I(n2180), .Z(n2162) );
  BUFFD1 U1694 ( .I(n2179), .Z(n2163) );
  BUFFD1 U1695 ( .I(n2179), .Z(n2164) );
  BUFFD1 U1696 ( .I(n2179), .Z(n2165) );
  BUFFD1 U1697 ( .I(n2179), .Z(n2166) );
  BUFFD1 U1698 ( .I(n2178), .Z(n2167) );
  BUFFD1 U1699 ( .I(n2178), .Z(n2168) );
  BUFFD1 U1700 ( .I(n2178), .Z(n2169) );
  BUFFD1 U1701 ( .I(n2178), .Z(n2170) );
  BUFFD1 U1702 ( .I(n2177), .Z(n2171) );
  BUFFD1 U1703 ( .I(n2177), .Z(n2172) );
  BUFFD1 U1704 ( .I(n2177), .Z(n2173) );
  BUFFD1 U1705 ( .I(n2177), .Z(n2174) );
  BUFFD1 U1706 ( .I(n2150), .Z(n2176) );
  BUFFD1 U1707 ( .I(n2137), .Z(n2140) );
  BUFFD1 U1708 ( .I(n2137), .Z(n2139) );
  BUFFD1 U1709 ( .I(n2136), .Z(n2141) );
  BUFFD1 U1710 ( .I(n2136), .Z(n2142) );
  BUFFD1 U1711 ( .I(n2135), .Z(n2144) );
  BUFFD1 U1712 ( .I(n2135), .Z(n2145) );
  BUFFD1 U1713 ( .I(n2141), .Z(n2146) );
  BUFFD1 U1714 ( .I(n2135), .Z(n2143) );
  BUFFD1 U1715 ( .I(n2137), .Z(n2138) );
  BUFFD1 U1716 ( .I(N45), .Z(n2127) );
  BUFFD1 U1717 ( .I(n2129), .Z(n2128) );
  BUFFD1 U1718 ( .I(n2125), .Z(n2129) );
  BUFFD1 U1719 ( .I(n2125), .Z(n2130) );
  BUFFD1 U1720 ( .I(n2125), .Z(n2131) );
  BUFFD1 U1721 ( .I(n2124), .Z(n2132) );
  BUFFD1 U1722 ( .I(N45), .Z(n2126) );
  BUFFD1 U1723 ( .I(n2230), .Z(n2229) );
  BUFFD1 U1724 ( .I(n2230), .Z(n2228) );
  BUFFD1 U1725 ( .I(n2231), .Z(n2227) );
  BUFFD1 U1726 ( .I(n2231), .Z(n2226) );
  BUFFD1 U1727 ( .I(n2232), .Z(n2225) );
  BUFFD1 U1728 ( .I(n2232), .Z(n2224) );
  BUFFD1 U1729 ( .I(n2224), .Z(n2223) );
  BUFFD1 U1730 ( .I(n2224), .Z(n2222) );
  BUFFD1 U1731 ( .I(n2233), .Z(n2221) );
  BUFFD1 U1732 ( .I(n2233), .Z(n2220) );
  BUFFD1 U1733 ( .I(n2234), .Z(n2219) );
  BUFFD1 U1734 ( .I(n2234), .Z(n2218) );
  BUFFD1 U1735 ( .I(n2235), .Z(n2217) );
  BUFFD1 U1736 ( .I(n2235), .Z(n2216) );
  BUFFD1 U1737 ( .I(n2236), .Z(n2215) );
  BUFFD1 U1738 ( .I(n2236), .Z(n2214) );
  BUFFD1 U1739 ( .I(n2237), .Z(n2213) );
  BUFFD1 U1740 ( .I(n2237), .Z(n2212) );
  BUFFD1 U1741 ( .I(n2238), .Z(n2211) );
  BUFFD1 U1742 ( .I(n2238), .Z(n2210) );
  BUFFD1 U1743 ( .I(n2239), .Z(n2209) );
  BUFFD1 U1744 ( .I(n2239), .Z(n2208) );
  BUFFD1 U1745 ( .I(n2240), .Z(n2207) );
  BUFFD1 U1746 ( .I(n2240), .Z(n2206) );
  BUFFD1 U1747 ( .I(n2241), .Z(n2205) );
  BUFFD1 U1748 ( .I(n2241), .Z(n2204) );
  BUFFD1 U1749 ( .I(n2242), .Z(n2203) );
  BUFFD1 U1750 ( .I(n2242), .Z(n2202) );
  BUFFD1 U1751 ( .I(n2243), .Z(n2201) );
  BUFFD1 U1752 ( .I(n2243), .Z(n2200) );
  BUFFD1 U1753 ( .I(n2244), .Z(n2199) );
  BUFFD1 U1754 ( .I(n2244), .Z(n2198) );
  BUFFD1 U1755 ( .I(n2245), .Z(n2197) );
  BUFFD1 U1756 ( .I(n2245), .Z(n2196) );
  BUFFD1 U1757 ( .I(n2246), .Z(n2195) );
  BUFFD1 U1758 ( .I(n2246), .Z(n2194) );
  BUFFD1 U1759 ( .I(n2247), .Z(n2193) );
  BUFFD1 U1760 ( .I(n2247), .Z(n2192) );
  BUFFD1 U1761 ( .I(n2248), .Z(n2191) );
  BUFFD1 U1762 ( .I(n2248), .Z(n2190) );
  BUFFD1 U1763 ( .I(n2249), .Z(n2189) );
  BUFFD1 U1764 ( .I(n2249), .Z(n2188) );
  BUFFD1 U1765 ( .I(n2183), .Z(n2181) );
  BUFFD1 U1766 ( .I(n2184), .Z(n2180) );
  BUFFD1 U1767 ( .I(n2184), .Z(n2179) );
  BUFFD1 U1768 ( .I(n2185), .Z(n2178) );
  BUFFD1 U1769 ( .I(n2185), .Z(n2177) );
  BUFFD1 U1770 ( .I(n2183), .Z(n2182) );
  BUFFD1 U1771 ( .I(N45), .Z(n2125) );
  BUFFD1 U1772 ( .I(N45), .Z(n2124) );
  BUFFD1 U1773 ( .I(n2133), .Z(n2137) );
  BUFFD1 U1774 ( .I(n2223), .Z(n2230) );
  BUFFD1 U1775 ( .I(n2222), .Z(n2231) );
  BUFFD1 U1776 ( .I(n2255), .Z(n2232) );
  BUFFD1 U1777 ( .I(n2216), .Z(n2233) );
  BUFFD1 U1778 ( .I(n2189), .Z(n2234) );
  BUFFD1 U1779 ( .I(n2254), .Z(n2235) );
  BUFFD1 U1780 ( .I(n2254), .Z(n2236) );
  BUFFD1 U1781 ( .I(n2254), .Z(n2237) );
  BUFFD1 U1782 ( .I(n2253), .Z(n2238) );
  BUFFD1 U1783 ( .I(n2253), .Z(n2239) );
  BUFFD1 U1784 ( .I(n2253), .Z(n2240) );
  BUFFD1 U1785 ( .I(n2252), .Z(n2241) );
  BUFFD1 U1786 ( .I(n2252), .Z(n2242) );
  BUFFD1 U1787 ( .I(n2252), .Z(n2243) );
  BUFFD1 U1788 ( .I(n2251), .Z(n2244) );
  BUFFD1 U1789 ( .I(n2251), .Z(n2245) );
  BUFFD1 U1790 ( .I(n2251), .Z(n2246) );
  BUFFD1 U1791 ( .I(n2250), .Z(n2247) );
  BUFFD1 U1792 ( .I(n2250), .Z(n2248) );
  BUFFD1 U1793 ( .I(n2250), .Z(n2249) );
  BUFFD1 U1794 ( .I(n2148), .Z(n2184) );
  BUFFD1 U1795 ( .I(n2148), .Z(n2185) );
  BUFFD1 U1796 ( .I(n2148), .Z(n2183) );
  BUFFD1 U1797 ( .I(n2118), .Z(n2122) );
  BUFFD1 U1798 ( .I(n2118), .Z(n2123) );
  BUFFD1 U1799 ( .I(n2120), .Z(n2121) );
  BUFFD1 U1800 ( .I(n2119), .Z(n2120) );
  BUFFD1 U1801 ( .I(n2257), .Z(n2117) );
  BUFFD1 U1802 ( .I(n2257), .Z(n2116) );
  BUFFD1 U1803 ( .I(N44), .Z(n2134) );
  BUFFD1 U1804 ( .I(N44), .Z(n2133) );
  BUFFD1 U1805 ( .I(n2201), .Z(n2255) );
  BUFFD1 U1806 ( .I(n2255), .Z(n2254) );
  BUFFD1 U1807 ( .I(n2186), .Z(n2253) );
  BUFFD1 U1808 ( .I(n2186), .Z(n2252) );
  BUFFD1 U1809 ( .I(n2221), .Z(n2251) );
  BUFFD1 U1810 ( .I(n2217), .Z(n2250) );
  BUFFD1 U1811 ( .I(n108), .Z(n2150) );
  XOR3D1 U1812 ( .A1(n96), .A2(n558), .A3(n257), .Z(n95) );
  BUFFD1 U1813 ( .I(N46), .Z(n2119) );
  INVD1 U1814 ( .I(n2114), .ZN(n2115) );
  XOR3D1 U1815 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n73), .Z(N85) );
  XOR3D1 U1816 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n73), .Z(n2147) );
  XOR3D1 U1817 ( .A1(DataI[0]), .A2(n74), .A3(n75), .Z(n73) );
  XOR3D1 U1818 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n76), .Z(n75) );
  XOR3D1 U1819 ( .A1(n77), .A2(DataI[3]), .A3(n78), .Z(n76) );
  XOR3D1 U1820 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n79), .Z(n78) );
  XOR3D1 U1821 ( .A1(n80), .A2(DataI[10]), .A3(n81), .Z(n79) );
  XOR3D1 U1822 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n82), .Z(n81) );
  XOR3D1 U1823 ( .A1(n83), .A2(DataI[17]), .A3(n84), .Z(n82) );
  BUFFD1 U1824 ( .I(n2187), .Z(n2186) );
  INVD1 U1825 ( .I(Reset), .ZN(n108) );
  BUFFD1 U1826 ( .I(N48), .Z(n2258) );
  ND3D1 U1827 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U1828 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  INVD1 U1829 ( .I(AddrW[2]), .ZN(n105) );
  BUFFD1 U1830 ( .I(ClockW), .Z(n2187) );
  MUX4ND0 U1831 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n2142), .S1(n2125), 
        .ZN(n2104) );
  MUX4ND0 U1832 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n2142), .S1(n2126), .ZN(
        n1714) );
  MUX4ND0 U1833 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n2138), .S1(n2124), .ZN(
        n1740) );
  MUX4ND0 U1834 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n2142), .S1(N45), .ZN(
        n1753) );
  MUX4ND0 U1835 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n2138), .S1(N45), .ZN(
        n1766) );
  MUX4ND0 U1836 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n2138), .S1(n2127), .ZN(
        n1779) );
  MUX4ND0 U1837 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n2142), .S1(n2130), 
        .ZN(n1818) );
  MUX4ND0 U1838 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n2142), .S1(n2127), 
        .ZN(n1831) );
  MUX4ND0 U1839 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n2142), .S1(n2124), 
        .ZN(n1844) );
  MUX4ND0 U1840 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n2141), .S1(n2125), 
        .ZN(n1857) );
  MUX4ND0 U1841 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n2141), .S1(n2129), 
        .ZN(n1870) );
  MUX4ND0 U1842 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n2141), .S1(n2126), 
        .ZN(n1883) );
  MUX4ND0 U1843 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n2141), .S1(n2128), 
        .ZN(n1896) );
  MUX4ND0 U1844 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n2141), .S1(n2124), 
        .ZN(n1909) );
  MUX4ND0 U1845 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n2141), .S1(n2124), 
        .ZN(n1922) );
  MUX4ND0 U1846 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n2141), .S1(n2132), 
        .ZN(n1935) );
  MUX4ND0 U1847 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n2141), .S1(N45), .ZN(
        n1948) );
  MUX4ND0 U1848 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n2141), .S1(n2126), 
        .ZN(n1961) );
  MUX4ND0 U1849 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n2141), .S1(n2124), 
        .ZN(n1974) );
  MUX4ND0 U1850 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n2141), .S1(n2126), 
        .ZN(n1987) );
  MUX4ND0 U1851 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n2141), .S1(n2132), 
        .ZN(n2000) );
  MUX4ND0 U1852 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n2141), .S1(n2130), 
        .ZN(n2013) );
  MUX4ND0 U1853 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n2142), .S1(n2126), .ZN(
        n1688) );
  MUX4ND0 U1854 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n2138), .S1(n2126), .ZN(
        n1701) );
  MUX4ND0 U1855 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n2141), .S1(n2131), 
        .ZN(n2026) );
  MUX4ND0 U1856 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n2142), .S1(n2125), 
        .ZN(n2039) );
  MUX4ND0 U1857 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n2142), .S1(N45), .ZN(
        n2052) );
  MUX4ND0 U1858 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n2142), .S1(n2124), 
        .ZN(n2065) );
  MUX4ND0 U1859 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n2142), .S1(n2124), 
        .ZN(n2078) );
  MUX4ND0 U1860 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n2142), .S1(N45), .ZN(
        n2091) );
  MUX4D0 U1861 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n2142), .S1(n2132), 
        .Z(n2105) );
  MUX4D0 U1862 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n2134), .S1(n2128), .Z(
        n1689) );
  MUX4D0 U1863 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n2144), .S1(n2132), .Z(
        n1702) );
  MUX4D0 U1864 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n2144), .S1(n2124), .Z(
        n1715) );
  MUX4D0 U1865 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n2145), .S1(n2126), .Z(
        n1741) );
  MUX4D0 U1866 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n2146), .S1(n2127), .Z(
        n1780) );
  MUX4D0 U1867 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n2146), .S1(n2124), 
        .Z(n1819) );
  MUX4D0 U1868 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n2145), .S1(n2126), 
        .Z(n1832) );
  MUX4D0 U1869 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(N44), .S1(n2125), .Z(
        n1845) );
  MUX4D0 U1870 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(N44), .S1(n2124), .Z(
        n1858) );
  MUX4D0 U1871 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(N44), .S1(n2125), .Z(
        n1871) );
  MUX4D0 U1872 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n2143), .S1(n2130), 
        .Z(n1884) );
  MUX4D0 U1873 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n2141), .S1(N45), .Z(
        n1897) );
  MUX4D0 U1874 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n2145), .S1(N45), .Z(
        n1910) );
  MUX4D0 U1875 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n2137), .S1(n2126), 
        .Z(n1923) );
  MUX4D0 U1876 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n2134), .S1(n2126), 
        .Z(n1936) );
  MUX4D0 U1877 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n2136), .S1(n2127), 
        .Z(n1949) );
  MUX4D0 U1878 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n2137), .S1(n2127), 
        .Z(n1962) );
  MUX4D0 U1879 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n2145), .S1(n2128), 
        .Z(n1975) );
  MUX4D0 U1880 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n2144), .S1(n2128), 
        .Z(n1988) );
  MUX4D0 U1881 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n2133), .S1(n2129), 
        .Z(n2001) );
  MUX4D0 U1882 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n2143), .S1(n2129), 
        .Z(n2014) );
  MUX4D0 U1883 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n2137), .S1(n2130), 
        .Z(n2027) );
  MUX4D0 U1884 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n2136), .S1(n2130), 
        .Z(n2040) );
  MUX4D0 U1885 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n2137), .S1(n2131), 
        .Z(n2053) );
  MUX4D0 U1886 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n2134), .S1(n2131), 
        .Z(n2066) );
  MUX4D0 U1887 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n2133), .S1(n2131), 
        .Z(n2079) );
  MUX4D0 U1888 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n2134), .S1(n2132), 
        .Z(n2092) );
  MUX4D0 U1889 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n2142), .S1(n2130), .Z(
        n2109) );
  MUX4D0 U1890 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n2142), .S1(n2129), 
        .Z(n2107) );
  MUX4D0 U1891 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n2143), .S1(n2132), .Z(
        n1693) );
  MUX4D0 U1892 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n2143), .S1(n2131), .Z(
        n1691) );
  MUX4D0 U1893 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n2144), .S1(n2129), .Z(
        n1706) );
  MUX4D0 U1894 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n2144), .S1(n2132), .Z(
        n1704) );
  MUX4D0 U1895 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n2144), .S1(n2125), .Z(
        n1719) );
  MUX4D0 U1896 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n2144), .S1(n2124), .Z(
        n1717) );
  MUX4D0 U1897 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n2145), .S1(n2132), .Z(
        n1745) );
  MUX4D0 U1898 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n2145), .S1(n2124), .Z(
        n1743) );
  MUX4D0 U1899 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(N44), .S1(n2128), .Z(n1758) );
  MUX4D0 U1900 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n2134), .S1(n2130), .Z(
        n1771) );
  MUX4D0 U1901 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n2133), .S1(n2127), .Z(
        n1769) );
  MUX4D0 U1902 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n2134), .S1(n2125), .Z(
        n1784) );
  MUX4D0 U1903 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n2146), .S1(n2126), .Z(
        n1782) );
  MUX4D0 U1904 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n2146), .S1(n2127), .Z(
        n1823) );
  MUX4D0 U1905 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n2146), .S1(N45), .Z(
        n1821) );
  MUX4D0 U1906 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(N44), .S1(n2126), .Z(
        n1836) );
  MUX4D0 U1907 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(N44), .S1(n2127), .Z(
        n1834) );
  MUX4D0 U1908 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(N44), .S1(n2124), .Z(
        n1849) );
  MUX4D0 U1909 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(N44), .S1(n2124), .Z(
        n1847) );
  MUX4D0 U1910 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n2136), .S1(n2125), .Z(
        n1862) );
  MUX4D0 U1911 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n2133), .S1(n2125), 
        .Z(n1860) );
  MUX4D0 U1912 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(N44), .S1(n2125), .Z(
        n1875) );
  MUX4D0 U1913 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n2133), .S1(n2124), 
        .Z(n1873) );
  MUX4D0 U1914 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n2135), .S1(n2124), .Z(
        n1888) );
  MUX4D0 U1915 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n2143), .S1(n2125), 
        .Z(n1886) );
  MUX4D0 U1916 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n2141), .S1(n2132), .Z(
        n1901) );
  MUX4D0 U1917 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n2135), .S1(n2130), 
        .Z(n1899) );
  MUX4D0 U1918 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n2139), .S1(n2127), .Z(
        n1914) );
  MUX4D0 U1919 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n2137), .S1(N45), .Z(
        n1912) );
  MUX4D0 U1920 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n2144), .S1(n2126), .Z(
        n1927) );
  MUX4D0 U1921 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n2144), .S1(n2126), 
        .Z(n1925) );
  MUX4D0 U1922 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n2145), .S1(n2127), .Z(
        n1940) );
  MUX4D0 U1923 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n2136), .S1(n2126), 
        .Z(n1938) );
  MUX4D0 U1924 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n2137), .S1(n2127), .Z(
        n1953) );
  MUX4D0 U1925 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n2137), .S1(n2127), 
        .Z(n1951) );
  MUX4D0 U1926 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n2144), .S1(n2128), .Z(
        n1966) );
  MUX4D0 U1927 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n2145), .S1(n2127), 
        .Z(n1964) );
  MUX4D0 U1928 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n2141), .S1(n2128), .Z(
        n1979) );
  MUX4D0 U1929 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n2136), .S1(n2128), 
        .Z(n1977) );
  MUX4D0 U1930 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n2140), .S1(n2128), .Z(
        n1992) );
  MUX4D0 U1931 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n2141), .S1(n2128), 
        .Z(n1990) );
  MUX4D0 U1932 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n2143), .S1(n2129), .Z(
        n2005) );
  MUX4D0 U1933 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n2143), .S1(n2129), 
        .Z(n2003) );
  MUX4D0 U1934 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n2143), .S1(n2129), .Z(
        n2018) );
  MUX4D0 U1935 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n2143), .S1(n2129), 
        .Z(n2016) );
  MUX4D0 U1936 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n2133), .S1(n2130), .Z(
        n2031) );
  MUX4D0 U1937 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n2133), .S1(n2130), 
        .Z(n2029) );
  MUX4D0 U1938 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n2133), .S1(n2130), .Z(
        n2044) );
  MUX4D0 U1939 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n2133), .S1(n2130), 
        .Z(n2042) );
  MUX4D0 U1940 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n2137), .S1(n2131), .Z(
        n2057) );
  MUX4D0 U1941 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n2137), .S1(n2131), 
        .Z(n2055) );
  MUX4D0 U1942 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n2134), .S1(n2131), .Z(
        n2070) );
  MUX4D0 U1943 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n2134), .S1(n2131), 
        .Z(n2068) );
  MUX4D0 U1944 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n2133), .S1(n2132), .Z(
        n2083) );
  MUX4D0 U1945 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n2137), .S1(n2132), 
        .Z(n2081) );
  MUX4D0 U1946 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n2133), .S1(n2132), .Z(
        n2096) );
  MUX4D0 U1947 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n2133), .S1(n2132), 
        .Z(n2094) );
  MUX4D0 U1948 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n2142), .S1(n2132), 
        .Z(n2106) );
  MUX4D0 U1949 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n2146), .S1(n2132), .Z(
        n1690) );
  MUX4D0 U1950 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n2144), .S1(n2125), .Z(
        n1703) );
  MUX4D0 U1951 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n2144), .S1(n2125), .Z(
        n1716) );
  MUX4D0 U1952 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n2145), .S1(N45), .Z(
        n1742) );
  MUX4D0 U1953 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n2134), .S1(N45), .Z(
        n1755) );
  MUX4D0 U1954 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n2134), .S1(N45), .Z(
        n1768) );
  MUX4D0 U1955 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n2133), .S1(n2132), .Z(
        n1781) );
  MUX4D0 U1956 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n2146), .S1(n2128), 
        .Z(n1820) );
  MUX4D0 U1957 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n2144), .S1(n2127), 
        .Z(n1833) );
  MUX4D0 U1958 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(N44), .S1(n2126), .Z(
        n1846) );
  MUX4D0 U1959 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n2134), .S1(n2125), 
        .Z(n1859) );
  MUX4D0 U1960 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(N44), .S1(n2127), .Z(
        n1872) );
  MUX4D0 U1961 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n2135), .S1(n2130), 
        .Z(n1885) );
  MUX4D0 U1962 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n2135), .S1(n2128), 
        .Z(n1898) );
  MUX4D0 U1963 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n2137), .S1(n2124), 
        .Z(n1911) );
  MUX4D0 U1964 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n2136), .S1(n2126), 
        .Z(n1924) );
  MUX4D0 U1965 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n2144), .S1(n2126), 
        .Z(n1937) );
  MUX4D0 U1966 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n2145), .S1(n2127), 
        .Z(n1950) );
  MUX4D0 U1967 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n2141), .S1(n2127), 
        .Z(n1963) );
  MUX4D0 U1968 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n2139), .S1(n2128), 
        .Z(n1976) );
  MUX4D0 U1969 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n2143), .S1(n2128), 
        .Z(n1989) );
  MUX4D0 U1970 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n2143), .S1(n2129), 
        .Z(n2002) );
  MUX4D0 U1971 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n2143), .S1(n2129), 
        .Z(n2015) );
  MUX4D0 U1972 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n2133), .S1(n2130), 
        .Z(n2028) );
  MUX4D0 U1973 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n2137), .S1(n2130), 
        .Z(n2041) );
  MUX4D0 U1974 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n2137), .S1(n2131), 
        .Z(n2054) );
  MUX4D0 U1975 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n2134), .S1(n2131), 
        .Z(n2067) );
  MUX4D0 U1976 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n2134), .S1(n2132), 
        .Z(n2080) );
  MUX4D0 U1977 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n2134), .S1(n2132), 
        .Z(n2093) );
  MUX4D0 U1978 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n2142), .S1(n2132), .Z(
        n2110) );
  MUX4D0 U1979 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n2142), .S1(n2132), 
        .Z(n2108) );
  MUX4D0 U1980 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n2143), .S1(n2125), .Z(
        n1694) );
  MUX4D0 U1981 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n2143), .S1(n2129), .Z(
        n1692) );
  MUX4D0 U1982 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n2144), .S1(n2124), .Z(
        n1707) );
  MUX4D0 U1983 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n2144), .S1(n2125), .Z(
        n1705) );
  MUX4D0 U1984 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n2144), .S1(n2130), .Z(
        n1720) );
  MUX4D0 U1985 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n2144), .S1(n2131), .Z(
        n1718) );
  MUX4D0 U1986 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n2145), .S1(n2125), .Z(
        n1746) );
  MUX4D0 U1987 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n2145), .S1(N45), .Z(
        n1744) );
  MUX4D0 U1988 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n2140), .S1(n2124), .Z(
        n1759) );
  MUX4D0 U1989 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n2137), .S1(n2125), .Z(
        n1757) );
  MUX4D0 U1990 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n2146), .S1(n2130), .Z(
        n1772) );
  MUX4D0 U1991 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n2133), .S1(n2128), .Z(
        n1770) );
  MUX4D0 U1992 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n2146), .S1(n2126), .Z(
        n1785) );
  MUX4D0 U1993 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n2146), .S1(n2132), .Z(
        n1783) );
  MUX4D0 U1994 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n2146), .S1(n2126), .Z(
        n1824) );
  MUX4D0 U1995 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n2146), .S1(n2128), 
        .Z(n1822) );
  MUX4D0 U1996 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n2145), .S1(n2128), .Z(
        n1837) );
  MUX4D0 U1997 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n2144), .S1(n2128), 
        .Z(n1835) );
  MUX4D0 U1998 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n2137), .S1(n2124), .Z(
        n1850) );
  MUX4D0 U1999 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n2133), .S1(n2124), 
        .Z(n1848) );
  MUX4D0 U2000 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n2137), .S1(n2125), .Z(
        n1863) );
  MUX4D0 U2001 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n2134), .S1(n2125), 
        .Z(n1861) );
  MUX4D0 U2002 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n2141), .S1(n2124), .Z(
        n1876) );
  MUX4D0 U2003 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(N44), .S1(n2124), .Z(
        n1874) );
  MUX4D0 U2004 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n2135), .S1(n2131), .Z(
        n1889) );
  MUX4D0 U2005 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n2135), .S1(n2131), 
        .Z(n1887) );
  MUX4D0 U2006 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n2143), .S1(n2131), .Z(
        n1902) );
  MUX4D0 U2007 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n2135), .S1(n2124), 
        .Z(n1900) );
  MUX4D0 U2008 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n2136), .S1(n2126), .Z(
        n1915) );
  MUX4D0 U2009 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n2141), .S1(n2128), 
        .Z(n1913) );
  MUX4D0 U2010 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n2145), .S1(n2126), .Z(
        n1928) );
  MUX4D0 U2011 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n2143), .S1(n2126), 
        .Z(n1926) );
  MUX4D0 U2012 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n2139), .S1(n2127), .Z(
        n1941) );
  MUX4D0 U2013 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n2144), .S1(n2127), 
        .Z(n1939) );
  MUX4D0 U2014 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n2142), .S1(n2127), .Z(
        n1954) );
  MUX4D0 U2015 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n2144), .S1(n2127), 
        .Z(n1952) );
  MUX4D0 U2016 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n2138), .S1(n2128), .Z(
        n1967) );
  MUX4D0 U2017 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n2137), .S1(n2127), 
        .Z(n1965) );
  MUX4D0 U2018 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n2135), .S1(n2128), .Z(
        n1980) );
  MUX4D0 U2019 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n2134), .S1(n2128), 
        .Z(n1978) );
  MUX4D0 U2020 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n2134), .S1(n2129), .Z(
        n1993) );
  MUX4D0 U2021 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n2145), .S1(n2128), 
        .Z(n1991) );
  MUX4D0 U2022 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n2143), .S1(n2129), .Z(
        n2006) );
  MUX4D0 U2023 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n2143), .S1(n2129), 
        .Z(n2004) );
  MUX4D0 U2024 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n2143), .S1(n2130), .Z(
        n2019) );
  MUX4D0 U2025 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n2143), .S1(n2129), 
        .Z(n2017) );
  MUX4D0 U2026 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n2137), .S1(n2130), .Z(
        n2032) );
  MUX4D0 U2027 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n2136), .S1(n2130), 
        .Z(n2030) );
  MUX4D0 U2028 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n2133), .S1(n2130), .Z(
        n2045) );
  MUX4D0 U2029 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n2133), .S1(n2130), 
        .Z(n2043) );
  MUX4D0 U2030 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n2137), .S1(n2131), .Z(
        n2058) );
  MUX4D0 U2031 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n2138), .S1(n2131), 
        .Z(n2056) );
  MUX4D0 U2032 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n2134), .S1(n2131), .Z(
        n2071) );
  MUX4D0 U2033 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n2134), .S1(n2131), 
        .Z(n2069) );
  MUX4D0 U2034 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n2137), .S1(n2132), .Z(
        n2084) );
  MUX4D0 U2035 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n2136), .S1(n2132), 
        .Z(n2082) );
  MUX4D0 U2036 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n2133), .S1(n2132), .Z(
        n2097) );
  MUX4D0 U2037 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n2134), .S1(n2132), 
        .Z(n2095) );
  MUX4ND0 U2038 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n2138), .S1(n2125), .ZN(
        n1727) );
  MUX4ND0 U2039 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n2142), .S1(n2131), .ZN(
        n1792) );
  MUX4ND0 U2040 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n2138), .S1(n2125), .ZN(
        n1805) );
  MUX4D0 U2041 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n2145), .S1(n2124), .Z(
        n1728) );
  MUX4D0 U2042 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n2140), .S1(n2129), .Z(
        n1754) );
  MUX4D0 U2043 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n2133), .S1(n2126), .Z(
        n1767) );
  MUX4D0 U2044 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n2146), .S1(N45), .Z(
        n1793) );
  MUX4D0 U2045 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n2146), .S1(n2130), .Z(
        n1806) );
  MUX4D0 U2046 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n2145), .S1(n2125), .Z(
        n1732) );
  MUX4D0 U2047 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n2145), .S1(n2124), .Z(
        n1730) );
  MUX4D0 U2048 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(N44), .S1(N45), .Z(n1756) );
  MUX4D0 U2049 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n2146), .S1(N45), .Z(n1797) );
  MUX4D0 U2050 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n2146), .S1(n2129), .Z(
        n1795) );
  MUX4D0 U2051 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n2146), .S1(n2127), .Z(
        n1810) );
  MUX4D0 U2052 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n2146), .S1(n2129), .Z(
        n1808) );
  MUX4D0 U2053 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n2145), .S1(n2125), .Z(
        n1729) );
  MUX4D0 U2054 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n2143), .S1(n2125), .Z(
        n1794) );
  MUX4D0 U2055 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n2146), .S1(n2124), .Z(
        n1807) );
  MUX4D0 U2056 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n2145), .S1(N45), .Z(n1733) );
  MUX4D0 U2057 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n2145), .S1(n2124), .Z(
        n1731) );
  MUX4D0 U2058 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(N44), .S1(N45), .Z(n1798)
         );
  MUX4D0 U2059 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n2135), .S1(n2126), .Z(
        n1796) );
  MUX4D0 U2060 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n2146), .S1(n2125), .Z(
        n1811) );
  MUX4D0 U2061 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n2146), .S1(n2128), .Z(
        n1809) );
  ND3D1 U2062 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U2063 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U2064 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U2065 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U2066 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U2067 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U2068 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U2069 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  ND3D1 U2070 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U2071 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U2072 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U2073 ( .I(AddrW[1]), .ZN(n106) );
  INVD1 U2074 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U2075 ( .I(AddrW[4]), .ZN(n102) );
  AN2D1 U2076 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  CKAN2D0 U2077 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX3ND0 U2078 ( .I0(n1686), .I1(n1687), .I2(n1688), .S0(n2125), .S1(n2120), 
        .ZN(n1685) );
  MUX3ND0 U2079 ( .I0(n1699), .I1(n1700), .I2(n1701), .S0(n2126), .S1(N46), 
        .ZN(n1698) );
  MUX3ND0 U2080 ( .I0(n1712), .I1(n1713), .I2(n1714), .S0(n2127), .S1(n2120), 
        .ZN(n1711) );
  MUX3ND0 U2081 ( .I0(n1725), .I1(n1726), .I2(n1727), .S0(n2131), .S1(n2120), 
        .ZN(n1724) );
  MUX3ND0 U2082 ( .I0(n1738), .I1(n1739), .I2(n1740), .S0(n2124), .S1(n2120), 
        .ZN(n1737) );
  MUX3ND0 U2083 ( .I0(n1751), .I1(n1752), .I2(n1753), .S0(n2128), .S1(n2120), 
        .ZN(n1750) );
  MUX3ND0 U2084 ( .I0(n1764), .I1(n1765), .I2(n1766), .S0(n2127), .S1(n2120), 
        .ZN(n1763) );
  MUX3ND0 U2085 ( .I0(n1777), .I1(n1778), .I2(n1779), .S0(n2126), .S1(n2120), 
        .ZN(n1776) );
  MUX3ND0 U2086 ( .I0(n1790), .I1(n1791), .I2(n1792), .S0(n2130), .S1(n2120), 
        .ZN(n1789) );
  MUX3ND0 U2087 ( .I0(n1803), .I1(n1804), .I2(n1805), .S0(n2127), .S1(n2120), 
        .ZN(n1802) );
  MUX3ND0 U2088 ( .I0(n1816), .I1(n1817), .I2(n1818), .S0(n2130), .S1(n2120), 
        .ZN(n1815) );
  MUX3ND0 U2089 ( .I0(n1829), .I1(n1830), .I2(n1831), .S0(n2128), .S1(n2120), 
        .ZN(n1828) );
  MUX3ND0 U2090 ( .I0(n1842), .I1(n1843), .I2(n1844), .S0(n2127), .S1(n2120), 
        .ZN(n1841) );
  MUX3ND0 U2091 ( .I0(n1855), .I1(n1856), .I2(n1857), .S0(n2128), .S1(n2120), 
        .ZN(n1854) );
  MUX3ND0 U2092 ( .I0(n1868), .I1(n1869), .I2(n1870), .S0(n2125), .S1(n2120), 
        .ZN(n1867) );
  MUX3ND0 U2093 ( .I0(n1881), .I1(n1882), .I2(n1883), .S0(n2126), .S1(n2118), 
        .ZN(n1880) );
  MUX3ND0 U2094 ( .I0(n1894), .I1(n1895), .I2(n1896), .S0(n2124), .S1(n2119), 
        .ZN(n1893) );
  MUX3ND0 U2095 ( .I0(n1907), .I1(n1908), .I2(n1909), .S0(n2129), .S1(n2119), 
        .ZN(n1906) );
  MUX3ND0 U2096 ( .I0(n1920), .I1(n1921), .I2(n1922), .S0(n2126), .S1(n2119), 
        .ZN(n1919) );
  MUX3ND0 U2097 ( .I0(n1933), .I1(n1934), .I2(n1935), .S0(n2126), .S1(n2119), 
        .ZN(n1932) );
  MUX3ND0 U2098 ( .I0(n1946), .I1(n1947), .I2(n1948), .S0(n2127), .S1(n2118), 
        .ZN(n1945) );
  MUX3ND0 U2099 ( .I0(n1959), .I1(n1960), .I2(n1961), .S0(n2128), .S1(n2118), 
        .ZN(n1958) );
  MUX3ND0 U2100 ( .I0(n1972), .I1(n1973), .I2(n1974), .S0(n2127), .S1(n2119), 
        .ZN(n1971) );
  MUX3ND0 U2101 ( .I0(n1985), .I1(n1986), .I2(n1987), .S0(n2128), .S1(n2118), 
        .ZN(n1984) );
  MUX3ND0 U2102 ( .I0(n1998), .I1(n1999), .I2(n2000), .S0(n2127), .S1(n2122), 
        .ZN(n1997) );
  MUX3ND0 U2103 ( .I0(n2011), .I1(n2012), .I2(n2013), .S0(n2129), .S1(n2119), 
        .ZN(n2010) );
  MUX3ND0 U2104 ( .I0(n2024), .I1(n2025), .I2(n2026), .S0(n2129), .S1(n2119), 
        .ZN(n2023) );
  MUX3ND0 U2105 ( .I0(n2037), .I1(n2038), .I2(n2039), .S0(n2129), .S1(n2119), 
        .ZN(n2036) );
  MUX3ND0 U2106 ( .I0(n2050), .I1(n2051), .I2(n2052), .S0(n2129), .S1(n2122), 
        .ZN(n2049) );
  MUX3ND0 U2107 ( .I0(n2063), .I1(n2064), .I2(n2065), .S0(N45), .S1(N46), .ZN(
        n2062) );
  MUX3ND0 U2108 ( .I0(n2076), .I1(n2077), .I2(n2078), .S0(n2129), .S1(n2119), 
        .ZN(n2075) );
  MUX3ND0 U2109 ( .I0(n2089), .I1(n2090), .I2(n2091), .S0(n2130), .S1(n2119), 
        .ZN(n2088) );
  MUX3ND0 U2110 ( .I0(n2102), .I1(n2103), .I2(n2104), .S0(n2128), .S1(n2120), 
        .ZN(n2101) );
  MUX3ND0 U2111 ( .I0(n2111), .I1(n2112), .I2(n2113), .S0(N47), .S1(n2115), 
        .ZN(N50) );
  MUX2ND0 U2112 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n2138), 
        .ZN(n1687) );
  MUX2ND0 U2113 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n2138), 
        .ZN(n1686) );
  MUX3ND0 U2114 ( .I0(n1690), .I1(n1689), .I2(n1685), .S0(n2123), .S1(N47), 
        .ZN(n1697) );
  MUX2ND0 U2115 ( .I0(n1692), .I1(n1691), .S(n2121), .ZN(n1696) );
  MUX2ND0 U2116 ( .I0(n1694), .I1(n1693), .S(n2121), .ZN(n1695) );
  MUX2ND0 U2117 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n2138), 
        .ZN(n1700) );
  MUX2ND0 U2118 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n2138), 
        .ZN(n1699) );
  MUX3ND0 U2119 ( .I0(n1703), .I1(n1702), .I2(n1698), .S0(n2123), .S1(n2257), 
        .ZN(n1710) );
  MUX2ND0 U2120 ( .I0(n1705), .I1(n1704), .S(n2120), .ZN(n1709) );
  MUX2ND0 U2121 ( .I0(n1707), .I1(n1706), .S(n2121), .ZN(n1708) );
  MUX2ND0 U2122 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n2138), 
        .ZN(n1713) );
  MUX2ND0 U2123 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n2139), 
        .ZN(n1712) );
  MUX3ND0 U2124 ( .I0(n1716), .I1(n1715), .I2(n1711), .S0(n2123), .S1(N47), 
        .ZN(n1723) );
  MUX2ND0 U2125 ( .I0(n1718), .I1(n1717), .S(n2121), .ZN(n1722) );
  MUX2ND0 U2126 ( .I0(n1720), .I1(n1719), .S(n2121), .ZN(n1721) );
  MUX2ND0 U2127 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n2139), 
        .ZN(n1726) );
  MUX2ND0 U2128 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n2139), 
        .ZN(n1725) );
  MUX3ND0 U2129 ( .I0(n1729), .I1(n1728), .I2(n1724), .S0(n2123), .S1(N47), 
        .ZN(n1736) );
  MUX2ND0 U2130 ( .I0(n1731), .I1(n1730), .S(n2121), .ZN(n1735) );
  MUX2ND0 U2131 ( .I0(n1733), .I1(n1732), .S(n2121), .ZN(n1734) );
  MUX2ND0 U2132 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n2139), 
        .ZN(n1739) );
  MUX2ND0 U2133 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n2139), 
        .ZN(n1738) );
  MUX3ND0 U2134 ( .I0(n1742), .I1(n1741), .I2(n1737), .S0(n2123), .S1(N47), 
        .ZN(n1749) );
  MUX2ND0 U2135 ( .I0(n1744), .I1(n1743), .S(n2121), .ZN(n1748) );
  MUX2ND0 U2136 ( .I0(n1746), .I1(n1745), .S(n2121), .ZN(n1747) );
  MUX2ND0 U2137 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n2139), 
        .ZN(n1752) );
  MUX2ND0 U2138 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n2140), 
        .ZN(n1751) );
  MUX3ND0 U2139 ( .I0(n1755), .I1(n1754), .I2(n1750), .S0(n2122), .S1(N47), 
        .ZN(n1762) );
  MUX2ND0 U2140 ( .I0(n1757), .I1(n1756), .S(n2121), .ZN(n1761) );
  MUX2ND0 U2141 ( .I0(n1759), .I1(n1758), .S(n2121), .ZN(n1760) );
  MUX2ND0 U2142 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n2140), 
        .ZN(n1765) );
  MUX2ND0 U2143 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n2140), 
        .ZN(n1764) );
  MUX3ND0 U2144 ( .I0(n1768), .I1(n1767), .I2(n1763), .S0(n2122), .S1(n2116), 
        .ZN(n1775) );
  MUX2ND0 U2145 ( .I0(n1770), .I1(n1769), .S(n2121), .ZN(n1774) );
  MUX2ND0 U2146 ( .I0(n1772), .I1(n1771), .S(n2121), .ZN(n1773) );
  MUX2ND0 U2147 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n2140), 
        .ZN(n1778) );
  MUX2ND0 U2148 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n2140), 
        .ZN(n1777) );
  MUX3ND0 U2149 ( .I0(n1781), .I1(n1780), .I2(n1776), .S0(n2121), .S1(n2257), 
        .ZN(n1788) );
  MUX2ND0 U2150 ( .I0(n1783), .I1(n1782), .S(n2121), .ZN(n1787) );
  MUX2ND0 U2151 ( .I0(n1785), .I1(n1784), .S(n2121), .ZN(n1786) );
  MUX2ND0 U2152 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n2142), 
        .ZN(n1791) );
  MUX2ND0 U2153 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n2140), 
        .ZN(n1790) );
  MUX3ND0 U2154 ( .I0(n1794), .I1(n1793), .I2(n1789), .S0(n2123), .S1(n2116), 
        .ZN(n1801) );
  MUX2ND0 U2155 ( .I0(n1796), .I1(n1795), .S(n2121), .ZN(n1800) );
  MUX2ND0 U2156 ( .I0(n1798), .I1(n1797), .S(n2121), .ZN(n1799) );
  MUX2ND0 U2157 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n2140), 
        .ZN(n1804) );
  MUX2ND0 U2158 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n2142), 
        .ZN(n1803) );
  MUX3ND0 U2159 ( .I0(n1807), .I1(n1806), .I2(n1802), .S0(n2122), .S1(n2116), 
        .ZN(n1814) );
  MUX2ND0 U2160 ( .I0(n1809), .I1(n1808), .S(n2121), .ZN(n1813) );
  MUX2ND0 U2161 ( .I0(n1811), .I1(n1810), .S(n2120), .ZN(n1812) );
  MUX2ND0 U2162 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(N44), 
        .ZN(n1817) );
  MUX2ND0 U2163 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n2140), 
        .ZN(n1816) );
  MUX3ND0 U2164 ( .I0(n1820), .I1(n1819), .I2(n1815), .S0(n2121), .S1(n2117), 
        .ZN(n1827) );
  MUX2ND0 U2165 ( .I0(n1822), .I1(n1821), .S(n2120), .ZN(n1826) );
  MUX2ND0 U2166 ( .I0(n1824), .I1(n1823), .S(n2120), .ZN(n1825) );
  MUX2ND0 U2167 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n2140), 
        .ZN(n1830) );
  MUX2ND0 U2168 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n2140), 
        .ZN(n1829) );
  MUX3ND0 U2169 ( .I0(n1833), .I1(n1832), .I2(n1828), .S0(n2121), .S1(n2257), 
        .ZN(n1840) );
  MUX2ND0 U2170 ( .I0(n1835), .I1(n1834), .S(n2121), .ZN(n1839) );
  MUX2ND0 U2171 ( .I0(n1837), .I1(n1836), .S(n2120), .ZN(n1838) );
  MUX2ND0 U2172 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n2140), 
        .ZN(n1843) );
  MUX2ND0 U2173 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n2140), 
        .ZN(n1842) );
  MUX3ND0 U2174 ( .I0(n1846), .I1(n1845), .I2(n1841), .S0(n2122), .S1(n2116), 
        .ZN(n1853) );
  MUX2ND0 U2175 ( .I0(n1848), .I1(n1847), .S(n2121), .ZN(n1852) );
  MUX2ND0 U2176 ( .I0(n1850), .I1(n1849), .S(n2120), .ZN(n1851) );
  MUX2ND0 U2177 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n2140), 
        .ZN(n1856) );
  MUX2ND0 U2178 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n2140), 
        .ZN(n1855) );
  MUX3ND0 U2179 ( .I0(n1859), .I1(n1858), .I2(n1854), .S0(n2122), .S1(n2257), 
        .ZN(n1866) );
  MUX2ND0 U2180 ( .I0(n1861), .I1(n1860), .S(n2121), .ZN(n1865) );
  MUX2ND0 U2181 ( .I0(n1863), .I1(n1862), .S(n2121), .ZN(n1864) );
  MUX2ND0 U2182 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n2140), 
        .ZN(n1869) );
  MUX2ND0 U2183 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n2140), 
        .ZN(n1868) );
  MUX3ND0 U2184 ( .I0(n1872), .I1(n1871), .I2(n1867), .S0(n2121), .S1(n2117), 
        .ZN(n1879) );
  MUX2ND0 U2185 ( .I0(n1874), .I1(n1873), .S(n2120), .ZN(n1878) );
  MUX2ND0 U2186 ( .I0(n1876), .I1(n1875), .S(n2120), .ZN(n1877) );
  MUX2ND0 U2187 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n2140), 
        .ZN(n1882) );
  MUX2ND0 U2188 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n2140), 
        .ZN(n1881) );
  MUX3ND0 U2189 ( .I0(n1885), .I1(n1884), .I2(n1880), .S0(n2120), .S1(n2117), 
        .ZN(n1892) );
  MUX2ND0 U2190 ( .I0(n1887), .I1(n1886), .S(n2120), .ZN(n1891) );
  MUX2ND0 U2191 ( .I0(n1889), .I1(n1888), .S(n2118), .ZN(n1890) );
  MUX2ND0 U2192 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n2140), 
        .ZN(n1895) );
  MUX2ND0 U2193 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n2140), 
        .ZN(n1894) );
  MUX3ND0 U2194 ( .I0(n1898), .I1(n1897), .I2(n1893), .S0(n2122), .S1(n2257), 
        .ZN(n1905) );
  MUX2ND0 U2195 ( .I0(n1900), .I1(n1899), .S(n2119), .ZN(n1904) );
  MUX2ND0 U2196 ( .I0(n1902), .I1(n1901), .S(n2118), .ZN(n1903) );
  MUX2ND0 U2197 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n2139), 
        .ZN(n1908) );
  MUX2ND0 U2198 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n2140), 
        .ZN(n1907) );
  MUX3ND0 U2199 ( .I0(n1911), .I1(n1910), .I2(n1906), .S0(n2122), .S1(n2117), 
        .ZN(n1918) );
  MUX2ND0 U2200 ( .I0(n1913), .I1(n1912), .S(n2119), .ZN(n1917) );
  MUX2ND0 U2201 ( .I0(n1915), .I1(n1914), .S(n2118), .ZN(n1916) );
  MUX2ND0 U2202 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n2140), 
        .ZN(n1921) );
  MUX2ND0 U2203 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n2139), 
        .ZN(n1920) );
  MUX3ND0 U2204 ( .I0(n1924), .I1(n1923), .I2(n1919), .S0(n2122), .S1(n2116), 
        .ZN(n1931) );
  MUX2ND0 U2205 ( .I0(n1926), .I1(n1925), .S(n2118), .ZN(n1930) );
  MUX2ND0 U2206 ( .I0(n1928), .I1(n1927), .S(n2118), .ZN(n1929) );
  MUX2ND0 U2207 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n2139), 
        .ZN(n1934) );
  MUX2ND0 U2208 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n2139), 
        .ZN(n1933) );
  MUX3ND0 U2209 ( .I0(n1937), .I1(n1936), .I2(n1932), .S0(n2119), .S1(n2116), 
        .ZN(n1944) );
  MUX2ND0 U2210 ( .I0(n1939), .I1(n1938), .S(n2119), .ZN(n1943) );
  MUX2ND0 U2211 ( .I0(n1941), .I1(n1940), .S(n2119), .ZN(n1942) );
  MUX2ND0 U2212 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n2139), 
        .ZN(n1947) );
  MUX2ND0 U2213 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n2139), 
        .ZN(n1946) );
  MUX3ND0 U2214 ( .I0(n1950), .I1(n1949), .I2(n1945), .S0(n2122), .S1(N47), 
        .ZN(n1957) );
  MUX2ND0 U2215 ( .I0(n1952), .I1(n1951), .S(n2119), .ZN(n1956) );
  MUX2ND0 U2216 ( .I0(n1954), .I1(n1953), .S(n2119), .ZN(n1955) );
  MUX2ND0 U2217 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n2139), 
        .ZN(n1960) );
  MUX2ND0 U2218 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n2139), 
        .ZN(n1959) );
  MUX3ND0 U2219 ( .I0(n1963), .I1(n1962), .I2(n1958), .S0(n2120), .S1(N47), 
        .ZN(n1970) );
  MUX2ND0 U2220 ( .I0(n1965), .I1(n1964), .S(n2119), .ZN(n1969) );
  MUX2ND0 U2221 ( .I0(n1967), .I1(n1966), .S(n2119), .ZN(n1968) );
  MUX2ND0 U2222 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n2139), 
        .ZN(n1973) );
  MUX2ND0 U2223 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n2139), 
        .ZN(n1972) );
  MUX3ND0 U2224 ( .I0(n1976), .I1(n1975), .I2(n1971), .S0(n2123), .S1(n2116), 
        .ZN(n1983) );
  MUX2ND0 U2225 ( .I0(n1978), .I1(n1977), .S(n2122), .ZN(n1982) );
  MUX2ND0 U2226 ( .I0(n1980), .I1(n1979), .S(n2122), .ZN(n1981) );
  MUX2ND0 U2227 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n2139), 
        .ZN(n1986) );
  MUX2ND0 U2228 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n2139), 
        .ZN(n1985) );
  MUX3ND0 U2229 ( .I0(n1989), .I1(n1988), .I2(n1984), .S0(n2122), .S1(N47), 
        .ZN(n1996) );
  MUX2ND0 U2230 ( .I0(n1991), .I1(n1990), .S(n2118), .ZN(n1995) );
  MUX2ND0 U2231 ( .I0(n1993), .I1(n1992), .S(n2119), .ZN(n1994) );
  MUX2ND0 U2232 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n2139), 
        .ZN(n1999) );
  MUX2ND0 U2233 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n2139), 
        .ZN(n1998) );
  MUX3ND0 U2234 ( .I0(n2002), .I1(n2001), .I2(n1997), .S0(n2122), .S1(N47), 
        .ZN(n2009) );
  MUX2ND0 U2235 ( .I0(n2004), .I1(n2003), .S(n2119), .ZN(n2008) );
  MUX2ND0 U2236 ( .I0(n2006), .I1(n2005), .S(n2119), .ZN(n2007) );
  MUX2ND0 U2237 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n2139), 
        .ZN(n2012) );
  MUX2ND0 U2238 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n2139), 
        .ZN(n2011) );
  MUX3ND0 U2239 ( .I0(n2015), .I1(n2014), .I2(n2010), .S0(n2122), .S1(n2117), 
        .ZN(n2022) );
  MUX2ND0 U2240 ( .I0(n2017), .I1(n2016), .S(n2122), .ZN(n2021) );
  MUX2ND0 U2241 ( .I0(n2019), .I1(n2018), .S(n2122), .ZN(n2020) );
  MUX2ND0 U2242 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n2139), 
        .ZN(n2025) );
  MUX2ND0 U2243 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n2138), 
        .ZN(n2024) );
  MUX3ND0 U2244 ( .I0(n2028), .I1(n2027), .I2(n2023), .S0(n2123), .S1(N47), 
        .ZN(n2035) );
  MUX2ND0 U2245 ( .I0(n2030), .I1(n2029), .S(n2122), .ZN(n2034) );
  MUX2ND0 U2246 ( .I0(n2032), .I1(n2031), .S(n2122), .ZN(n2033) );
  MUX2ND0 U2247 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n2138), 
        .ZN(n2038) );
  MUX2ND0 U2248 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n2138), 
        .ZN(n2037) );
  MUX3ND0 U2249 ( .I0(n2041), .I1(n2040), .I2(n2036), .S0(n2122), .S1(n2116), 
        .ZN(n2048) );
  MUX2ND0 U2250 ( .I0(n2043), .I1(n2042), .S(n2122), .ZN(n2047) );
  MUX2ND0 U2251 ( .I0(n2045), .I1(n2044), .S(n2122), .ZN(n2046) );
  MUX2ND0 U2252 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n2138), 
        .ZN(n2051) );
  MUX2ND0 U2253 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n2138), 
        .ZN(n2050) );
  MUX3ND0 U2254 ( .I0(n2054), .I1(n2053), .I2(n2049), .S0(n2123), .S1(n2117), 
        .ZN(n2061) );
  MUX2ND0 U2255 ( .I0(n2056), .I1(n2055), .S(n2122), .ZN(n2060) );
  MUX2ND0 U2256 ( .I0(n2058), .I1(n2057), .S(n2122), .ZN(n2059) );
  MUX2ND0 U2257 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n2138), 
        .ZN(n2064) );
  MUX2ND0 U2258 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n2138), 
        .ZN(n2063) );
  MUX3ND0 U2259 ( .I0(n2067), .I1(n2066), .I2(n2062), .S0(n2123), .S1(n2116), 
        .ZN(n2074) );
  MUX2ND0 U2260 ( .I0(n2069), .I1(n2068), .S(n2119), .ZN(n2073) );
  MUX2ND0 U2261 ( .I0(n2071), .I1(n2070), .S(n2118), .ZN(n2072) );
  MUX2ND0 U2262 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n2138), 
        .ZN(n2077) );
  MUX2ND0 U2263 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n2138), 
        .ZN(n2076) );
  MUX3ND0 U2264 ( .I0(n2080), .I1(n2079), .I2(n2075), .S0(n2123), .S1(n2116), 
        .ZN(n2087) );
  MUX2ND0 U2265 ( .I0(n2082), .I1(n2081), .S(n2119), .ZN(n2086) );
  MUX2ND0 U2266 ( .I0(n2084), .I1(n2083), .S(n2119), .ZN(n2085) );
  MUX2ND0 U2267 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n2138), 
        .ZN(n2090) );
  MUX2ND0 U2268 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n2138), 
        .ZN(n2089) );
  MUX3ND0 U2269 ( .I0(n2093), .I1(n2092), .I2(n2088), .S0(n2123), .S1(n2116), 
        .ZN(n2100) );
  MUX2ND0 U2270 ( .I0(n2095), .I1(n2094), .S(n2123), .ZN(n2099) );
  MUX2ND0 U2271 ( .I0(n2097), .I1(n2096), .S(n2119), .ZN(n2098) );
  MUX2ND0 U2272 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n2138), 
        .ZN(n2103) );
  MUX2ND0 U2273 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n2140), 
        .ZN(n2102) );
  MUX3ND0 U2274 ( .I0(n2106), .I1(n2105), .I2(n2101), .S0(n2123), .S1(n2117), 
        .ZN(n2113) );
  MUX2ND0 U2275 ( .I0(n2108), .I1(n2107), .S(n2122), .ZN(n2112) );
  MUX2ND0 U2276 ( .I0(n2110), .I1(n2109), .S(N46), .ZN(n2111) );
endmodule


module PLLTop ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(Reset) );
  VFO VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(Reset) );
  MultiCounter MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(Reset)
         );
endmodule


module ClockComparator ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   N5, N6, N7, N8, N9, N19, N20, n2, n3, n4, n5, n6, n7, n1, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47;
  wire   [1:0] ClockInN;
  wire   [1:0] CounterClockN;

  MOAI22D1 U5 ( .A1(n4), .A2(n5), .B1(n6), .B2(ClockInN[1]), .ZN(N20) );
  MOAI22D1 U8 ( .A1(CounterClockN[1]), .A2(n7), .B1(n6), .B2(N9), .ZN(N19) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n3), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n2), .Q(
        CounterClockN[1]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n3), .Q(
        AdjustFreq[1]) );
  DFCNQD1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n2), .Q(
        CounterClockN[0]) );
  DFCNQD1 \ClockInN_reg[1]  ( .D(n8), .CP(ClockIn), .CDN(n2), .Q(ClockInN[1])
         );
  DFCNQD1 \ClockInN_reg[0]  ( .D(n21), .CP(ClockIn), .CDN(n2), .Q(ClockInN[0])
         );
  DFSND1 ZeroCounters_reg ( .D(n33), .CP(ClockIn), .SDN(n3), .QN(n2) );
  INVD8 U3 ( .I(n1), .ZN(n8) );
  INVD0 U4 ( .I(n15), .ZN(n1) );
  INVD0 U6 ( .I(n9), .ZN(n10) );
  CKNXD16 U7 ( .I(N6), .ZN(n9) );
  CKXOR2D0 U9 ( .A1(n11), .A2(n29), .Z(N6) );
  CKBD0 U10 ( .CLK(ClockInN[1]), .C(n11) );
  INVD0 U11 ( .I(n12), .ZN(n13) );
  CKNXD16 U12 ( .I(n10), .ZN(n12) );
  CKNXD16 U13 ( .I(n14), .ZN(n15) );
  INVD0 U14 ( .I(n17), .ZN(n14) );
  INVD0 U15 ( .I(n18), .ZN(n19) );
  CKNXD16 U16 ( .I(n16), .ZN(n17) );
  INVD0 U17 ( .I(n19), .ZN(n16) );
  CKNXD16 U18 ( .I(n13), .ZN(n18) );
  CKNXD16 U19 ( .I(n23), .ZN(n20) );
  INVD1 U20 ( .I(n20), .ZN(n21) );
  INVD0 U21 ( .I(n22), .ZN(n23) );
  CKNXD16 U22 ( .I(n25), .ZN(n22) );
  INVD0 U23 ( .I(N5), .ZN(n30) );
  INVD0 U24 ( .I(n24), .ZN(n25) );
  CKNXD16 U25 ( .I(n28), .ZN(n24) );
  CKBXD0 U26 ( .I(n31), .Z(n28) );
  BUFFD0 U27 ( .I(n27), .Z(n29) );
  INVD0 U28 ( .I(ClockInN[0]), .ZN(n26) );
  CKNXD16 U29 ( .I(n26), .ZN(n27) );
  CKNXD16 U30 ( .I(n30), .ZN(n31) );
  CKNXD16 U31 ( .I(n29), .ZN(N5) );
  INVD16 U32 ( .I(n42), .ZN(n43) );
  INVD0 U33 ( .I(n45), .ZN(n42) );
  CKNXD0 U34 ( .I(n46), .ZN(n47) );
  CKNXD16 U35 ( .I(n32), .ZN(n46) );
  BUFFD0 U36 ( .I(N9), .Z(n32) );
  CKBD0 U37 ( .CLK(n35), .C(n33) );
  CKNXD16 U38 ( .I(n34), .ZN(n35) );
  CKNXD0 U39 ( .I(n37), .ZN(n34) );
  INVD0 U40 ( .I(n47), .ZN(n44) );
  CKNXD16 U41 ( .I(n36), .ZN(n37) );
  CKNXD0 U42 ( .I(n39), .ZN(n36) );
  CKNXD16 U43 ( .I(n38), .ZN(n39) );
  CKNXD0 U44 ( .I(n41), .ZN(n38) );
  CKNXD16 U45 ( .I(n40), .ZN(n41) );
  CKNXD0 U46 ( .I(n43), .ZN(n40) );
  CKNXD16 U47 ( .I(n44), .ZN(n45) );
  AN2D8 U48 ( .A1(n11), .A2(ClockInN[0]), .Z(N9) );
  INVD1 U49 ( .I(Reset), .ZN(n3) );
  XOR2D1 U50 ( .A1(CounterClockN[1]), .A2(CounterClockN[0]), .Z(n5) );
  AOI21D1 U51 ( .A1(ClockInN[0]), .A2(n6), .B(N9), .ZN(n4) );
  INR3D0 U52 ( .A1(CounterClockN[0]), .B1(ClockInN[1]), .B2(ClockInN[0]), .ZN(
        n7) );
  ND2D1 U53 ( .A1(CounterClockN[1]), .A2(CounterClockN[0]), .ZN(n6) );
  XOR2D1 U54 ( .A1(CounterClockN[1]), .A2(CounterClockN[0]), .Z(N8) );
  INVD1 U55 ( .I(CounterClockN[0]), .ZN(N7) );
endmodule


module VFO ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N8, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20,
         N21, N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N41,
         N54, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n1,
         n2, n4, n5, n6, n7, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay83ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay83ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay83ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay83ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay83ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_DW01_dec_0 \Sampler/sub_183  ( .A({n27, n23, n29, n38, n19, n60}), .SUM(
        {N40, N39, N38, N37, N36, N35}) );
  VFO_DW01_inc_0 \Sampler/add_180  ( .A({n27, n23, n29, n38, n19, n60}), .SUM(
        {N32, N31, N30, N29, N28, N27}) );
  VFO_DW01_inc_1 \ClockOutGen/add_161  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  VFO_DW01_cmp2_2 \ClockOutGen/lt_160  ( .A(FastDivvy), .B(DivideFactor), 
        .LEQ(n3), .TC(n3), .LT_LE(N8) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[5]) );
  ND2D1 U30 ( .A1(WireD[5]), .A2(n20), .ZN(WireD[0]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[3]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n20), .Q(
        FastDivvy[1]) );
  DFCNQD1 ClockOutReg_reg ( .D(n17), .CP(FastClock), .CDN(n20), .Q(ClockOut)
         );
  DFSNQD1 \DivideFactor_reg[0]  ( .D(n1), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[0]) );
  DFSNQD1 \DivideFactor_reg[1]  ( .D(n7), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[1]) );
  DFSNQD1 \DivideFactor_reg[4]  ( .D(n21), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[4]) );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(n25), .E(n39), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[3]  ( .D(n104), .E(n39), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[3]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(n30), .E(n39), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[2]) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n4), .Z(n2) );
  BUFFD0 U5 ( .I(n5), .Z(n4) );
  BUFFD0 U6 ( .I(n6), .Z(n5) );
  BUFFD0 U7 ( .I(n48), .Z(n6) );
  AN2D0 U8 ( .A1(n125), .A2(n11), .Z(n9) );
  BUFFD0 U9 ( .I(n61), .Z(n7) );
  BUFFD0 U10 ( .I(n37), .Z(n19) );
  BUFFD0 U11 ( .I(n75), .Z(n21) );
  BUFFD0 U12 ( .I(n40), .Z(n22) );
  BUFFD0 U13 ( .I(n88), .Z(n23) );
  BUFFD0 U14 ( .I(n22), .Z(n24) );
  INVD4 U15 ( .I(n44), .ZN(n89) );
  BUFFD0 U16 ( .I(n26), .Z(n25) );
  BUFFD0 U17 ( .I(n91), .Z(n26) );
  BUFFD0 U18 ( .I(n28), .Z(n27) );
  BUFFD0 U19 ( .I(DivideFactor[5]), .Z(n28) );
  CKND12 U20 ( .CLK(n113), .CN(n114) );
  INVD16 U21 ( .I(n43), .ZN(n102) );
  BUFFD0 U22 ( .I(DivideFactor[3]), .Z(n29) );
  BUFFD10 U23 ( .I(n121), .Z(n124) );
  BUFFD0 U24 ( .I(n31), .Z(n30) );
  BUFFD0 U25 ( .I(n32), .Z(n31) );
  BUFFD0 U26 ( .I(n33), .Z(n32) );
  BUFFD0 U27 ( .I(n34), .Z(n33) );
  BUFFD0 U28 ( .I(n35), .Z(n34) );
  BUFFD0 U29 ( .I(n36), .Z(n35) );
  BUFFD0 U31 ( .I(n116), .Z(n36) );
  BUFFD0 U32 ( .I(DivideFactor[1]), .Z(n37) );
  BUFFD0 U33 ( .I(DivideFactor[2]), .Z(n38) );
  BUFFD0 U34 ( .I(n127), .Z(n39) );
  AO222D1 U35 ( .A1(N39), .A2(n8), .B1(N31), .B2(n9), .C1(n23), .C2(n126), .Z(
        n40) );
  AN3D1 U36 ( .A1(n42), .A2(n38), .A3(n29), .Z(n41) );
  AN3D1 U37 ( .A1(n27), .A2(n23), .A3(n19), .Z(n42) );
  AOI22D0 U38 ( .A1(N38), .A2(n12), .B1(N30), .B2(n11), .ZN(n43) );
  AOI22D0 U39 ( .A1(N40), .A2(n12), .B1(N32), .B2(n11), .ZN(n44) );
  AOI222D0 U40 ( .A1(N36), .A2(n8), .B1(N28), .B2(n9), .C1(n19), .C2(n126), 
        .ZN(n45) );
  INVD1 U41 ( .I(n45), .ZN(n18) );
  AOI222D0 U42 ( .A1(N35), .A2(n8), .B1(N27), .B2(n9), .C1(n60), .C2(n126), 
        .ZN(n46) );
  AOI22D0 U43 ( .A1(N37), .A2(n12), .B1(N29), .B2(n11), .ZN(n47) );
  CKND12 U44 ( .CLK(n55), .CN(n56) );
  BUFFD0 U45 ( .I(n50), .Z(n48) );
  CKNXD16 U46 ( .I(n49), .ZN(n50) );
  CKNXD0 U47 ( .I(n52), .ZN(n49) );
  CKNXD16 U48 ( .I(n51), .ZN(n52) );
  CKNXD0 U49 ( .I(n54), .ZN(n51) );
  CKNXD16 U50 ( .I(n53), .ZN(n54) );
  CKNXD0 U51 ( .I(n56), .ZN(n53) );
  CKNXD0 U52 ( .I(n58), .ZN(n55) );
  CKNXD16 U53 ( .I(n57), .ZN(n58) );
  INVD0 U54 ( .I(n59), .ZN(n57) );
  INVD0 U55 ( .I(n46), .ZN(n59) );
  CKBXD0 U56 ( .I(DivideFactor[0]), .Z(n60) );
  CKBD12 U57 ( .CLK(n74), .C(n72) );
  BUFFD0 U58 ( .I(n63), .Z(n61) );
  CKNXD16 U59 ( .I(n62), .ZN(n63) );
  CKNXD0 U60 ( .I(n65), .ZN(n62) );
  CKNXD16 U61 ( .I(n64), .ZN(n65) );
  CKNXD0 U62 ( .I(n67), .ZN(n64) );
  CKNXD16 U63 ( .I(n66), .ZN(n67) );
  CKNXD0 U64 ( .I(n69), .ZN(n66) );
  CKNXD16 U65 ( .I(n68), .ZN(n69) );
  INVD0 U66 ( .I(n71), .ZN(n68) );
  CKNXD16 U67 ( .I(n70), .ZN(n71) );
  INVD0 U68 ( .I(n72), .ZN(n70) );
  INVD0 U69 ( .I(n73), .ZN(n74) );
  CKNXD16 U70 ( .I(n18), .ZN(n73) );
  BUFFD0 U71 ( .I(n77), .Z(n75) );
  CKNXD16 U72 ( .I(n76), .ZN(n77) );
  CKNXD0 U73 ( .I(n79), .ZN(n76) );
  CKNXD16 U74 ( .I(n78), .ZN(n79) );
  CKNXD0 U75 ( .I(n81), .ZN(n78) );
  CKNXD16 U76 ( .I(n80), .ZN(n81) );
  CKNXD0 U77 ( .I(n83), .ZN(n80) );
  CKNXD16 U78 ( .I(n82), .ZN(n83) );
  CKNXD0 U79 ( .I(n85), .ZN(n82) );
  CKNXD16 U80 ( .I(n84), .ZN(n85) );
  INVD0 U81 ( .I(n87), .ZN(n84) );
  CKNXD0 U82 ( .I(n24), .ZN(n86) );
  CKNXD16 U83 ( .I(n86), .ZN(n87) );
  BUFFD0 U84 ( .I(DivideFactor[4]), .Z(n88) );
  CKNXD16 U85 ( .I(n90), .ZN(n91) );
  CKNXD0 U86 ( .I(n93), .ZN(n90) );
  CKNXD16 U87 ( .I(n92), .ZN(n93) );
  CKNXD0 U88 ( .I(n95), .ZN(n92) );
  CKNXD16 U89 ( .I(n94), .ZN(n95) );
  CKNXD0 U90 ( .I(n97), .ZN(n94) );
  CKNXD16 U91 ( .I(n96), .ZN(n97) );
  CKNXD0 U92 ( .I(n99), .ZN(n96) );
  CKNXD16 U93 ( .I(n98), .ZN(n99) );
  CKNXD0 U94 ( .I(n101), .ZN(n98) );
  CKNXD16 U95 ( .I(n100), .ZN(n101) );
  INVD0 U96 ( .I(n89), .ZN(n100) );
  CKNXD16 U97 ( .I(n103), .ZN(n104) );
  CKNXD0 U98 ( .I(n106), .ZN(n103) );
  CKNXD16 U99 ( .I(n105), .ZN(n106) );
  CKNXD0 U100 ( .I(n108), .ZN(n105) );
  CKNXD16 U101 ( .I(n107), .ZN(n108) );
  CKNXD0 U102 ( .I(n110), .ZN(n107) );
  CKNXD16 U103 ( .I(n109), .ZN(n110) );
  CKNXD0 U104 ( .I(n112), .ZN(n109) );
  CKNXD16 U105 ( .I(n111), .ZN(n112) );
  CKNXD0 U106 ( .I(n114), .ZN(n111) );
  INVD0 U107 ( .I(n102), .ZN(n113) );
  CKNXD16 U108 ( .I(n115), .ZN(n116) );
  INVD0 U109 ( .I(n119), .ZN(n115) );
  INVD0 U110 ( .I(n47), .ZN(n117) );
  CKNXD16 U111 ( .I(n118), .ZN(n119) );
  INVD0 U112 ( .I(n123), .ZN(n118) );
  INVD0 U113 ( .I(n120), .ZN(n121) );
  CKNXD16 U114 ( .I(n117), .ZN(n120) );
  CKNXD16 U115 ( .I(n122), .ZN(n123) );
  INVD0 U116 ( .I(n124), .ZN(n122) );
  INVD0 U117 ( .I(n41), .ZN(n125) );
  BUFFD0 U118 ( .I(n128), .Z(n126) );
  BUFFD0 U119 ( .I(n129), .Z(n127) );
  BUFFD0 U120 ( .I(n130), .Z(n128) );
  BUFFD0 U121 ( .I(n131), .Z(n129) );
  BUFFD0 U122 ( .I(n132), .Z(n130) );
  BUFFD0 U123 ( .I(n133), .Z(n131) );
  BUFFD0 U124 ( .I(n134), .Z(n132) );
  BUFFD0 U125 ( .I(n135), .Z(n133) );
  BUFFD0 U126 ( .I(n136), .Z(n134) );
  BUFFD0 U127 ( .I(n137), .Z(n135) );
  BUFFD0 U128 ( .I(n138), .Z(n136) );
  BUFFD0 U129 ( .I(n139), .Z(n137) );
  BUFFD0 U130 ( .I(n140), .Z(n138) );
  BUFFD0 U131 ( .I(n141), .Z(n139) );
  BUFFD0 U132 ( .I(n142), .Z(n140) );
  BUFFD0 U133 ( .I(n143), .Z(n141) );
  BUFFD0 U134 ( .I(n10), .Z(n142) );
  BUFFD0 U135 ( .I(n144), .Z(n143) );
  BUFFD0 U136 ( .I(n145), .Z(n144) );
  BUFFD0 U137 ( .I(n146), .Z(n145) );
  BUFFD0 U138 ( .I(n147), .Z(n146) );
  BUFFD0 U139 ( .I(n148), .Z(n147) );
  BUFFD0 U140 ( .I(n149), .Z(n148) );
  BUFFD0 U141 ( .I(n150), .Z(n149) );
  BUFFD0 U142 ( .I(n151), .Z(n150) );
  BUFFD0 U143 ( .I(n152), .Z(n151) );
  BUFFD0 U144 ( .I(n153), .Z(n152) );
  BUFFD0 U145 ( .I(N54), .Z(n153) );
  OAI21D0 U146 ( .A1(n13), .A2(n14), .B(n15), .ZN(n10) );
  INVD1 U147 ( .I(n126), .ZN(N54) );
  AN2D1 U148 ( .A1(N41), .A2(n12), .Z(n8) );
  NR2D1 U149 ( .A1(n16), .A2(n14), .ZN(n12) );
  INVD1 U150 ( .I(Reset), .ZN(n20) );
  AN2D1 U151 ( .A1(N13), .A2(N8), .Z(N20) );
  AN2D1 U152 ( .A1(N12), .A2(N8), .Z(N19) );
  AN2D1 U153 ( .A1(N11), .A2(N8), .Z(N18) );
  AN2D1 U154 ( .A1(N10), .A2(N8), .Z(N17) );
  IOA21D1 U155 ( .A1(n16), .A2(n125), .B(n14), .ZN(n15) );
  AN2D1 U156 ( .A1(N41), .A2(AdjustFreq[1]), .Z(n13) );
  INVD1 U157 ( .I(WireD[0]), .ZN(FastClock) );
  INVD1 U158 ( .I(AdjustFreq[0]), .ZN(n14) );
  NR2D1 U159 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n11) );
  XNR2D1 U160 ( .A1(ClockOut), .A2(N8), .ZN(n17) );
  INVD1 U161 ( .I(AdjustFreq[1]), .ZN(n16) );
  AN2D1 U162 ( .A1(N14), .A2(N8), .Z(N21) );
  AN2D1 U163 ( .A1(N9), .A2(N8), .Z(N16) );
  TIEL U164 ( .ZN(n3) );
  AN3D0 U165 ( .A1(n29), .A2(n38), .A3(n19), .Z(n154) );
  OR3D0 U166 ( .A1(n27), .A2(n23), .A3(n154), .Z(N41) );
endmodule


module MultiCounter ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1, n2, n3, n4;
  wire   [3:0] Ctr;

  MultiCounter_DW01_inc_0 add_16 ( .A({CarryOut, Ctr[3:1], n2}), .SUM({N4, N5, 
        N3, N2, N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  CKBXD0 U3 ( .I(n4), .Z(n2) );
  INVD16 U4 ( .I(n3), .ZN(n4) );
  INVD0 U5 ( .I(Ctr[0]), .ZN(n3) );
  INVD1 U6 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n10, n11, n12, \carry[4] , \carry[3] , \carry[2] , n2, n3, n5, n7, n9
;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n10) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(n12) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n11) );
  CKBD0 U1 ( .CLK(n9), .C(SUM[4]) );
  INVD8 U2 ( .I(n2), .ZN(n9) );
  XNR2D0 U3 ( .A1(\carry[4] ), .A2(A[4]), .ZN(n2) );
  CKNXD16 U4 ( .I(n3), .ZN(SUM[1]) );
  INVD0 U5 ( .I(n12), .ZN(n3) );
  CKNXD16 U6 ( .I(n5), .ZN(SUM[2]) );
  INVD0 U7 ( .I(n11), .ZN(n5) );
  CKNXD16 U8 ( .I(n7), .ZN(SUM[3]) );
  INVD0 U9 ( .I(n10), .ZN(n7) );
  CKND0 U10 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKNXD16 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CKXOR2D0 U2 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
endmodule


module VFO_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_cmp2_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [5:0] A;
  input [5:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  OAI21D0 U1 ( .A1(A[5]), .A2(n1), .B(n2), .ZN(LT_LE) );
  IOA21D0 U2 ( .A1(n1), .A2(A[5]), .B(n3), .ZN(n2) );
  IOA21D0 U3 ( .A1(n4), .A2(B[4]), .B(n5), .ZN(n3) );
  OAI221D0 U4 ( .A1(B[3]), .A2(n6), .B1(B[4]), .B2(n4), .C(n7), .ZN(n5) );
  AO221D0 U5 ( .A1(n8), .A2(B[2]), .B1(n6), .B2(B[3]), .C(n9), .Z(n7) );
  OA222D0 U6 ( .A1(n10), .A2(n11), .B1(B[1]), .B2(n12), .C1(B[2]), .C2(n8), 
        .Z(n9) );
  INR2D0 U7 ( .A1(n10), .B1(A[1]), .ZN(n12) );
  CKND0 U8 ( .CLK(A[1]), .CN(n11) );
  INR2D0 U9 ( .A1(B[0]), .B1(A[0]), .ZN(n10) );
  CKND0 U10 ( .CLK(A[2]), .CN(n8) );
  CKND0 U11 ( .CLK(A[3]), .CN(n6) );
  CKND0 U12 ( .CLK(A[4]), .CN(n4) );
  CKND0 U13 ( .CLK(B[5]), .CN(n1) );
endmodule


module DesDecoder_DWid32_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n3, \carry[4] , \carry[3] , \carry[2] , n2;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  XOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  INVD3 U2 ( .I(A[0]), .ZN(n3) );
  BUFFD0 U3 ( .I(n2), .Z(SUM[0]) );
  CKBD0 U4 ( .CLK(n3), .C(n2) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n10, n11, \carry[4] , \carry[3] , \carry[2] , n1, n3, n4, n5, n7, n8;

  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(n11) );
  HA1D4 U1_1_1 ( .A(A[1]), .B(n7), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(n10) );
  INVD1 U1 ( .I(n5), .ZN(SUM[3]) );
  CKNXD0 U2 ( .I(n1), .ZN(SUM[2]) );
  CKNXD16 U3 ( .I(n4), .ZN(n1) );
  INVD0 U4 ( .I(n3), .ZN(n4) );
  CKNXD16 U5 ( .I(n11), .ZN(n3) );
  INVD0 U6 ( .I(n10), .ZN(n5) );
  CKNXD16 U7 ( .I(n7), .ZN(SUM[0]) );
  INVD0 U8 ( .I(n8), .ZN(n7) );
  CKNXD16 U9 ( .I(A[0]), .ZN(n8) );
  CKXOR2D0 U10 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
endmodule

