library verilog;
use verilog.vl_types.all;
entity block_nonblock_tb is
end block_nonblock_tb;
