
`ifndef RKV_I2C_USER_TESTS_SVH
`define RKV_I2C_USER_TESTS_SVH

`endif // RKV_I2C_USER_TESTS_SVH

