library verilog;
use verilog.vl_types.all;
entity uvm_pkg_sv_unit is
end uvm_pkg_sv_unit;
