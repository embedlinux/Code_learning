
module CondGenerate ( Result, ArgA, ArgB, Sel, Enable );
  output [31:0] Result;
  input [31:0] ArgA;
  input [31:0] ArgB;
  input Sel, Enable;
  wire   n11, n12, n13, n1, n3, n5, n7, n8, n9, n10;

  Mux32Bit Mux1 ( .Out({Result[31:25], n11, n12, Result[22:10], n13, 
        Result[8:0]}), .A(ArgA), .B(ArgB), .Sel(n10), .unused(Enable) );
  CKBD0 U1 ( .CLK(n8), .C(n1) );
  CKNXD16 U2 ( .I(n1), .ZN(Result[23]) );
  CKBD0 U3 ( .CLK(n7), .C(n3) );
  CKNXD16 U4 ( .I(n3), .ZN(Result[9]) );
  CKBD0 U5 ( .CLK(n9), .C(n5) );
  CKNXD16 U6 ( .I(n5), .ZN(Result[24]) );
  BUFFD1 U7 ( .I(Sel), .Z(n10) );
  CKND0 U8 ( .CLK(n13), .CN(n7) );
  CKND0 U9 ( .CLK(n12), .CN(n8) );
  CKND0 U10 ( .CLK(n11), .CN(n9) );
endmodule


module Mux32Bit ( Out, A, B, Sel, unused );
  output [31:0] Out;
  input [31:0] A;
  input [31:0] B;
  input Sel, unused;
  wire   n194, n1, n2, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, n22,
         n24, n26, n28, n30, n32, n33, n34, n35, n36, n37, n39, n41, n42, n44,
         n46, n47, n49, n51, n53, n55, n56, n58, n60, n62, n64, n66, n68, n70,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193;

  OAI22D0 U1 ( .A1(n179), .A2(n108), .B1(n180), .B2(n169), .ZN(n1) );
  INVD1 U2 ( .I(n1), .ZN(n178) );
  OAI22D0 U3 ( .A1(n176), .A2(n159), .B1(n177), .B2(n147), .ZN(n2) );
  INVD1 U4 ( .I(n2), .ZN(n175) );
  MAOI22D0 U5 ( .A1(B[22]), .A2(n121), .B1(n188), .B2(n192), .ZN(n3) );
  OAI22D0 U6 ( .A1(n190), .A2(n115), .B1(n191), .B2(n121), .ZN(n4) );
  INVD1 U7 ( .I(n4), .ZN(n189) );
  OAI22D0 U8 ( .A1(n183), .A2(n123), .B1(n184), .B2(n147), .ZN(n5) );
  INVD1 U9 ( .I(n5), .ZN(n182) );
  AOI22D0 U10 ( .A1(B[1]), .A2(n169), .B1(A[1]), .B2(n193), .ZN(n112) );
  AOI22D0 U11 ( .A1(B[6]), .A2(n135), .B1(A[6]), .B2(Sel), .ZN(n98) );
  AOI22D0 U12 ( .A1(B[7]), .A2(n169), .B1(A[7]), .B2(n149), .ZN(n105) );
  AOI22D0 U13 ( .A1(A[20]), .A2(n193), .B1(B[20]), .B2(n121), .ZN(n128) );
  AOI22D0 U14 ( .A1(B[25]), .A2(n121), .B1(A[25]), .B2(Sel), .ZN(n119) );
  AOI22D0 U15 ( .A1(B[26]), .A2(n192), .B1(A[26]), .B2(Sel), .ZN(n127) );
  CKBD0 U16 ( .CLK(n178), .C(n6) );
  CKNXD16 U17 ( .I(n6), .ZN(Out[8]) );
  CKBD0 U18 ( .CLK(n189), .C(n8) );
  CKNXD16 U19 ( .I(n8), .ZN(Out[30]) );
  CKBD0 U20 ( .CLK(n41), .C(n10) );
  CKNXD16 U21 ( .I(n10), .ZN(Out[21]) );
  CKBD0 U22 ( .CLK(n46), .C(n12) );
  CKNXD16 U23 ( .I(n12), .ZN(Out[28]) );
  CKBD0 U24 ( .CLK(n32), .C(n14) );
  CKNXD16 U25 ( .I(n14), .ZN(Out[6]) );
  CKBD0 U26 ( .CLK(n55), .C(n16) );
  CKNXD16 U27 ( .I(n16), .ZN(Out[20]) );
  CKBD0 U28 ( .CLK(n182), .C(n18) );
  CKNXD16 U29 ( .I(n18), .ZN(Out[31]) );
  CKBD0 U30 ( .CLK(n175), .C(n20) );
  CKNXD16 U31 ( .I(n20), .ZN(Out[19]) );
  CKBD0 U32 ( .CLK(n35), .C(n22) );
  CKNXD16 U33 ( .I(n22), .ZN(Out[25]) );
  CKBD0 U34 ( .CLK(n36), .C(n24) );
  CKNXD16 U35 ( .I(n24), .ZN(Out[26]) );
  CKBD0 U36 ( .CLK(n34), .C(n26) );
  CKNXD16 U37 ( .I(n26), .ZN(Out[1]) );
  CKBD0 U38 ( .CLK(n33), .C(n28) );
  CKNXD16 U39 ( .I(n28), .ZN(Out[7]) );
  CKBD0 U40 ( .CLK(n87), .C(n30) );
  CKNXD16 U41 ( .I(n30), .ZN(Out[5]) );
  CKBD0 U42 ( .CLK(n98), .C(n32) );
  CKBD0 U43 ( .CLK(n105), .C(n33) );
  CKBXD0 U44 ( .I(n112), .Z(n34) );
  CKBXD0 U45 ( .I(n119), .Z(n35) );
  CKBXD0 U46 ( .I(n127), .Z(n36) );
  CKBD0 U47 ( .CLK(n129), .C(n37) );
  CKNXD16 U48 ( .I(n37), .ZN(Out[27]) );
  CKBD0 U49 ( .CLK(n141), .C(n39) );
  CKNXD16 U50 ( .I(n39), .ZN(Out[29]) );
  CKBD0 U51 ( .CLK(n153), .C(n41) );
  CKBD0 U52 ( .CLK(n163), .C(n42) );
  CKNXD16 U53 ( .I(n42), .ZN(Out[16]) );
  CKBD0 U54 ( .CLK(n3), .C(n44) );
  CKNXD16 U55 ( .I(n44), .ZN(Out[22]) );
  CKBD0 U56 ( .CLK(n186), .C(n46) );
  CKBD0 U57 ( .CLK(n168), .C(n47) );
  CKNXD16 U58 ( .I(n47), .ZN(Out[15]) );
  CKBD0 U59 ( .CLK(n157), .C(n49) );
  CKNXD16 U60 ( .I(n49), .ZN(Out[0]) );
  CKBD0 U61 ( .CLK(n146), .C(n51) );
  CKNXD16 U62 ( .I(n51), .ZN(Out[17]) );
  CKBD0 U63 ( .CLK(n134), .C(n53) );
  CKNXD16 U64 ( .I(n53), .ZN(Out[18]) );
  CKBXD0 U65 ( .I(n128), .Z(n55) );
  CKBD0 U66 ( .CLK(n120), .C(n56) );
  CKNXD16 U67 ( .I(n56), .ZN(Out[10]) );
  CKBD0 U68 ( .CLK(n113), .C(n58) );
  CKNXD16 U69 ( .I(n58), .ZN(Out[11]) );
  CKBD0 U70 ( .CLK(n106), .C(n60) );
  CKNXD16 U71 ( .I(n60), .ZN(Out[12]) );
  CKBD0 U72 ( .CLK(n99), .C(n62) );
  CKNXD16 U73 ( .I(n62), .ZN(Out[13]) );
  CKBD0 U74 ( .CLK(n92), .C(n64) );
  CKNXD16 U75 ( .I(n64), .ZN(Out[14]) );
  CKBD0 U76 ( .CLK(n72), .C(n66) );
  CKNXD16 U77 ( .I(n66), .ZN(Out[3]) );
  CKBD0 U78 ( .CLK(n77), .C(n68) );
  CKNXD16 U79 ( .I(n68), .ZN(Out[4]) );
  CKBD0 U80 ( .CLK(n82), .C(n70) );
  CKNXD16 U81 ( .I(n70), .ZN(Out[2]) );
  CKND0 U82 ( .CLK(A[3]), .CN(n73) );
  INVD1 U83 ( .I(B[3]), .ZN(n74) );
  NR2D0 U84 ( .A1(n169), .A2(n73), .ZN(n75) );
  NR2D0 U85 ( .A1(n101), .A2(n74), .ZN(n76) );
  NR2XD0 U86 ( .A1(n75), .A2(n76), .ZN(n72) );
  CKND0 U87 ( .CLK(A[4]), .CN(n78) );
  CKND0 U88 ( .CLK(B[4]), .CN(n79) );
  NR2D0 U89 ( .A1(n147), .A2(n78), .ZN(n80) );
  NR2D0 U90 ( .A1(n94), .A2(n79), .ZN(n81) );
  NR2XD0 U91 ( .A1(n80), .A2(n81), .ZN(n77) );
  CKND0 U92 ( .CLK(A[2]), .CN(n83) );
  CKND0 U93 ( .CLK(B[2]), .CN(n84) );
  NR2D1 U94 ( .A1(n147), .A2(n83), .ZN(n85) );
  NR2D0 U95 ( .A1(n101), .A2(n84), .ZN(n86) );
  NR2XD0 U96 ( .A1(n85), .A2(n86), .ZN(n82) );
  CKND0 U97 ( .CLK(A[5]), .CN(n88) );
  CKND0 U98 ( .CLK(B[5]), .CN(n89) );
  NR2D0 U99 ( .A1(n147), .A2(n88), .ZN(n90) );
  NR2D0 U100 ( .A1(n94), .A2(n89), .ZN(n91) );
  NR2XD0 U101 ( .A1(n90), .A2(n91), .ZN(n87) );
  CKND0 U102 ( .CLK(A[14]), .CN(n93) );
  CKND0 U103 ( .CLK(n192), .CN(n94) );
  CKND0 U104 ( .CLK(B[14]), .CN(n95) );
  NR2D0 U105 ( .A1(n147), .A2(n93), .ZN(n96) );
  NR2D0 U106 ( .A1(n94), .A2(n95), .ZN(n97) );
  NR2XD0 U107 ( .A1(n96), .A2(n97), .ZN(n92) );
  CKND0 U108 ( .CLK(A[13]), .CN(n100) );
  CKND0 U109 ( .CLK(n192), .CN(n101) );
  CKND0 U110 ( .CLK(B[13]), .CN(n102) );
  NR2D0 U111 ( .A1(n121), .A2(n100), .ZN(n103) );
  NR2D0 U112 ( .A1(n101), .A2(n102), .ZN(n104) );
  NR2XD0 U113 ( .A1(n103), .A2(n104), .ZN(n99) );
  CKND0 U114 ( .CLK(A[12]), .CN(n107) );
  CKND0 U115 ( .CLK(n192), .CN(n108) );
  CKND0 U116 ( .CLK(B[12]), .CN(n109) );
  NR2D0 U117 ( .A1(n192), .A2(n107), .ZN(n110) );
  NR2D0 U118 ( .A1(n108), .A2(n109), .ZN(n111) );
  NR2XD0 U119 ( .A1(n110), .A2(n111), .ZN(n106) );
  CKND0 U120 ( .CLK(A[11]), .CN(n114) );
  CKND0 U121 ( .CLK(n192), .CN(n115) );
  CKND0 U122 ( .CLK(B[11]), .CN(n116) );
  NR2D0 U123 ( .A1(n147), .A2(n114), .ZN(n117) );
  NR2D0 U124 ( .A1(n115), .A2(n116), .ZN(n118) );
  NR2XD0 U125 ( .A1(n117), .A2(n118), .ZN(n113) );
  INVD0 U126 ( .I(Sel), .ZN(n121) );
  CKND0 U127 ( .CLK(A[10]), .CN(n122) );
  CKND0 U128 ( .CLK(n192), .CN(n123) );
  CKND0 U129 ( .CLK(B[10]), .CN(n124) );
  NR2D0 U130 ( .A1(n121), .A2(n122), .ZN(n125) );
  NR2D0 U131 ( .A1(n123), .A2(n124), .ZN(n126) );
  NR2XD0 U132 ( .A1(n125), .A2(n126), .ZN(n120) );
  INVD1 U133 ( .I(n193), .ZN(n192) );
  INVD0 U134 ( .I(A[27]), .ZN(n130) );
  CKND0 U135 ( .CLK(B[27]), .CN(n131) );
  NR2D1 U136 ( .A1(n121), .A2(n130), .ZN(n132) );
  NR2D0 U137 ( .A1(n101), .A2(n131), .ZN(n133) );
  NR2XD0 U138 ( .A1(n132), .A2(n133), .ZN(n129) );
  INVD0 U139 ( .I(n193), .ZN(n135) );
  INVD0 U140 ( .I(A[18]), .ZN(n136) );
  INVD0 U141 ( .I(n192), .ZN(n137) );
  CKND0 U142 ( .CLK(B[18]), .CN(n138) );
  NR2D1 U143 ( .A1(n135), .A2(n136), .ZN(n139) );
  NR2D0 U144 ( .A1(n137), .A2(n138), .ZN(n140) );
  NR2XD0 U145 ( .A1(n139), .A2(n140), .ZN(n134) );
  INVD0 U146 ( .I(A[29]), .ZN(n142) );
  CKND0 U147 ( .CLK(B[29]), .CN(n143) );
  NR2D1 U148 ( .A1(n147), .A2(n142), .ZN(n144) );
  NR2D0 U149 ( .A1(n94), .A2(n143), .ZN(n145) );
  NR2XD0 U150 ( .A1(n144), .A2(n145), .ZN(n141) );
  INVD0 U151 ( .I(n193), .ZN(n147) );
  CKND0 U152 ( .CLK(A[17]), .CN(n148) );
  INVD0 U153 ( .I(n192), .ZN(n149) );
  CKND0 U154 ( .CLK(B[17]), .CN(n150) );
  NR2D0 U155 ( .A1(n147), .A2(n148), .ZN(n151) );
  NR2D0 U156 ( .A1(n149), .A2(n150), .ZN(n152) );
  NR2XD0 U157 ( .A1(n151), .A2(n152), .ZN(n146) );
  BUFFD0 U158 ( .I(Sel), .Z(n193) );
  CKND0 U159 ( .CLK(A[21]), .CN(n154) );
  NR2D0 U160 ( .A1(n147), .A2(n154), .ZN(n155) );
  NR2D0 U161 ( .A1(n185), .A2(n115), .ZN(n156) );
  NR2XD0 U162 ( .A1(n155), .A2(n156), .ZN(n153) );
  INVD1 U163 ( .I(B[21]), .ZN(n185) );
  CKND0 U164 ( .CLK(A[0]), .CN(n158) );
  CKND0 U165 ( .CLK(n192), .CN(n159) );
  CKND0 U166 ( .CLK(B[0]), .CN(n160) );
  NR2D0 U167 ( .A1(n121), .A2(n158), .ZN(n161) );
  NR2D0 U168 ( .A1(n159), .A2(n160), .ZN(n162) );
  NR2XD0 U169 ( .A1(n161), .A2(n162), .ZN(n157) );
  INVD0 U170 ( .I(n192), .ZN(n164) );
  CKND0 U171 ( .CLK(B[16]), .CN(n165) );
  NR2D0 U172 ( .A1(n164), .A2(n165), .ZN(n166) );
  NR2D0 U173 ( .A1(n181), .A2(n192), .ZN(n167) );
  NR2XD0 U174 ( .A1(n166), .A2(n167), .ZN(n163) );
  INVD1 U175 ( .I(A[16]), .ZN(n181) );
  INVD0 U176 ( .I(n193), .ZN(n169) );
  CKND0 U177 ( .CLK(A[15]), .CN(n170) );
  INVD0 U178 ( .I(n192), .ZN(n171) );
  INVD1 U179 ( .I(B[15]), .ZN(n172) );
  NR2D0 U180 ( .A1(n169), .A2(n170), .ZN(n173) );
  NR2D0 U181 ( .A1(n171), .A2(n172), .ZN(n174) );
  NR2XD0 U182 ( .A1(n173), .A2(n174), .ZN(n168) );
  INVD1 U183 ( .I(B[8]), .ZN(n179) );
  INVD1 U184 ( .I(A[8]), .ZN(n180) );
  INVD1 U185 ( .I(B[19]), .ZN(n176) );
  INVD1 U186 ( .I(A[19]), .ZN(n177) );
  INVD1 U187 ( .I(B[30]), .ZN(n190) );
  INVD1 U188 ( .I(A[30]), .ZN(n191) );
  INVD1 U189 ( .I(B[31]), .ZN(n183) );
  INVD1 U190 ( .I(A[31]), .ZN(n184) );
  INVD1 U191 ( .I(A[22]), .ZN(n188) );
  INVD1 U192 ( .I(A[28]), .ZN(n187) );
  CKND0 U193 ( .CLK(n194), .CN(n186) );
  IOA22D0 U194 ( .B1(n187), .B2(n121), .A1(B[28]), .A2(n121), .ZN(n194) );
  AO22D0 U195 ( .A1(B[9]), .A2(n121), .B1(n164), .B2(A[9]), .Z(Out[9]) );
  AO22D0 U196 ( .A1(B[23]), .A2(n121), .B1(A[23]), .B2(n171), .Z(Out[23]) );
  AO22D0 U197 ( .A1(B[24]), .A2(n121), .B1(A[24]), .B2(n137), .Z(Out[24]) );
endmodule

