
module FIFO_Top ( Dout, Din, ReadIn, WriteIn, Clocker, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, Clocker, Reseter;
  wire   E_FIFO, F_FIFO, Mem_Enable, ReadWire, WriteWire, _0_net_, n4, n5;
  wire   [4:0] SM_MemAddr;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(E_FIFO), .FullFIFO(F_FIFO), .ReadCmd(ReadWire), .WriteCmd(
        WriteWire), .ReadReq(ReadIn), .WriteReq(WriteIn), .Clk(Clocker), 
        .Reset(Reseter) );
  Mem1kx32gen RegFile1 ( .DataO(Dout), .DataI(Din), .Addr(SM_MemAddr), 
        .ClockIn(_0_net_), .ChipEna(Mem_Enable), .Read(ReadWire), .Write(
        WriteWire) );
  INVD1 U10 ( .I(n5), .ZN(n4) );
  INR2D1 U11 ( .A1(ReadWire), .B1(WriteWire), .ZN(n5) );
  AO22D0 U12 ( .A1(SM_WriteAddr[2]), .A2(n4), .B1(SM_ReadAddr[2]), .B2(n5), 
        .Z(SM_MemAddr[2]) );
  AO22D0 U13 ( .A1(SM_WriteAddr[4]), .A2(n4), .B1(SM_ReadAddr[4]), .B2(n5), 
        .Z(SM_MemAddr[4]) );
  AO22D0 U14 ( .A1(SM_WriteAddr[0]), .A2(n4), .B1(SM_ReadAddr[0]), .B2(n5), 
        .Z(SM_MemAddr[0]) );
  AO22D0 U15 ( .A1(SM_WriteAddr[3]), .A2(n4), .B1(SM_ReadAddr[3]), .B2(n5), 
        .Z(SM_MemAddr[3]) );
  AO22D0 U16 ( .A1(SM_WriteAddr[1]), .A2(n4), .B1(SM_ReadAddr[1]), .B2(n5), 
        .Z(SM_MemAddr[1]) );
  AOI211D1 U17 ( .A1(WriteWire), .A2(ReadWire), .B(F_FIFO), .C(E_FIFO), .ZN(
        Mem_Enable) );
  INVD1 U18 ( .I(Clocker), .ZN(_0_net_) );
endmodule


module FIFOStateM ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, Clk, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, Clk, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N72, N73, N74, N75, N76, N88, N89, N90, N91, N92,
         N93, N95, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N144, N146, N148, N150, N152, N155,
         N158, N161, N164, N167, N169, N172, N175, N178, N181, N184, N186,
         N187, N190, N191, N200, N201, N202, N211, N212, N213, N214, N217,
         N220, N223, N226, N229, N232, N235, N238, N241, n2, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n1, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n73, n74, n75,
         n76;
  wire   [2:0] CurState;
  wire   [2:0] NextState;

  LHQD1 \WriteCount_tri_enable_reg[0]  ( .E(N200), .D(N201), .Q(N9) );
  LHQD1 \NextState_reg[0]  ( .E(N190), .D(N144), .Q(NextState[0]) );
  LHQD1 \WriteCount_reg[1]  ( .E(N200), .D(N155), .Q(N238) );
  LHQD1 \ReadCount_reg[1]  ( .E(N211), .D(N172), .Q(N223) );
  LHQD1 \NextState_reg[1]  ( .E(N190), .D(N146), .Q(NextState[1]) );
  LHQD1 \NextState_reg[2]  ( .E(N190), .D(N148), .Q(NextState[2]) );
  LHQD1 EmptyFIFOReg_reg ( .E(N213), .D(N184), .Q(EmptyFIFO) );
  LHQD1 WriteCmdReg_reg ( .E(N202), .D(N167), .Q(WriteCmd) );
  LHQD1 FullFIFOReg_reg ( .E(N191), .D(N150), .Q(FullFIFO) );
  LHQD1 \WriteCount_tri_enable_reg[4]  ( .E(N200), .D(N201), .Q(N5) );
  LHQD1 \WriteCount_tri_enable_reg[2]  ( .E(N200), .D(N201), .Q(N7) );
  LHQD1 \WriteCount_tri_enable_reg[1]  ( .E(N200), .D(N201), .Q(N8) );
  LHQD1 \WriteCount_tri_enable_reg[3]  ( .E(N200), .D(N201), .Q(N6) );
  LHQD1 \ReadCount_tri_enable_reg[4]  ( .E(N211), .D(N212), .Q(N0) );
  LHQD1 \ReadCount_tri_enable_reg[2]  ( .E(N211), .D(N212), .Q(N2) );
  LHQD1 \ReadCount_tri_enable_reg[0]  ( .E(N211), .D(N212), .Q(N4) );
  LHQD1 \ReadCount_tri_enable_reg[1]  ( .E(N211), .D(N212), .Q(N3) );
  LHQD1 \ReadCount_tri_enable_reg[3]  ( .E(N211), .D(N212), .Q(N1) );
  LHQD1 ReadCmdReg_reg ( .E(N187), .D(N186), .Q(ReadCmd) );
  LHQD1 \ReadCount_reg[0]  ( .E(N211), .D(N169), .Q(N226) );
  LHQD1 \ReadCount_reg[4]  ( .E(N211), .D(N181), .Q(N214) );
  LHQD1 \WriteCount_reg[4]  ( .E(N200), .D(N164), .Q(N229) );
  LHQD1 \WriteCount_reg[3]  ( .E(N200), .D(N161), .Q(N232) );
  LHQD1 \WriteCount_reg[2]  ( .E(N200), .D(N158), .Q(N235) );
  LHQD1 \ReadCount_reg[2]  ( .E(N211), .D(N175), .Q(N220) );
  LHQD1 \ReadCount_reg[3]  ( .E(N211), .D(N178), .Q(N217) );
  LHQD1 \WriteCount_reg[0]  ( .E(N200), .D(N152), .Q(N241) );
  BUFTD1 \WriteCount_tri[0]  ( .I(N241), .OE(n70), .Z(WriteAddr[0]) );
  BUFTD1 \WriteCount_tri[1]  ( .I(N238), .OE(n69), .Z(WriteAddr[1]) );
  BUFTD1 \WriteCount_tri[2]  ( .I(N235), .OE(n68), .Z(WriteAddr[2]) );
  BUFTD1 \WriteCount_tri[3]  ( .I(N232), .OE(n67), .Z(WriteAddr[3]) );
  BUFTD1 \WriteCount_tri[4]  ( .I(N229), .OE(n66), .Z(WriteAddr[4]) );
  BUFTD1 \ReadCount_tri[0]  ( .I(N226), .OE(n65), .Z(ReadAddr[0]) );
  BUFTD1 \ReadCount_tri[1]  ( .I(N223), .OE(n64), .Z(ReadAddr[1]) );
  BUFTD1 \ReadCount_tri[2]  ( .I(N220), .OE(n63), .Z(ReadAddr[2]) );
  BUFTD1 \ReadCount_tri[3]  ( .I(N217), .OE(n62), .Z(ReadAddr[3]) );
  BUFTD1 \ReadCount_tri[4]  ( .I(N214), .OE(n61), .Z(ReadAddr[4]) );
  MOAI22D1 U25 ( .A1(Clk), .A2(n26), .B1(n20), .B2(N213), .ZN(N200) );
  OA21D1 U27 ( .A1(n29), .A2(n21), .B(n30), .Z(n26) );
  AO222D1 U60 ( .A1(ReadAddr[4]), .A2(n33), .B1(N54), .B2(n43), .C1(N76), .C2(
        n52), .Z(N164) );
  AO222D1 U61 ( .A1(ReadAddr[3]), .A2(n33), .B1(N53), .B2(n43), .C1(N75), .C2(
        n52), .Z(N161) );
  AO222D1 U62 ( .A1(ReadAddr[2]), .A2(n33), .B1(N52), .B2(n43), .C1(N74), .C2(
        n52), .Z(N158) );
  AO222D1 U63 ( .A1(ReadAddr[1]), .A2(n33), .B1(N51), .B2(n43), .C1(N73), .C2(
        n52), .Z(N155) );
  AO222D1 U64 ( .A1(ReadAddr[0]), .A2(n33), .B1(N50), .B2(n43), .C1(N72), .C2(
        n52), .Z(N152) );
  FIFOStateM_DW01_inc_0 add_210 ( .A({n2, N105, N104, N103, N102, N101}), 
        .SUM({N111, N110, N109, N108, N107, N106}) );
  FIFOStateM_DW01_inc_1 add_198 ( .A({n2, N76, N75, N74, N73, N72}), .SUM({N93, 
        N92, N91, N90, N89, N88}) );
  FIFOStateM_DW01_inc_2 add_110_C147 ( .A({N45, N46, N47, N48, N49}), .SUM({
        N54, N53, N52, N51, N50}) );
  FIFOStateM_DW01_inc_3 r109 ( .A(ReadAddr), .SUM({N105, N104, N103, N102, 
        N101}) );
  FIFOStateM_DW01_inc_4 r106 ( .A(WriteAddr), .SUM({N76, N75, N74, N73, N72})
         );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(Clk), .CDN(n71), .Q(n58), 
        .QN(n72) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(Clk), .CDN(n71), .Q(
        CurState[2]), .QN(n36) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(Clk), .CDN(n71), .Q(
        CurState[0]), .QN(n41) );
  NR3D0 U3 ( .A1(n41), .A2(n72), .A3(n36), .ZN(n33) );
  INVD1 U4 ( .I(n47), .ZN(n42) );
  INVD1 U5 ( .I(n43), .ZN(n51) );
  NR2D1 U6 ( .A1(n27), .A2(n21), .ZN(n43) );
  INVD1 U7 ( .I(n53), .ZN(n52) );
  INVD1 U8 ( .I(n50), .ZN(n31) );
  NR2D1 U9 ( .A1(n52), .A2(n50), .ZN(n47) );
  OAI21D1 U10 ( .A1(n47), .A2(n46), .B(n51), .ZN(N167) );
  NR2D1 U11 ( .A1(n54), .A2(n46), .ZN(N150) );
  INVD1 U12 ( .I(n25), .ZN(N186) );
  INVD1 U13 ( .I(n38), .ZN(n48) );
  INVD1 U14 ( .I(n23), .ZN(N211) );
  NR3D0 U15 ( .A1(n41), .A2(n58), .A3(n36), .ZN(n50) );
  AOI21D1 U16 ( .A1(n42), .A2(n46), .B(n33), .ZN(n25) );
  OAI221D0 U17 ( .A1(n46), .A2(n53), .B1(N112), .B2(n29), .C(n59), .ZN(N144)
         );
  NR2D1 U18 ( .A1(n33), .A2(n50), .ZN(n59) );
  INVD1 U19 ( .I(n32), .ZN(n27) );
  OAI21D1 U20 ( .A1(n46), .A2(n55), .B(n54), .ZN(N148) );
  AOI21D1 U21 ( .A1(N95), .A2(n49), .B(n50), .ZN(n55) );
  INVD1 U22 ( .I(n49), .ZN(n29) );
  NR2D1 U23 ( .A1(n40), .A2(n49), .ZN(n53) );
  INVD1 U24 ( .I(n33), .ZN(n54) );
  NR2D1 U26 ( .A1(n27), .A2(n20), .ZN(N184) );
  ND3D1 U28 ( .A1(n51), .A2(n31), .A3(n56), .ZN(N146) );
  AOI22D0 U29 ( .A1(n49), .A2(n57), .B1(n40), .B2(n39), .ZN(n56) );
  ND2D1 U30 ( .A1(N95), .A2(n39), .ZN(n57) );
  AN2D1 U31 ( .A1(N150), .A2(n22), .Z(N201) );
  AN2D1 U32 ( .A1(N184), .A2(n22), .Z(N212) );
  AO22D0 U33 ( .A1(n32), .A2(N45), .B1(N105), .B2(n48), .Z(N181) );
  AO22D0 U34 ( .A1(n32), .A2(N49), .B1(N101), .B2(n48), .Z(N169) );
  AO22D0 U35 ( .A1(n32), .A2(N48), .B1(N102), .B2(n48), .Z(N172) );
  AO22D0 U36 ( .A1(n32), .A2(N46), .B1(N104), .B2(n48), .Z(N178) );
  AO22D0 U37 ( .A1(n32), .A2(N47), .B1(N103), .B2(n48), .Z(N175) );
  NR3D0 U38 ( .A1(n33), .A2(n49), .A3(n50), .ZN(n38) );
  INVD1 U39 ( .I(n39), .ZN(n46) );
  INVD1 U40 ( .I(n20), .ZN(n21) );
  OAI21D1 U41 ( .A1(n45), .A2(n32), .B(n22), .ZN(n23) );
  NR2D1 U42 ( .A1(n38), .A2(n39), .ZN(n45) );
  INVD1 U43 ( .I(n40), .ZN(n28) );
  INVD1 U44 ( .I(N0), .ZN(n61) );
  INVD1 U45 ( .I(N1), .ZN(n62) );
  INVD1 U46 ( .I(N2), .ZN(n63) );
  INVD1 U47 ( .I(N3), .ZN(n64) );
  INVD1 U48 ( .I(N4), .ZN(n65) );
  INVD1 U49 ( .I(N5), .ZN(n66) );
  INVD1 U50 ( .I(N6), .ZN(n67) );
  INVD1 U51 ( .I(N7), .ZN(n68) );
  INVD1 U52 ( .I(N8), .ZN(n69) );
  INVD1 U53 ( .I(N9), .ZN(n70) );
  NR3D0 U54 ( .A1(CurState[2]), .A2(n72), .A3(n41), .ZN(n49) );
  NR3D0 U55 ( .A1(CurState[2]), .A2(n72), .A3(CurState[0]), .ZN(n40) );
  NR3D0 U56 ( .A1(CurState[0]), .A2(CurState[2]), .A3(n58), .ZN(n32) );
  INR2D1 U57 ( .A1(WriteAddr[1]), .B1(Reset), .ZN(N48) );
  INR2D1 U58 ( .A1(WriteAddr[2]), .B1(Reset), .ZN(N47) );
  INR2D1 U59 ( .A1(WriteAddr[3]), .B1(Reset), .ZN(N46) );
  INR2D1 U65 ( .A1(WriteAddr[4]), .B1(Reset), .ZN(N45) );
  AO22D0 U66 ( .A1(n20), .A2(N73), .B1(n21), .B2(WriteAddr[1]), .Z(N99) );
  AN2D1 U67 ( .A1(WriteAddr[0]), .A2(n71), .Z(N49) );
  AO22D0 U68 ( .A1(n21), .A2(WriteAddr[0]), .B1(n20), .B2(N72), .Z(N100) );
  INVD1 U69 ( .I(Clk), .ZN(n22) );
  XNR2D1 U70 ( .A1(n1), .A2(N109), .ZN(n73) );
  AOI22D0 U71 ( .A1(n20), .A2(N75), .B1(n21), .B2(WriteAddr[3]), .ZN(n1) );
  AO22D0 U72 ( .A1(n20), .A2(N74), .B1(n21), .B2(WriteAddr[2]), .Z(N98) );
  XNR2D1 U73 ( .A1(n3), .A2(N110), .ZN(n75) );
  AOI22D0 U74 ( .A1(n20), .A2(N76), .B1(n21), .B2(WriteAddr[4]), .ZN(n3) );
  ND2D1 U75 ( .A1(ReadReq), .A2(n60), .ZN(n39) );
  NR2D1 U76 ( .A1(n60), .A2(ReadReq), .ZN(n20) );
  INVD1 U77 ( .I(WriteReq), .ZN(n60) );
  INVD1 U78 ( .I(Reset), .ZN(n71) );
  AOI221D0 U79 ( .A1(n42), .A2(n20), .B1(Reset), .B2(n32), .C(n43), .ZN(n24)
         );
  AOI21D1 U80 ( .A1(Reset), .A2(n32), .B(n33), .ZN(n30) );
  AOI31D0 U81 ( .A1(n24), .A2(n34), .A3(n35), .B(Clk), .ZN(N190) );
  ND2D1 U82 ( .A1(CurState[2]), .A2(n41), .ZN(n34) );
  AOI31D0 U83 ( .A1(n72), .A2(n36), .A3(CurState[0]), .B(n37), .ZN(n35) );
  AOI21D1 U84 ( .A1(n38), .A2(n28), .B(n39), .ZN(n37) );
  AOI21D1 U85 ( .A1(n27), .A2(n28), .B(Clk), .ZN(N213) );
  OAI21D1 U86 ( .A1(Clk), .A2(n44), .B(n23), .ZN(N187) );
  AOI22D0 U87 ( .A1(n20), .A2(n42), .B1(n40), .B2(n46), .ZN(n44) );
  AOI21D1 U88 ( .A1(n30), .A2(n31), .B(Clk), .ZN(N191) );
  AOI21D1 U89 ( .A1(n24), .A2(n25), .B(Clk), .ZN(N202) );
  TIEL U90 ( .ZN(n2) );
  INR2D0 U91 ( .A1(N88), .B1(ReadAddr[0]), .ZN(n5) );
  CKND0 U92 ( .CLK(ReadAddr[1]), .CN(n4) );
  OAI22D0 U93 ( .A1(n5), .A2(n4), .B1(N89), .B2(n5), .ZN(n9) );
  INR2D0 U94 ( .A1(ReadAddr[0]), .B1(N88), .ZN(n7) );
  CKND0 U95 ( .CLK(N89), .CN(n6) );
  OAI22D0 U96 ( .A1(ReadAddr[1]), .A2(n7), .B1(n7), .B2(n6), .ZN(n8) );
  IND3D0 U97 ( .A1(N93), .B1(n9), .B2(n8), .ZN(n13) );
  CKXOR2D0 U98 ( .A1(N92), .A2(ReadAddr[4]), .Z(n12) );
  CKXOR2D0 U99 ( .A1(N90), .A2(ReadAddr[2]), .Z(n11) );
  CKXOR2D0 U100 ( .A1(N91), .A2(ReadAddr[3]), .Z(n10) );
  NR4D0 U101 ( .A1(n13), .A2(n12), .A3(n11), .A4(n10), .ZN(N95) );
  INR2D0 U102 ( .A1(N106), .B1(N100), .ZN(n15) );
  CKND0 U103 ( .CLK(N99), .CN(n14) );
  OAI22D0 U104 ( .A1(N107), .A2(n15), .B1(n15), .B2(n14), .ZN(n19) );
  INR2D0 U105 ( .A1(N100), .B1(N106), .ZN(n17) );
  CKND0 U106 ( .CLK(N107), .CN(n16) );
  OAI22D0 U107 ( .A1(n17), .A2(n16), .B1(N99), .B2(n17), .ZN(n18) );
  IND3D0 U108 ( .A1(N111), .B1(n19), .B2(n18), .ZN(n76) );
  CKXOR2D0 U109 ( .A1(N98), .A2(N108), .Z(n74) );
  NR4D0 U110 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N112) );
endmodule


module Mem1kx32gen ( Dready, ParityErr, DataO, DataI, Addr, ClockIn, ChipEna, 
        Read, Write );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] Addr;
  input ClockIn, ChipEna, Read, Write;
  output Dready, ParityErr;
  wire   ChipClock, \WordArray[0].Word[0].QWire , \WordArray[0].Word[1].QWire ,
         \WordArray[0].Word[2].QWire , \WordArray[0].Word[3].QWire ,
         \WordArray[0].Word[4].QWire , \WordArray[0].Word[5].QWire ,
         \WordArray[0].Word[6].QWire , \WordArray[0].Word[7].QWire ,
         \WordArray[0].Word[8].QWire , \WordArray[0].Word[9].QWire , _9_net_,
         \WordArray[0].Word[10].QWire , \WordArray[0].Word[11].QWire ,
         \WordArray[0].Word[12].QWire , \WordArray[0].Word[13].QWire ,
         \WordArray[0].Word[14].QWire , \WordArray[0].Word[15].QWire ,
         \WordArray[0].Word[16].QWire , \WordArray[0].Word[17].QWire ,
         \WordArray[0].Word[18].QWire , \WordArray[0].Word[19].QWire ,
         \WordArray[0].Word[20].QWire , \WordArray[0].Word[21].QWire ,
         \WordArray[0].Word[22].QWire , \WordArray[0].Word[23].QWire ,
         \WordArray[0].Word[24].QWire , \WordArray[0].Word[25].QWire ,
         \WordArray[0].Word[26].QWire , \WordArray[0].Word[27].QWire ,
         \WordArray[0].Word[28].QWire , \WordArray[0].Word[29].QWire ,
         \WordArray[0].Word[30].QWire , \WordArray[0].Word[31].QWire ,
         \WordArray[1].Word[0].QWire , \WordArray[1].Word[1].QWire ,
         \WordArray[1].Word[2].QWire , \WordArray[1].Word[3].QWire ,
         \WordArray[1].Word[4].QWire , \WordArray[1].Word[5].QWire ,
         \WordArray[1].Word[6].QWire , \WordArray[1].Word[7].QWire ,
         \WordArray[1].Word[8].QWire , \WordArray[1].Word[9].QWire ,
         \WordArray[1].Word[10].QWire , \WordArray[1].Word[11].QWire ,
         \WordArray[1].Word[12].QWire , \WordArray[1].Word[13].QWire ,
         \WordArray[1].Word[14].QWire , \WordArray[1].Word[15].QWire ,
         \WordArray[1].Word[16].QWire , \WordArray[1].Word[17].QWire ,
         \WordArray[1].Word[18].QWire , \WordArray[1].Word[19].QWire ,
         \WordArray[1].Word[20].QWire , \WordArray[1].Word[21].QWire ,
         \WordArray[1].Word[22].QWire , \WordArray[1].Word[23].QWire ,
         \WordArray[1].Word[24].QWire , \WordArray[1].Word[25].QWire ,
         \WordArray[1].Word[26].QWire , \WordArray[1].Word[27].QWire ,
         \WordArray[1].Word[28].QWire , \WordArray[1].Word[29].QWire ,
         \WordArray[1].Word[30].QWire , \WordArray[1].Word[31].QWire ,
         _65_net_, \WordArray[2].Word[0].QWire , \WordArray[2].Word[1].QWire ,
         \WordArray[2].Word[2].QWire , \WordArray[2].Word[3].QWire ,
         \WordArray[2].Word[4].QWire , \WordArray[2].Word[5].QWire ,
         \WordArray[2].Word[6].QWire , \WordArray[2].Word[7].QWire ,
         \WordArray[2].Word[8].QWire , \WordArray[2].Word[9].QWire ,
         \WordArray[2].Word[10].QWire , \WordArray[2].Word[11].QWire ,
         \WordArray[2].Word[12].QWire , \WordArray[2].Word[13].QWire ,
         \WordArray[2].Word[14].QWire , \WordArray[2].Word[15].QWire ,
         \WordArray[2].Word[16].QWire , \WordArray[2].Word[17].QWire ,
         \WordArray[2].Word[18].QWire , \WordArray[2].Word[19].QWire ,
         \WordArray[2].Word[20].QWire , \WordArray[2].Word[21].QWire ,
         \WordArray[2].Word[22].QWire , \WordArray[2].Word[23].QWire ,
         \WordArray[2].Word[24].QWire , \WordArray[2].Word[25].QWire ,
         \WordArray[2].Word[26].QWire , \WordArray[2].Word[27].QWire ,
         \WordArray[2].Word[28].QWire , \WordArray[2].Word[29].QWire ,
         \WordArray[2].Word[30].QWire , \WordArray[2].Word[31].QWire ,
         _98_net_, \WordArray[3].Word[0].QWire , _99_net_,
         \WordArray[3].Word[1].QWire , \WordArray[3].Word[2].QWire ,
         \WordArray[3].Word[3].QWire , \WordArray[3].Word[4].QWire ,
         \WordArray[3].Word[5].QWire , \WordArray[3].Word[6].QWire ,
         \WordArray[3].Word[7].QWire , \WordArray[3].Word[8].QWire ,
         \WordArray[3].Word[9].QWire , \WordArray[3].Word[10].QWire ,
         \WordArray[3].Word[11].QWire , \WordArray[3].Word[12].QWire ,
         \WordArray[3].Word[13].QWire , \WordArray[3].Word[14].QWire ,
         \WordArray[3].Word[15].QWire , \WordArray[3].Word[16].QWire ,
         \WordArray[3].Word[17].QWire , \WordArray[3].Word[18].QWire ,
         \WordArray[3].Word[19].QWire , \WordArray[3].Word[20].QWire ,
         \WordArray[3].Word[21].QWire , \WordArray[3].Word[22].QWire ,
         \WordArray[3].Word[23].QWire , \WordArray[3].Word[24].QWire ,
         \WordArray[3].Word[25].QWire , \WordArray[3].Word[26].QWire ,
         \WordArray[3].Word[27].QWire , \WordArray[3].Word[28].QWire ,
         \WordArray[3].Word[29].QWire , \WordArray[3].Word[30].QWire ,
         \WordArray[3].Word[31].QWire , \WordArray[4].Word[0].QWire ,
         \WordArray[4].Word[1].QWire , \WordArray[4].Word[2].QWire ,
         \WordArray[4].Word[3].QWire , \WordArray[4].Word[4].QWire ,
         \WordArray[4].Word[5].QWire , \WordArray[4].Word[6].QWire ,
         \WordArray[4].Word[7].QWire , \WordArray[4].Word[8].QWire ,
         \WordArray[4].Word[9].QWire , \WordArray[4].Word[10].QWire ,
         \WordArray[4].Word[11].QWire , \WordArray[4].Word[12].QWire ,
         \WordArray[4].Word[13].QWire , \WordArray[4].Word[14].QWire ,
         \WordArray[4].Word[15].QWire , \WordArray[4].Word[16].QWire ,
         \WordArray[4].Word[17].QWire , \WordArray[4].Word[18].QWire ,
         \WordArray[4].Word[19].QWire , \WordArray[4].Word[20].QWire ,
         \WordArray[4].Word[21].QWire , \WordArray[4].Word[22].QWire ,
         \WordArray[4].Word[23].QWire , \WordArray[4].Word[24].QWire ,
         \WordArray[4].Word[25].QWire , \WordArray[4].Word[26].QWire ,
         \WordArray[4].Word[27].QWire , \WordArray[4].Word[28].QWire ,
         \WordArray[4].Word[29].QWire , \WordArray[4].Word[30].QWire ,
         \WordArray[4].Word[31].QWire , _164_net_,
         \WordArray[5].Word[0].QWire , \WordArray[5].Word[1].QWire ,
         \WordArray[5].Word[2].QWire , \WordArray[5].Word[3].QWire ,
         \WordArray[5].Word[4].QWire , \WordArray[5].Word[5].QWire ,
         \WordArray[5].Word[6].QWire , \WordArray[5].Word[7].QWire ,
         \WordArray[5].Word[8].QWire , \WordArray[5].Word[9].QWire ,
         \WordArray[5].Word[10].QWire , \WordArray[5].Word[11].QWire ,
         \WordArray[5].Word[12].QWire , \WordArray[5].Word[13].QWire ,
         \WordArray[5].Word[14].QWire , \WordArray[5].Word[15].QWire ,
         \WordArray[5].Word[16].QWire , \WordArray[5].Word[17].QWire ,
         \WordArray[5].Word[18].QWire , \WordArray[5].Word[19].QWire ,
         \WordArray[5].Word[20].QWire , \WordArray[5].Word[21].QWire ,
         \WordArray[5].Word[22].QWire , \WordArray[5].Word[23].QWire ,
         \WordArray[5].Word[24].QWire , \WordArray[5].Word[25].QWire ,
         \WordArray[5].Word[26].QWire , \WordArray[5].Word[27].QWire ,
         \WordArray[5].Word[28].QWire , \WordArray[5].Word[29].QWire ,
         \WordArray[5].Word[30].QWire , \WordArray[5].Word[31].QWire ,
         _197_net_, \WordArray[6].Word[0].QWire , \WordArray[6].Word[1].QWire ,
         \WordArray[6].Word[2].QWire , \WordArray[6].Word[3].QWire ,
         \WordArray[6].Word[4].QWire , \WordArray[6].Word[5].QWire ,
         \WordArray[6].Word[6].QWire , \WordArray[6].Word[7].QWire ,
         \WordArray[6].Word[8].QWire , \WordArray[6].Word[9].QWire ,
         \WordArray[6].Word[10].QWire , \WordArray[6].Word[11].QWire ,
         \WordArray[6].Word[12].QWire , \WordArray[6].Word[13].QWire ,
         \WordArray[6].Word[14].QWire , \WordArray[6].Word[15].QWire ,
         \WordArray[6].Word[16].QWire , \WordArray[6].Word[17].QWire ,
         \WordArray[6].Word[18].QWire , \WordArray[6].Word[19].QWire ,
         \WordArray[6].Word[20].QWire , \WordArray[6].Word[21].QWire ,
         \WordArray[6].Word[22].QWire , \WordArray[6].Word[23].QWire ,
         \WordArray[6].Word[24].QWire , \WordArray[6].Word[25].QWire ,
         \WordArray[6].Word[26].QWire , \WordArray[6].Word[27].QWire ,
         \WordArray[6].Word[28].QWire , \WordArray[6].Word[29].QWire ,
         \WordArray[6].Word[30].QWire , \WordArray[6].Word[31].QWire ,
         _230_net_, \WordArray[7].Word[0].QWire , \WordArray[7].Word[1].QWire ,
         \WordArray[7].Word[2].QWire , \WordArray[7].Word[3].QWire ,
         \WordArray[7].Word[4].QWire , \WordArray[7].Word[5].QWire ,
         \WordArray[7].Word[6].QWire , \WordArray[7].Word[7].QWire ,
         \WordArray[7].Word[8].QWire , \WordArray[7].Word[9].QWire ,
         \WordArray[7].Word[10].QWire , \WordArray[7].Word[11].QWire ,
         \WordArray[7].Word[12].QWire , \WordArray[7].Word[13].QWire ,
         \WordArray[7].Word[14].QWire , \WordArray[7].Word[15].QWire ,
         \WordArray[7].Word[16].QWire , \WordArray[7].Word[17].QWire ,
         \WordArray[7].Word[18].QWire , \WordArray[7].Word[19].QWire ,
         \WordArray[7].Word[20].QWire , \WordArray[7].Word[21].QWire ,
         \WordArray[7].Word[22].QWire , \WordArray[7].Word[23].QWire ,
         \WordArray[7].Word[24].QWire , \WordArray[7].Word[25].QWire ,
         \WordArray[7].Word[26].QWire , \WordArray[7].Word[27].QWire ,
         \WordArray[7].Word[28].QWire , \WordArray[7].Word[29].QWire ,
         \WordArray[7].Word[30].QWire , \WordArray[7].Word[31].QWire ,
         _263_net_, \WordArray[8].Word[0].QWire , \WordArray[8].Word[1].QWire ,
         \WordArray[8].Word[2].QWire , \WordArray[8].Word[3].QWire ,
         \WordArray[8].Word[4].QWire , \WordArray[8].Word[5].QWire ,
         \WordArray[8].Word[6].QWire , \WordArray[8].Word[7].QWire ,
         \WordArray[8].Word[8].QWire , \WordArray[8].Word[9].QWire ,
         \WordArray[8].Word[10].QWire , \WordArray[8].Word[11].QWire ,
         \WordArray[8].Word[12].QWire , \WordArray[8].Word[13].QWire ,
         \WordArray[8].Word[14].QWire , \WordArray[8].Word[15].QWire ,
         \WordArray[8].Word[16].QWire , \WordArray[8].Word[17].QWire ,
         \WordArray[8].Word[18].QWire , \WordArray[8].Word[19].QWire ,
         \WordArray[8].Word[20].QWire , \WordArray[8].Word[21].QWire ,
         \WordArray[8].Word[22].QWire , \WordArray[8].Word[23].QWire ,
         \WordArray[8].Word[24].QWire , \WordArray[8].Word[25].QWire ,
         \WordArray[8].Word[26].QWire , \WordArray[8].Word[27].QWire ,
         \WordArray[8].Word[28].QWire , \WordArray[8].Word[29].QWire ,
         \WordArray[8].Word[30].QWire , \WordArray[8].Word[31].QWire ,
         _296_net_, \WordArray[9].Word[0].QWire , \WordArray[9].CoreIn[32] ,
         \WordArray[9].Word[1].QWire , \WordArray[9].Word[2].QWire ,
         \WordArray[9].Word[3].QWire , \WordArray[9].Word[4].QWire ,
         \WordArray[9].Word[5].QWire , \WordArray[9].Word[6].QWire ,
         \WordArray[9].Word[7].QWire , \WordArray[9].Word[8].QWire ,
         \WordArray[9].Word[9].QWire , \WordArray[9].Word[10].QWire ,
         \WordArray[9].Word[11].QWire , \WordArray[9].Word[12].QWire ,
         \WordArray[9].Word[13].QWire , \WordArray[9].Word[14].QWire ,
         \WordArray[9].Word[15].QWire , \WordArray[9].Word[16].QWire ,
         \WordArray[9].Word[17].QWire , \WordArray[9].Word[18].QWire ,
         \WordArray[9].Word[19].QWire , \WordArray[9].Word[20].QWire ,
         \WordArray[9].Word[21].QWire , \WordArray[9].Word[22].QWire ,
         \WordArray[9].Word[23].QWire , \WordArray[9].Word[24].QWire ,
         \WordArray[9].Word[25].QWire , \WordArray[9].Word[26].QWire ,
         \WordArray[9].Word[27].QWire , \WordArray[9].Word[28].QWire ,
         \WordArray[9].Word[29].QWire , \WordArray[9].Word[30].QWire ,
         \WordArray[9].Word[31].QWire , _329_net_,
         \WordArray[10].Word[0].QWire , \WordArray[10].Word[1].QWire ,
         \WordArray[10].Word[2].QWire , \WordArray[10].Word[3].QWire ,
         \WordArray[10].Word[4].QWire , \WordArray[10].Word[5].QWire ,
         \WordArray[10].Word[6].QWire , \WordArray[10].Word[7].QWire ,
         \WordArray[10].Word[8].QWire , \WordArray[10].Word[9].QWire ,
         \WordArray[10].Word[10].QWire , \WordArray[10].Word[11].QWire ,
         \WordArray[10].Word[12].QWire , \WordArray[10].Word[13].QWire ,
         \WordArray[10].Word[14].QWire , \WordArray[10].Word[15].QWire ,
         \WordArray[10].Word[16].QWire , \WordArray[10].Word[17].QWire ,
         \WordArray[10].Word[18].QWire , \WordArray[10].Word[19].QWire ,
         \WordArray[10].Word[20].QWire , \WordArray[10].Word[21].QWire ,
         \WordArray[10].Word[22].QWire , \WordArray[10].Word[23].QWire ,
         \WordArray[10].Word[24].QWire , \WordArray[10].Word[25].QWire ,
         \WordArray[10].Word[26].QWire , \WordArray[10].Word[27].QWire ,
         \WordArray[10].Word[28].QWire , \WordArray[10].Word[29].QWire ,
         \WordArray[10].Word[30].QWire , \WordArray[10].Word[31].QWire ,
         _362_net_, \WordArray[11].Word[0].QWire ,
         \WordArray[11].Word[1].QWire , \WordArray[11].Word[2].QWire ,
         \WordArray[11].Word[3].QWire , \WordArray[11].Word[4].QWire ,
         \WordArray[11].Word[5].QWire , \WordArray[11].Word[6].QWire ,
         \WordArray[11].Word[7].QWire , \WordArray[11].Word[8].QWire ,
         \WordArray[11].Word[9].QWire , \WordArray[11].Word[10].QWire ,
         \WordArray[11].Word[11].QWire , \WordArray[11].Word[12].QWire ,
         \WordArray[11].Word[13].QWire , \WordArray[11].Word[14].QWire ,
         \WordArray[11].Word[15].QWire , \WordArray[11].Word[16].QWire ,
         \WordArray[11].Word[17].QWire , \WordArray[11].Word[18].QWire ,
         \WordArray[11].Word[19].QWire , \WordArray[11].Word[20].QWire ,
         \WordArray[11].Word[21].QWire , \WordArray[11].Word[22].QWire ,
         \WordArray[11].Word[23].QWire , \WordArray[11].Word[24].QWire ,
         \WordArray[11].Word[25].QWire , \WordArray[11].Word[26].QWire ,
         \WordArray[11].Word[27].QWire , \WordArray[11].Word[28].QWire ,
         \WordArray[11].Word[29].QWire , \WordArray[11].Word[30].QWire ,
         \WordArray[11].Word[31].QWire , _395_net_,
         \WordArray[12].Word[0].QWire , \WordArray[12].Word[1].QWire ,
         \WordArray[12].Word[2].QWire , \WordArray[12].Word[3].QWire ,
         \WordArray[12].Word[4].QWire , \WordArray[12].Word[5].QWire ,
         \WordArray[12].Word[6].QWire , \WordArray[12].Word[7].QWire ,
         \WordArray[12].Word[8].QWire , \WordArray[12].Word[9].QWire ,
         \WordArray[12].Word[10].QWire , \WordArray[12].Word[11].QWire ,
         \WordArray[12].Word[12].QWire , \WordArray[12].Word[13].QWire ,
         \WordArray[12].Word[14].QWire , \WordArray[12].Word[15].QWire ,
         \WordArray[12].Word[16].QWire , \WordArray[12].Word[17].QWire ,
         \WordArray[12].Word[18].QWire , \WordArray[12].Word[19].QWire ,
         \WordArray[12].Word[20].QWire , \WordArray[12].Word[21].QWire ,
         \WordArray[12].Word[22].QWire , \WordArray[12].Word[23].QWire ,
         \WordArray[12].Word[24].QWire , \WordArray[12].Word[25].QWire ,
         \WordArray[12].Word[26].QWire , \WordArray[12].Word[27].QWire ,
         \WordArray[12].Word[28].QWire , \WordArray[12].Word[29].QWire ,
         \WordArray[12].Word[30].QWire , \WordArray[12].Word[31].QWire ,
         _428_net_, \WordArray[13].Word[0].QWire ,
         \WordArray[13].Word[1].QWire , \WordArray[13].Word[2].QWire ,
         \WordArray[13].Word[3].QWire , \WordArray[13].Word[4].QWire ,
         \WordArray[13].Word[5].QWire , \WordArray[13].Word[6].QWire ,
         \WordArray[13].Word[7].QWire , \WordArray[13].Word[8].QWire ,
         \WordArray[13].Word[9].QWire , \WordArray[13].Word[10].QWire ,
         \WordArray[13].Word[11].QWire , \WordArray[13].Word[12].QWire ,
         \WordArray[13].Word[13].QWire , \WordArray[13].Word[14].QWire ,
         \WordArray[13].Word[15].QWire , \WordArray[13].Word[16].QWire ,
         \WordArray[13].Word[17].QWire , \WordArray[13].Word[18].QWire ,
         \WordArray[13].Word[19].QWire , \WordArray[13].Word[20].QWire ,
         \WordArray[13].Word[21].QWire , \WordArray[13].Word[22].QWire ,
         \WordArray[13].Word[23].QWire , \WordArray[13].Word[24].QWire ,
         \WordArray[13].Word[25].QWire , \WordArray[13].Word[26].QWire ,
         \WordArray[13].Word[27].QWire , \WordArray[13].Word[28].QWire ,
         \WordArray[13].Word[29].QWire , \WordArray[13].Word[30].QWire ,
         \WordArray[13].Word[31].QWire , _461_net_,
         \WordArray[14].Word[0].QWire , \WordArray[14].Word[1].QWire ,
         \WordArray[14].Word[2].QWire , \WordArray[14].Word[3].QWire ,
         \WordArray[14].Word[4].QWire , \WordArray[14].Word[5].QWire ,
         \WordArray[14].Word[6].QWire , \WordArray[14].Word[7].QWire ,
         \WordArray[14].Word[8].QWire , \WordArray[14].Word[9].QWire ,
         \WordArray[14].Word[10].QWire , \WordArray[14].Word[11].QWire ,
         \WordArray[14].Word[12].QWire , \WordArray[14].Word[13].QWire ,
         \WordArray[14].Word[14].QWire , \WordArray[14].Word[15].QWire ,
         \WordArray[14].Word[16].QWire , \WordArray[14].Word[17].QWire ,
         \WordArray[14].Word[18].QWire , \WordArray[14].Word[19].QWire ,
         \WordArray[14].Word[20].QWire , \WordArray[14].Word[21].QWire ,
         \WordArray[14].Word[22].QWire , \WordArray[14].Word[23].QWire ,
         \WordArray[14].Word[24].QWire , \WordArray[14].Word[25].QWire ,
         \WordArray[14].Word[26].QWire , \WordArray[14].Word[27].QWire ,
         \WordArray[14].Word[28].QWire , \WordArray[14].Word[29].QWire ,
         \WordArray[14].Word[30].QWire , \WordArray[14].Word[31].QWire ,
         _494_net_, \WordArray[15].Word[0].QWire ,
         \WordArray[15].Word[1].QWire , \WordArray[15].Word[2].QWire ,
         \WordArray[15].Word[3].QWire , \WordArray[15].Word[4].QWire ,
         \WordArray[15].Word[5].QWire , \WordArray[15].Word[6].QWire ,
         \WordArray[15].Word[7].QWire , \WordArray[15].Word[8].QWire ,
         \WordArray[15].Word[9].QWire , \WordArray[15].Word[10].QWire ,
         \WordArray[15].Word[11].QWire , \WordArray[15].Word[12].QWire ,
         \WordArray[15].Word[13].QWire , \WordArray[15].Word[14].QWire ,
         \WordArray[15].Word[15].QWire , \WordArray[15].Word[16].QWire ,
         \WordArray[15].Word[17].QWire , \WordArray[15].Word[18].QWire ,
         \WordArray[15].Word[19].QWire , \WordArray[15].Word[20].QWire ,
         \WordArray[15].Word[21].QWire , \WordArray[15].Word[22].QWire ,
         \WordArray[15].Word[23].QWire , \WordArray[15].Word[24].QWire ,
         \WordArray[15].Word[25].QWire , \WordArray[15].Word[26].QWire ,
         \WordArray[15].Word[27].QWire , \WordArray[15].Word[28].QWire ,
         \WordArray[15].Word[29].QWire , \WordArray[15].Word[30].QWire ,
         \WordArray[15].Word[31].QWire , _527_net_,
         \WordArray[16].Word[0].QWire , \WordArray[16].Word[1].QWire ,
         \WordArray[16].Word[2].QWire , \WordArray[16].Word[3].QWire ,
         \WordArray[16].Word[4].QWire , \WordArray[16].Word[5].QWire ,
         \WordArray[16].Word[6].QWire , \WordArray[16].Word[7].QWire ,
         \WordArray[16].Word[8].QWire , \WordArray[16].Word[9].QWire ,
         \WordArray[16].Word[10].QWire , \WordArray[16].Word[11].QWire ,
         \WordArray[16].Word[12].QWire , \WordArray[16].Word[13].QWire ,
         \WordArray[16].Word[14].QWire , \WordArray[16].Word[15].QWire ,
         \WordArray[16].Word[16].QWire , \WordArray[16].Word[17].QWire ,
         \WordArray[16].Word[18].QWire , \WordArray[16].Word[19].QWire ,
         \WordArray[16].Word[20].QWire , \WordArray[16].Word[21].QWire ,
         \WordArray[16].Word[22].QWire , \WordArray[16].Word[23].QWire ,
         \WordArray[16].Word[24].QWire , \WordArray[16].Word[25].QWire ,
         \WordArray[16].Word[26].QWire , \WordArray[16].Word[27].QWire ,
         \WordArray[16].Word[28].QWire , \WordArray[16].Word[29].QWire ,
         \WordArray[16].Word[30].QWire , \WordArray[16].Word[31].QWire ,
         _560_net_, \WordArray[17].Word[0].QWire ,
         \WordArray[17].Word[1].QWire , \WordArray[17].Word[2].QWire ,
         \WordArray[17].Word[3].QWire , \WordArray[17].Word[4].QWire ,
         \WordArray[17].Word[5].QWire , \WordArray[17].Word[6].QWire ,
         \WordArray[17].Word[7].QWire , \WordArray[17].Word[8].QWire ,
         \WordArray[17].Word[9].QWire , \WordArray[17].Word[10].QWire ,
         \WordArray[17].Word[11].QWire , \WordArray[17].Word[12].QWire ,
         \WordArray[17].Word[13].QWire , \WordArray[17].Word[14].QWire ,
         \WordArray[17].Word[15].QWire , \WordArray[17].Word[16].QWire ,
         \WordArray[17].Word[17].QWire , \WordArray[17].Word[18].QWire ,
         \WordArray[17].Word[19].QWire , \WordArray[17].Word[20].QWire ,
         \WordArray[17].Word[21].QWire , \WordArray[17].Word[22].QWire ,
         \WordArray[17].Word[23].QWire , \WordArray[17].Word[24].QWire ,
         \WordArray[17].Word[25].QWire , \WordArray[17].Word[26].QWire ,
         \WordArray[17].Word[27].QWire , \WordArray[17].Word[28].QWire ,
         \WordArray[17].Word[29].QWire , \WordArray[17].Word[30].QWire ,
         \WordArray[17].Word[31].QWire , _593_net_,
         \WordArray[18].Word[0].QWire , \WordArray[18].Word[1].QWire ,
         \WordArray[18].Word[2].QWire , \WordArray[18].Word[3].QWire ,
         \WordArray[18].Word[4].QWire , \WordArray[18].Word[5].QWire ,
         \WordArray[18].Word[6].QWire , \WordArray[18].Word[7].QWire ,
         \WordArray[18].Word[8].QWire , \WordArray[18].Word[9].QWire ,
         \WordArray[18].Word[10].QWire , \WordArray[18].Word[11].QWire ,
         \WordArray[18].Word[12].QWire , \WordArray[18].Word[13].QWire ,
         \WordArray[18].Word[14].QWire , \WordArray[18].Word[15].QWire ,
         \WordArray[18].Word[16].QWire , \WordArray[18].Word[17].QWire ,
         \WordArray[18].Word[18].QWire , \WordArray[18].Word[19].QWire ,
         \WordArray[18].Word[20].QWire , \WordArray[18].Word[21].QWire ,
         \WordArray[18].Word[22].QWire , \WordArray[18].Word[23].QWire ,
         \WordArray[18].Word[24].QWire , \WordArray[18].Word[25].QWire ,
         \WordArray[18].Word[26].QWire , \WordArray[18].Word[27].QWire ,
         \WordArray[18].Word[28].QWire , \WordArray[18].Word[29].QWire ,
         \WordArray[18].Word[30].QWire , \WordArray[18].Word[31].QWire ,
         _626_net_, \WordArray[19].Word[0].QWire ,
         \WordArray[19].Word[1].QWire , \WordArray[19].Word[2].QWire ,
         \WordArray[19].Word[3].QWire , \WordArray[19].Word[4].QWire ,
         \WordArray[19].Word[5].QWire , \WordArray[19].Word[6].QWire ,
         \WordArray[19].Word[7].QWire , \WordArray[19].Word[8].QWire ,
         \WordArray[19].Word[9].QWire , \WordArray[19].Word[10].QWire ,
         \WordArray[19].Word[11].QWire , \WordArray[19].Word[12].QWire ,
         \WordArray[19].Word[13].QWire , \WordArray[19].Word[14].QWire ,
         \WordArray[19].Word[15].QWire , \WordArray[19].Word[16].QWire ,
         \WordArray[19].Word[17].QWire , \WordArray[19].Word[18].QWire ,
         \WordArray[19].Word[19].QWire , \WordArray[19].Word[20].QWire ,
         \WordArray[19].Word[21].QWire , \WordArray[19].Word[22].QWire ,
         \WordArray[19].Word[23].QWire , \WordArray[19].Word[24].QWire ,
         \WordArray[19].Word[25].QWire , \WordArray[19].Word[26].QWire ,
         \WordArray[19].Word[27].QWire , \WordArray[19].Word[28].QWire ,
         \WordArray[19].Word[29].QWire , \WordArray[19].Word[30].QWire ,
         \WordArray[19].Word[31].QWire , _659_net_,
         \WordArray[20].Word[0].QWire , \WordArray[20].Word[1].QWire ,
         \WordArray[20].Word[2].QWire , \WordArray[20].Word[3].QWire ,
         \WordArray[20].Word[4].QWire , \WordArray[20].Word[5].QWire ,
         \WordArray[20].Word[6].QWire , \WordArray[20].Word[7].QWire ,
         \WordArray[20].Word[8].QWire , \WordArray[20].Word[9].QWire ,
         \WordArray[20].Word[10].QWire , \WordArray[20].Word[11].QWire ,
         \WordArray[20].Word[12].QWire , \WordArray[20].Word[13].QWire ,
         \WordArray[20].Word[14].QWire , \WordArray[20].Word[15].QWire ,
         \WordArray[20].Word[16].QWire , \WordArray[20].Word[17].QWire ,
         \WordArray[20].Word[18].QWire , \WordArray[20].Word[19].QWire ,
         \WordArray[20].Word[20].QWire , \WordArray[20].Word[21].QWire ,
         \WordArray[20].Word[22].QWire , \WordArray[20].Word[23].QWire ,
         \WordArray[20].Word[24].QWire , \WordArray[20].Word[25].QWire ,
         \WordArray[20].Word[26].QWire , \WordArray[20].Word[27].QWire ,
         \WordArray[20].Word[28].QWire , \WordArray[20].Word[29].QWire ,
         \WordArray[20].Word[30].QWire , \WordArray[20].Word[31].QWire ,
         _692_net_, \WordArray[21].Word[0].QWire ,
         \WordArray[21].Word[1].QWire , \WordArray[21].Word[2].QWire ,
         \WordArray[21].Word[3].QWire , \WordArray[21].Word[4].QWire ,
         \WordArray[21].Word[5].QWire , \WordArray[21].Word[6].QWire ,
         \WordArray[21].Word[7].QWire , \WordArray[21].Word[8].QWire ,
         \WordArray[21].Word[9].QWire , \WordArray[21].Word[10].QWire ,
         \WordArray[21].Word[11].QWire , \WordArray[21].Word[12].QWire ,
         \WordArray[21].Word[13].QWire , \WordArray[21].Word[14].QWire ,
         \WordArray[21].Word[15].QWire , \WordArray[21].Word[16].QWire ,
         \WordArray[21].Word[17].QWire , \WordArray[21].Word[18].QWire ,
         \WordArray[21].Word[19].QWire , \WordArray[21].Word[20].QWire ,
         \WordArray[21].Word[21].QWire , \WordArray[21].Word[22].QWire ,
         \WordArray[21].Word[23].QWire , \WordArray[21].Word[24].QWire ,
         \WordArray[21].Word[25].QWire , \WordArray[21].Word[26].QWire ,
         \WordArray[21].Word[27].QWire , \WordArray[21].Word[28].QWire ,
         \WordArray[21].Word[29].QWire , \WordArray[21].Word[30].QWire ,
         \WordArray[21].Word[31].QWire , _725_net_,
         \WordArray[22].Word[0].QWire , \WordArray[22].Word[1].QWire ,
         \WordArray[22].Word[2].QWire , \WordArray[22].Word[3].QWire ,
         \WordArray[22].Word[4].QWire , \WordArray[22].Word[5].QWire ,
         \WordArray[22].Word[6].QWire , \WordArray[22].Word[7].QWire ,
         \WordArray[22].Word[8].QWire , \WordArray[22].Word[9].QWire ,
         \WordArray[22].Word[10].QWire , \WordArray[22].Word[11].QWire ,
         \WordArray[22].Word[12].QWire , \WordArray[22].Word[13].QWire ,
         \WordArray[22].Word[14].QWire , \WordArray[22].Word[15].QWire ,
         \WordArray[22].Word[16].QWire , \WordArray[22].Word[17].QWire ,
         \WordArray[22].Word[18].QWire , \WordArray[22].Word[19].QWire ,
         \WordArray[22].Word[20].QWire , \WordArray[22].Word[21].QWire ,
         \WordArray[22].Word[22].QWire , \WordArray[22].Word[23].QWire ,
         \WordArray[22].Word[24].QWire , \WordArray[22].Word[25].QWire ,
         \WordArray[22].Word[26].QWire , \WordArray[22].Word[27].QWire ,
         \WordArray[22].Word[28].QWire , \WordArray[22].Word[29].QWire ,
         \WordArray[22].Word[30].QWire , \WordArray[22].Word[31].QWire ,
         _758_net_, \WordArray[23].Word[0].QWire ,
         \WordArray[23].Word[1].QWire , \WordArray[23].Word[2].QWire ,
         \WordArray[23].Word[3].QWire , \WordArray[23].Word[4].QWire ,
         \WordArray[23].Word[5].QWire , \WordArray[23].Word[6].QWire ,
         \WordArray[23].Word[7].QWire , \WordArray[23].Word[8].QWire ,
         \WordArray[23].Word[9].QWire , \WordArray[23].Word[10].QWire ,
         \WordArray[23].Word[11].QWire , \WordArray[23].Word[12].QWire ,
         \WordArray[23].Word[13].QWire , \WordArray[23].Word[14].QWire ,
         \WordArray[23].Word[15].QWire , \WordArray[23].Word[16].QWire ,
         \WordArray[23].Word[17].QWire , \WordArray[23].Word[18].QWire ,
         \WordArray[23].Word[19].QWire , \WordArray[23].Word[20].QWire ,
         \WordArray[23].Word[21].QWire , \WordArray[23].Word[22].QWire ,
         \WordArray[23].Word[23].QWire , \WordArray[23].Word[24].QWire ,
         \WordArray[23].Word[25].QWire , \WordArray[23].Word[26].QWire ,
         \WordArray[23].Word[27].QWire , \WordArray[23].Word[28].QWire ,
         \WordArray[23].Word[29].QWire , \WordArray[23].Word[30].QWire ,
         \WordArray[23].Word[31].QWire , _791_net_,
         \WordArray[24].Word[0].QWire , \WordArray[24].Word[1].QWire ,
         \WordArray[24].Word[2].QWire , \WordArray[24].Word[3].QWire ,
         \WordArray[24].Word[4].QWire , \WordArray[24].Word[5].QWire ,
         \WordArray[24].Word[6].QWire , \WordArray[24].Word[7].QWire ,
         \WordArray[24].Word[8].QWire , \WordArray[24].Word[9].QWire ,
         \WordArray[24].Word[10].QWire , \WordArray[24].Word[11].QWire ,
         \WordArray[24].Word[12].QWire , \WordArray[24].Word[13].QWire ,
         \WordArray[24].Word[14].QWire , \WordArray[24].Word[15].QWire ,
         \WordArray[24].Word[16].QWire , \WordArray[24].Word[17].QWire ,
         \WordArray[24].Word[18].QWire , \WordArray[24].Word[19].QWire ,
         \WordArray[24].Word[20].QWire , \WordArray[24].Word[21].QWire ,
         \WordArray[24].Word[22].QWire , \WordArray[24].Word[23].QWire ,
         \WordArray[24].Word[24].QWire , \WordArray[24].Word[25].QWire ,
         \WordArray[24].Word[26].QWire , \WordArray[24].Word[27].QWire ,
         \WordArray[24].Word[28].QWire , \WordArray[24].Word[29].QWire ,
         \WordArray[24].Word[30].QWire , \WordArray[24].Word[31].QWire ,
         _824_net_, \WordArray[25].Word[0].QWire ,
         \WordArray[25].Word[1].QWire , \WordArray[25].Word[2].QWire ,
         \WordArray[25].Word[3].QWire , \WordArray[25].Word[4].QWire ,
         \WordArray[25].Word[5].QWire , \WordArray[25].Word[6].QWire ,
         \WordArray[25].Word[7].QWire , \WordArray[25].Word[8].QWire ,
         \WordArray[25].Word[9].QWire , \WordArray[25].Word[10].QWire ,
         \WordArray[25].Word[11].QWire , \WordArray[25].Word[12].QWire ,
         \WordArray[25].Word[13].QWire , \WordArray[25].Word[14].QWire ,
         \WordArray[25].Word[15].QWire , \WordArray[25].Word[16].QWire ,
         \WordArray[25].Word[17].QWire , \WordArray[25].Word[18].QWire ,
         \WordArray[25].Word[19].QWire , \WordArray[25].Word[20].QWire ,
         \WordArray[25].Word[21].QWire , \WordArray[25].Word[22].QWire ,
         \WordArray[25].Word[23].QWire , \WordArray[25].Word[24].QWire ,
         \WordArray[25].Word[25].QWire , \WordArray[25].Word[26].QWire ,
         \WordArray[25].Word[27].QWire , \WordArray[25].Word[28].QWire ,
         \WordArray[25].Word[29].QWire , \WordArray[25].Word[30].QWire ,
         \WordArray[25].Word[31].QWire , _857_net_,
         \WordArray[26].Word[0].QWire , \WordArray[26].Word[1].QWire ,
         \WordArray[26].Word[2].QWire , \WordArray[26].Word[3].QWire ,
         \WordArray[26].Word[4].QWire , \WordArray[26].Word[5].QWire ,
         \WordArray[26].Word[6].QWire , \WordArray[26].Word[7].QWire ,
         \WordArray[26].Word[8].QWire , \WordArray[26].Word[9].QWire ,
         \WordArray[26].Word[10].QWire , \WordArray[26].Word[11].QWire ,
         \WordArray[26].Word[12].QWire , \WordArray[26].Word[13].QWire ,
         \WordArray[26].Word[14].QWire , \WordArray[26].Word[15].QWire ,
         \WordArray[26].Word[16].QWire , \WordArray[26].Word[17].QWire ,
         \WordArray[26].Word[18].QWire , \WordArray[26].Word[19].QWire ,
         \WordArray[26].Word[20].QWire , \WordArray[26].Word[21].QWire ,
         \WordArray[26].Word[22].QWire , \WordArray[26].Word[23].QWire ,
         \WordArray[26].Word[24].QWire , \WordArray[26].Word[25].QWire ,
         \WordArray[26].Word[26].QWire , \WordArray[26].Word[27].QWire ,
         \WordArray[26].Word[28].QWire , \WordArray[26].Word[29].QWire ,
         \WordArray[26].Word[30].QWire , \WordArray[26].Word[31].QWire ,
         _890_net_, \WordArray[27].Word[0].QWire ,
         \WordArray[27].Word[1].QWire , \WordArray[27].Word[2].QWire ,
         \WordArray[27].Word[3].QWire , \WordArray[27].Word[4].QWire ,
         \WordArray[27].Word[5].QWire , \WordArray[27].Word[6].QWire ,
         \WordArray[27].Word[7].QWire , \WordArray[27].Word[8].QWire ,
         \WordArray[27].Word[9].QWire , \WordArray[27].Word[10].QWire ,
         \WordArray[27].Word[11].QWire , \WordArray[27].Word[12].QWire ,
         \WordArray[27].Word[13].QWire , \WordArray[27].Word[14].QWire ,
         \WordArray[27].Word[15].QWire , \WordArray[27].Word[16].QWire ,
         \WordArray[27].Word[17].QWire , \WordArray[27].Word[18].QWire ,
         \WordArray[27].Word[19].QWire , \WordArray[27].Word[20].QWire ,
         \WordArray[27].Word[21].QWire , \WordArray[27].Word[22].QWire ,
         \WordArray[27].Word[23].QWire , \WordArray[27].Word[24].QWire ,
         \WordArray[27].Word[25].QWire , \WordArray[27].Word[26].QWire ,
         \WordArray[27].Word[27].QWire , \WordArray[27].Word[28].QWire ,
         \WordArray[27].Word[29].QWire , \WordArray[27].Word[30].QWire ,
         \WordArray[27].Word[31].QWire , _923_net_,
         \WordArray[28].Word[0].QWire , \WordArray[28].Word[1].QWire ,
         \WordArray[28].Word[2].QWire , \WordArray[28].Word[3].QWire ,
         \WordArray[28].Word[4].QWire , \WordArray[28].Word[5].QWire ,
         \WordArray[28].Word[6].QWire , \WordArray[28].Word[7].QWire ,
         \WordArray[28].Word[8].QWire , \WordArray[28].Word[9].QWire ,
         \WordArray[28].Word[10].QWire , \WordArray[28].Word[11].QWire ,
         \WordArray[28].Word[12].QWire , \WordArray[28].Word[13].QWire ,
         \WordArray[28].Word[14].QWire , \WordArray[28].Word[15].QWire ,
         \WordArray[28].Word[16].QWire , \WordArray[28].Word[17].QWire ,
         \WordArray[28].Word[18].QWire , \WordArray[28].Word[19].QWire ,
         \WordArray[28].Word[20].QWire , \WordArray[28].Word[21].QWire ,
         \WordArray[28].Word[22].QWire , \WordArray[28].Word[23].QWire ,
         \WordArray[28].Word[24].QWire , \WordArray[28].Word[25].QWire ,
         \WordArray[28].Word[26].QWire , \WordArray[28].Word[27].QWire ,
         \WordArray[28].Word[28].QWire , \WordArray[28].Word[29].QWire ,
         \WordArray[28].Word[30].QWire , \WordArray[28].Word[31].QWire ,
         _956_net_, \WordArray[29].Word[0].QWire ,
         \WordArray[29].Word[1].QWire , \WordArray[29].Word[2].QWire ,
         \WordArray[29].Word[3].QWire , \WordArray[29].Word[4].QWire ,
         \WordArray[29].Word[5].QWire , \WordArray[29].Word[6].QWire ,
         \WordArray[29].Word[7].QWire , \WordArray[29].Word[8].QWire ,
         \WordArray[29].Word[9].QWire , \WordArray[29].Word[10].QWire ,
         \WordArray[29].Word[11].QWire , \WordArray[29].Word[12].QWire ,
         \WordArray[29].Word[13].QWire , \WordArray[29].Word[14].QWire ,
         \WordArray[29].Word[15].QWire , \WordArray[29].Word[16].QWire ,
         \WordArray[29].Word[17].QWire , \WordArray[29].Word[18].QWire ,
         \WordArray[29].Word[19].QWire , \WordArray[29].Word[20].QWire ,
         \WordArray[29].Word[21].QWire , \WordArray[29].Word[22].QWire ,
         \WordArray[29].Word[23].QWire , \WordArray[29].Word[24].QWire ,
         \WordArray[29].Word[25].QWire , \WordArray[29].Word[26].QWire ,
         \WordArray[29].Word[27].QWire , \WordArray[29].Word[28].QWire ,
         \WordArray[29].Word[29].QWire , \WordArray[29].Word[30].QWire ,
         \WordArray[29].Word[31].QWire , _989_net_,
         \WordArray[30].Word[0].QWire , \WordArray[30].Word[1].QWire ,
         \WordArray[30].Word[2].QWire , \WordArray[30].Word[3].QWire ,
         \WordArray[30].Word[4].QWire , \WordArray[30].Word[5].QWire ,
         \WordArray[30].Word[6].QWire , \WordArray[30].Word[7].QWire ,
         \WordArray[30].Word[8].QWire , \WordArray[30].Word[9].QWire ,
         _999_net_, \WordArray[30].Word[10].QWire ,
         \WordArray[30].Word[11].QWire , \WordArray[30].Word[12].QWire ,
         \WordArray[30].Word[13].QWire , \WordArray[30].Word[14].QWire ,
         \WordArray[30].Word[15].QWire , \WordArray[30].Word[16].QWire ,
         \WordArray[30].Word[17].QWire , \WordArray[30].Word[18].QWire ,
         \WordArray[30].Word[19].QWire , \WordArray[30].Word[20].QWire ,
         \WordArray[30].Word[21].QWire , \WordArray[30].Word[22].QWire ,
         \WordArray[30].Word[23].QWire , \WordArray[30].Word[24].QWire ,
         \WordArray[30].Word[25].QWire , \WordArray[30].Word[26].QWire ,
         \WordArray[30].Word[27].QWire , \WordArray[30].Word[28].QWire ,
         \WordArray[30].Word[29].QWire , \WordArray[30].Word[30].QWire ,
         \WordArray[30].Word[31].QWire , \WordArray[31].Word[0].QWire ,
         \WordArray[31].Word[1].QWire , \WordArray[31].Word[2].QWire ,
         \WordArray[31].Word[3].QWire , \WordArray[31].Word[4].QWire ,
         \WordArray[31].Word[5].QWire , \WordArray[31].Word[6].QWire ,
         \WordArray[31].Word[7].QWire , \WordArray[31].Word[8].QWire ,
         \WordArray[31].Word[9].QWire , \WordArray[31].Word[10].QWire ,
         \WordArray[31].Word[11].QWire , \WordArray[31].Word[12].QWire ,
         \WordArray[31].Word[13].QWire , \WordArray[31].Word[14].QWire ,
         \WordArray[31].Word[15].QWire , \WordArray[31].Word[16].QWire ,
         \WordArray[31].Word[17].QWire , \WordArray[31].Word[18].QWire ,
         \WordArray[31].Word[19].QWire , \WordArray[31].Word[20].QWire ,
         \WordArray[31].Word[21].QWire , \WordArray[31].Word[22].QWire ,
         \WordArray[31].Word[23].QWire , \WordArray[31].Word[24].QWire ,
         \WordArray[31].Word[25].QWire , \WordArray[31].Word[26].QWire ,
         \WordArray[31].Word[27].QWire , \WordArray[31].Word[28].QWire ,
         \WordArray[31].Word[29].QWire , \WordArray[31].Word[30].QWire ,
         \WordArray[31].Word[31].QWire , _1055_net_, N1127, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166;
  wire   [31:0] DataRead;

  BUFTD1 \WordArray[31].Word[31].Buf  ( .I(\WordArray[31].Word[31].QWire ), 
        .OE(n36), .Z(DataRead[31]) );
  BUFTD1 \WordArray[31].Word[30].Buf  ( .I(\WordArray[31].Word[30].QWire ), 
        .OE(n36), .Z(DataRead[30]) );
  BUFTD1 \WordArray[31].Word[29].Buf  ( .I(\WordArray[31].Word[29].QWire ), 
        .OE(n36), .Z(DataRead[29]) );
  BUFTD1 \WordArray[31].Word[28].Buf  ( .I(\WordArray[31].Word[28].QWire ), 
        .OE(n35), .Z(DataRead[28]) );
  BUFTD1 \WordArray[31].Word[27].Buf  ( .I(\WordArray[31].Word[27].QWire ), 
        .OE(n36), .Z(DataRead[27]) );
  BUFTD1 \WordArray[31].Word[26].Buf  ( .I(\WordArray[31].Word[26].QWire ), 
        .OE(n35), .Z(DataRead[26]) );
  BUFTD1 \WordArray[31].Word[25].Buf  ( .I(\WordArray[31].Word[25].QWire ), 
        .OE(n36), .Z(DataRead[25]) );
  BUFTD1 \WordArray[31].Word[24].Buf  ( .I(\WordArray[31].Word[24].QWire ), 
        .OE(n36), .Z(DataRead[24]) );
  BUFTD1 \WordArray[31].Word[23].Buf  ( .I(\WordArray[31].Word[23].QWire ), 
        .OE(n36), .Z(DataRead[23]) );
  BUFTD1 \WordArray[31].Word[22].Buf  ( .I(\WordArray[31].Word[22].QWire ), 
        .OE(n35), .Z(DataRead[22]) );
  BUFTD1 \WordArray[31].Word[21].Buf  ( .I(\WordArray[31].Word[21].QWire ), 
        .OE(n36), .Z(DataRead[21]) );
  BUFTD1 \WordArray[31].Word[20].Buf  ( .I(\WordArray[31].Word[20].QWire ), 
        .OE(n36), .Z(DataRead[20]) );
  BUFTD1 \WordArray[31].Word[19].Buf  ( .I(\WordArray[31].Word[19].QWire ), 
        .OE(n35), .Z(DataRead[19]) );
  BUFTD1 \WordArray[31].Word[18].Buf  ( .I(\WordArray[31].Word[18].QWire ), 
        .OE(n35), .Z(DataRead[18]) );
  BUFTD1 \WordArray[31].Word[17].Buf  ( .I(\WordArray[31].Word[17].QWire ), 
        .OE(n35), .Z(DataRead[17]) );
  BUFTD1 \WordArray[31].Word[16].Buf  ( .I(\WordArray[31].Word[16].QWire ), 
        .OE(n35), .Z(DataRead[16]) );
  BUFTD1 \WordArray[31].Word[15].Buf  ( .I(\WordArray[31].Word[15].QWire ), 
        .OE(n35), .Z(DataRead[15]) );
  BUFTD1 \WordArray[31].Word[14].Buf  ( .I(\WordArray[31].Word[14].QWire ), 
        .OE(n35), .Z(DataRead[14]) );
  BUFTD1 \WordArray[31].Word[13].Buf  ( .I(\WordArray[31].Word[13].QWire ), 
        .OE(n35), .Z(DataRead[13]) );
  BUFTD1 \WordArray[31].Word[12].Buf  ( .I(\WordArray[31].Word[12].QWire ), 
        .OE(n35), .Z(DataRead[12]) );
  BUFTD1 \WordArray[31].Word[11].Buf  ( .I(\WordArray[31].Word[11].QWire ), 
        .OE(n35), .Z(DataRead[11]) );
  BUFTD1 \WordArray[31].Word[10].Buf  ( .I(\WordArray[31].Word[10].QWire ), 
        .OE(n35), .Z(DataRead[10]) );
  BUFTD1 \WordArray[31].Word[9].Buf  ( .I(\WordArray[31].Word[9].QWire ), .OE(
        n36), .Z(DataRead[9]) );
  BUFTD1 \WordArray[31].Word[8].Buf  ( .I(\WordArray[31].Word[8].QWire ), .OE(
        n36), .Z(DataRead[8]) );
  BUFTD1 \WordArray[31].Word[7].Buf  ( .I(\WordArray[31].Word[7].QWire ), .OE(
        n36), .Z(DataRead[7]) );
  BUFTD1 \WordArray[31].Word[6].Buf  ( .I(\WordArray[31].Word[6].QWire ), .OE(
        n36), .Z(DataRead[6]) );
  BUFTD1 \WordArray[31].Word[5].Buf  ( .I(\WordArray[31].Word[5].QWire ), .OE(
        n36), .Z(DataRead[5]) );
  BUFTD1 \WordArray[31].Word[4].Buf  ( .I(\WordArray[31].Word[4].QWire ), .OE(
        n35), .Z(DataRead[4]) );
  BUFTD1 \WordArray[31].Word[3].Buf  ( .I(\WordArray[31].Word[3].QWire ), .OE(
        n36), .Z(DataRead[3]) );
  BUFTD1 \WordArray[31].Word[2].Buf  ( .I(\WordArray[31].Word[2].QWire ), .OE(
        n35), .Z(DataRead[2]) );
  BUFTD1 \WordArray[31].Word[1].Buf  ( .I(\WordArray[31].Word[1].QWire ), .OE(
        n36), .Z(DataRead[1]) );
  BUFTD1 \WordArray[31].Word[0].Buf  ( .I(\WordArray[31].Word[0].QWire ), .OE(
        n35), .Z(DataRead[0]) );
  BUFTD1 \WordArray[30].Word[31].Buf  ( .I(\WordArray[30].Word[31].QWire ), 
        .OE(n38), .Z(DataRead[31]) );
  BUFTD1 \WordArray[30].Word[30].Buf  ( .I(\WordArray[30].Word[30].QWire ), 
        .OE(n38), .Z(DataRead[30]) );
  BUFTD1 \WordArray[30].Word[29].Buf  ( .I(\WordArray[30].Word[29].QWire ), 
        .OE(n38), .Z(DataRead[29]) );
  BUFTD1 \WordArray[30].Word[28].Buf  ( .I(\WordArray[30].Word[28].QWire ), 
        .OE(n37), .Z(DataRead[28]) );
  BUFTD1 \WordArray[30].Word[27].Buf  ( .I(\WordArray[30].Word[27].QWire ), 
        .OE(n38), .Z(DataRead[27]) );
  BUFTD1 \WordArray[30].Word[26].Buf  ( .I(\WordArray[30].Word[26].QWire ), 
        .OE(n37), .Z(DataRead[26]) );
  BUFTD1 \WordArray[30].Word[25].Buf  ( .I(\WordArray[30].Word[25].QWire ), 
        .OE(n38), .Z(DataRead[25]) );
  BUFTD1 \WordArray[30].Word[24].Buf  ( .I(\WordArray[30].Word[24].QWire ), 
        .OE(n38), .Z(DataRead[24]) );
  BUFTD1 \WordArray[30].Word[23].Buf  ( .I(\WordArray[30].Word[23].QWire ), 
        .OE(n38), .Z(DataRead[23]) );
  BUFTD1 \WordArray[30].Word[22].Buf  ( .I(\WordArray[30].Word[22].QWire ), 
        .OE(n37), .Z(DataRead[22]) );
  BUFTD1 \WordArray[30].Word[21].Buf  ( .I(\WordArray[30].Word[21].QWire ), 
        .OE(n38), .Z(DataRead[21]) );
  BUFTD1 \WordArray[30].Word[20].Buf  ( .I(\WordArray[30].Word[20].QWire ), 
        .OE(n38), .Z(DataRead[20]) );
  BUFTD1 \WordArray[30].Word[19].Buf  ( .I(\WordArray[30].Word[19].QWire ), 
        .OE(n37), .Z(DataRead[19]) );
  BUFTD1 \WordArray[30].Word[18].Buf  ( .I(\WordArray[30].Word[18].QWire ), 
        .OE(n37), .Z(DataRead[18]) );
  BUFTD1 \WordArray[30].Word[17].Buf  ( .I(\WordArray[30].Word[17].QWire ), 
        .OE(n37), .Z(DataRead[17]) );
  BUFTD1 \WordArray[30].Word[16].Buf  ( .I(\WordArray[30].Word[16].QWire ), 
        .OE(n37), .Z(DataRead[16]) );
  BUFTD1 \WordArray[30].Word[15].Buf  ( .I(\WordArray[30].Word[15].QWire ), 
        .OE(n37), .Z(DataRead[15]) );
  BUFTD1 \WordArray[30].Word[14].Buf  ( .I(\WordArray[30].Word[14].QWire ), 
        .OE(n37), .Z(DataRead[14]) );
  BUFTD1 \WordArray[30].Word[13].Buf  ( .I(\WordArray[30].Word[13].QWire ), 
        .OE(n37), .Z(DataRead[13]) );
  BUFTD1 \WordArray[30].Word[12].Buf  ( .I(\WordArray[30].Word[12].QWire ), 
        .OE(n37), .Z(DataRead[12]) );
  BUFTD1 \WordArray[30].Word[11].Buf  ( .I(\WordArray[30].Word[11].QWire ), 
        .OE(n37), .Z(DataRead[11]) );
  BUFTD1 \WordArray[30].Word[10].Buf  ( .I(\WordArray[30].Word[10].QWire ), 
        .OE(n37), .Z(DataRead[10]) );
  BUFTD1 \WordArray[30].Word[9].Buf  ( .I(\WordArray[30].Word[9].QWire ), .OE(
        n38), .Z(DataRead[9]) );
  BUFTD1 \WordArray[30].Word[8].Buf  ( .I(\WordArray[30].Word[8].QWire ), .OE(
        n38), .Z(DataRead[8]) );
  BUFTD1 \WordArray[30].Word[7].Buf  ( .I(\WordArray[30].Word[7].QWire ), .OE(
        n38), .Z(DataRead[7]) );
  BUFTD1 \WordArray[30].Word[6].Buf  ( .I(\WordArray[30].Word[6].QWire ), .OE(
        n38), .Z(DataRead[6]) );
  BUFTD1 \WordArray[30].Word[5].Buf  ( .I(\WordArray[30].Word[5].QWire ), .OE(
        n38), .Z(DataRead[5]) );
  BUFTD1 \WordArray[30].Word[4].Buf  ( .I(\WordArray[30].Word[4].QWire ), .OE(
        n37), .Z(DataRead[4]) );
  BUFTD1 \WordArray[30].Word[3].Buf  ( .I(\WordArray[30].Word[3].QWire ), .OE(
        n38), .Z(DataRead[3]) );
  BUFTD1 \WordArray[30].Word[2].Buf  ( .I(\WordArray[30].Word[2].QWire ), .OE(
        n37), .Z(DataRead[2]) );
  BUFTD1 \WordArray[30].Word[1].Buf  ( .I(\WordArray[30].Word[1].QWire ), .OE(
        n38), .Z(DataRead[1]) );
  BUFTD1 \WordArray[30].Word[0].Buf  ( .I(\WordArray[30].Word[0].QWire ), .OE(
        n37), .Z(DataRead[0]) );
  BUFTD1 \WordArray[29].Word[31].Buf  ( .I(\WordArray[29].Word[31].QWire ), 
        .OE(n40), .Z(DataRead[31]) );
  BUFTD1 \WordArray[29].Word[30].Buf  ( .I(\WordArray[29].Word[30].QWire ), 
        .OE(n40), .Z(DataRead[30]) );
  BUFTD1 \WordArray[29].Word[29].Buf  ( .I(\WordArray[29].Word[29].QWire ), 
        .OE(n40), .Z(DataRead[29]) );
  BUFTD1 \WordArray[29].Word[28].Buf  ( .I(\WordArray[29].Word[28].QWire ), 
        .OE(n39), .Z(DataRead[28]) );
  BUFTD1 \WordArray[29].Word[27].Buf  ( .I(\WordArray[29].Word[27].QWire ), 
        .OE(n40), .Z(DataRead[27]) );
  BUFTD1 \WordArray[29].Word[26].Buf  ( .I(\WordArray[29].Word[26].QWire ), 
        .OE(n39), .Z(DataRead[26]) );
  BUFTD1 \WordArray[29].Word[25].Buf  ( .I(\WordArray[29].Word[25].QWire ), 
        .OE(n40), .Z(DataRead[25]) );
  BUFTD1 \WordArray[29].Word[24].Buf  ( .I(\WordArray[29].Word[24].QWire ), 
        .OE(n40), .Z(DataRead[24]) );
  BUFTD1 \WordArray[29].Word[23].Buf  ( .I(\WordArray[29].Word[23].QWire ), 
        .OE(n40), .Z(DataRead[23]) );
  BUFTD1 \WordArray[29].Word[22].Buf  ( .I(\WordArray[29].Word[22].QWire ), 
        .OE(n39), .Z(DataRead[22]) );
  BUFTD1 \WordArray[29].Word[21].Buf  ( .I(\WordArray[29].Word[21].QWire ), 
        .OE(n40), .Z(DataRead[21]) );
  BUFTD1 \WordArray[29].Word[20].Buf  ( .I(\WordArray[29].Word[20].QWire ), 
        .OE(n40), .Z(DataRead[20]) );
  BUFTD1 \WordArray[29].Word[19].Buf  ( .I(\WordArray[29].Word[19].QWire ), 
        .OE(n39), .Z(DataRead[19]) );
  BUFTD1 \WordArray[29].Word[18].Buf  ( .I(\WordArray[29].Word[18].QWire ), 
        .OE(n39), .Z(DataRead[18]) );
  BUFTD1 \WordArray[29].Word[17].Buf  ( .I(\WordArray[29].Word[17].QWire ), 
        .OE(n39), .Z(DataRead[17]) );
  BUFTD1 \WordArray[29].Word[16].Buf  ( .I(\WordArray[29].Word[16].QWire ), 
        .OE(n39), .Z(DataRead[16]) );
  BUFTD1 \WordArray[29].Word[15].Buf  ( .I(\WordArray[29].Word[15].QWire ), 
        .OE(n39), .Z(DataRead[15]) );
  BUFTD1 \WordArray[29].Word[14].Buf  ( .I(\WordArray[29].Word[14].QWire ), 
        .OE(n39), .Z(DataRead[14]) );
  BUFTD1 \WordArray[29].Word[13].Buf  ( .I(\WordArray[29].Word[13].QWire ), 
        .OE(n39), .Z(DataRead[13]) );
  BUFTD1 \WordArray[29].Word[12].Buf  ( .I(\WordArray[29].Word[12].QWire ), 
        .OE(n39), .Z(DataRead[12]) );
  BUFTD1 \WordArray[29].Word[11].Buf  ( .I(\WordArray[29].Word[11].QWire ), 
        .OE(n39), .Z(DataRead[11]) );
  BUFTD1 \WordArray[29].Word[10].Buf  ( .I(\WordArray[29].Word[10].QWire ), 
        .OE(n39), .Z(DataRead[10]) );
  BUFTD1 \WordArray[29].Word[9].Buf  ( .I(\WordArray[29].Word[9].QWire ), .OE(
        n40), .Z(DataRead[9]) );
  BUFTD1 \WordArray[29].Word[8].Buf  ( .I(\WordArray[29].Word[8].QWire ), .OE(
        n40), .Z(DataRead[8]) );
  BUFTD1 \WordArray[29].Word[7].Buf  ( .I(\WordArray[29].Word[7].QWire ), .OE(
        n40), .Z(DataRead[7]) );
  BUFTD1 \WordArray[29].Word[6].Buf  ( .I(\WordArray[29].Word[6].QWire ), .OE(
        n40), .Z(DataRead[6]) );
  BUFTD1 \WordArray[29].Word[5].Buf  ( .I(\WordArray[29].Word[5].QWire ), .OE(
        n40), .Z(DataRead[5]) );
  BUFTD1 \WordArray[29].Word[4].Buf  ( .I(\WordArray[29].Word[4].QWire ), .OE(
        n39), .Z(DataRead[4]) );
  BUFTD1 \WordArray[29].Word[3].Buf  ( .I(\WordArray[29].Word[3].QWire ), .OE(
        n40), .Z(DataRead[3]) );
  BUFTD1 \WordArray[29].Word[2].Buf  ( .I(\WordArray[29].Word[2].QWire ), .OE(
        n39), .Z(DataRead[2]) );
  BUFTD1 \WordArray[29].Word[1].Buf  ( .I(\WordArray[29].Word[1].QWire ), .OE(
        n40), .Z(DataRead[1]) );
  BUFTD1 \WordArray[29].Word[0].Buf  ( .I(\WordArray[29].Word[0].QWire ), .OE(
        n39), .Z(DataRead[0]) );
  BUFTD1 \WordArray[28].Word[31].Buf  ( .I(\WordArray[28].Word[31].QWire ), 
        .OE(n42), .Z(DataRead[31]) );
  BUFTD1 \WordArray[28].Word[30].Buf  ( .I(\WordArray[28].Word[30].QWire ), 
        .OE(n42), .Z(DataRead[30]) );
  BUFTD1 \WordArray[28].Word[29].Buf  ( .I(\WordArray[28].Word[29].QWire ), 
        .OE(n42), .Z(DataRead[29]) );
  BUFTD1 \WordArray[28].Word[28].Buf  ( .I(\WordArray[28].Word[28].QWire ), 
        .OE(n41), .Z(DataRead[28]) );
  BUFTD1 \WordArray[28].Word[27].Buf  ( .I(\WordArray[28].Word[27].QWire ), 
        .OE(n42), .Z(DataRead[27]) );
  BUFTD1 \WordArray[28].Word[26].Buf  ( .I(\WordArray[28].Word[26].QWire ), 
        .OE(n41), .Z(DataRead[26]) );
  BUFTD1 \WordArray[28].Word[25].Buf  ( .I(\WordArray[28].Word[25].QWire ), 
        .OE(n42), .Z(DataRead[25]) );
  BUFTD1 \WordArray[28].Word[24].Buf  ( .I(\WordArray[28].Word[24].QWire ), 
        .OE(n42), .Z(DataRead[24]) );
  BUFTD1 \WordArray[28].Word[23].Buf  ( .I(\WordArray[28].Word[23].QWire ), 
        .OE(n42), .Z(DataRead[23]) );
  BUFTD1 \WordArray[28].Word[22].Buf  ( .I(\WordArray[28].Word[22].QWire ), 
        .OE(n41), .Z(DataRead[22]) );
  BUFTD1 \WordArray[28].Word[21].Buf  ( .I(\WordArray[28].Word[21].QWire ), 
        .OE(n42), .Z(DataRead[21]) );
  BUFTD1 \WordArray[28].Word[20].Buf  ( .I(\WordArray[28].Word[20].QWire ), 
        .OE(n42), .Z(DataRead[20]) );
  BUFTD1 \WordArray[28].Word[19].Buf  ( .I(\WordArray[28].Word[19].QWire ), 
        .OE(n41), .Z(DataRead[19]) );
  BUFTD1 \WordArray[28].Word[18].Buf  ( .I(\WordArray[28].Word[18].QWire ), 
        .OE(n41), .Z(DataRead[18]) );
  BUFTD1 \WordArray[28].Word[17].Buf  ( .I(\WordArray[28].Word[17].QWire ), 
        .OE(n41), .Z(DataRead[17]) );
  BUFTD1 \WordArray[28].Word[16].Buf  ( .I(\WordArray[28].Word[16].QWire ), 
        .OE(n41), .Z(DataRead[16]) );
  BUFTD1 \WordArray[28].Word[15].Buf  ( .I(\WordArray[28].Word[15].QWire ), 
        .OE(n41), .Z(DataRead[15]) );
  BUFTD1 \WordArray[28].Word[14].Buf  ( .I(\WordArray[28].Word[14].QWire ), 
        .OE(n41), .Z(DataRead[14]) );
  BUFTD1 \WordArray[28].Word[13].Buf  ( .I(\WordArray[28].Word[13].QWire ), 
        .OE(n41), .Z(DataRead[13]) );
  BUFTD1 \WordArray[28].Word[12].Buf  ( .I(\WordArray[28].Word[12].QWire ), 
        .OE(n41), .Z(DataRead[12]) );
  BUFTD1 \WordArray[28].Word[11].Buf  ( .I(\WordArray[28].Word[11].QWire ), 
        .OE(n41), .Z(DataRead[11]) );
  BUFTD1 \WordArray[28].Word[10].Buf  ( .I(\WordArray[28].Word[10].QWire ), 
        .OE(n41), .Z(DataRead[10]) );
  BUFTD1 \WordArray[28].Word[9].Buf  ( .I(\WordArray[28].Word[9].QWire ), .OE(
        n42), .Z(DataRead[9]) );
  BUFTD1 \WordArray[28].Word[8].Buf  ( .I(\WordArray[28].Word[8].QWire ), .OE(
        n42), .Z(DataRead[8]) );
  BUFTD1 \WordArray[28].Word[7].Buf  ( .I(\WordArray[28].Word[7].QWire ), .OE(
        n42), .Z(DataRead[7]) );
  BUFTD1 \WordArray[28].Word[6].Buf  ( .I(\WordArray[28].Word[6].QWire ), .OE(
        n42), .Z(DataRead[6]) );
  BUFTD1 \WordArray[28].Word[5].Buf  ( .I(\WordArray[28].Word[5].QWire ), .OE(
        n42), .Z(DataRead[5]) );
  BUFTD1 \WordArray[28].Word[4].Buf  ( .I(\WordArray[28].Word[4].QWire ), .OE(
        n41), .Z(DataRead[4]) );
  BUFTD1 \WordArray[28].Word[3].Buf  ( .I(\WordArray[28].Word[3].QWire ), .OE(
        n42), .Z(DataRead[3]) );
  BUFTD1 \WordArray[28].Word[2].Buf  ( .I(\WordArray[28].Word[2].QWire ), .OE(
        n41), .Z(DataRead[2]) );
  BUFTD1 \WordArray[28].Word[1].Buf  ( .I(\WordArray[28].Word[1].QWire ), .OE(
        n42), .Z(DataRead[1]) );
  BUFTD1 \WordArray[28].Word[0].Buf  ( .I(\WordArray[28].Word[0].QWire ), .OE(
        n41), .Z(DataRead[0]) );
  BUFTD1 \WordArray[27].Word[31].Buf  ( .I(\WordArray[27].Word[31].QWire ), 
        .OE(n44), .Z(DataRead[31]) );
  BUFTD1 \WordArray[27].Word[30].Buf  ( .I(\WordArray[27].Word[30].QWire ), 
        .OE(n44), .Z(DataRead[30]) );
  BUFTD1 \WordArray[27].Word[29].Buf  ( .I(\WordArray[27].Word[29].QWire ), 
        .OE(n44), .Z(DataRead[29]) );
  BUFTD1 \WordArray[27].Word[28].Buf  ( .I(\WordArray[27].Word[28].QWire ), 
        .OE(n43), .Z(DataRead[28]) );
  BUFTD1 \WordArray[27].Word[27].Buf  ( .I(\WordArray[27].Word[27].QWire ), 
        .OE(n44), .Z(DataRead[27]) );
  BUFTD1 \WordArray[27].Word[26].Buf  ( .I(\WordArray[27].Word[26].QWire ), 
        .OE(n43), .Z(DataRead[26]) );
  BUFTD1 \WordArray[27].Word[25].Buf  ( .I(\WordArray[27].Word[25].QWire ), 
        .OE(n44), .Z(DataRead[25]) );
  BUFTD1 \WordArray[27].Word[24].Buf  ( .I(\WordArray[27].Word[24].QWire ), 
        .OE(n44), .Z(DataRead[24]) );
  BUFTD1 \WordArray[27].Word[23].Buf  ( .I(\WordArray[27].Word[23].QWire ), 
        .OE(n44), .Z(DataRead[23]) );
  BUFTD1 \WordArray[27].Word[22].Buf  ( .I(\WordArray[27].Word[22].QWire ), 
        .OE(n43), .Z(DataRead[22]) );
  BUFTD1 \WordArray[27].Word[21].Buf  ( .I(\WordArray[27].Word[21].QWire ), 
        .OE(n44), .Z(DataRead[21]) );
  BUFTD1 \WordArray[27].Word[20].Buf  ( .I(\WordArray[27].Word[20].QWire ), 
        .OE(n44), .Z(DataRead[20]) );
  BUFTD1 \WordArray[27].Word[19].Buf  ( .I(\WordArray[27].Word[19].QWire ), 
        .OE(n43), .Z(DataRead[19]) );
  BUFTD1 \WordArray[27].Word[18].Buf  ( .I(\WordArray[27].Word[18].QWire ), 
        .OE(n43), .Z(DataRead[18]) );
  BUFTD1 \WordArray[27].Word[17].Buf  ( .I(\WordArray[27].Word[17].QWire ), 
        .OE(n43), .Z(DataRead[17]) );
  BUFTD1 \WordArray[27].Word[16].Buf  ( .I(\WordArray[27].Word[16].QWire ), 
        .OE(n43), .Z(DataRead[16]) );
  BUFTD1 \WordArray[27].Word[15].Buf  ( .I(\WordArray[27].Word[15].QWire ), 
        .OE(n43), .Z(DataRead[15]) );
  BUFTD1 \WordArray[27].Word[14].Buf  ( .I(\WordArray[27].Word[14].QWire ), 
        .OE(n43), .Z(DataRead[14]) );
  BUFTD1 \WordArray[27].Word[13].Buf  ( .I(\WordArray[27].Word[13].QWire ), 
        .OE(n43), .Z(DataRead[13]) );
  BUFTD1 \WordArray[27].Word[12].Buf  ( .I(\WordArray[27].Word[12].QWire ), 
        .OE(n43), .Z(DataRead[12]) );
  BUFTD1 \WordArray[27].Word[11].Buf  ( .I(\WordArray[27].Word[11].QWire ), 
        .OE(n43), .Z(DataRead[11]) );
  BUFTD1 \WordArray[27].Word[10].Buf  ( .I(\WordArray[27].Word[10].QWire ), 
        .OE(n43), .Z(DataRead[10]) );
  BUFTD1 \WordArray[27].Word[9].Buf  ( .I(\WordArray[27].Word[9].QWire ), .OE(
        n44), .Z(DataRead[9]) );
  BUFTD1 \WordArray[27].Word[8].Buf  ( .I(\WordArray[27].Word[8].QWire ), .OE(
        n44), .Z(DataRead[8]) );
  BUFTD1 \WordArray[27].Word[7].Buf  ( .I(\WordArray[27].Word[7].QWire ), .OE(
        n44), .Z(DataRead[7]) );
  BUFTD1 \WordArray[27].Word[6].Buf  ( .I(\WordArray[27].Word[6].QWire ), .OE(
        n44), .Z(DataRead[6]) );
  BUFTD1 \WordArray[27].Word[5].Buf  ( .I(\WordArray[27].Word[5].QWire ), .OE(
        n44), .Z(DataRead[5]) );
  BUFTD1 \WordArray[27].Word[4].Buf  ( .I(\WordArray[27].Word[4].QWire ), .OE(
        n43), .Z(DataRead[4]) );
  BUFTD1 \WordArray[27].Word[3].Buf  ( .I(\WordArray[27].Word[3].QWire ), .OE(
        n44), .Z(DataRead[3]) );
  BUFTD1 \WordArray[27].Word[2].Buf  ( .I(\WordArray[27].Word[2].QWire ), .OE(
        n43), .Z(DataRead[2]) );
  BUFTD1 \WordArray[27].Word[1].Buf  ( .I(\WordArray[27].Word[1].QWire ), .OE(
        n44), .Z(DataRead[1]) );
  BUFTD1 \WordArray[27].Word[0].Buf  ( .I(\WordArray[27].Word[0].QWire ), .OE(
        n43), .Z(DataRead[0]) );
  BUFTD1 \WordArray[26].Word[31].Buf  ( .I(\WordArray[26].Word[31].QWire ), 
        .OE(n46), .Z(DataRead[31]) );
  BUFTD1 \WordArray[26].Word[30].Buf  ( .I(\WordArray[26].Word[30].QWire ), 
        .OE(n46), .Z(DataRead[30]) );
  BUFTD1 \WordArray[26].Word[29].Buf  ( .I(\WordArray[26].Word[29].QWire ), 
        .OE(n46), .Z(DataRead[29]) );
  BUFTD1 \WordArray[26].Word[28].Buf  ( .I(\WordArray[26].Word[28].QWire ), 
        .OE(n45), .Z(DataRead[28]) );
  BUFTD1 \WordArray[26].Word[27].Buf  ( .I(\WordArray[26].Word[27].QWire ), 
        .OE(n46), .Z(DataRead[27]) );
  BUFTD1 \WordArray[26].Word[26].Buf  ( .I(\WordArray[26].Word[26].QWire ), 
        .OE(n45), .Z(DataRead[26]) );
  BUFTD1 \WordArray[26].Word[25].Buf  ( .I(\WordArray[26].Word[25].QWire ), 
        .OE(n46), .Z(DataRead[25]) );
  BUFTD1 \WordArray[26].Word[24].Buf  ( .I(\WordArray[26].Word[24].QWire ), 
        .OE(n46), .Z(DataRead[24]) );
  BUFTD1 \WordArray[26].Word[23].Buf  ( .I(\WordArray[26].Word[23].QWire ), 
        .OE(n46), .Z(DataRead[23]) );
  BUFTD1 \WordArray[26].Word[22].Buf  ( .I(\WordArray[26].Word[22].QWire ), 
        .OE(n45), .Z(DataRead[22]) );
  BUFTD1 \WordArray[26].Word[21].Buf  ( .I(\WordArray[26].Word[21].QWire ), 
        .OE(n46), .Z(DataRead[21]) );
  BUFTD1 \WordArray[26].Word[20].Buf  ( .I(\WordArray[26].Word[20].QWire ), 
        .OE(n46), .Z(DataRead[20]) );
  BUFTD1 \WordArray[26].Word[19].Buf  ( .I(\WordArray[26].Word[19].QWire ), 
        .OE(n45), .Z(DataRead[19]) );
  BUFTD1 \WordArray[26].Word[18].Buf  ( .I(\WordArray[26].Word[18].QWire ), 
        .OE(n45), .Z(DataRead[18]) );
  BUFTD1 \WordArray[26].Word[17].Buf  ( .I(\WordArray[26].Word[17].QWire ), 
        .OE(n45), .Z(DataRead[17]) );
  BUFTD1 \WordArray[26].Word[16].Buf  ( .I(\WordArray[26].Word[16].QWire ), 
        .OE(n45), .Z(DataRead[16]) );
  BUFTD1 \WordArray[26].Word[15].Buf  ( .I(\WordArray[26].Word[15].QWire ), 
        .OE(n45), .Z(DataRead[15]) );
  BUFTD1 \WordArray[26].Word[14].Buf  ( .I(\WordArray[26].Word[14].QWire ), 
        .OE(n45), .Z(DataRead[14]) );
  BUFTD1 \WordArray[26].Word[13].Buf  ( .I(\WordArray[26].Word[13].QWire ), 
        .OE(n45), .Z(DataRead[13]) );
  BUFTD1 \WordArray[26].Word[12].Buf  ( .I(\WordArray[26].Word[12].QWire ), 
        .OE(n45), .Z(DataRead[12]) );
  BUFTD1 \WordArray[26].Word[11].Buf  ( .I(\WordArray[26].Word[11].QWire ), 
        .OE(n45), .Z(DataRead[11]) );
  BUFTD1 \WordArray[26].Word[10].Buf  ( .I(\WordArray[26].Word[10].QWire ), 
        .OE(n45), .Z(DataRead[10]) );
  BUFTD1 \WordArray[26].Word[9].Buf  ( .I(\WordArray[26].Word[9].QWire ), .OE(
        n46), .Z(DataRead[9]) );
  BUFTD1 \WordArray[26].Word[8].Buf  ( .I(\WordArray[26].Word[8].QWire ), .OE(
        n46), .Z(DataRead[8]) );
  BUFTD1 \WordArray[26].Word[7].Buf  ( .I(\WordArray[26].Word[7].QWire ), .OE(
        n46), .Z(DataRead[7]) );
  BUFTD1 \WordArray[26].Word[6].Buf  ( .I(\WordArray[26].Word[6].QWire ), .OE(
        n46), .Z(DataRead[6]) );
  BUFTD1 \WordArray[26].Word[5].Buf  ( .I(\WordArray[26].Word[5].QWire ), .OE(
        n46), .Z(DataRead[5]) );
  BUFTD1 \WordArray[26].Word[4].Buf  ( .I(\WordArray[26].Word[4].QWire ), .OE(
        n45), .Z(DataRead[4]) );
  BUFTD1 \WordArray[26].Word[3].Buf  ( .I(\WordArray[26].Word[3].QWire ), .OE(
        n46), .Z(DataRead[3]) );
  BUFTD1 \WordArray[26].Word[2].Buf  ( .I(\WordArray[26].Word[2].QWire ), .OE(
        n45), .Z(DataRead[2]) );
  BUFTD1 \WordArray[26].Word[1].Buf  ( .I(\WordArray[26].Word[1].QWire ), .OE(
        n46), .Z(DataRead[1]) );
  BUFTD1 \WordArray[26].Word[0].Buf  ( .I(\WordArray[26].Word[0].QWire ), .OE(
        n45), .Z(DataRead[0]) );
  BUFTD1 \WordArray[25].Word[31].Buf  ( .I(\WordArray[25].Word[31].QWire ), 
        .OE(n48), .Z(DataRead[31]) );
  BUFTD1 \WordArray[25].Word[30].Buf  ( .I(\WordArray[25].Word[30].QWire ), 
        .OE(n48), .Z(DataRead[30]) );
  BUFTD1 \WordArray[25].Word[29].Buf  ( .I(\WordArray[25].Word[29].QWire ), 
        .OE(n48), .Z(DataRead[29]) );
  BUFTD1 \WordArray[25].Word[28].Buf  ( .I(\WordArray[25].Word[28].QWire ), 
        .OE(n47), .Z(DataRead[28]) );
  BUFTD1 \WordArray[25].Word[27].Buf  ( .I(\WordArray[25].Word[27].QWire ), 
        .OE(n48), .Z(DataRead[27]) );
  BUFTD1 \WordArray[25].Word[26].Buf  ( .I(\WordArray[25].Word[26].QWire ), 
        .OE(n47), .Z(DataRead[26]) );
  BUFTD1 \WordArray[25].Word[25].Buf  ( .I(\WordArray[25].Word[25].QWire ), 
        .OE(n48), .Z(DataRead[25]) );
  BUFTD1 \WordArray[25].Word[24].Buf  ( .I(\WordArray[25].Word[24].QWire ), 
        .OE(n48), .Z(DataRead[24]) );
  BUFTD1 \WordArray[25].Word[23].Buf  ( .I(\WordArray[25].Word[23].QWire ), 
        .OE(n48), .Z(DataRead[23]) );
  BUFTD1 \WordArray[25].Word[22].Buf  ( .I(\WordArray[25].Word[22].QWire ), 
        .OE(n47), .Z(DataRead[22]) );
  BUFTD1 \WordArray[25].Word[21].Buf  ( .I(\WordArray[25].Word[21].QWire ), 
        .OE(n48), .Z(DataRead[21]) );
  BUFTD1 \WordArray[25].Word[20].Buf  ( .I(\WordArray[25].Word[20].QWire ), 
        .OE(n48), .Z(DataRead[20]) );
  BUFTD1 \WordArray[25].Word[19].Buf  ( .I(\WordArray[25].Word[19].QWire ), 
        .OE(n47), .Z(DataRead[19]) );
  BUFTD1 \WordArray[25].Word[18].Buf  ( .I(\WordArray[25].Word[18].QWire ), 
        .OE(n47), .Z(DataRead[18]) );
  BUFTD1 \WordArray[25].Word[17].Buf  ( .I(\WordArray[25].Word[17].QWire ), 
        .OE(n47), .Z(DataRead[17]) );
  BUFTD1 \WordArray[25].Word[16].Buf  ( .I(\WordArray[25].Word[16].QWire ), 
        .OE(n47), .Z(DataRead[16]) );
  BUFTD1 \WordArray[25].Word[15].Buf  ( .I(\WordArray[25].Word[15].QWire ), 
        .OE(n47), .Z(DataRead[15]) );
  BUFTD1 \WordArray[25].Word[14].Buf  ( .I(\WordArray[25].Word[14].QWire ), 
        .OE(n47), .Z(DataRead[14]) );
  BUFTD1 \WordArray[25].Word[13].Buf  ( .I(\WordArray[25].Word[13].QWire ), 
        .OE(n47), .Z(DataRead[13]) );
  BUFTD1 \WordArray[25].Word[12].Buf  ( .I(\WordArray[25].Word[12].QWire ), 
        .OE(n47), .Z(DataRead[12]) );
  BUFTD1 \WordArray[25].Word[11].Buf  ( .I(\WordArray[25].Word[11].QWire ), 
        .OE(n47), .Z(DataRead[11]) );
  BUFTD1 \WordArray[25].Word[10].Buf  ( .I(\WordArray[25].Word[10].QWire ), 
        .OE(n47), .Z(DataRead[10]) );
  BUFTD1 \WordArray[25].Word[9].Buf  ( .I(\WordArray[25].Word[9].QWire ), .OE(
        n48), .Z(DataRead[9]) );
  BUFTD1 \WordArray[25].Word[8].Buf  ( .I(\WordArray[25].Word[8].QWire ), .OE(
        n48), .Z(DataRead[8]) );
  BUFTD1 \WordArray[25].Word[7].Buf  ( .I(\WordArray[25].Word[7].QWire ), .OE(
        n48), .Z(DataRead[7]) );
  BUFTD1 \WordArray[25].Word[6].Buf  ( .I(\WordArray[25].Word[6].QWire ), .OE(
        n48), .Z(DataRead[6]) );
  BUFTD1 \WordArray[25].Word[5].Buf  ( .I(\WordArray[25].Word[5].QWire ), .OE(
        n48), .Z(DataRead[5]) );
  BUFTD1 \WordArray[25].Word[4].Buf  ( .I(\WordArray[25].Word[4].QWire ), .OE(
        n47), .Z(DataRead[4]) );
  BUFTD1 \WordArray[25].Word[3].Buf  ( .I(\WordArray[25].Word[3].QWire ), .OE(
        n48), .Z(DataRead[3]) );
  BUFTD1 \WordArray[25].Word[2].Buf  ( .I(\WordArray[25].Word[2].QWire ), .OE(
        n47), .Z(DataRead[2]) );
  BUFTD1 \WordArray[25].Word[1].Buf  ( .I(\WordArray[25].Word[1].QWire ), .OE(
        n48), .Z(DataRead[1]) );
  BUFTD1 \WordArray[25].Word[0].Buf  ( .I(\WordArray[25].Word[0].QWire ), .OE(
        n47), .Z(DataRead[0]) );
  BUFTD1 \WordArray[24].Word[31].Buf  ( .I(\WordArray[24].Word[31].QWire ), 
        .OE(n50), .Z(DataRead[31]) );
  BUFTD1 \WordArray[24].Word[30].Buf  ( .I(\WordArray[24].Word[30].QWire ), 
        .OE(n50), .Z(DataRead[30]) );
  BUFTD1 \WordArray[24].Word[29].Buf  ( .I(\WordArray[24].Word[29].QWire ), 
        .OE(n50), .Z(DataRead[29]) );
  BUFTD1 \WordArray[24].Word[28].Buf  ( .I(\WordArray[24].Word[28].QWire ), 
        .OE(n49), .Z(DataRead[28]) );
  BUFTD1 \WordArray[24].Word[27].Buf  ( .I(\WordArray[24].Word[27].QWire ), 
        .OE(n50), .Z(DataRead[27]) );
  BUFTD1 \WordArray[24].Word[26].Buf  ( .I(\WordArray[24].Word[26].QWire ), 
        .OE(n49), .Z(DataRead[26]) );
  BUFTD1 \WordArray[24].Word[25].Buf  ( .I(\WordArray[24].Word[25].QWire ), 
        .OE(n50), .Z(DataRead[25]) );
  BUFTD1 \WordArray[24].Word[24].Buf  ( .I(\WordArray[24].Word[24].QWire ), 
        .OE(n50), .Z(DataRead[24]) );
  BUFTD1 \WordArray[24].Word[23].Buf  ( .I(\WordArray[24].Word[23].QWire ), 
        .OE(n50), .Z(DataRead[23]) );
  BUFTD1 \WordArray[24].Word[22].Buf  ( .I(\WordArray[24].Word[22].QWire ), 
        .OE(n49), .Z(DataRead[22]) );
  BUFTD1 \WordArray[24].Word[21].Buf  ( .I(\WordArray[24].Word[21].QWire ), 
        .OE(n50), .Z(DataRead[21]) );
  BUFTD1 \WordArray[24].Word[20].Buf  ( .I(\WordArray[24].Word[20].QWire ), 
        .OE(n50), .Z(DataRead[20]) );
  BUFTD1 \WordArray[24].Word[19].Buf  ( .I(\WordArray[24].Word[19].QWire ), 
        .OE(n49), .Z(DataRead[19]) );
  BUFTD1 \WordArray[24].Word[18].Buf  ( .I(\WordArray[24].Word[18].QWire ), 
        .OE(n49), .Z(DataRead[18]) );
  BUFTD1 \WordArray[24].Word[17].Buf  ( .I(\WordArray[24].Word[17].QWire ), 
        .OE(n49), .Z(DataRead[17]) );
  BUFTD1 \WordArray[24].Word[16].Buf  ( .I(\WordArray[24].Word[16].QWire ), 
        .OE(n49), .Z(DataRead[16]) );
  BUFTD1 \WordArray[24].Word[15].Buf  ( .I(\WordArray[24].Word[15].QWire ), 
        .OE(n49), .Z(DataRead[15]) );
  BUFTD1 \WordArray[24].Word[14].Buf  ( .I(\WordArray[24].Word[14].QWire ), 
        .OE(n49), .Z(DataRead[14]) );
  BUFTD1 \WordArray[24].Word[13].Buf  ( .I(\WordArray[24].Word[13].QWire ), 
        .OE(n49), .Z(DataRead[13]) );
  BUFTD1 \WordArray[24].Word[12].Buf  ( .I(\WordArray[24].Word[12].QWire ), 
        .OE(n49), .Z(DataRead[12]) );
  BUFTD1 \WordArray[24].Word[11].Buf  ( .I(\WordArray[24].Word[11].QWire ), 
        .OE(n49), .Z(DataRead[11]) );
  BUFTD1 \WordArray[24].Word[10].Buf  ( .I(\WordArray[24].Word[10].QWire ), 
        .OE(n49), .Z(DataRead[10]) );
  BUFTD1 \WordArray[24].Word[9].Buf  ( .I(\WordArray[24].Word[9].QWire ), .OE(
        n50), .Z(DataRead[9]) );
  BUFTD1 \WordArray[24].Word[8].Buf  ( .I(\WordArray[24].Word[8].QWire ), .OE(
        n50), .Z(DataRead[8]) );
  BUFTD1 \WordArray[24].Word[7].Buf  ( .I(\WordArray[24].Word[7].QWire ), .OE(
        n50), .Z(DataRead[7]) );
  BUFTD1 \WordArray[24].Word[6].Buf  ( .I(\WordArray[24].Word[6].QWire ), .OE(
        n50), .Z(DataRead[6]) );
  BUFTD1 \WordArray[24].Word[5].Buf  ( .I(\WordArray[24].Word[5].QWire ), .OE(
        n50), .Z(DataRead[5]) );
  BUFTD1 \WordArray[24].Word[4].Buf  ( .I(\WordArray[24].Word[4].QWire ), .OE(
        n49), .Z(DataRead[4]) );
  BUFTD1 \WordArray[24].Word[3].Buf  ( .I(\WordArray[24].Word[3].QWire ), .OE(
        n50), .Z(DataRead[3]) );
  BUFTD1 \WordArray[24].Word[2].Buf  ( .I(\WordArray[24].Word[2].QWire ), .OE(
        n49), .Z(DataRead[2]) );
  BUFTD1 \WordArray[24].Word[1].Buf  ( .I(\WordArray[24].Word[1].QWire ), .OE(
        n50), .Z(DataRead[1]) );
  BUFTD1 \WordArray[24].Word[0].Buf  ( .I(\WordArray[24].Word[0].QWire ), .OE(
        n49), .Z(DataRead[0]) );
  BUFTD1 \WordArray[23].Word[31].Buf  ( .I(\WordArray[23].Word[31].QWire ), 
        .OE(n52), .Z(DataRead[31]) );
  BUFTD1 \WordArray[23].Word[30].Buf  ( .I(\WordArray[23].Word[30].QWire ), 
        .OE(n52), .Z(DataRead[30]) );
  BUFTD1 \WordArray[23].Word[29].Buf  ( .I(\WordArray[23].Word[29].QWire ), 
        .OE(n52), .Z(DataRead[29]) );
  BUFTD1 \WordArray[23].Word[28].Buf  ( .I(\WordArray[23].Word[28].QWire ), 
        .OE(n51), .Z(DataRead[28]) );
  BUFTD1 \WordArray[23].Word[27].Buf  ( .I(\WordArray[23].Word[27].QWire ), 
        .OE(n52), .Z(DataRead[27]) );
  BUFTD1 \WordArray[23].Word[26].Buf  ( .I(\WordArray[23].Word[26].QWire ), 
        .OE(n51), .Z(DataRead[26]) );
  BUFTD1 \WordArray[23].Word[25].Buf  ( .I(\WordArray[23].Word[25].QWire ), 
        .OE(n52), .Z(DataRead[25]) );
  BUFTD1 \WordArray[23].Word[24].Buf  ( .I(\WordArray[23].Word[24].QWire ), 
        .OE(n52), .Z(DataRead[24]) );
  BUFTD1 \WordArray[23].Word[23].Buf  ( .I(\WordArray[23].Word[23].QWire ), 
        .OE(n52), .Z(DataRead[23]) );
  BUFTD1 \WordArray[23].Word[22].Buf  ( .I(\WordArray[23].Word[22].QWire ), 
        .OE(n51), .Z(DataRead[22]) );
  BUFTD1 \WordArray[23].Word[21].Buf  ( .I(\WordArray[23].Word[21].QWire ), 
        .OE(n52), .Z(DataRead[21]) );
  BUFTD1 \WordArray[23].Word[20].Buf  ( .I(\WordArray[23].Word[20].QWire ), 
        .OE(n52), .Z(DataRead[20]) );
  BUFTD1 \WordArray[23].Word[19].Buf  ( .I(\WordArray[23].Word[19].QWire ), 
        .OE(n51), .Z(DataRead[19]) );
  BUFTD1 \WordArray[23].Word[18].Buf  ( .I(\WordArray[23].Word[18].QWire ), 
        .OE(n51), .Z(DataRead[18]) );
  BUFTD1 \WordArray[23].Word[17].Buf  ( .I(\WordArray[23].Word[17].QWire ), 
        .OE(n51), .Z(DataRead[17]) );
  BUFTD1 \WordArray[23].Word[16].Buf  ( .I(\WordArray[23].Word[16].QWire ), 
        .OE(n51), .Z(DataRead[16]) );
  BUFTD1 \WordArray[23].Word[15].Buf  ( .I(\WordArray[23].Word[15].QWire ), 
        .OE(n51), .Z(DataRead[15]) );
  BUFTD1 \WordArray[23].Word[14].Buf  ( .I(\WordArray[23].Word[14].QWire ), 
        .OE(n51), .Z(DataRead[14]) );
  BUFTD1 \WordArray[23].Word[13].Buf  ( .I(\WordArray[23].Word[13].QWire ), 
        .OE(n51), .Z(DataRead[13]) );
  BUFTD1 \WordArray[23].Word[12].Buf  ( .I(\WordArray[23].Word[12].QWire ), 
        .OE(n51), .Z(DataRead[12]) );
  BUFTD1 \WordArray[23].Word[11].Buf  ( .I(\WordArray[23].Word[11].QWire ), 
        .OE(n51), .Z(DataRead[11]) );
  BUFTD1 \WordArray[23].Word[10].Buf  ( .I(\WordArray[23].Word[10].QWire ), 
        .OE(n51), .Z(DataRead[10]) );
  BUFTD1 \WordArray[23].Word[9].Buf  ( .I(\WordArray[23].Word[9].QWire ), .OE(
        n52), .Z(DataRead[9]) );
  BUFTD1 \WordArray[23].Word[8].Buf  ( .I(\WordArray[23].Word[8].QWire ), .OE(
        n52), .Z(DataRead[8]) );
  BUFTD1 \WordArray[23].Word[7].Buf  ( .I(\WordArray[23].Word[7].QWire ), .OE(
        n52), .Z(DataRead[7]) );
  BUFTD1 \WordArray[23].Word[6].Buf  ( .I(\WordArray[23].Word[6].QWire ), .OE(
        n52), .Z(DataRead[6]) );
  BUFTD1 \WordArray[23].Word[5].Buf  ( .I(\WordArray[23].Word[5].QWire ), .OE(
        n52), .Z(DataRead[5]) );
  BUFTD1 \WordArray[23].Word[4].Buf  ( .I(\WordArray[23].Word[4].QWire ), .OE(
        n51), .Z(DataRead[4]) );
  BUFTD1 \WordArray[23].Word[3].Buf  ( .I(\WordArray[23].Word[3].QWire ), .OE(
        n52), .Z(DataRead[3]) );
  BUFTD1 \WordArray[23].Word[2].Buf  ( .I(\WordArray[23].Word[2].QWire ), .OE(
        n51), .Z(DataRead[2]) );
  BUFTD1 \WordArray[23].Word[1].Buf  ( .I(\WordArray[23].Word[1].QWire ), .OE(
        n52), .Z(DataRead[1]) );
  BUFTD1 \WordArray[23].Word[0].Buf  ( .I(\WordArray[23].Word[0].QWire ), .OE(
        n51), .Z(DataRead[0]) );
  BUFTD1 \WordArray[22].Word[31].Buf  ( .I(\WordArray[22].Word[31].QWire ), 
        .OE(n54), .Z(DataRead[31]) );
  BUFTD1 \WordArray[22].Word[30].Buf  ( .I(\WordArray[22].Word[30].QWire ), 
        .OE(n54), .Z(DataRead[30]) );
  BUFTD1 \WordArray[22].Word[29].Buf  ( .I(\WordArray[22].Word[29].QWire ), 
        .OE(n54), .Z(DataRead[29]) );
  BUFTD1 \WordArray[22].Word[28].Buf  ( .I(\WordArray[22].Word[28].QWire ), 
        .OE(n53), .Z(DataRead[28]) );
  BUFTD1 \WordArray[22].Word[27].Buf  ( .I(\WordArray[22].Word[27].QWire ), 
        .OE(n54), .Z(DataRead[27]) );
  BUFTD1 \WordArray[22].Word[26].Buf  ( .I(\WordArray[22].Word[26].QWire ), 
        .OE(n53), .Z(DataRead[26]) );
  BUFTD1 \WordArray[22].Word[25].Buf  ( .I(\WordArray[22].Word[25].QWire ), 
        .OE(n54), .Z(DataRead[25]) );
  BUFTD1 \WordArray[22].Word[24].Buf  ( .I(\WordArray[22].Word[24].QWire ), 
        .OE(n54), .Z(DataRead[24]) );
  BUFTD1 \WordArray[22].Word[23].Buf  ( .I(\WordArray[22].Word[23].QWire ), 
        .OE(n54), .Z(DataRead[23]) );
  BUFTD1 \WordArray[22].Word[22].Buf  ( .I(\WordArray[22].Word[22].QWire ), 
        .OE(n53), .Z(DataRead[22]) );
  BUFTD1 \WordArray[22].Word[21].Buf  ( .I(\WordArray[22].Word[21].QWire ), 
        .OE(n54), .Z(DataRead[21]) );
  BUFTD1 \WordArray[22].Word[20].Buf  ( .I(\WordArray[22].Word[20].QWire ), 
        .OE(n54), .Z(DataRead[20]) );
  BUFTD1 \WordArray[22].Word[19].Buf  ( .I(\WordArray[22].Word[19].QWire ), 
        .OE(n53), .Z(DataRead[19]) );
  BUFTD1 \WordArray[22].Word[18].Buf  ( .I(\WordArray[22].Word[18].QWire ), 
        .OE(n53), .Z(DataRead[18]) );
  BUFTD1 \WordArray[22].Word[17].Buf  ( .I(\WordArray[22].Word[17].QWire ), 
        .OE(n53), .Z(DataRead[17]) );
  BUFTD1 \WordArray[22].Word[16].Buf  ( .I(\WordArray[22].Word[16].QWire ), 
        .OE(n53), .Z(DataRead[16]) );
  BUFTD1 \WordArray[22].Word[15].Buf  ( .I(\WordArray[22].Word[15].QWire ), 
        .OE(n53), .Z(DataRead[15]) );
  BUFTD1 \WordArray[22].Word[14].Buf  ( .I(\WordArray[22].Word[14].QWire ), 
        .OE(n53), .Z(DataRead[14]) );
  BUFTD1 \WordArray[22].Word[13].Buf  ( .I(\WordArray[22].Word[13].QWire ), 
        .OE(n53), .Z(DataRead[13]) );
  BUFTD1 \WordArray[22].Word[12].Buf  ( .I(\WordArray[22].Word[12].QWire ), 
        .OE(n53), .Z(DataRead[12]) );
  BUFTD1 \WordArray[22].Word[11].Buf  ( .I(\WordArray[22].Word[11].QWire ), 
        .OE(n53), .Z(DataRead[11]) );
  BUFTD1 \WordArray[22].Word[10].Buf  ( .I(\WordArray[22].Word[10].QWire ), 
        .OE(n53), .Z(DataRead[10]) );
  BUFTD1 \WordArray[22].Word[9].Buf  ( .I(\WordArray[22].Word[9].QWire ), .OE(
        n54), .Z(DataRead[9]) );
  BUFTD1 \WordArray[22].Word[8].Buf  ( .I(\WordArray[22].Word[8].QWire ), .OE(
        n54), .Z(DataRead[8]) );
  BUFTD1 \WordArray[22].Word[7].Buf  ( .I(\WordArray[22].Word[7].QWire ), .OE(
        n54), .Z(DataRead[7]) );
  BUFTD1 \WordArray[22].Word[6].Buf  ( .I(\WordArray[22].Word[6].QWire ), .OE(
        n54), .Z(DataRead[6]) );
  BUFTD1 \WordArray[22].Word[5].Buf  ( .I(\WordArray[22].Word[5].QWire ), .OE(
        n54), .Z(DataRead[5]) );
  BUFTD1 \WordArray[22].Word[4].Buf  ( .I(\WordArray[22].Word[4].QWire ), .OE(
        n53), .Z(DataRead[4]) );
  BUFTD1 \WordArray[22].Word[3].Buf  ( .I(\WordArray[22].Word[3].QWire ), .OE(
        n54), .Z(DataRead[3]) );
  BUFTD1 \WordArray[22].Word[2].Buf  ( .I(\WordArray[22].Word[2].QWire ), .OE(
        n53), .Z(DataRead[2]) );
  BUFTD1 \WordArray[22].Word[1].Buf  ( .I(\WordArray[22].Word[1].QWire ), .OE(
        n54), .Z(DataRead[1]) );
  BUFTD1 \WordArray[22].Word[0].Buf  ( .I(\WordArray[22].Word[0].QWire ), .OE(
        n53), .Z(DataRead[0]) );
  BUFTD1 \WordArray[21].Word[31].Buf  ( .I(\WordArray[21].Word[31].QWire ), 
        .OE(n56), .Z(DataRead[31]) );
  BUFTD1 \WordArray[21].Word[30].Buf  ( .I(\WordArray[21].Word[30].QWire ), 
        .OE(n56), .Z(DataRead[30]) );
  BUFTD1 \WordArray[21].Word[29].Buf  ( .I(\WordArray[21].Word[29].QWire ), 
        .OE(n56), .Z(DataRead[29]) );
  BUFTD1 \WordArray[21].Word[28].Buf  ( .I(\WordArray[21].Word[28].QWire ), 
        .OE(n55), .Z(DataRead[28]) );
  BUFTD1 \WordArray[21].Word[27].Buf  ( .I(\WordArray[21].Word[27].QWire ), 
        .OE(n56), .Z(DataRead[27]) );
  BUFTD1 \WordArray[21].Word[26].Buf  ( .I(\WordArray[21].Word[26].QWire ), 
        .OE(n55), .Z(DataRead[26]) );
  BUFTD1 \WordArray[21].Word[25].Buf  ( .I(\WordArray[21].Word[25].QWire ), 
        .OE(n56), .Z(DataRead[25]) );
  BUFTD1 \WordArray[21].Word[24].Buf  ( .I(\WordArray[21].Word[24].QWire ), 
        .OE(n56), .Z(DataRead[24]) );
  BUFTD1 \WordArray[21].Word[23].Buf  ( .I(\WordArray[21].Word[23].QWire ), 
        .OE(n56), .Z(DataRead[23]) );
  BUFTD1 \WordArray[21].Word[22].Buf  ( .I(\WordArray[21].Word[22].QWire ), 
        .OE(n55), .Z(DataRead[22]) );
  BUFTD1 \WordArray[21].Word[21].Buf  ( .I(\WordArray[21].Word[21].QWire ), 
        .OE(n56), .Z(DataRead[21]) );
  BUFTD1 \WordArray[21].Word[20].Buf  ( .I(\WordArray[21].Word[20].QWire ), 
        .OE(n56), .Z(DataRead[20]) );
  BUFTD1 \WordArray[21].Word[19].Buf  ( .I(\WordArray[21].Word[19].QWire ), 
        .OE(n55), .Z(DataRead[19]) );
  BUFTD1 \WordArray[21].Word[18].Buf  ( .I(\WordArray[21].Word[18].QWire ), 
        .OE(n55), .Z(DataRead[18]) );
  BUFTD1 \WordArray[21].Word[17].Buf  ( .I(\WordArray[21].Word[17].QWire ), 
        .OE(n55), .Z(DataRead[17]) );
  BUFTD1 \WordArray[21].Word[16].Buf  ( .I(\WordArray[21].Word[16].QWire ), 
        .OE(n55), .Z(DataRead[16]) );
  BUFTD1 \WordArray[21].Word[15].Buf  ( .I(\WordArray[21].Word[15].QWire ), 
        .OE(n55), .Z(DataRead[15]) );
  BUFTD1 \WordArray[21].Word[14].Buf  ( .I(\WordArray[21].Word[14].QWire ), 
        .OE(n55), .Z(DataRead[14]) );
  BUFTD1 \WordArray[21].Word[13].Buf  ( .I(\WordArray[21].Word[13].QWire ), 
        .OE(n55), .Z(DataRead[13]) );
  BUFTD1 \WordArray[21].Word[12].Buf  ( .I(\WordArray[21].Word[12].QWire ), 
        .OE(n55), .Z(DataRead[12]) );
  BUFTD1 \WordArray[21].Word[11].Buf  ( .I(\WordArray[21].Word[11].QWire ), 
        .OE(n55), .Z(DataRead[11]) );
  BUFTD1 \WordArray[21].Word[10].Buf  ( .I(\WordArray[21].Word[10].QWire ), 
        .OE(n55), .Z(DataRead[10]) );
  BUFTD1 \WordArray[21].Word[9].Buf  ( .I(\WordArray[21].Word[9].QWire ), .OE(
        n56), .Z(DataRead[9]) );
  BUFTD1 \WordArray[21].Word[8].Buf  ( .I(\WordArray[21].Word[8].QWire ), .OE(
        n56), .Z(DataRead[8]) );
  BUFTD1 \WordArray[21].Word[7].Buf  ( .I(\WordArray[21].Word[7].QWire ), .OE(
        n56), .Z(DataRead[7]) );
  BUFTD1 \WordArray[21].Word[6].Buf  ( .I(\WordArray[21].Word[6].QWire ), .OE(
        n56), .Z(DataRead[6]) );
  BUFTD1 \WordArray[21].Word[5].Buf  ( .I(\WordArray[21].Word[5].QWire ), .OE(
        n56), .Z(DataRead[5]) );
  BUFTD1 \WordArray[21].Word[4].Buf  ( .I(\WordArray[21].Word[4].QWire ), .OE(
        n55), .Z(DataRead[4]) );
  BUFTD1 \WordArray[21].Word[3].Buf  ( .I(\WordArray[21].Word[3].QWire ), .OE(
        n56), .Z(DataRead[3]) );
  BUFTD1 \WordArray[21].Word[2].Buf  ( .I(\WordArray[21].Word[2].QWire ), .OE(
        n55), .Z(DataRead[2]) );
  BUFTD1 \WordArray[21].Word[1].Buf  ( .I(\WordArray[21].Word[1].QWire ), .OE(
        n56), .Z(DataRead[1]) );
  BUFTD1 \WordArray[21].Word[0].Buf  ( .I(\WordArray[21].Word[0].QWire ), .OE(
        n55), .Z(DataRead[0]) );
  BUFTD1 \WordArray[20].Word[31].Buf  ( .I(\WordArray[20].Word[31].QWire ), 
        .OE(n58), .Z(DataRead[31]) );
  BUFTD1 \WordArray[20].Word[30].Buf  ( .I(\WordArray[20].Word[30].QWire ), 
        .OE(n58), .Z(DataRead[30]) );
  BUFTD1 \WordArray[20].Word[29].Buf  ( .I(\WordArray[20].Word[29].QWire ), 
        .OE(n58), .Z(DataRead[29]) );
  BUFTD1 \WordArray[20].Word[28].Buf  ( .I(\WordArray[20].Word[28].QWire ), 
        .OE(n57), .Z(DataRead[28]) );
  BUFTD1 \WordArray[20].Word[27].Buf  ( .I(\WordArray[20].Word[27].QWire ), 
        .OE(n58), .Z(DataRead[27]) );
  BUFTD1 \WordArray[20].Word[26].Buf  ( .I(\WordArray[20].Word[26].QWire ), 
        .OE(n57), .Z(DataRead[26]) );
  BUFTD1 \WordArray[20].Word[25].Buf  ( .I(\WordArray[20].Word[25].QWire ), 
        .OE(n58), .Z(DataRead[25]) );
  BUFTD1 \WordArray[20].Word[24].Buf  ( .I(\WordArray[20].Word[24].QWire ), 
        .OE(n58), .Z(DataRead[24]) );
  BUFTD1 \WordArray[20].Word[23].Buf  ( .I(\WordArray[20].Word[23].QWire ), 
        .OE(n58), .Z(DataRead[23]) );
  BUFTD1 \WordArray[20].Word[22].Buf  ( .I(\WordArray[20].Word[22].QWire ), 
        .OE(n57), .Z(DataRead[22]) );
  BUFTD1 \WordArray[20].Word[21].Buf  ( .I(\WordArray[20].Word[21].QWire ), 
        .OE(n58), .Z(DataRead[21]) );
  BUFTD1 \WordArray[20].Word[20].Buf  ( .I(\WordArray[20].Word[20].QWire ), 
        .OE(n58), .Z(DataRead[20]) );
  BUFTD1 \WordArray[20].Word[19].Buf  ( .I(\WordArray[20].Word[19].QWire ), 
        .OE(n57), .Z(DataRead[19]) );
  BUFTD1 \WordArray[20].Word[18].Buf  ( .I(\WordArray[20].Word[18].QWire ), 
        .OE(n57), .Z(DataRead[18]) );
  BUFTD1 \WordArray[20].Word[17].Buf  ( .I(\WordArray[20].Word[17].QWire ), 
        .OE(n57), .Z(DataRead[17]) );
  BUFTD1 \WordArray[20].Word[16].Buf  ( .I(\WordArray[20].Word[16].QWire ), 
        .OE(n57), .Z(DataRead[16]) );
  BUFTD1 \WordArray[20].Word[15].Buf  ( .I(\WordArray[20].Word[15].QWire ), 
        .OE(n57), .Z(DataRead[15]) );
  BUFTD1 \WordArray[20].Word[14].Buf  ( .I(\WordArray[20].Word[14].QWire ), 
        .OE(n57), .Z(DataRead[14]) );
  BUFTD1 \WordArray[20].Word[13].Buf  ( .I(\WordArray[20].Word[13].QWire ), 
        .OE(n57), .Z(DataRead[13]) );
  BUFTD1 \WordArray[20].Word[12].Buf  ( .I(\WordArray[20].Word[12].QWire ), 
        .OE(n57), .Z(DataRead[12]) );
  BUFTD1 \WordArray[20].Word[11].Buf  ( .I(\WordArray[20].Word[11].QWire ), 
        .OE(n57), .Z(DataRead[11]) );
  BUFTD1 \WordArray[20].Word[10].Buf  ( .I(\WordArray[20].Word[10].QWire ), 
        .OE(n57), .Z(DataRead[10]) );
  BUFTD1 \WordArray[20].Word[9].Buf  ( .I(\WordArray[20].Word[9].QWire ), .OE(
        n58), .Z(DataRead[9]) );
  BUFTD1 \WordArray[20].Word[8].Buf  ( .I(\WordArray[20].Word[8].QWire ), .OE(
        n58), .Z(DataRead[8]) );
  BUFTD1 \WordArray[20].Word[7].Buf  ( .I(\WordArray[20].Word[7].QWire ), .OE(
        n58), .Z(DataRead[7]) );
  BUFTD1 \WordArray[20].Word[6].Buf  ( .I(\WordArray[20].Word[6].QWire ), .OE(
        n58), .Z(DataRead[6]) );
  BUFTD1 \WordArray[20].Word[5].Buf  ( .I(\WordArray[20].Word[5].QWire ), .OE(
        n58), .Z(DataRead[5]) );
  BUFTD1 \WordArray[20].Word[4].Buf  ( .I(\WordArray[20].Word[4].QWire ), .OE(
        n57), .Z(DataRead[4]) );
  BUFTD1 \WordArray[20].Word[3].Buf  ( .I(\WordArray[20].Word[3].QWire ), .OE(
        n58), .Z(DataRead[3]) );
  BUFTD1 \WordArray[20].Word[2].Buf  ( .I(\WordArray[20].Word[2].QWire ), .OE(
        n57), .Z(DataRead[2]) );
  BUFTD1 \WordArray[20].Word[1].Buf  ( .I(\WordArray[20].Word[1].QWire ), .OE(
        n58), .Z(DataRead[1]) );
  BUFTD1 \WordArray[20].Word[0].Buf  ( .I(\WordArray[20].Word[0].QWire ), .OE(
        n57), .Z(DataRead[0]) );
  BUFTD1 \WordArray[19].Word[31].Buf  ( .I(\WordArray[19].Word[31].QWire ), 
        .OE(n60), .Z(DataRead[31]) );
  BUFTD1 \WordArray[19].Word[30].Buf  ( .I(\WordArray[19].Word[30].QWire ), 
        .OE(n60), .Z(DataRead[30]) );
  BUFTD1 \WordArray[19].Word[29].Buf  ( .I(\WordArray[19].Word[29].QWire ), 
        .OE(n60), .Z(DataRead[29]) );
  BUFTD1 \WordArray[19].Word[28].Buf  ( .I(\WordArray[19].Word[28].QWire ), 
        .OE(n59), .Z(DataRead[28]) );
  BUFTD1 \WordArray[19].Word[27].Buf  ( .I(\WordArray[19].Word[27].QWire ), 
        .OE(n60), .Z(DataRead[27]) );
  BUFTD1 \WordArray[19].Word[26].Buf  ( .I(\WordArray[19].Word[26].QWire ), 
        .OE(n59), .Z(DataRead[26]) );
  BUFTD1 \WordArray[19].Word[25].Buf  ( .I(\WordArray[19].Word[25].QWire ), 
        .OE(n60), .Z(DataRead[25]) );
  BUFTD1 \WordArray[19].Word[24].Buf  ( .I(\WordArray[19].Word[24].QWire ), 
        .OE(n60), .Z(DataRead[24]) );
  BUFTD1 \WordArray[19].Word[23].Buf  ( .I(\WordArray[19].Word[23].QWire ), 
        .OE(n60), .Z(DataRead[23]) );
  BUFTD1 \WordArray[19].Word[22].Buf  ( .I(\WordArray[19].Word[22].QWire ), 
        .OE(n59), .Z(DataRead[22]) );
  BUFTD1 \WordArray[19].Word[21].Buf  ( .I(\WordArray[19].Word[21].QWire ), 
        .OE(n60), .Z(DataRead[21]) );
  BUFTD1 \WordArray[19].Word[20].Buf  ( .I(\WordArray[19].Word[20].QWire ), 
        .OE(n60), .Z(DataRead[20]) );
  BUFTD1 \WordArray[19].Word[19].Buf  ( .I(\WordArray[19].Word[19].QWire ), 
        .OE(n59), .Z(DataRead[19]) );
  BUFTD1 \WordArray[19].Word[18].Buf  ( .I(\WordArray[19].Word[18].QWire ), 
        .OE(n59), .Z(DataRead[18]) );
  BUFTD1 \WordArray[19].Word[17].Buf  ( .I(\WordArray[19].Word[17].QWire ), 
        .OE(n59), .Z(DataRead[17]) );
  BUFTD1 \WordArray[19].Word[16].Buf  ( .I(\WordArray[19].Word[16].QWire ), 
        .OE(n59), .Z(DataRead[16]) );
  BUFTD1 \WordArray[19].Word[15].Buf  ( .I(\WordArray[19].Word[15].QWire ), 
        .OE(n59), .Z(DataRead[15]) );
  BUFTD1 \WordArray[19].Word[14].Buf  ( .I(\WordArray[19].Word[14].QWire ), 
        .OE(n59), .Z(DataRead[14]) );
  BUFTD1 \WordArray[19].Word[13].Buf  ( .I(\WordArray[19].Word[13].QWire ), 
        .OE(n59), .Z(DataRead[13]) );
  BUFTD1 \WordArray[19].Word[12].Buf  ( .I(\WordArray[19].Word[12].QWire ), 
        .OE(n59), .Z(DataRead[12]) );
  BUFTD1 \WordArray[19].Word[11].Buf  ( .I(\WordArray[19].Word[11].QWire ), 
        .OE(n59), .Z(DataRead[11]) );
  BUFTD1 \WordArray[19].Word[10].Buf  ( .I(\WordArray[19].Word[10].QWire ), 
        .OE(n59), .Z(DataRead[10]) );
  BUFTD1 \WordArray[19].Word[9].Buf  ( .I(\WordArray[19].Word[9].QWire ), .OE(
        n60), .Z(DataRead[9]) );
  BUFTD1 \WordArray[19].Word[8].Buf  ( .I(\WordArray[19].Word[8].QWire ), .OE(
        n60), .Z(DataRead[8]) );
  BUFTD1 \WordArray[19].Word[7].Buf  ( .I(\WordArray[19].Word[7].QWire ), .OE(
        n60), .Z(DataRead[7]) );
  BUFTD1 \WordArray[19].Word[6].Buf  ( .I(\WordArray[19].Word[6].QWire ), .OE(
        n60), .Z(DataRead[6]) );
  BUFTD1 \WordArray[19].Word[5].Buf  ( .I(\WordArray[19].Word[5].QWire ), .OE(
        n60), .Z(DataRead[5]) );
  BUFTD1 \WordArray[19].Word[4].Buf  ( .I(\WordArray[19].Word[4].QWire ), .OE(
        n59), .Z(DataRead[4]) );
  BUFTD1 \WordArray[19].Word[3].Buf  ( .I(\WordArray[19].Word[3].QWire ), .OE(
        n60), .Z(DataRead[3]) );
  BUFTD1 \WordArray[19].Word[2].Buf  ( .I(\WordArray[19].Word[2].QWire ), .OE(
        n59), .Z(DataRead[2]) );
  BUFTD1 \WordArray[19].Word[1].Buf  ( .I(\WordArray[19].Word[1].QWire ), .OE(
        n60), .Z(DataRead[1]) );
  BUFTD1 \WordArray[19].Word[0].Buf  ( .I(\WordArray[19].Word[0].QWire ), .OE(
        n59), .Z(DataRead[0]) );
  BUFTD1 \WordArray[18].Word[31].Buf  ( .I(\WordArray[18].Word[31].QWire ), 
        .OE(n62), .Z(DataRead[31]) );
  BUFTD1 \WordArray[18].Word[30].Buf  ( .I(\WordArray[18].Word[30].QWire ), 
        .OE(n62), .Z(DataRead[30]) );
  BUFTD1 \WordArray[18].Word[29].Buf  ( .I(\WordArray[18].Word[29].QWire ), 
        .OE(n62), .Z(DataRead[29]) );
  BUFTD1 \WordArray[18].Word[28].Buf  ( .I(\WordArray[18].Word[28].QWire ), 
        .OE(n61), .Z(DataRead[28]) );
  BUFTD1 \WordArray[18].Word[27].Buf  ( .I(\WordArray[18].Word[27].QWire ), 
        .OE(n62), .Z(DataRead[27]) );
  BUFTD1 \WordArray[18].Word[26].Buf  ( .I(\WordArray[18].Word[26].QWire ), 
        .OE(n61), .Z(DataRead[26]) );
  BUFTD1 \WordArray[18].Word[25].Buf  ( .I(\WordArray[18].Word[25].QWire ), 
        .OE(n62), .Z(DataRead[25]) );
  BUFTD1 \WordArray[18].Word[24].Buf  ( .I(\WordArray[18].Word[24].QWire ), 
        .OE(n62), .Z(DataRead[24]) );
  BUFTD1 \WordArray[18].Word[23].Buf  ( .I(\WordArray[18].Word[23].QWire ), 
        .OE(n62), .Z(DataRead[23]) );
  BUFTD1 \WordArray[18].Word[22].Buf  ( .I(\WordArray[18].Word[22].QWire ), 
        .OE(n61), .Z(DataRead[22]) );
  BUFTD1 \WordArray[18].Word[21].Buf  ( .I(\WordArray[18].Word[21].QWire ), 
        .OE(n62), .Z(DataRead[21]) );
  BUFTD1 \WordArray[18].Word[20].Buf  ( .I(\WordArray[18].Word[20].QWire ), 
        .OE(n62), .Z(DataRead[20]) );
  BUFTD1 \WordArray[18].Word[19].Buf  ( .I(\WordArray[18].Word[19].QWire ), 
        .OE(n61), .Z(DataRead[19]) );
  BUFTD1 \WordArray[18].Word[18].Buf  ( .I(\WordArray[18].Word[18].QWire ), 
        .OE(n61), .Z(DataRead[18]) );
  BUFTD1 \WordArray[18].Word[17].Buf  ( .I(\WordArray[18].Word[17].QWire ), 
        .OE(n61), .Z(DataRead[17]) );
  BUFTD1 \WordArray[18].Word[16].Buf  ( .I(\WordArray[18].Word[16].QWire ), 
        .OE(n61), .Z(DataRead[16]) );
  BUFTD1 \WordArray[18].Word[15].Buf  ( .I(\WordArray[18].Word[15].QWire ), 
        .OE(n61), .Z(DataRead[15]) );
  BUFTD1 \WordArray[18].Word[14].Buf  ( .I(\WordArray[18].Word[14].QWire ), 
        .OE(n61), .Z(DataRead[14]) );
  BUFTD1 \WordArray[18].Word[13].Buf  ( .I(\WordArray[18].Word[13].QWire ), 
        .OE(n61), .Z(DataRead[13]) );
  BUFTD1 \WordArray[18].Word[12].Buf  ( .I(\WordArray[18].Word[12].QWire ), 
        .OE(n61), .Z(DataRead[12]) );
  BUFTD1 \WordArray[18].Word[11].Buf  ( .I(\WordArray[18].Word[11].QWire ), 
        .OE(n61), .Z(DataRead[11]) );
  BUFTD1 \WordArray[18].Word[10].Buf  ( .I(\WordArray[18].Word[10].QWire ), 
        .OE(n61), .Z(DataRead[10]) );
  BUFTD1 \WordArray[18].Word[9].Buf  ( .I(\WordArray[18].Word[9].QWire ), .OE(
        n62), .Z(DataRead[9]) );
  BUFTD1 \WordArray[18].Word[8].Buf  ( .I(\WordArray[18].Word[8].QWire ), .OE(
        n62), .Z(DataRead[8]) );
  BUFTD1 \WordArray[18].Word[7].Buf  ( .I(\WordArray[18].Word[7].QWire ), .OE(
        n62), .Z(DataRead[7]) );
  BUFTD1 \WordArray[18].Word[6].Buf  ( .I(\WordArray[18].Word[6].QWire ), .OE(
        n62), .Z(DataRead[6]) );
  BUFTD1 \WordArray[18].Word[5].Buf  ( .I(\WordArray[18].Word[5].QWire ), .OE(
        n62), .Z(DataRead[5]) );
  BUFTD1 \WordArray[18].Word[4].Buf  ( .I(\WordArray[18].Word[4].QWire ), .OE(
        n61), .Z(DataRead[4]) );
  BUFTD1 \WordArray[18].Word[3].Buf  ( .I(\WordArray[18].Word[3].QWire ), .OE(
        n62), .Z(DataRead[3]) );
  BUFTD1 \WordArray[18].Word[2].Buf  ( .I(\WordArray[18].Word[2].QWire ), .OE(
        n61), .Z(DataRead[2]) );
  BUFTD1 \WordArray[18].Word[1].Buf  ( .I(\WordArray[18].Word[1].QWire ), .OE(
        n62), .Z(DataRead[1]) );
  BUFTD1 \WordArray[18].Word[0].Buf  ( .I(\WordArray[18].Word[0].QWire ), .OE(
        n61), .Z(DataRead[0]) );
  BUFTD1 \WordArray[17].Word[31].Buf  ( .I(\WordArray[17].Word[31].QWire ), 
        .OE(n64), .Z(DataRead[31]) );
  BUFTD1 \WordArray[17].Word[30].Buf  ( .I(\WordArray[17].Word[30].QWire ), 
        .OE(n64), .Z(DataRead[30]) );
  BUFTD1 \WordArray[17].Word[29].Buf  ( .I(\WordArray[17].Word[29].QWire ), 
        .OE(n64), .Z(DataRead[29]) );
  BUFTD1 \WordArray[17].Word[28].Buf  ( .I(\WordArray[17].Word[28].QWire ), 
        .OE(n63), .Z(DataRead[28]) );
  BUFTD1 \WordArray[17].Word[27].Buf  ( .I(\WordArray[17].Word[27].QWire ), 
        .OE(n64), .Z(DataRead[27]) );
  BUFTD1 \WordArray[17].Word[26].Buf  ( .I(\WordArray[17].Word[26].QWire ), 
        .OE(n63), .Z(DataRead[26]) );
  BUFTD1 \WordArray[17].Word[25].Buf  ( .I(\WordArray[17].Word[25].QWire ), 
        .OE(n64), .Z(DataRead[25]) );
  BUFTD1 \WordArray[17].Word[24].Buf  ( .I(\WordArray[17].Word[24].QWire ), 
        .OE(n64), .Z(DataRead[24]) );
  BUFTD1 \WordArray[17].Word[23].Buf  ( .I(\WordArray[17].Word[23].QWire ), 
        .OE(n64), .Z(DataRead[23]) );
  BUFTD1 \WordArray[17].Word[22].Buf  ( .I(\WordArray[17].Word[22].QWire ), 
        .OE(n63), .Z(DataRead[22]) );
  BUFTD1 \WordArray[17].Word[21].Buf  ( .I(\WordArray[17].Word[21].QWire ), 
        .OE(n64), .Z(DataRead[21]) );
  BUFTD1 \WordArray[17].Word[20].Buf  ( .I(\WordArray[17].Word[20].QWire ), 
        .OE(n64), .Z(DataRead[20]) );
  BUFTD1 \WordArray[17].Word[19].Buf  ( .I(\WordArray[17].Word[19].QWire ), 
        .OE(n63), .Z(DataRead[19]) );
  BUFTD1 \WordArray[17].Word[18].Buf  ( .I(\WordArray[17].Word[18].QWire ), 
        .OE(n63), .Z(DataRead[18]) );
  BUFTD1 \WordArray[17].Word[17].Buf  ( .I(\WordArray[17].Word[17].QWire ), 
        .OE(n63), .Z(DataRead[17]) );
  BUFTD1 \WordArray[17].Word[16].Buf  ( .I(\WordArray[17].Word[16].QWire ), 
        .OE(n63), .Z(DataRead[16]) );
  BUFTD1 \WordArray[17].Word[15].Buf  ( .I(\WordArray[17].Word[15].QWire ), 
        .OE(n63), .Z(DataRead[15]) );
  BUFTD1 \WordArray[17].Word[14].Buf  ( .I(\WordArray[17].Word[14].QWire ), 
        .OE(n63), .Z(DataRead[14]) );
  BUFTD1 \WordArray[17].Word[13].Buf  ( .I(\WordArray[17].Word[13].QWire ), 
        .OE(n63), .Z(DataRead[13]) );
  BUFTD1 \WordArray[17].Word[12].Buf  ( .I(\WordArray[17].Word[12].QWire ), 
        .OE(n63), .Z(DataRead[12]) );
  BUFTD1 \WordArray[17].Word[11].Buf  ( .I(\WordArray[17].Word[11].QWire ), 
        .OE(n63), .Z(DataRead[11]) );
  BUFTD1 \WordArray[17].Word[10].Buf  ( .I(\WordArray[17].Word[10].QWire ), 
        .OE(n63), .Z(DataRead[10]) );
  BUFTD1 \WordArray[17].Word[9].Buf  ( .I(\WordArray[17].Word[9].QWire ), .OE(
        n64), .Z(DataRead[9]) );
  BUFTD1 \WordArray[17].Word[8].Buf  ( .I(\WordArray[17].Word[8].QWire ), .OE(
        n64), .Z(DataRead[8]) );
  BUFTD1 \WordArray[17].Word[7].Buf  ( .I(\WordArray[17].Word[7].QWire ), .OE(
        n64), .Z(DataRead[7]) );
  BUFTD1 \WordArray[17].Word[6].Buf  ( .I(\WordArray[17].Word[6].QWire ), .OE(
        n64), .Z(DataRead[6]) );
  BUFTD1 \WordArray[17].Word[5].Buf  ( .I(\WordArray[17].Word[5].QWire ), .OE(
        n64), .Z(DataRead[5]) );
  BUFTD1 \WordArray[17].Word[4].Buf  ( .I(\WordArray[17].Word[4].QWire ), .OE(
        n63), .Z(DataRead[4]) );
  BUFTD1 \WordArray[17].Word[3].Buf  ( .I(\WordArray[17].Word[3].QWire ), .OE(
        n64), .Z(DataRead[3]) );
  BUFTD1 \WordArray[17].Word[2].Buf  ( .I(\WordArray[17].Word[2].QWire ), .OE(
        n63), .Z(DataRead[2]) );
  BUFTD1 \WordArray[17].Word[1].Buf  ( .I(\WordArray[17].Word[1].QWire ), .OE(
        n64), .Z(DataRead[1]) );
  BUFTD1 \WordArray[17].Word[0].Buf  ( .I(\WordArray[17].Word[0].QWire ), .OE(
        n63), .Z(DataRead[0]) );
  BUFTD1 \WordArray[16].Word[31].Buf  ( .I(\WordArray[16].Word[31].QWire ), 
        .OE(n66), .Z(DataRead[31]) );
  BUFTD1 \WordArray[16].Word[30].Buf  ( .I(\WordArray[16].Word[30].QWire ), 
        .OE(n66), .Z(DataRead[30]) );
  BUFTD1 \WordArray[16].Word[29].Buf  ( .I(\WordArray[16].Word[29].QWire ), 
        .OE(n66), .Z(DataRead[29]) );
  BUFTD1 \WordArray[16].Word[28].Buf  ( .I(\WordArray[16].Word[28].QWire ), 
        .OE(n65), .Z(DataRead[28]) );
  BUFTD1 \WordArray[16].Word[27].Buf  ( .I(\WordArray[16].Word[27].QWire ), 
        .OE(n66), .Z(DataRead[27]) );
  BUFTD1 \WordArray[16].Word[26].Buf  ( .I(\WordArray[16].Word[26].QWire ), 
        .OE(n65), .Z(DataRead[26]) );
  BUFTD1 \WordArray[16].Word[25].Buf  ( .I(\WordArray[16].Word[25].QWire ), 
        .OE(n66), .Z(DataRead[25]) );
  BUFTD1 \WordArray[16].Word[24].Buf  ( .I(\WordArray[16].Word[24].QWire ), 
        .OE(n66), .Z(DataRead[24]) );
  BUFTD1 \WordArray[16].Word[23].Buf  ( .I(\WordArray[16].Word[23].QWire ), 
        .OE(n66), .Z(DataRead[23]) );
  BUFTD1 \WordArray[16].Word[22].Buf  ( .I(\WordArray[16].Word[22].QWire ), 
        .OE(n65), .Z(DataRead[22]) );
  BUFTD1 \WordArray[16].Word[21].Buf  ( .I(\WordArray[16].Word[21].QWire ), 
        .OE(n66), .Z(DataRead[21]) );
  BUFTD1 \WordArray[16].Word[20].Buf  ( .I(\WordArray[16].Word[20].QWire ), 
        .OE(n66), .Z(DataRead[20]) );
  BUFTD1 \WordArray[16].Word[19].Buf  ( .I(\WordArray[16].Word[19].QWire ), 
        .OE(n65), .Z(DataRead[19]) );
  BUFTD1 \WordArray[16].Word[18].Buf  ( .I(\WordArray[16].Word[18].QWire ), 
        .OE(n65), .Z(DataRead[18]) );
  BUFTD1 \WordArray[16].Word[17].Buf  ( .I(\WordArray[16].Word[17].QWire ), 
        .OE(n65), .Z(DataRead[17]) );
  BUFTD1 \WordArray[16].Word[16].Buf  ( .I(\WordArray[16].Word[16].QWire ), 
        .OE(n65), .Z(DataRead[16]) );
  BUFTD1 \WordArray[16].Word[15].Buf  ( .I(\WordArray[16].Word[15].QWire ), 
        .OE(n65), .Z(DataRead[15]) );
  BUFTD1 \WordArray[16].Word[14].Buf  ( .I(\WordArray[16].Word[14].QWire ), 
        .OE(n65), .Z(DataRead[14]) );
  BUFTD1 \WordArray[16].Word[13].Buf  ( .I(\WordArray[16].Word[13].QWire ), 
        .OE(n65), .Z(DataRead[13]) );
  BUFTD1 \WordArray[16].Word[12].Buf  ( .I(\WordArray[16].Word[12].QWire ), 
        .OE(n65), .Z(DataRead[12]) );
  BUFTD1 \WordArray[16].Word[11].Buf  ( .I(\WordArray[16].Word[11].QWire ), 
        .OE(n65), .Z(DataRead[11]) );
  BUFTD1 \WordArray[16].Word[10].Buf  ( .I(\WordArray[16].Word[10].QWire ), 
        .OE(n65), .Z(DataRead[10]) );
  BUFTD1 \WordArray[16].Word[9].Buf  ( .I(\WordArray[16].Word[9].QWire ), .OE(
        n66), .Z(DataRead[9]) );
  BUFTD1 \WordArray[16].Word[8].Buf  ( .I(\WordArray[16].Word[8].QWire ), .OE(
        n66), .Z(DataRead[8]) );
  BUFTD1 \WordArray[16].Word[7].Buf  ( .I(\WordArray[16].Word[7].QWire ), .OE(
        n66), .Z(DataRead[7]) );
  BUFTD1 \WordArray[16].Word[6].Buf  ( .I(\WordArray[16].Word[6].QWire ), .OE(
        n66), .Z(DataRead[6]) );
  BUFTD1 \WordArray[16].Word[5].Buf  ( .I(\WordArray[16].Word[5].QWire ), .OE(
        n66), .Z(DataRead[5]) );
  BUFTD1 \WordArray[16].Word[4].Buf  ( .I(\WordArray[16].Word[4].QWire ), .OE(
        n65), .Z(DataRead[4]) );
  BUFTD1 \WordArray[16].Word[3].Buf  ( .I(\WordArray[16].Word[3].QWire ), .OE(
        n66), .Z(DataRead[3]) );
  BUFTD1 \WordArray[16].Word[2].Buf  ( .I(\WordArray[16].Word[2].QWire ), .OE(
        n65), .Z(DataRead[2]) );
  BUFTD1 \WordArray[16].Word[1].Buf  ( .I(\WordArray[16].Word[1].QWire ), .OE(
        n66), .Z(DataRead[1]) );
  BUFTD1 \WordArray[16].Word[0].Buf  ( .I(\WordArray[16].Word[0].QWire ), .OE(
        n65), .Z(DataRead[0]) );
  BUFTD1 \WordArray[15].Word[31].Buf  ( .I(\WordArray[15].Word[31].QWire ), 
        .OE(n68), .Z(DataRead[31]) );
  BUFTD1 \WordArray[15].Word[30].Buf  ( .I(\WordArray[15].Word[30].QWire ), 
        .OE(n68), .Z(DataRead[30]) );
  BUFTD1 \WordArray[15].Word[29].Buf  ( .I(\WordArray[15].Word[29].QWire ), 
        .OE(n68), .Z(DataRead[29]) );
  BUFTD1 \WordArray[15].Word[28].Buf  ( .I(\WordArray[15].Word[28].QWire ), 
        .OE(n67), .Z(DataRead[28]) );
  BUFTD1 \WordArray[15].Word[27].Buf  ( .I(\WordArray[15].Word[27].QWire ), 
        .OE(n68), .Z(DataRead[27]) );
  BUFTD1 \WordArray[15].Word[26].Buf  ( .I(\WordArray[15].Word[26].QWire ), 
        .OE(n67), .Z(DataRead[26]) );
  BUFTD1 \WordArray[15].Word[25].Buf  ( .I(\WordArray[15].Word[25].QWire ), 
        .OE(n68), .Z(DataRead[25]) );
  BUFTD1 \WordArray[15].Word[24].Buf  ( .I(\WordArray[15].Word[24].QWire ), 
        .OE(n68), .Z(DataRead[24]) );
  BUFTD1 \WordArray[15].Word[23].Buf  ( .I(\WordArray[15].Word[23].QWire ), 
        .OE(n68), .Z(DataRead[23]) );
  BUFTD1 \WordArray[15].Word[22].Buf  ( .I(\WordArray[15].Word[22].QWire ), 
        .OE(n67), .Z(DataRead[22]) );
  BUFTD1 \WordArray[15].Word[21].Buf  ( .I(\WordArray[15].Word[21].QWire ), 
        .OE(n68), .Z(DataRead[21]) );
  BUFTD1 \WordArray[15].Word[20].Buf  ( .I(\WordArray[15].Word[20].QWire ), 
        .OE(n68), .Z(DataRead[20]) );
  BUFTD1 \WordArray[15].Word[19].Buf  ( .I(\WordArray[15].Word[19].QWire ), 
        .OE(n67), .Z(DataRead[19]) );
  BUFTD1 \WordArray[15].Word[18].Buf  ( .I(\WordArray[15].Word[18].QWire ), 
        .OE(n67), .Z(DataRead[18]) );
  BUFTD1 \WordArray[15].Word[17].Buf  ( .I(\WordArray[15].Word[17].QWire ), 
        .OE(n67), .Z(DataRead[17]) );
  BUFTD1 \WordArray[15].Word[16].Buf  ( .I(\WordArray[15].Word[16].QWire ), 
        .OE(n67), .Z(DataRead[16]) );
  BUFTD1 \WordArray[15].Word[15].Buf  ( .I(\WordArray[15].Word[15].QWire ), 
        .OE(n67), .Z(DataRead[15]) );
  BUFTD1 \WordArray[15].Word[14].Buf  ( .I(\WordArray[15].Word[14].QWire ), 
        .OE(n67), .Z(DataRead[14]) );
  BUFTD1 \WordArray[15].Word[13].Buf  ( .I(\WordArray[15].Word[13].QWire ), 
        .OE(n67), .Z(DataRead[13]) );
  BUFTD1 \WordArray[15].Word[12].Buf  ( .I(\WordArray[15].Word[12].QWire ), 
        .OE(n67), .Z(DataRead[12]) );
  BUFTD1 \WordArray[15].Word[11].Buf  ( .I(\WordArray[15].Word[11].QWire ), 
        .OE(n67), .Z(DataRead[11]) );
  BUFTD1 \WordArray[15].Word[10].Buf  ( .I(\WordArray[15].Word[10].QWire ), 
        .OE(n67), .Z(DataRead[10]) );
  BUFTD1 \WordArray[15].Word[9].Buf  ( .I(\WordArray[15].Word[9].QWire ), .OE(
        n68), .Z(DataRead[9]) );
  BUFTD1 \WordArray[15].Word[8].Buf  ( .I(\WordArray[15].Word[8].QWire ), .OE(
        n68), .Z(DataRead[8]) );
  BUFTD1 \WordArray[15].Word[7].Buf  ( .I(\WordArray[15].Word[7].QWire ), .OE(
        n68), .Z(DataRead[7]) );
  BUFTD1 \WordArray[15].Word[6].Buf  ( .I(\WordArray[15].Word[6].QWire ), .OE(
        n68), .Z(DataRead[6]) );
  BUFTD1 \WordArray[15].Word[5].Buf  ( .I(\WordArray[15].Word[5].QWire ), .OE(
        n68), .Z(DataRead[5]) );
  BUFTD1 \WordArray[15].Word[4].Buf  ( .I(\WordArray[15].Word[4].QWire ), .OE(
        n67), .Z(DataRead[4]) );
  BUFTD1 \WordArray[15].Word[3].Buf  ( .I(\WordArray[15].Word[3].QWire ), .OE(
        n68), .Z(DataRead[3]) );
  BUFTD1 \WordArray[15].Word[2].Buf  ( .I(\WordArray[15].Word[2].QWire ), .OE(
        n67), .Z(DataRead[2]) );
  BUFTD1 \WordArray[15].Word[1].Buf  ( .I(\WordArray[15].Word[1].QWire ), .OE(
        n68), .Z(DataRead[1]) );
  BUFTD1 \WordArray[15].Word[0].Buf  ( .I(\WordArray[15].Word[0].QWire ), .OE(
        n67), .Z(DataRead[0]) );
  BUFTD1 \WordArray[14].Word[31].Buf  ( .I(\WordArray[14].Word[31].QWire ), 
        .OE(n70), .Z(DataRead[31]) );
  BUFTD1 \WordArray[14].Word[30].Buf  ( .I(\WordArray[14].Word[30].QWire ), 
        .OE(n70), .Z(DataRead[30]) );
  BUFTD1 \WordArray[14].Word[29].Buf  ( .I(\WordArray[14].Word[29].QWire ), 
        .OE(n70), .Z(DataRead[29]) );
  BUFTD1 \WordArray[14].Word[28].Buf  ( .I(\WordArray[14].Word[28].QWire ), 
        .OE(n69), .Z(DataRead[28]) );
  BUFTD1 \WordArray[14].Word[27].Buf  ( .I(\WordArray[14].Word[27].QWire ), 
        .OE(n70), .Z(DataRead[27]) );
  BUFTD1 \WordArray[14].Word[26].Buf  ( .I(\WordArray[14].Word[26].QWire ), 
        .OE(n69), .Z(DataRead[26]) );
  BUFTD1 \WordArray[14].Word[25].Buf  ( .I(\WordArray[14].Word[25].QWire ), 
        .OE(n70), .Z(DataRead[25]) );
  BUFTD1 \WordArray[14].Word[24].Buf  ( .I(\WordArray[14].Word[24].QWire ), 
        .OE(n70), .Z(DataRead[24]) );
  BUFTD1 \WordArray[14].Word[23].Buf  ( .I(\WordArray[14].Word[23].QWire ), 
        .OE(n70), .Z(DataRead[23]) );
  BUFTD1 \WordArray[14].Word[22].Buf  ( .I(\WordArray[14].Word[22].QWire ), 
        .OE(n69), .Z(DataRead[22]) );
  BUFTD1 \WordArray[14].Word[21].Buf  ( .I(\WordArray[14].Word[21].QWire ), 
        .OE(n70), .Z(DataRead[21]) );
  BUFTD1 \WordArray[14].Word[20].Buf  ( .I(\WordArray[14].Word[20].QWire ), 
        .OE(n70), .Z(DataRead[20]) );
  BUFTD1 \WordArray[14].Word[19].Buf  ( .I(\WordArray[14].Word[19].QWire ), 
        .OE(n69), .Z(DataRead[19]) );
  BUFTD1 \WordArray[14].Word[18].Buf  ( .I(\WordArray[14].Word[18].QWire ), 
        .OE(n69), .Z(DataRead[18]) );
  BUFTD1 \WordArray[14].Word[17].Buf  ( .I(\WordArray[14].Word[17].QWire ), 
        .OE(n69), .Z(DataRead[17]) );
  BUFTD1 \WordArray[14].Word[16].Buf  ( .I(\WordArray[14].Word[16].QWire ), 
        .OE(n69), .Z(DataRead[16]) );
  BUFTD1 \WordArray[14].Word[15].Buf  ( .I(\WordArray[14].Word[15].QWire ), 
        .OE(n69), .Z(DataRead[15]) );
  BUFTD1 \WordArray[14].Word[14].Buf  ( .I(\WordArray[14].Word[14].QWire ), 
        .OE(n69), .Z(DataRead[14]) );
  BUFTD1 \WordArray[14].Word[13].Buf  ( .I(\WordArray[14].Word[13].QWire ), 
        .OE(n69), .Z(DataRead[13]) );
  BUFTD1 \WordArray[14].Word[12].Buf  ( .I(\WordArray[14].Word[12].QWire ), 
        .OE(n69), .Z(DataRead[12]) );
  BUFTD1 \WordArray[14].Word[11].Buf  ( .I(\WordArray[14].Word[11].QWire ), 
        .OE(n69), .Z(DataRead[11]) );
  BUFTD1 \WordArray[14].Word[10].Buf  ( .I(\WordArray[14].Word[10].QWire ), 
        .OE(n69), .Z(DataRead[10]) );
  BUFTD1 \WordArray[14].Word[9].Buf  ( .I(\WordArray[14].Word[9].QWire ), .OE(
        n70), .Z(DataRead[9]) );
  BUFTD1 \WordArray[14].Word[8].Buf  ( .I(\WordArray[14].Word[8].QWire ), .OE(
        n70), .Z(DataRead[8]) );
  BUFTD1 \WordArray[14].Word[7].Buf  ( .I(\WordArray[14].Word[7].QWire ), .OE(
        n70), .Z(DataRead[7]) );
  BUFTD1 \WordArray[14].Word[6].Buf  ( .I(\WordArray[14].Word[6].QWire ), .OE(
        n70), .Z(DataRead[6]) );
  BUFTD1 \WordArray[14].Word[5].Buf  ( .I(\WordArray[14].Word[5].QWire ), .OE(
        n70), .Z(DataRead[5]) );
  BUFTD1 \WordArray[14].Word[4].Buf  ( .I(\WordArray[14].Word[4].QWire ), .OE(
        n69), .Z(DataRead[4]) );
  BUFTD1 \WordArray[14].Word[3].Buf  ( .I(\WordArray[14].Word[3].QWire ), .OE(
        n70), .Z(DataRead[3]) );
  BUFTD1 \WordArray[14].Word[2].Buf  ( .I(\WordArray[14].Word[2].QWire ), .OE(
        n69), .Z(DataRead[2]) );
  BUFTD1 \WordArray[14].Word[1].Buf  ( .I(\WordArray[14].Word[1].QWire ), .OE(
        n70), .Z(DataRead[1]) );
  BUFTD1 \WordArray[14].Word[0].Buf  ( .I(\WordArray[14].Word[0].QWire ), .OE(
        n69), .Z(DataRead[0]) );
  BUFTD1 \WordArray[13].Word[31].Buf  ( .I(\WordArray[13].Word[31].QWire ), 
        .OE(n72), .Z(DataRead[31]) );
  BUFTD1 \WordArray[13].Word[30].Buf  ( .I(\WordArray[13].Word[30].QWire ), 
        .OE(n72), .Z(DataRead[30]) );
  BUFTD1 \WordArray[13].Word[29].Buf  ( .I(\WordArray[13].Word[29].QWire ), 
        .OE(n72), .Z(DataRead[29]) );
  BUFTD1 \WordArray[13].Word[28].Buf  ( .I(\WordArray[13].Word[28].QWire ), 
        .OE(n71), .Z(DataRead[28]) );
  BUFTD1 \WordArray[13].Word[27].Buf  ( .I(\WordArray[13].Word[27].QWire ), 
        .OE(n72), .Z(DataRead[27]) );
  BUFTD1 \WordArray[13].Word[26].Buf  ( .I(\WordArray[13].Word[26].QWire ), 
        .OE(n71), .Z(DataRead[26]) );
  BUFTD1 \WordArray[13].Word[25].Buf  ( .I(\WordArray[13].Word[25].QWire ), 
        .OE(n72), .Z(DataRead[25]) );
  BUFTD1 \WordArray[13].Word[24].Buf  ( .I(\WordArray[13].Word[24].QWire ), 
        .OE(n72), .Z(DataRead[24]) );
  BUFTD1 \WordArray[13].Word[23].Buf  ( .I(\WordArray[13].Word[23].QWire ), 
        .OE(n72), .Z(DataRead[23]) );
  BUFTD1 \WordArray[13].Word[22].Buf  ( .I(\WordArray[13].Word[22].QWire ), 
        .OE(n71), .Z(DataRead[22]) );
  BUFTD1 \WordArray[13].Word[21].Buf  ( .I(\WordArray[13].Word[21].QWire ), 
        .OE(n72), .Z(DataRead[21]) );
  BUFTD1 \WordArray[13].Word[20].Buf  ( .I(\WordArray[13].Word[20].QWire ), 
        .OE(n72), .Z(DataRead[20]) );
  BUFTD1 \WordArray[13].Word[19].Buf  ( .I(\WordArray[13].Word[19].QWire ), 
        .OE(n71), .Z(DataRead[19]) );
  BUFTD1 \WordArray[13].Word[18].Buf  ( .I(\WordArray[13].Word[18].QWire ), 
        .OE(n71), .Z(DataRead[18]) );
  BUFTD1 \WordArray[13].Word[17].Buf  ( .I(\WordArray[13].Word[17].QWire ), 
        .OE(n71), .Z(DataRead[17]) );
  BUFTD1 \WordArray[13].Word[16].Buf  ( .I(\WordArray[13].Word[16].QWire ), 
        .OE(n71), .Z(DataRead[16]) );
  BUFTD1 \WordArray[13].Word[15].Buf  ( .I(\WordArray[13].Word[15].QWire ), 
        .OE(n71), .Z(DataRead[15]) );
  BUFTD1 \WordArray[13].Word[14].Buf  ( .I(\WordArray[13].Word[14].QWire ), 
        .OE(n71), .Z(DataRead[14]) );
  BUFTD1 \WordArray[13].Word[13].Buf  ( .I(\WordArray[13].Word[13].QWire ), 
        .OE(n71), .Z(DataRead[13]) );
  BUFTD1 \WordArray[13].Word[12].Buf  ( .I(\WordArray[13].Word[12].QWire ), 
        .OE(n71), .Z(DataRead[12]) );
  BUFTD1 \WordArray[13].Word[11].Buf  ( .I(\WordArray[13].Word[11].QWire ), 
        .OE(n71), .Z(DataRead[11]) );
  BUFTD1 \WordArray[13].Word[10].Buf  ( .I(\WordArray[13].Word[10].QWire ), 
        .OE(n71), .Z(DataRead[10]) );
  BUFTD1 \WordArray[13].Word[9].Buf  ( .I(\WordArray[13].Word[9].QWire ), .OE(
        n72), .Z(DataRead[9]) );
  BUFTD1 \WordArray[13].Word[8].Buf  ( .I(\WordArray[13].Word[8].QWire ), .OE(
        n72), .Z(DataRead[8]) );
  BUFTD1 \WordArray[13].Word[7].Buf  ( .I(\WordArray[13].Word[7].QWire ), .OE(
        n72), .Z(DataRead[7]) );
  BUFTD1 \WordArray[13].Word[6].Buf  ( .I(\WordArray[13].Word[6].QWire ), .OE(
        n72), .Z(DataRead[6]) );
  BUFTD1 \WordArray[13].Word[5].Buf  ( .I(\WordArray[13].Word[5].QWire ), .OE(
        n72), .Z(DataRead[5]) );
  BUFTD1 \WordArray[13].Word[4].Buf  ( .I(\WordArray[13].Word[4].QWire ), .OE(
        n71), .Z(DataRead[4]) );
  BUFTD1 \WordArray[13].Word[3].Buf  ( .I(\WordArray[13].Word[3].QWire ), .OE(
        n72), .Z(DataRead[3]) );
  BUFTD1 \WordArray[13].Word[2].Buf  ( .I(\WordArray[13].Word[2].QWire ), .OE(
        n71), .Z(DataRead[2]) );
  BUFTD1 \WordArray[13].Word[1].Buf  ( .I(\WordArray[13].Word[1].QWire ), .OE(
        n72), .Z(DataRead[1]) );
  BUFTD1 \WordArray[13].Word[0].Buf  ( .I(\WordArray[13].Word[0].QWire ), .OE(
        n71), .Z(DataRead[0]) );
  BUFTD1 \WordArray[12].Word[31].Buf  ( .I(\WordArray[12].Word[31].QWire ), 
        .OE(n74), .Z(DataRead[31]) );
  BUFTD1 \WordArray[12].Word[30].Buf  ( .I(\WordArray[12].Word[30].QWire ), 
        .OE(n74), .Z(DataRead[30]) );
  BUFTD1 \WordArray[12].Word[29].Buf  ( .I(\WordArray[12].Word[29].QWire ), 
        .OE(n74), .Z(DataRead[29]) );
  BUFTD1 \WordArray[12].Word[28].Buf  ( .I(\WordArray[12].Word[28].QWire ), 
        .OE(n73), .Z(DataRead[28]) );
  BUFTD1 \WordArray[12].Word[27].Buf  ( .I(\WordArray[12].Word[27].QWire ), 
        .OE(n74), .Z(DataRead[27]) );
  BUFTD1 \WordArray[12].Word[26].Buf  ( .I(\WordArray[12].Word[26].QWire ), 
        .OE(n73), .Z(DataRead[26]) );
  BUFTD1 \WordArray[12].Word[25].Buf  ( .I(\WordArray[12].Word[25].QWire ), 
        .OE(n74), .Z(DataRead[25]) );
  BUFTD1 \WordArray[12].Word[24].Buf  ( .I(\WordArray[12].Word[24].QWire ), 
        .OE(n74), .Z(DataRead[24]) );
  BUFTD1 \WordArray[12].Word[23].Buf  ( .I(\WordArray[12].Word[23].QWire ), 
        .OE(n74), .Z(DataRead[23]) );
  BUFTD1 \WordArray[12].Word[22].Buf  ( .I(\WordArray[12].Word[22].QWire ), 
        .OE(n73), .Z(DataRead[22]) );
  BUFTD1 \WordArray[12].Word[21].Buf  ( .I(\WordArray[12].Word[21].QWire ), 
        .OE(n74), .Z(DataRead[21]) );
  BUFTD1 \WordArray[12].Word[20].Buf  ( .I(\WordArray[12].Word[20].QWire ), 
        .OE(n74), .Z(DataRead[20]) );
  BUFTD1 \WordArray[12].Word[19].Buf  ( .I(\WordArray[12].Word[19].QWire ), 
        .OE(n73), .Z(DataRead[19]) );
  BUFTD1 \WordArray[12].Word[18].Buf  ( .I(\WordArray[12].Word[18].QWire ), 
        .OE(n73), .Z(DataRead[18]) );
  BUFTD1 \WordArray[12].Word[17].Buf  ( .I(\WordArray[12].Word[17].QWire ), 
        .OE(n73), .Z(DataRead[17]) );
  BUFTD1 \WordArray[12].Word[16].Buf  ( .I(\WordArray[12].Word[16].QWire ), 
        .OE(n73), .Z(DataRead[16]) );
  BUFTD1 \WordArray[12].Word[15].Buf  ( .I(\WordArray[12].Word[15].QWire ), 
        .OE(n73), .Z(DataRead[15]) );
  BUFTD1 \WordArray[12].Word[14].Buf  ( .I(\WordArray[12].Word[14].QWire ), 
        .OE(n73), .Z(DataRead[14]) );
  BUFTD1 \WordArray[12].Word[13].Buf  ( .I(\WordArray[12].Word[13].QWire ), 
        .OE(n73), .Z(DataRead[13]) );
  BUFTD1 \WordArray[12].Word[12].Buf  ( .I(\WordArray[12].Word[12].QWire ), 
        .OE(n73), .Z(DataRead[12]) );
  BUFTD1 \WordArray[12].Word[11].Buf  ( .I(\WordArray[12].Word[11].QWire ), 
        .OE(n73), .Z(DataRead[11]) );
  BUFTD1 \WordArray[12].Word[10].Buf  ( .I(\WordArray[12].Word[10].QWire ), 
        .OE(n73), .Z(DataRead[10]) );
  BUFTD1 \WordArray[12].Word[9].Buf  ( .I(\WordArray[12].Word[9].QWire ), .OE(
        n74), .Z(DataRead[9]) );
  BUFTD1 \WordArray[12].Word[8].Buf  ( .I(\WordArray[12].Word[8].QWire ), .OE(
        n74), .Z(DataRead[8]) );
  BUFTD1 \WordArray[12].Word[7].Buf  ( .I(\WordArray[12].Word[7].QWire ), .OE(
        n74), .Z(DataRead[7]) );
  BUFTD1 \WordArray[12].Word[6].Buf  ( .I(\WordArray[12].Word[6].QWire ), .OE(
        n74), .Z(DataRead[6]) );
  BUFTD1 \WordArray[12].Word[5].Buf  ( .I(\WordArray[12].Word[5].QWire ), .OE(
        n74), .Z(DataRead[5]) );
  BUFTD1 \WordArray[12].Word[4].Buf  ( .I(\WordArray[12].Word[4].QWire ), .OE(
        n73), .Z(DataRead[4]) );
  BUFTD1 \WordArray[12].Word[3].Buf  ( .I(\WordArray[12].Word[3].QWire ), .OE(
        n74), .Z(DataRead[3]) );
  BUFTD1 \WordArray[12].Word[2].Buf  ( .I(\WordArray[12].Word[2].QWire ), .OE(
        n73), .Z(DataRead[2]) );
  BUFTD1 \WordArray[12].Word[1].Buf  ( .I(\WordArray[12].Word[1].QWire ), .OE(
        n74), .Z(DataRead[1]) );
  BUFTD1 \WordArray[12].Word[0].Buf  ( .I(\WordArray[12].Word[0].QWire ), .OE(
        n73), .Z(DataRead[0]) );
  BUFTD1 \WordArray[11].Word[31].Buf  ( .I(\WordArray[11].Word[31].QWire ), 
        .OE(n76), .Z(DataRead[31]) );
  BUFTD1 \WordArray[11].Word[30].Buf  ( .I(\WordArray[11].Word[30].QWire ), 
        .OE(n76), .Z(DataRead[30]) );
  BUFTD1 \WordArray[11].Word[29].Buf  ( .I(\WordArray[11].Word[29].QWire ), 
        .OE(n76), .Z(DataRead[29]) );
  BUFTD1 \WordArray[11].Word[28].Buf  ( .I(\WordArray[11].Word[28].QWire ), 
        .OE(n75), .Z(DataRead[28]) );
  BUFTD1 \WordArray[11].Word[27].Buf  ( .I(\WordArray[11].Word[27].QWire ), 
        .OE(n76), .Z(DataRead[27]) );
  BUFTD1 \WordArray[11].Word[26].Buf  ( .I(\WordArray[11].Word[26].QWire ), 
        .OE(n75), .Z(DataRead[26]) );
  BUFTD1 \WordArray[11].Word[25].Buf  ( .I(\WordArray[11].Word[25].QWire ), 
        .OE(n76), .Z(DataRead[25]) );
  BUFTD1 \WordArray[11].Word[24].Buf  ( .I(\WordArray[11].Word[24].QWire ), 
        .OE(n76), .Z(DataRead[24]) );
  BUFTD1 \WordArray[11].Word[23].Buf  ( .I(\WordArray[11].Word[23].QWire ), 
        .OE(n76), .Z(DataRead[23]) );
  BUFTD1 \WordArray[11].Word[22].Buf  ( .I(\WordArray[11].Word[22].QWire ), 
        .OE(n75), .Z(DataRead[22]) );
  BUFTD1 \WordArray[11].Word[21].Buf  ( .I(\WordArray[11].Word[21].QWire ), 
        .OE(n76), .Z(DataRead[21]) );
  BUFTD1 \WordArray[11].Word[20].Buf  ( .I(\WordArray[11].Word[20].QWire ), 
        .OE(n76), .Z(DataRead[20]) );
  BUFTD1 \WordArray[11].Word[19].Buf  ( .I(\WordArray[11].Word[19].QWire ), 
        .OE(n75), .Z(DataRead[19]) );
  BUFTD1 \WordArray[11].Word[18].Buf  ( .I(\WordArray[11].Word[18].QWire ), 
        .OE(n75), .Z(DataRead[18]) );
  BUFTD1 \WordArray[11].Word[17].Buf  ( .I(\WordArray[11].Word[17].QWire ), 
        .OE(n75), .Z(DataRead[17]) );
  BUFTD1 \WordArray[11].Word[16].Buf  ( .I(\WordArray[11].Word[16].QWire ), 
        .OE(n75), .Z(DataRead[16]) );
  BUFTD1 \WordArray[11].Word[15].Buf  ( .I(\WordArray[11].Word[15].QWire ), 
        .OE(n75), .Z(DataRead[15]) );
  BUFTD1 \WordArray[11].Word[14].Buf  ( .I(\WordArray[11].Word[14].QWire ), 
        .OE(n75), .Z(DataRead[14]) );
  BUFTD1 \WordArray[11].Word[13].Buf  ( .I(\WordArray[11].Word[13].QWire ), 
        .OE(n75), .Z(DataRead[13]) );
  BUFTD1 \WordArray[11].Word[12].Buf  ( .I(\WordArray[11].Word[12].QWire ), 
        .OE(n75), .Z(DataRead[12]) );
  BUFTD1 \WordArray[11].Word[11].Buf  ( .I(\WordArray[11].Word[11].QWire ), 
        .OE(n75), .Z(DataRead[11]) );
  BUFTD1 \WordArray[11].Word[10].Buf  ( .I(\WordArray[11].Word[10].QWire ), 
        .OE(n75), .Z(DataRead[10]) );
  BUFTD1 \WordArray[11].Word[9].Buf  ( .I(\WordArray[11].Word[9].QWire ), .OE(
        n76), .Z(DataRead[9]) );
  BUFTD1 \WordArray[11].Word[8].Buf  ( .I(\WordArray[11].Word[8].QWire ), .OE(
        n76), .Z(DataRead[8]) );
  BUFTD1 \WordArray[11].Word[7].Buf  ( .I(\WordArray[11].Word[7].QWire ), .OE(
        n76), .Z(DataRead[7]) );
  BUFTD1 \WordArray[11].Word[6].Buf  ( .I(\WordArray[11].Word[6].QWire ), .OE(
        n76), .Z(DataRead[6]) );
  BUFTD1 \WordArray[11].Word[5].Buf  ( .I(\WordArray[11].Word[5].QWire ), .OE(
        n76), .Z(DataRead[5]) );
  BUFTD1 \WordArray[11].Word[4].Buf  ( .I(\WordArray[11].Word[4].QWire ), .OE(
        n75), .Z(DataRead[4]) );
  BUFTD1 \WordArray[11].Word[3].Buf  ( .I(\WordArray[11].Word[3].QWire ), .OE(
        n76), .Z(DataRead[3]) );
  BUFTD1 \WordArray[11].Word[2].Buf  ( .I(\WordArray[11].Word[2].QWire ), .OE(
        n75), .Z(DataRead[2]) );
  BUFTD1 \WordArray[11].Word[1].Buf  ( .I(\WordArray[11].Word[1].QWire ), .OE(
        n76), .Z(DataRead[1]) );
  BUFTD1 \WordArray[11].Word[0].Buf  ( .I(\WordArray[11].Word[0].QWire ), .OE(
        n75), .Z(DataRead[0]) );
  BUFTD1 \WordArray[10].Word[31].Buf  ( .I(\WordArray[10].Word[31].QWire ), 
        .OE(n78), .Z(DataRead[31]) );
  BUFTD1 \WordArray[10].Word[30].Buf  ( .I(\WordArray[10].Word[30].QWire ), 
        .OE(n78), .Z(DataRead[30]) );
  BUFTD1 \WordArray[10].Word[29].Buf  ( .I(\WordArray[10].Word[29].QWire ), 
        .OE(n78), .Z(DataRead[29]) );
  BUFTD1 \WordArray[10].Word[28].Buf  ( .I(\WordArray[10].Word[28].QWire ), 
        .OE(n77), .Z(DataRead[28]) );
  BUFTD1 \WordArray[10].Word[27].Buf  ( .I(\WordArray[10].Word[27].QWire ), 
        .OE(n78), .Z(DataRead[27]) );
  BUFTD1 \WordArray[10].Word[26].Buf  ( .I(\WordArray[10].Word[26].QWire ), 
        .OE(n77), .Z(DataRead[26]) );
  BUFTD1 \WordArray[10].Word[25].Buf  ( .I(\WordArray[10].Word[25].QWire ), 
        .OE(n78), .Z(DataRead[25]) );
  BUFTD1 \WordArray[10].Word[24].Buf  ( .I(\WordArray[10].Word[24].QWire ), 
        .OE(n78), .Z(DataRead[24]) );
  BUFTD1 \WordArray[10].Word[23].Buf  ( .I(\WordArray[10].Word[23].QWire ), 
        .OE(n78), .Z(DataRead[23]) );
  BUFTD1 \WordArray[10].Word[22].Buf  ( .I(\WordArray[10].Word[22].QWire ), 
        .OE(n77), .Z(DataRead[22]) );
  BUFTD1 \WordArray[10].Word[21].Buf  ( .I(\WordArray[10].Word[21].QWire ), 
        .OE(n78), .Z(DataRead[21]) );
  BUFTD1 \WordArray[10].Word[20].Buf  ( .I(\WordArray[10].Word[20].QWire ), 
        .OE(n78), .Z(DataRead[20]) );
  BUFTD1 \WordArray[10].Word[19].Buf  ( .I(\WordArray[10].Word[19].QWire ), 
        .OE(n77), .Z(DataRead[19]) );
  BUFTD1 \WordArray[10].Word[18].Buf  ( .I(\WordArray[10].Word[18].QWire ), 
        .OE(n77), .Z(DataRead[18]) );
  BUFTD1 \WordArray[10].Word[17].Buf  ( .I(\WordArray[10].Word[17].QWire ), 
        .OE(n77), .Z(DataRead[17]) );
  BUFTD1 \WordArray[10].Word[16].Buf  ( .I(\WordArray[10].Word[16].QWire ), 
        .OE(n77), .Z(DataRead[16]) );
  BUFTD1 \WordArray[10].Word[15].Buf  ( .I(\WordArray[10].Word[15].QWire ), 
        .OE(n77), .Z(DataRead[15]) );
  BUFTD1 \WordArray[10].Word[14].Buf  ( .I(\WordArray[10].Word[14].QWire ), 
        .OE(n77), .Z(DataRead[14]) );
  BUFTD1 \WordArray[10].Word[13].Buf  ( .I(\WordArray[10].Word[13].QWire ), 
        .OE(n77), .Z(DataRead[13]) );
  BUFTD1 \WordArray[10].Word[12].Buf  ( .I(\WordArray[10].Word[12].QWire ), 
        .OE(n77), .Z(DataRead[12]) );
  BUFTD1 \WordArray[10].Word[11].Buf  ( .I(\WordArray[10].Word[11].QWire ), 
        .OE(n77), .Z(DataRead[11]) );
  BUFTD1 \WordArray[10].Word[10].Buf  ( .I(\WordArray[10].Word[10].QWire ), 
        .OE(n77), .Z(DataRead[10]) );
  BUFTD1 \WordArray[10].Word[9].Buf  ( .I(\WordArray[10].Word[9].QWire ), .OE(
        n78), .Z(DataRead[9]) );
  BUFTD1 \WordArray[10].Word[8].Buf  ( .I(\WordArray[10].Word[8].QWire ), .OE(
        n78), .Z(DataRead[8]) );
  BUFTD1 \WordArray[10].Word[7].Buf  ( .I(\WordArray[10].Word[7].QWire ), .OE(
        n78), .Z(DataRead[7]) );
  BUFTD1 \WordArray[10].Word[6].Buf  ( .I(\WordArray[10].Word[6].QWire ), .OE(
        n78), .Z(DataRead[6]) );
  BUFTD1 \WordArray[10].Word[5].Buf  ( .I(\WordArray[10].Word[5].QWire ), .OE(
        n78), .Z(DataRead[5]) );
  BUFTD1 \WordArray[10].Word[4].Buf  ( .I(\WordArray[10].Word[4].QWire ), .OE(
        n77), .Z(DataRead[4]) );
  BUFTD1 \WordArray[10].Word[3].Buf  ( .I(\WordArray[10].Word[3].QWire ), .OE(
        n78), .Z(DataRead[3]) );
  BUFTD1 \WordArray[10].Word[2].Buf  ( .I(\WordArray[10].Word[2].QWire ), .OE(
        n77), .Z(DataRead[2]) );
  BUFTD1 \WordArray[10].Word[1].Buf  ( .I(\WordArray[10].Word[1].QWire ), .OE(
        n78), .Z(DataRead[1]) );
  BUFTD1 \WordArray[10].Word[0].Buf  ( .I(\WordArray[10].Word[0].QWire ), .OE(
        n77), .Z(DataRead[0]) );
  BUFTD1 \WordArray[9].Word[31].Buf  ( .I(\WordArray[9].Word[31].QWire ), .OE(
        n80), .Z(DataRead[31]) );
  BUFTD1 \WordArray[9].Word[30].Buf  ( .I(\WordArray[9].Word[30].QWire ), .OE(
        n80), .Z(DataRead[30]) );
  BUFTD1 \WordArray[9].Word[29].Buf  ( .I(\WordArray[9].Word[29].QWire ), .OE(
        n80), .Z(DataRead[29]) );
  BUFTD1 \WordArray[9].Word[28].Buf  ( .I(\WordArray[9].Word[28].QWire ), .OE(
        n79), .Z(DataRead[28]) );
  BUFTD1 \WordArray[9].Word[27].Buf  ( .I(\WordArray[9].Word[27].QWire ), .OE(
        n80), .Z(DataRead[27]) );
  BUFTD1 \WordArray[9].Word[26].Buf  ( .I(\WordArray[9].Word[26].QWire ), .OE(
        n79), .Z(DataRead[26]) );
  BUFTD1 \WordArray[9].Word[25].Buf  ( .I(\WordArray[9].Word[25].QWire ), .OE(
        n80), .Z(DataRead[25]) );
  BUFTD1 \WordArray[9].Word[24].Buf  ( .I(\WordArray[9].Word[24].QWire ), .OE(
        n80), .Z(DataRead[24]) );
  BUFTD1 \WordArray[9].Word[23].Buf  ( .I(\WordArray[9].Word[23].QWire ), .OE(
        n80), .Z(DataRead[23]) );
  BUFTD1 \WordArray[9].Word[22].Buf  ( .I(\WordArray[9].Word[22].QWire ), .OE(
        n79), .Z(DataRead[22]) );
  BUFTD1 \WordArray[9].Word[21].Buf  ( .I(\WordArray[9].Word[21].QWire ), .OE(
        n80), .Z(DataRead[21]) );
  BUFTD1 \WordArray[9].Word[20].Buf  ( .I(\WordArray[9].Word[20].QWire ), .OE(
        n80), .Z(DataRead[20]) );
  BUFTD1 \WordArray[9].Word[19].Buf  ( .I(\WordArray[9].Word[19].QWire ), .OE(
        n79), .Z(DataRead[19]) );
  BUFTD1 \WordArray[9].Word[18].Buf  ( .I(\WordArray[9].Word[18].QWire ), .OE(
        n79), .Z(DataRead[18]) );
  BUFTD1 \WordArray[9].Word[17].Buf  ( .I(\WordArray[9].Word[17].QWire ), .OE(
        n79), .Z(DataRead[17]) );
  BUFTD1 \WordArray[9].Word[16].Buf  ( .I(\WordArray[9].Word[16].QWire ), .OE(
        n79), .Z(DataRead[16]) );
  BUFTD1 \WordArray[9].Word[15].Buf  ( .I(\WordArray[9].Word[15].QWire ), .OE(
        n79), .Z(DataRead[15]) );
  BUFTD1 \WordArray[9].Word[14].Buf  ( .I(\WordArray[9].Word[14].QWire ), .OE(
        n79), .Z(DataRead[14]) );
  BUFTD1 \WordArray[9].Word[13].Buf  ( .I(\WordArray[9].Word[13].QWire ), .OE(
        n79), .Z(DataRead[13]) );
  BUFTD1 \WordArray[9].Word[12].Buf  ( .I(\WordArray[9].Word[12].QWire ), .OE(
        n79), .Z(DataRead[12]) );
  BUFTD1 \WordArray[9].Word[11].Buf  ( .I(\WordArray[9].Word[11].QWire ), .OE(
        n79), .Z(DataRead[11]) );
  BUFTD1 \WordArray[9].Word[10].Buf  ( .I(\WordArray[9].Word[10].QWire ), .OE(
        n79), .Z(DataRead[10]) );
  BUFTD1 \WordArray[9].Word[9].Buf  ( .I(\WordArray[9].Word[9].QWire ), .OE(
        n80), .Z(DataRead[9]) );
  BUFTD1 \WordArray[9].Word[8].Buf  ( .I(\WordArray[9].Word[8].QWire ), .OE(
        n80), .Z(DataRead[8]) );
  BUFTD1 \WordArray[9].Word[7].Buf  ( .I(\WordArray[9].Word[7].QWire ), .OE(
        n80), .Z(DataRead[7]) );
  BUFTD1 \WordArray[9].Word[6].Buf  ( .I(\WordArray[9].Word[6].QWire ), .OE(
        n80), .Z(DataRead[6]) );
  BUFTD1 \WordArray[9].Word[5].Buf  ( .I(\WordArray[9].Word[5].QWire ), .OE(
        n80), .Z(DataRead[5]) );
  BUFTD1 \WordArray[9].Word[4].Buf  ( .I(\WordArray[9].Word[4].QWire ), .OE(
        n79), .Z(DataRead[4]) );
  BUFTD1 \WordArray[9].Word[3].Buf  ( .I(\WordArray[9].Word[3].QWire ), .OE(
        n80), .Z(DataRead[3]) );
  BUFTD1 \WordArray[9].Word[2].Buf  ( .I(\WordArray[9].Word[2].QWire ), .OE(
        n79), .Z(DataRead[2]) );
  BUFTD1 \WordArray[9].Word[1].Buf  ( .I(\WordArray[9].Word[1].QWire ), .OE(
        n80), .Z(DataRead[1]) );
  BUFTD1 \WordArray[9].Word[0].Buf  ( .I(\WordArray[9].Word[0].QWire ), .OE(
        n79), .Z(DataRead[0]) );
  BUFTD1 \WordArray[8].Word[31].Buf  ( .I(\WordArray[8].Word[31].QWire ), .OE(
        n82), .Z(DataRead[31]) );
  BUFTD1 \WordArray[8].Word[30].Buf  ( .I(\WordArray[8].Word[30].QWire ), .OE(
        n82), .Z(DataRead[30]) );
  BUFTD1 \WordArray[8].Word[29].Buf  ( .I(\WordArray[8].Word[29].QWire ), .OE(
        n82), .Z(DataRead[29]) );
  BUFTD1 \WordArray[8].Word[28].Buf  ( .I(\WordArray[8].Word[28].QWire ), .OE(
        n81), .Z(DataRead[28]) );
  BUFTD1 \WordArray[8].Word[27].Buf  ( .I(\WordArray[8].Word[27].QWire ), .OE(
        n82), .Z(DataRead[27]) );
  BUFTD1 \WordArray[8].Word[26].Buf  ( .I(\WordArray[8].Word[26].QWire ), .OE(
        n81), .Z(DataRead[26]) );
  BUFTD1 \WordArray[8].Word[25].Buf  ( .I(\WordArray[8].Word[25].QWire ), .OE(
        n82), .Z(DataRead[25]) );
  BUFTD1 \WordArray[8].Word[24].Buf  ( .I(\WordArray[8].Word[24].QWire ), .OE(
        n82), .Z(DataRead[24]) );
  BUFTD1 \WordArray[8].Word[23].Buf  ( .I(\WordArray[8].Word[23].QWire ), .OE(
        n82), .Z(DataRead[23]) );
  BUFTD1 \WordArray[8].Word[22].Buf  ( .I(\WordArray[8].Word[22].QWire ), .OE(
        n81), .Z(DataRead[22]) );
  BUFTD1 \WordArray[8].Word[21].Buf  ( .I(\WordArray[8].Word[21].QWire ), .OE(
        n82), .Z(DataRead[21]) );
  BUFTD1 \WordArray[8].Word[20].Buf  ( .I(\WordArray[8].Word[20].QWire ), .OE(
        n82), .Z(DataRead[20]) );
  BUFTD1 \WordArray[8].Word[19].Buf  ( .I(\WordArray[8].Word[19].QWire ), .OE(
        n81), .Z(DataRead[19]) );
  BUFTD1 \WordArray[8].Word[18].Buf  ( .I(\WordArray[8].Word[18].QWire ), .OE(
        n81), .Z(DataRead[18]) );
  BUFTD1 \WordArray[8].Word[17].Buf  ( .I(\WordArray[8].Word[17].QWire ), .OE(
        n81), .Z(DataRead[17]) );
  BUFTD1 \WordArray[8].Word[16].Buf  ( .I(\WordArray[8].Word[16].QWire ), .OE(
        n81), .Z(DataRead[16]) );
  BUFTD1 \WordArray[8].Word[15].Buf  ( .I(\WordArray[8].Word[15].QWire ), .OE(
        n81), .Z(DataRead[15]) );
  BUFTD1 \WordArray[8].Word[14].Buf  ( .I(\WordArray[8].Word[14].QWire ), .OE(
        n81), .Z(DataRead[14]) );
  BUFTD1 \WordArray[8].Word[13].Buf  ( .I(\WordArray[8].Word[13].QWire ), .OE(
        n81), .Z(DataRead[13]) );
  BUFTD1 \WordArray[8].Word[12].Buf  ( .I(\WordArray[8].Word[12].QWire ), .OE(
        n81), .Z(DataRead[12]) );
  BUFTD1 \WordArray[8].Word[11].Buf  ( .I(\WordArray[8].Word[11].QWire ), .OE(
        n81), .Z(DataRead[11]) );
  BUFTD1 \WordArray[8].Word[10].Buf  ( .I(\WordArray[8].Word[10].QWire ), .OE(
        n81), .Z(DataRead[10]) );
  BUFTD1 \WordArray[8].Word[9].Buf  ( .I(\WordArray[8].Word[9].QWire ), .OE(
        n82), .Z(DataRead[9]) );
  BUFTD1 \WordArray[8].Word[8].Buf  ( .I(\WordArray[8].Word[8].QWire ), .OE(
        n82), .Z(DataRead[8]) );
  BUFTD1 \WordArray[8].Word[7].Buf  ( .I(\WordArray[8].Word[7].QWire ), .OE(
        n82), .Z(DataRead[7]) );
  BUFTD1 \WordArray[8].Word[6].Buf  ( .I(\WordArray[8].Word[6].QWire ), .OE(
        n82), .Z(DataRead[6]) );
  BUFTD1 \WordArray[8].Word[5].Buf  ( .I(\WordArray[8].Word[5].QWire ), .OE(
        n82), .Z(DataRead[5]) );
  BUFTD1 \WordArray[8].Word[4].Buf  ( .I(\WordArray[8].Word[4].QWire ), .OE(
        n81), .Z(DataRead[4]) );
  BUFTD1 \WordArray[8].Word[3].Buf  ( .I(\WordArray[8].Word[3].QWire ), .OE(
        n82), .Z(DataRead[3]) );
  BUFTD1 \WordArray[8].Word[2].Buf  ( .I(\WordArray[8].Word[2].QWire ), .OE(
        n81), .Z(DataRead[2]) );
  BUFTD1 \WordArray[8].Word[1].Buf  ( .I(\WordArray[8].Word[1].QWire ), .OE(
        n82), .Z(DataRead[1]) );
  BUFTD1 \WordArray[8].Word[0].Buf  ( .I(\WordArray[8].Word[0].QWire ), .OE(
        n81), .Z(DataRead[0]) );
  BUFTD1 \WordArray[7].Word[31].Buf  ( .I(\WordArray[7].Word[31].QWire ), .OE(
        n84), .Z(DataRead[31]) );
  BUFTD1 \WordArray[7].Word[30].Buf  ( .I(\WordArray[7].Word[30].QWire ), .OE(
        n84), .Z(DataRead[30]) );
  BUFTD1 \WordArray[7].Word[29].Buf  ( .I(\WordArray[7].Word[29].QWire ), .OE(
        n84), .Z(DataRead[29]) );
  BUFTD1 \WordArray[7].Word[28].Buf  ( .I(\WordArray[7].Word[28].QWire ), .OE(
        n83), .Z(DataRead[28]) );
  BUFTD1 \WordArray[7].Word[27].Buf  ( .I(\WordArray[7].Word[27].QWire ), .OE(
        n84), .Z(DataRead[27]) );
  BUFTD1 \WordArray[7].Word[26].Buf  ( .I(\WordArray[7].Word[26].QWire ), .OE(
        n83), .Z(DataRead[26]) );
  BUFTD1 \WordArray[7].Word[25].Buf  ( .I(\WordArray[7].Word[25].QWire ), .OE(
        n84), .Z(DataRead[25]) );
  BUFTD1 \WordArray[7].Word[24].Buf  ( .I(\WordArray[7].Word[24].QWire ), .OE(
        n84), .Z(DataRead[24]) );
  BUFTD1 \WordArray[7].Word[23].Buf  ( .I(\WordArray[7].Word[23].QWire ), .OE(
        n84), .Z(DataRead[23]) );
  BUFTD1 \WordArray[7].Word[22].Buf  ( .I(\WordArray[7].Word[22].QWire ), .OE(
        n83), .Z(DataRead[22]) );
  BUFTD1 \WordArray[7].Word[21].Buf  ( .I(\WordArray[7].Word[21].QWire ), .OE(
        n84), .Z(DataRead[21]) );
  BUFTD1 \WordArray[7].Word[20].Buf  ( .I(\WordArray[7].Word[20].QWire ), .OE(
        n84), .Z(DataRead[20]) );
  BUFTD1 \WordArray[7].Word[19].Buf  ( .I(\WordArray[7].Word[19].QWire ), .OE(
        n83), .Z(DataRead[19]) );
  BUFTD1 \WordArray[7].Word[18].Buf  ( .I(\WordArray[7].Word[18].QWire ), .OE(
        n83), .Z(DataRead[18]) );
  BUFTD1 \WordArray[7].Word[17].Buf  ( .I(\WordArray[7].Word[17].QWire ), .OE(
        n83), .Z(DataRead[17]) );
  BUFTD1 \WordArray[7].Word[16].Buf  ( .I(\WordArray[7].Word[16].QWire ), .OE(
        n83), .Z(DataRead[16]) );
  BUFTD1 \WordArray[7].Word[15].Buf  ( .I(\WordArray[7].Word[15].QWire ), .OE(
        n83), .Z(DataRead[15]) );
  BUFTD1 \WordArray[7].Word[14].Buf  ( .I(\WordArray[7].Word[14].QWire ), .OE(
        n83), .Z(DataRead[14]) );
  BUFTD1 \WordArray[7].Word[13].Buf  ( .I(\WordArray[7].Word[13].QWire ), .OE(
        n83), .Z(DataRead[13]) );
  BUFTD1 \WordArray[7].Word[12].Buf  ( .I(\WordArray[7].Word[12].QWire ), .OE(
        n83), .Z(DataRead[12]) );
  BUFTD1 \WordArray[7].Word[11].Buf  ( .I(\WordArray[7].Word[11].QWire ), .OE(
        n83), .Z(DataRead[11]) );
  BUFTD1 \WordArray[7].Word[10].Buf  ( .I(\WordArray[7].Word[10].QWire ), .OE(
        n83), .Z(DataRead[10]) );
  BUFTD1 \WordArray[7].Word[9].Buf  ( .I(\WordArray[7].Word[9].QWire ), .OE(
        n84), .Z(DataRead[9]) );
  BUFTD1 \WordArray[7].Word[8].Buf  ( .I(\WordArray[7].Word[8].QWire ), .OE(
        n84), .Z(DataRead[8]) );
  BUFTD1 \WordArray[7].Word[7].Buf  ( .I(\WordArray[7].Word[7].QWire ), .OE(
        n84), .Z(DataRead[7]) );
  BUFTD1 \WordArray[7].Word[6].Buf  ( .I(\WordArray[7].Word[6].QWire ), .OE(
        n84), .Z(DataRead[6]) );
  BUFTD1 \WordArray[7].Word[5].Buf  ( .I(\WordArray[7].Word[5].QWire ), .OE(
        n84), .Z(DataRead[5]) );
  BUFTD1 \WordArray[7].Word[4].Buf  ( .I(\WordArray[7].Word[4].QWire ), .OE(
        n83), .Z(DataRead[4]) );
  BUFTD1 \WordArray[7].Word[3].Buf  ( .I(\WordArray[7].Word[3].QWire ), .OE(
        n84), .Z(DataRead[3]) );
  BUFTD1 \WordArray[7].Word[2].Buf  ( .I(\WordArray[7].Word[2].QWire ), .OE(
        n83), .Z(DataRead[2]) );
  BUFTD1 \WordArray[7].Word[1].Buf  ( .I(\WordArray[7].Word[1].QWire ), .OE(
        n84), .Z(DataRead[1]) );
  BUFTD1 \WordArray[7].Word[0].Buf  ( .I(\WordArray[7].Word[0].QWire ), .OE(
        n83), .Z(DataRead[0]) );
  BUFTD1 \WordArray[6].Word[31].Buf  ( .I(\WordArray[6].Word[31].QWire ), .OE(
        n86), .Z(DataRead[31]) );
  BUFTD1 \WordArray[6].Word[30].Buf  ( .I(\WordArray[6].Word[30].QWire ), .OE(
        n86), .Z(DataRead[30]) );
  BUFTD1 \WordArray[6].Word[29].Buf  ( .I(\WordArray[6].Word[29].QWire ), .OE(
        n86), .Z(DataRead[29]) );
  BUFTD1 \WordArray[6].Word[28].Buf  ( .I(\WordArray[6].Word[28].QWire ), .OE(
        n85), .Z(DataRead[28]) );
  BUFTD1 \WordArray[6].Word[27].Buf  ( .I(\WordArray[6].Word[27].QWire ), .OE(
        n86), .Z(DataRead[27]) );
  BUFTD1 \WordArray[6].Word[26].Buf  ( .I(\WordArray[6].Word[26].QWire ), .OE(
        n85), .Z(DataRead[26]) );
  BUFTD1 \WordArray[6].Word[25].Buf  ( .I(\WordArray[6].Word[25].QWire ), .OE(
        n86), .Z(DataRead[25]) );
  BUFTD1 \WordArray[6].Word[24].Buf  ( .I(\WordArray[6].Word[24].QWire ), .OE(
        n86), .Z(DataRead[24]) );
  BUFTD1 \WordArray[6].Word[23].Buf  ( .I(\WordArray[6].Word[23].QWire ), .OE(
        n86), .Z(DataRead[23]) );
  BUFTD1 \WordArray[6].Word[22].Buf  ( .I(\WordArray[6].Word[22].QWire ), .OE(
        n85), .Z(DataRead[22]) );
  BUFTD1 \WordArray[6].Word[21].Buf  ( .I(\WordArray[6].Word[21].QWire ), .OE(
        n86), .Z(DataRead[21]) );
  BUFTD1 \WordArray[6].Word[20].Buf  ( .I(\WordArray[6].Word[20].QWire ), .OE(
        n86), .Z(DataRead[20]) );
  BUFTD1 \WordArray[6].Word[19].Buf  ( .I(\WordArray[6].Word[19].QWire ), .OE(
        n85), .Z(DataRead[19]) );
  BUFTD1 \WordArray[6].Word[18].Buf  ( .I(\WordArray[6].Word[18].QWire ), .OE(
        n85), .Z(DataRead[18]) );
  BUFTD1 \WordArray[6].Word[17].Buf  ( .I(\WordArray[6].Word[17].QWire ), .OE(
        n85), .Z(DataRead[17]) );
  BUFTD1 \WordArray[6].Word[16].Buf  ( .I(\WordArray[6].Word[16].QWire ), .OE(
        n85), .Z(DataRead[16]) );
  BUFTD1 \WordArray[6].Word[15].Buf  ( .I(\WordArray[6].Word[15].QWire ), .OE(
        n85), .Z(DataRead[15]) );
  BUFTD1 \WordArray[6].Word[14].Buf  ( .I(\WordArray[6].Word[14].QWire ), .OE(
        n85), .Z(DataRead[14]) );
  BUFTD1 \WordArray[6].Word[13].Buf  ( .I(\WordArray[6].Word[13].QWire ), .OE(
        n85), .Z(DataRead[13]) );
  BUFTD1 \WordArray[6].Word[12].Buf  ( .I(\WordArray[6].Word[12].QWire ), .OE(
        n85), .Z(DataRead[12]) );
  BUFTD1 \WordArray[6].Word[11].Buf  ( .I(\WordArray[6].Word[11].QWire ), .OE(
        n85), .Z(DataRead[11]) );
  BUFTD1 \WordArray[6].Word[10].Buf  ( .I(\WordArray[6].Word[10].QWire ), .OE(
        n85), .Z(DataRead[10]) );
  BUFTD1 \WordArray[6].Word[9].Buf  ( .I(\WordArray[6].Word[9].QWire ), .OE(
        n86), .Z(DataRead[9]) );
  BUFTD1 \WordArray[6].Word[8].Buf  ( .I(\WordArray[6].Word[8].QWire ), .OE(
        n86), .Z(DataRead[8]) );
  BUFTD1 \WordArray[6].Word[7].Buf  ( .I(\WordArray[6].Word[7].QWire ), .OE(
        n86), .Z(DataRead[7]) );
  BUFTD1 \WordArray[6].Word[6].Buf  ( .I(\WordArray[6].Word[6].QWire ), .OE(
        n86), .Z(DataRead[6]) );
  BUFTD1 \WordArray[6].Word[5].Buf  ( .I(\WordArray[6].Word[5].QWire ), .OE(
        n86), .Z(DataRead[5]) );
  BUFTD1 \WordArray[6].Word[4].Buf  ( .I(\WordArray[6].Word[4].QWire ), .OE(
        n85), .Z(DataRead[4]) );
  BUFTD1 \WordArray[6].Word[3].Buf  ( .I(\WordArray[6].Word[3].QWire ), .OE(
        n86), .Z(DataRead[3]) );
  BUFTD1 \WordArray[6].Word[2].Buf  ( .I(\WordArray[6].Word[2].QWire ), .OE(
        n85), .Z(DataRead[2]) );
  BUFTD1 \WordArray[6].Word[1].Buf  ( .I(\WordArray[6].Word[1].QWire ), .OE(
        n86), .Z(DataRead[1]) );
  BUFTD1 \WordArray[6].Word[0].Buf  ( .I(\WordArray[6].Word[0].QWire ), .OE(
        n85), .Z(DataRead[0]) );
  BUFTD1 \WordArray[5].Word[31].Buf  ( .I(\WordArray[5].Word[31].QWire ), .OE(
        n88), .Z(DataRead[31]) );
  BUFTD1 \WordArray[5].Word[30].Buf  ( .I(\WordArray[5].Word[30].QWire ), .OE(
        n88), .Z(DataRead[30]) );
  BUFTD1 \WordArray[5].Word[29].Buf  ( .I(\WordArray[5].Word[29].QWire ), .OE(
        n88), .Z(DataRead[29]) );
  BUFTD1 \WordArray[5].Word[28].Buf  ( .I(\WordArray[5].Word[28].QWire ), .OE(
        n87), .Z(DataRead[28]) );
  BUFTD1 \WordArray[5].Word[27].Buf  ( .I(\WordArray[5].Word[27].QWire ), .OE(
        n88), .Z(DataRead[27]) );
  BUFTD1 \WordArray[5].Word[26].Buf  ( .I(\WordArray[5].Word[26].QWire ), .OE(
        n87), .Z(DataRead[26]) );
  BUFTD1 \WordArray[5].Word[25].Buf  ( .I(\WordArray[5].Word[25].QWire ), .OE(
        n88), .Z(DataRead[25]) );
  BUFTD1 \WordArray[5].Word[24].Buf  ( .I(\WordArray[5].Word[24].QWire ), .OE(
        n88), .Z(DataRead[24]) );
  BUFTD1 \WordArray[5].Word[23].Buf  ( .I(\WordArray[5].Word[23].QWire ), .OE(
        n88), .Z(DataRead[23]) );
  BUFTD1 \WordArray[5].Word[22].Buf  ( .I(\WordArray[5].Word[22].QWire ), .OE(
        n87), .Z(DataRead[22]) );
  BUFTD1 \WordArray[5].Word[21].Buf  ( .I(\WordArray[5].Word[21].QWire ), .OE(
        n88), .Z(DataRead[21]) );
  BUFTD1 \WordArray[5].Word[20].Buf  ( .I(\WordArray[5].Word[20].QWire ), .OE(
        n88), .Z(DataRead[20]) );
  BUFTD1 \WordArray[5].Word[19].Buf  ( .I(\WordArray[5].Word[19].QWire ), .OE(
        n87), .Z(DataRead[19]) );
  BUFTD1 \WordArray[5].Word[18].Buf  ( .I(\WordArray[5].Word[18].QWire ), .OE(
        n87), .Z(DataRead[18]) );
  BUFTD1 \WordArray[5].Word[17].Buf  ( .I(\WordArray[5].Word[17].QWire ), .OE(
        n87), .Z(DataRead[17]) );
  BUFTD1 \WordArray[5].Word[16].Buf  ( .I(\WordArray[5].Word[16].QWire ), .OE(
        n87), .Z(DataRead[16]) );
  BUFTD1 \WordArray[5].Word[15].Buf  ( .I(\WordArray[5].Word[15].QWire ), .OE(
        n87), .Z(DataRead[15]) );
  BUFTD1 \WordArray[5].Word[14].Buf  ( .I(\WordArray[5].Word[14].QWire ), .OE(
        n87), .Z(DataRead[14]) );
  BUFTD1 \WordArray[5].Word[13].Buf  ( .I(\WordArray[5].Word[13].QWire ), .OE(
        n87), .Z(DataRead[13]) );
  BUFTD1 \WordArray[5].Word[12].Buf  ( .I(\WordArray[5].Word[12].QWire ), .OE(
        n87), .Z(DataRead[12]) );
  BUFTD1 \WordArray[5].Word[11].Buf  ( .I(\WordArray[5].Word[11].QWire ), .OE(
        n87), .Z(DataRead[11]) );
  BUFTD1 \WordArray[5].Word[10].Buf  ( .I(\WordArray[5].Word[10].QWire ), .OE(
        n87), .Z(DataRead[10]) );
  BUFTD1 \WordArray[5].Word[9].Buf  ( .I(\WordArray[5].Word[9].QWire ), .OE(
        n88), .Z(DataRead[9]) );
  BUFTD1 \WordArray[5].Word[8].Buf  ( .I(\WordArray[5].Word[8].QWire ), .OE(
        n88), .Z(DataRead[8]) );
  BUFTD1 \WordArray[5].Word[7].Buf  ( .I(\WordArray[5].Word[7].QWire ), .OE(
        n88), .Z(DataRead[7]) );
  BUFTD1 \WordArray[5].Word[6].Buf  ( .I(\WordArray[5].Word[6].QWire ), .OE(
        n88), .Z(DataRead[6]) );
  BUFTD1 \WordArray[5].Word[5].Buf  ( .I(\WordArray[5].Word[5].QWire ), .OE(
        n88), .Z(DataRead[5]) );
  BUFTD1 \WordArray[5].Word[4].Buf  ( .I(\WordArray[5].Word[4].QWire ), .OE(
        n87), .Z(DataRead[4]) );
  BUFTD1 \WordArray[5].Word[3].Buf  ( .I(\WordArray[5].Word[3].QWire ), .OE(
        n88), .Z(DataRead[3]) );
  BUFTD1 \WordArray[5].Word[2].Buf  ( .I(\WordArray[5].Word[2].QWire ), .OE(
        n87), .Z(DataRead[2]) );
  BUFTD1 \WordArray[5].Word[1].Buf  ( .I(\WordArray[5].Word[1].QWire ), .OE(
        n88), .Z(DataRead[1]) );
  BUFTD1 \WordArray[5].Word[0].Buf  ( .I(\WordArray[5].Word[0].QWire ), .OE(
        n87), .Z(DataRead[0]) );
  BUFTD1 \WordArray[4].Word[31].Buf  ( .I(\WordArray[4].Word[31].QWire ), .OE(
        n90), .Z(DataRead[31]) );
  BUFTD1 \WordArray[4].Word[30].Buf  ( .I(\WordArray[4].Word[30].QWire ), .OE(
        n90), .Z(DataRead[30]) );
  BUFTD1 \WordArray[4].Word[29].Buf  ( .I(\WordArray[4].Word[29].QWire ), .OE(
        n90), .Z(DataRead[29]) );
  BUFTD1 \WordArray[4].Word[28].Buf  ( .I(\WordArray[4].Word[28].QWire ), .OE(
        n89), .Z(DataRead[28]) );
  BUFTD1 \WordArray[4].Word[27].Buf  ( .I(\WordArray[4].Word[27].QWire ), .OE(
        n90), .Z(DataRead[27]) );
  BUFTD1 \WordArray[4].Word[26].Buf  ( .I(\WordArray[4].Word[26].QWire ), .OE(
        n89), .Z(DataRead[26]) );
  BUFTD1 \WordArray[4].Word[25].Buf  ( .I(\WordArray[4].Word[25].QWire ), .OE(
        n90), .Z(DataRead[25]) );
  BUFTD1 \WordArray[4].Word[24].Buf  ( .I(\WordArray[4].Word[24].QWire ), .OE(
        n90), .Z(DataRead[24]) );
  BUFTD1 \WordArray[4].Word[23].Buf  ( .I(\WordArray[4].Word[23].QWire ), .OE(
        n90), .Z(DataRead[23]) );
  BUFTD1 \WordArray[4].Word[22].Buf  ( .I(\WordArray[4].Word[22].QWire ), .OE(
        n89), .Z(DataRead[22]) );
  BUFTD1 \WordArray[4].Word[21].Buf  ( .I(\WordArray[4].Word[21].QWire ), .OE(
        n90), .Z(DataRead[21]) );
  BUFTD1 \WordArray[4].Word[20].Buf  ( .I(\WordArray[4].Word[20].QWire ), .OE(
        n90), .Z(DataRead[20]) );
  BUFTD1 \WordArray[4].Word[19].Buf  ( .I(\WordArray[4].Word[19].QWire ), .OE(
        n89), .Z(DataRead[19]) );
  BUFTD1 \WordArray[4].Word[18].Buf  ( .I(\WordArray[4].Word[18].QWire ), .OE(
        n89), .Z(DataRead[18]) );
  BUFTD1 \WordArray[4].Word[17].Buf  ( .I(\WordArray[4].Word[17].QWire ), .OE(
        n89), .Z(DataRead[17]) );
  BUFTD1 \WordArray[4].Word[16].Buf  ( .I(\WordArray[4].Word[16].QWire ), .OE(
        n89), .Z(DataRead[16]) );
  BUFTD1 \WordArray[4].Word[15].Buf  ( .I(\WordArray[4].Word[15].QWire ), .OE(
        n89), .Z(DataRead[15]) );
  BUFTD1 \WordArray[4].Word[14].Buf  ( .I(\WordArray[4].Word[14].QWire ), .OE(
        n89), .Z(DataRead[14]) );
  BUFTD1 \WordArray[4].Word[13].Buf  ( .I(\WordArray[4].Word[13].QWire ), .OE(
        n89), .Z(DataRead[13]) );
  BUFTD1 \WordArray[4].Word[12].Buf  ( .I(\WordArray[4].Word[12].QWire ), .OE(
        n89), .Z(DataRead[12]) );
  BUFTD1 \WordArray[4].Word[11].Buf  ( .I(\WordArray[4].Word[11].QWire ), .OE(
        n89), .Z(DataRead[11]) );
  BUFTD1 \WordArray[4].Word[10].Buf  ( .I(\WordArray[4].Word[10].QWire ), .OE(
        n89), .Z(DataRead[10]) );
  BUFTD1 \WordArray[4].Word[9].Buf  ( .I(\WordArray[4].Word[9].QWire ), .OE(
        n90), .Z(DataRead[9]) );
  BUFTD1 \WordArray[4].Word[8].Buf  ( .I(\WordArray[4].Word[8].QWire ), .OE(
        n90), .Z(DataRead[8]) );
  BUFTD1 \WordArray[4].Word[7].Buf  ( .I(\WordArray[4].Word[7].QWire ), .OE(
        n90), .Z(DataRead[7]) );
  BUFTD1 \WordArray[4].Word[6].Buf  ( .I(\WordArray[4].Word[6].QWire ), .OE(
        n90), .Z(DataRead[6]) );
  BUFTD1 \WordArray[4].Word[5].Buf  ( .I(\WordArray[4].Word[5].QWire ), .OE(
        n90), .Z(DataRead[5]) );
  BUFTD1 \WordArray[4].Word[4].Buf  ( .I(\WordArray[4].Word[4].QWire ), .OE(
        n89), .Z(DataRead[4]) );
  BUFTD1 \WordArray[4].Word[3].Buf  ( .I(\WordArray[4].Word[3].QWire ), .OE(
        n90), .Z(DataRead[3]) );
  BUFTD1 \WordArray[4].Word[2].Buf  ( .I(\WordArray[4].Word[2].QWire ), .OE(
        n89), .Z(DataRead[2]) );
  BUFTD1 \WordArray[4].Word[1].Buf  ( .I(\WordArray[4].Word[1].QWire ), .OE(
        n90), .Z(DataRead[1]) );
  BUFTD1 \WordArray[4].Word[0].Buf  ( .I(\WordArray[4].Word[0].QWire ), .OE(
        n89), .Z(DataRead[0]) );
  BUFTD1 \WordArray[3].Word[31].Buf  ( .I(\WordArray[3].Word[31].QWire ), .OE(
        n92), .Z(DataRead[31]) );
  BUFTD1 \WordArray[3].Word[30].Buf  ( .I(\WordArray[3].Word[30].QWire ), .OE(
        n92), .Z(DataRead[30]) );
  BUFTD1 \WordArray[3].Word[29].Buf  ( .I(\WordArray[3].Word[29].QWire ), .OE(
        n92), .Z(DataRead[29]) );
  BUFTD1 \WordArray[3].Word[28].Buf  ( .I(\WordArray[3].Word[28].QWire ), .OE(
        n91), .Z(DataRead[28]) );
  BUFTD1 \WordArray[3].Word[27].Buf  ( .I(\WordArray[3].Word[27].QWire ), .OE(
        n92), .Z(DataRead[27]) );
  BUFTD1 \WordArray[3].Word[26].Buf  ( .I(\WordArray[3].Word[26].QWire ), .OE(
        n91), .Z(DataRead[26]) );
  BUFTD1 \WordArray[3].Word[25].Buf  ( .I(\WordArray[3].Word[25].QWire ), .OE(
        n92), .Z(DataRead[25]) );
  BUFTD1 \WordArray[3].Word[24].Buf  ( .I(\WordArray[3].Word[24].QWire ), .OE(
        n92), .Z(DataRead[24]) );
  BUFTD1 \WordArray[3].Word[23].Buf  ( .I(\WordArray[3].Word[23].QWire ), .OE(
        n92), .Z(DataRead[23]) );
  BUFTD1 \WordArray[3].Word[22].Buf  ( .I(\WordArray[3].Word[22].QWire ), .OE(
        n91), .Z(DataRead[22]) );
  BUFTD1 \WordArray[3].Word[21].Buf  ( .I(\WordArray[3].Word[21].QWire ), .OE(
        n92), .Z(DataRead[21]) );
  BUFTD1 \WordArray[3].Word[20].Buf  ( .I(\WordArray[3].Word[20].QWire ), .OE(
        n92), .Z(DataRead[20]) );
  BUFTD1 \WordArray[3].Word[19].Buf  ( .I(\WordArray[3].Word[19].QWire ), .OE(
        n91), .Z(DataRead[19]) );
  BUFTD1 \WordArray[3].Word[18].Buf  ( .I(\WordArray[3].Word[18].QWire ), .OE(
        n91), .Z(DataRead[18]) );
  BUFTD1 \WordArray[3].Word[17].Buf  ( .I(\WordArray[3].Word[17].QWire ), .OE(
        n91), .Z(DataRead[17]) );
  BUFTD1 \WordArray[3].Word[16].Buf  ( .I(\WordArray[3].Word[16].QWire ), .OE(
        n91), .Z(DataRead[16]) );
  BUFTD1 \WordArray[3].Word[15].Buf  ( .I(\WordArray[3].Word[15].QWire ), .OE(
        n91), .Z(DataRead[15]) );
  BUFTD1 \WordArray[3].Word[14].Buf  ( .I(\WordArray[3].Word[14].QWire ), .OE(
        n91), .Z(DataRead[14]) );
  BUFTD1 \WordArray[3].Word[13].Buf  ( .I(\WordArray[3].Word[13].QWire ), .OE(
        n91), .Z(DataRead[13]) );
  BUFTD1 \WordArray[3].Word[12].Buf  ( .I(\WordArray[3].Word[12].QWire ), .OE(
        n91), .Z(DataRead[12]) );
  BUFTD1 \WordArray[3].Word[11].Buf  ( .I(\WordArray[3].Word[11].QWire ), .OE(
        n91), .Z(DataRead[11]) );
  BUFTD1 \WordArray[3].Word[10].Buf  ( .I(\WordArray[3].Word[10].QWire ), .OE(
        n91), .Z(DataRead[10]) );
  BUFTD1 \WordArray[3].Word[9].Buf  ( .I(\WordArray[3].Word[9].QWire ), .OE(
        n92), .Z(DataRead[9]) );
  BUFTD1 \WordArray[3].Word[8].Buf  ( .I(\WordArray[3].Word[8].QWire ), .OE(
        n92), .Z(DataRead[8]) );
  BUFTD1 \WordArray[3].Word[7].Buf  ( .I(\WordArray[3].Word[7].QWire ), .OE(
        n92), .Z(DataRead[7]) );
  BUFTD1 \WordArray[3].Word[6].Buf  ( .I(\WordArray[3].Word[6].QWire ), .OE(
        n92), .Z(DataRead[6]) );
  BUFTD1 \WordArray[3].Word[5].Buf  ( .I(\WordArray[3].Word[5].QWire ), .OE(
        n92), .Z(DataRead[5]) );
  BUFTD1 \WordArray[3].Word[4].Buf  ( .I(\WordArray[3].Word[4].QWire ), .OE(
        n91), .Z(DataRead[4]) );
  BUFTD1 \WordArray[3].Word[3].Buf  ( .I(\WordArray[3].Word[3].QWire ), .OE(
        n92), .Z(DataRead[3]) );
  BUFTD1 \WordArray[3].Word[2].Buf  ( .I(\WordArray[3].Word[2].QWire ), .OE(
        n91), .Z(DataRead[2]) );
  BUFTD1 \WordArray[3].Word[1].Buf  ( .I(\WordArray[3].Word[1].QWire ), .OE(
        n92), .Z(DataRead[1]) );
  BUFTD1 \WordArray[3].Word[0].Buf  ( .I(\WordArray[3].Word[0].QWire ), .OE(
        n91), .Z(DataRead[0]) );
  BUFTD1 \WordArray[2].Word[31].Buf  ( .I(\WordArray[2].Word[31].QWire ), .OE(
        n94), .Z(DataRead[31]) );
  BUFTD1 \WordArray[2].Word[30].Buf  ( .I(\WordArray[2].Word[30].QWire ), .OE(
        n94), .Z(DataRead[30]) );
  BUFTD1 \WordArray[2].Word[29].Buf  ( .I(\WordArray[2].Word[29].QWire ), .OE(
        n94), .Z(DataRead[29]) );
  BUFTD1 \WordArray[2].Word[28].Buf  ( .I(\WordArray[2].Word[28].QWire ), .OE(
        n93), .Z(DataRead[28]) );
  BUFTD1 \WordArray[2].Word[27].Buf  ( .I(\WordArray[2].Word[27].QWire ), .OE(
        n94), .Z(DataRead[27]) );
  BUFTD1 \WordArray[2].Word[26].Buf  ( .I(\WordArray[2].Word[26].QWire ), .OE(
        n93), .Z(DataRead[26]) );
  BUFTD1 \WordArray[2].Word[25].Buf  ( .I(\WordArray[2].Word[25].QWire ), .OE(
        n94), .Z(DataRead[25]) );
  BUFTD1 \WordArray[2].Word[24].Buf  ( .I(\WordArray[2].Word[24].QWire ), .OE(
        n94), .Z(DataRead[24]) );
  BUFTD1 \WordArray[2].Word[23].Buf  ( .I(\WordArray[2].Word[23].QWire ), .OE(
        n94), .Z(DataRead[23]) );
  BUFTD1 \WordArray[2].Word[22].Buf  ( .I(\WordArray[2].Word[22].QWire ), .OE(
        n93), .Z(DataRead[22]) );
  BUFTD1 \WordArray[2].Word[21].Buf  ( .I(\WordArray[2].Word[21].QWire ), .OE(
        n94), .Z(DataRead[21]) );
  BUFTD1 \WordArray[2].Word[20].Buf  ( .I(\WordArray[2].Word[20].QWire ), .OE(
        n94), .Z(DataRead[20]) );
  BUFTD1 \WordArray[2].Word[19].Buf  ( .I(\WordArray[2].Word[19].QWire ), .OE(
        n93), .Z(DataRead[19]) );
  BUFTD1 \WordArray[2].Word[18].Buf  ( .I(\WordArray[2].Word[18].QWire ), .OE(
        n93), .Z(DataRead[18]) );
  BUFTD1 \WordArray[2].Word[17].Buf  ( .I(\WordArray[2].Word[17].QWire ), .OE(
        n93), .Z(DataRead[17]) );
  BUFTD1 \WordArray[2].Word[16].Buf  ( .I(\WordArray[2].Word[16].QWire ), .OE(
        n93), .Z(DataRead[16]) );
  BUFTD1 \WordArray[2].Word[15].Buf  ( .I(\WordArray[2].Word[15].QWire ), .OE(
        n93), .Z(DataRead[15]) );
  BUFTD1 \WordArray[2].Word[14].Buf  ( .I(\WordArray[2].Word[14].QWire ), .OE(
        n93), .Z(DataRead[14]) );
  BUFTD1 \WordArray[2].Word[13].Buf  ( .I(\WordArray[2].Word[13].QWire ), .OE(
        n93), .Z(DataRead[13]) );
  BUFTD1 \WordArray[2].Word[12].Buf  ( .I(\WordArray[2].Word[12].QWire ), .OE(
        n93), .Z(DataRead[12]) );
  BUFTD1 \WordArray[2].Word[11].Buf  ( .I(\WordArray[2].Word[11].QWire ), .OE(
        n93), .Z(DataRead[11]) );
  BUFTD1 \WordArray[2].Word[10].Buf  ( .I(\WordArray[2].Word[10].QWire ), .OE(
        n93), .Z(DataRead[10]) );
  BUFTD1 \WordArray[2].Word[9].Buf  ( .I(\WordArray[2].Word[9].QWire ), .OE(
        n94), .Z(DataRead[9]) );
  BUFTD1 \WordArray[2].Word[8].Buf  ( .I(\WordArray[2].Word[8].QWire ), .OE(
        n94), .Z(DataRead[8]) );
  BUFTD1 \WordArray[2].Word[7].Buf  ( .I(\WordArray[2].Word[7].QWire ), .OE(
        n94), .Z(DataRead[7]) );
  BUFTD1 \WordArray[2].Word[6].Buf  ( .I(\WordArray[2].Word[6].QWire ), .OE(
        n94), .Z(DataRead[6]) );
  BUFTD1 \WordArray[2].Word[5].Buf  ( .I(\WordArray[2].Word[5].QWire ), .OE(
        n94), .Z(DataRead[5]) );
  BUFTD1 \WordArray[2].Word[4].Buf  ( .I(\WordArray[2].Word[4].QWire ), .OE(
        n93), .Z(DataRead[4]) );
  BUFTD1 \WordArray[2].Word[3].Buf  ( .I(\WordArray[2].Word[3].QWire ), .OE(
        n94), .Z(DataRead[3]) );
  BUFTD1 \WordArray[2].Word[2].Buf  ( .I(\WordArray[2].Word[2].QWire ), .OE(
        n93), .Z(DataRead[2]) );
  BUFTD1 \WordArray[2].Word[1].Buf  ( .I(\WordArray[2].Word[1].QWire ), .OE(
        n94), .Z(DataRead[1]) );
  BUFTD1 \WordArray[2].Word[0].Buf  ( .I(\WordArray[2].Word[0].QWire ), .OE(
        n93), .Z(DataRead[0]) );
  BUFTD1 \WordArray[1].Word[31].Buf  ( .I(\WordArray[1].Word[31].QWire ), .OE(
        n96), .Z(DataRead[31]) );
  BUFTD1 \WordArray[1].Word[30].Buf  ( .I(\WordArray[1].Word[30].QWire ), .OE(
        n96), .Z(DataRead[30]) );
  BUFTD1 \WordArray[1].Word[29].Buf  ( .I(\WordArray[1].Word[29].QWire ), .OE(
        n96), .Z(DataRead[29]) );
  BUFTD1 \WordArray[1].Word[28].Buf  ( .I(\WordArray[1].Word[28].QWire ), .OE(
        n95), .Z(DataRead[28]) );
  BUFTD1 \WordArray[1].Word[27].Buf  ( .I(\WordArray[1].Word[27].QWire ), .OE(
        n96), .Z(DataRead[27]) );
  BUFTD1 \WordArray[1].Word[26].Buf  ( .I(\WordArray[1].Word[26].QWire ), .OE(
        n95), .Z(DataRead[26]) );
  BUFTD1 \WordArray[1].Word[25].Buf  ( .I(\WordArray[1].Word[25].QWire ), .OE(
        n96), .Z(DataRead[25]) );
  BUFTD1 \WordArray[1].Word[24].Buf  ( .I(\WordArray[1].Word[24].QWire ), .OE(
        n96), .Z(DataRead[24]) );
  BUFTD1 \WordArray[1].Word[23].Buf  ( .I(\WordArray[1].Word[23].QWire ), .OE(
        n96), .Z(DataRead[23]) );
  BUFTD1 \WordArray[1].Word[22].Buf  ( .I(\WordArray[1].Word[22].QWire ), .OE(
        n95), .Z(DataRead[22]) );
  BUFTD1 \WordArray[1].Word[21].Buf  ( .I(\WordArray[1].Word[21].QWire ), .OE(
        n96), .Z(DataRead[21]) );
  BUFTD1 \WordArray[1].Word[20].Buf  ( .I(\WordArray[1].Word[20].QWire ), .OE(
        n96), .Z(DataRead[20]) );
  BUFTD1 \WordArray[1].Word[19].Buf  ( .I(\WordArray[1].Word[19].QWire ), .OE(
        n95), .Z(DataRead[19]) );
  BUFTD1 \WordArray[1].Word[18].Buf  ( .I(\WordArray[1].Word[18].QWire ), .OE(
        n95), .Z(DataRead[18]) );
  BUFTD1 \WordArray[1].Word[17].Buf  ( .I(\WordArray[1].Word[17].QWire ), .OE(
        n95), .Z(DataRead[17]) );
  BUFTD1 \WordArray[1].Word[16].Buf  ( .I(\WordArray[1].Word[16].QWire ), .OE(
        n95), .Z(DataRead[16]) );
  BUFTD1 \WordArray[1].Word[15].Buf  ( .I(\WordArray[1].Word[15].QWire ), .OE(
        n95), .Z(DataRead[15]) );
  BUFTD1 \WordArray[1].Word[14].Buf  ( .I(\WordArray[1].Word[14].QWire ), .OE(
        n95), .Z(DataRead[14]) );
  BUFTD1 \WordArray[1].Word[13].Buf  ( .I(\WordArray[1].Word[13].QWire ), .OE(
        n95), .Z(DataRead[13]) );
  BUFTD1 \WordArray[1].Word[12].Buf  ( .I(\WordArray[1].Word[12].QWire ), .OE(
        n95), .Z(DataRead[12]) );
  BUFTD1 \WordArray[1].Word[11].Buf  ( .I(\WordArray[1].Word[11].QWire ), .OE(
        n95), .Z(DataRead[11]) );
  BUFTD1 \WordArray[1].Word[10].Buf  ( .I(\WordArray[1].Word[10].QWire ), .OE(
        n95), .Z(DataRead[10]) );
  BUFTD1 \WordArray[1].Word[9].Buf  ( .I(\WordArray[1].Word[9].QWire ), .OE(
        n96), .Z(DataRead[9]) );
  BUFTD1 \WordArray[1].Word[8].Buf  ( .I(\WordArray[1].Word[8].QWire ), .OE(
        n96), .Z(DataRead[8]) );
  BUFTD1 \WordArray[1].Word[7].Buf  ( .I(\WordArray[1].Word[7].QWire ), .OE(
        n96), .Z(DataRead[7]) );
  BUFTD1 \WordArray[1].Word[6].Buf  ( .I(\WordArray[1].Word[6].QWire ), .OE(
        n96), .Z(DataRead[6]) );
  BUFTD1 \WordArray[1].Word[5].Buf  ( .I(\WordArray[1].Word[5].QWire ), .OE(
        n96), .Z(DataRead[5]) );
  BUFTD1 \WordArray[1].Word[4].Buf  ( .I(\WordArray[1].Word[4].QWire ), .OE(
        n95), .Z(DataRead[4]) );
  BUFTD1 \WordArray[1].Word[3].Buf  ( .I(\WordArray[1].Word[3].QWire ), .OE(
        n96), .Z(DataRead[3]) );
  BUFTD1 \WordArray[1].Word[2].Buf  ( .I(\WordArray[1].Word[2].QWire ), .OE(
        n95), .Z(DataRead[2]) );
  BUFTD1 \WordArray[1].Word[1].Buf  ( .I(\WordArray[1].Word[1].QWire ), .OE(
        n96), .Z(DataRead[1]) );
  BUFTD1 \WordArray[1].Word[0].Buf  ( .I(\WordArray[1].Word[0].QWire ), .OE(
        n95), .Z(DataRead[0]) );
  BUFTD1 \WordArray[0].Word[31].Buf  ( .I(\WordArray[0].Word[31].QWire ), .OE(
        n97), .Z(DataRead[31]) );
  BUFTD1 \WordArray[0].Word[30].Buf  ( .I(\WordArray[0].Word[30].QWire ), .OE(
        n98), .Z(DataRead[30]) );
  BUFTD1 \WordArray[0].Word[29].Buf  ( .I(\WordArray[0].Word[29].QWire ), .OE(
        n97), .Z(DataRead[29]) );
  BUFTD1 \WordArray[0].Word[28].Buf  ( .I(\WordArray[0].Word[28].QWire ), .OE(
        n97), .Z(DataRead[28]) );
  BUFTD1 \WordArray[0].Word[27].Buf  ( .I(\WordArray[0].Word[27].QWire ), .OE(
        n97), .Z(DataRead[27]) );
  BUFTD1 \WordArray[0].Word[26].Buf  ( .I(\WordArray[0].Word[26].QWire ), .OE(
        n97), .Z(DataRead[26]) );
  BUFTD1 \WordArray[0].Word[25].Buf  ( .I(\WordArray[0].Word[25].QWire ), .OE(
        n97), .Z(DataRead[25]) );
  BUFTD1 \WordArray[0].Word[24].Buf  ( .I(\WordArray[0].Word[24].QWire ), .OE(
        n97), .Z(DataRead[24]) );
  BUFTD1 \WordArray[0].Word[23].Buf  ( .I(\WordArray[0].Word[23].QWire ), .OE(
        n97), .Z(DataRead[23]) );
  BUFTD1 \WordArray[0].Word[22].Buf  ( .I(\WordArray[0].Word[22].QWire ), .OE(
        n97), .Z(DataRead[22]) );
  BUFTD1 \WordArray[0].Word[21].Buf  ( .I(\WordArray[0].Word[21].QWire ), .OE(
        n98), .Z(DataRead[21]) );
  BUFTD1 \WordArray[0].Word[20].Buf  ( .I(\WordArray[0].Word[20].QWire ), .OE(
        n97), .Z(DataRead[20]) );
  BUFTD1 \WordArray[0].Word[19].Buf  ( .I(\WordArray[0].Word[19].QWire ), .OE(
        n97), .Z(DataRead[19]) );
  BUFTD1 \WordArray[0].Word[18].Buf  ( .I(\WordArray[0].Word[18].QWire ), .OE(
        n98), .Z(DataRead[18]) );
  BUFTD1 \WordArray[0].Word[17].Buf  ( .I(\WordArray[0].Word[17].QWire ), .OE(
        n98), .Z(DataRead[17]) );
  BUFTD1 \WordArray[0].Word[16].Buf  ( .I(\WordArray[0].Word[16].QWire ), .OE(
        n98), .Z(DataRead[16]) );
  BUFTD1 \WordArray[0].Word[15].Buf  ( .I(\WordArray[0].Word[15].QWire ), .OE(
        n98), .Z(DataRead[15]) );
  BUFTD1 \WordArray[0].Word[14].Buf  ( .I(\WordArray[0].Word[14].QWire ), .OE(
        n98), .Z(DataRead[14]) );
  BUFTD1 \WordArray[0].Word[13].Buf  ( .I(\WordArray[0].Word[13].QWire ), .OE(
        n98), .Z(DataRead[13]) );
  BUFTD1 \WordArray[0].Word[12].Buf  ( .I(\WordArray[0].Word[12].QWire ), .OE(
        n98), .Z(DataRead[12]) );
  BUFTD1 \WordArray[0].Word[11].Buf  ( .I(\WordArray[0].Word[11].QWire ), .OE(
        n98), .Z(DataRead[11]) );
  BUFTD1 \WordArray[0].Word[10].Buf  ( .I(\WordArray[0].Word[10].QWire ), .OE(
        n98), .Z(DataRead[10]) );
  BUFTD1 \WordArray[0].Word[9].Buf  ( .I(\WordArray[0].Word[9].QWire ), .OE(
        n97), .Z(DataRead[9]) );
  BUFTD1 \WordArray[0].Word[8].Buf  ( .I(\WordArray[0].Word[8].QWire ), .OE(
        n97), .Z(DataRead[8]) );
  BUFTD1 \WordArray[0].Word[7].Buf  ( .I(\WordArray[0].Word[7].QWire ), .OE(
        n98), .Z(DataRead[7]) );
  BUFTD1 \WordArray[0].Word[6].Buf  ( .I(\WordArray[0].Word[6].QWire ), .OE(
        n97), .Z(DataRead[6]) );
  BUFTD1 \WordArray[0].Word[5].Buf  ( .I(\WordArray[0].Word[5].QWire ), .OE(
        n98), .Z(DataRead[5]) );
  BUFTD1 \WordArray[0].Word[4].Buf  ( .I(\WordArray[0].Word[4].QWire ), .OE(
        n97), .Z(DataRead[4]) );
  BUFTD1 \WordArray[0].Word[3].Buf  ( .I(\WordArray[0].Word[3].QWire ), .OE(
        n98), .Z(DataRead[3]) );
  BUFTD1 \WordArray[0].Word[2].Buf  ( .I(\WordArray[0].Word[2].QWire ), .OE(
        n97), .Z(DataRead[2]) );
  BUFTD1 \WordArray[0].Word[1].Buf  ( .I(\WordArray[0].Word[1].QWire ), .OE(
        n98), .Z(DataRead[1]) );
  BUFTD1 \WordArray[0].Word[0].Buf  ( .I(\WordArray[0].Word[0].QWire ), .OE(
        n98), .Z(DataRead[0]) );
  BUFTD1 \DataO_tri[0]  ( .I(DataRead[0]), .OE(n101), .Z(DataO[0]) );
  BUFTD1 \DataO_tri[1]  ( .I(DataRead[1]), .OE(n101), .Z(DataO[1]) );
  BUFTD1 \DataO_tri[2]  ( .I(DataRead[2]), .OE(n102), .Z(DataO[2]) );
  BUFTD1 \DataO_tri[3]  ( .I(DataRead[3]), .OE(n102), .Z(DataO[3]) );
  BUFTD1 \DataO_tri[4]  ( .I(DataRead[4]), .OE(n102), .Z(DataO[4]) );
  BUFTD1 \DataO_tri[5]  ( .I(DataRead[5]), .OE(n102), .Z(DataO[5]) );
  BUFTD1 \DataO_tri[6]  ( .I(DataRead[6]), .OE(n102), .Z(DataO[6]) );
  BUFTD1 \DataO_tri[7]  ( .I(DataRead[7]), .OE(n102), .Z(DataO[7]) );
  BUFTD1 \DataO_tri[8]  ( .I(DataRead[8]), .OE(n102), .Z(DataO[8]) );
  BUFTD1 \DataO_tri[9]  ( .I(DataRead[9]), .OE(n102), .Z(DataO[9]) );
  BUFTD1 \DataO_tri[10]  ( .I(DataRead[10]), .OE(n101), .Z(DataO[10]) );
  BUFTD1 \DataO_tri[11]  ( .I(DataRead[11]), .OE(n101), .Z(DataO[11]) );
  BUFTD1 \DataO_tri[12]  ( .I(DataRead[12]), .OE(n101), .Z(DataO[12]) );
  BUFTD1 \DataO_tri[13]  ( .I(DataRead[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD1 \DataO_tri[14]  ( .I(DataRead[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD1 \DataO_tri[15]  ( .I(DataRead[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD1 \DataO_tri[16]  ( .I(DataRead[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD1 \DataO_tri[17]  ( .I(DataRead[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD1 \DataO_tri[18]  ( .I(DataRead[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD1 \DataO_tri[19]  ( .I(DataRead[19]), .OE(n101), .Z(DataO[19]) );
  BUFTD1 \DataO_tri[20]  ( .I(DataRead[20]), .OE(n101), .Z(DataO[20]) );
  BUFTD1 \DataO_tri[21]  ( .I(DataRead[21]), .OE(n101), .Z(DataO[21]) );
  BUFTD1 \DataO_tri[22]  ( .I(DataRead[22]), .OE(n101), .Z(DataO[22]) );
  BUFTD1 \DataO_tri[23]  ( .I(DataRead[23]), .OE(n101), .Z(DataO[23]) );
  BUFTD1 \DataO_tri[24]  ( .I(DataRead[24]), .OE(n101), .Z(DataO[24]) );
  BUFTD1 \DataO_tri[25]  ( .I(DataRead[25]), .OE(n101), .Z(DataO[25]) );
  BUFTD1 \DataO_tri[26]  ( .I(DataRead[26]), .OE(n101), .Z(DataO[26]) );
  BUFTD1 \DataO_tri[27]  ( .I(DataRead[27]), .OE(n101), .Z(DataO[27]) );
  BUFTD1 \DataO_tri[28]  ( .I(DataRead[28]), .OE(n101), .Z(DataO[28]) );
  BUFTD1 \DataO_tri[29]  ( .I(DataRead[29]), .OE(n101), .Z(DataO[29]) );
  BUFTD1 \DataO_tri[30]  ( .I(DataRead[30]), .OE(n102), .Z(DataO[30]) );
  BUFTD1 \DataO_tri[31]  ( .I(DataRead[31]), .OE(n102), .Z(DataO[31]) );
  XNR4D1 U43 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n2126) );
  XOR4D1 U44 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n2125) );
  XOR4D1 U45 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n2122) );
  XOR4D1 U46 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n2119) );
  XNR4D1 U47 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n2116) );
  XOR4D1 U49 ( .A1(n2129), .A2(DataRead[12]), .A3(n2130), .A4(DataRead[11]), 
        .Z(n2128) );
  XOR4D1 U50 ( .A1(DataRead[23]), .A2(DataRead[22]), .A3(DataRead[13]), .A4(
        DataRead[21]), .Z(n2130) );
  XOR4D1 U51 ( .A1(n2131), .A2(n2132), .A3(n2133), .A4(n2134), .Z(n2129) );
  XOR4D1 U52 ( .A1(n2135), .A2(n2136), .A3(DataRead[10]), .A4(DataRead[14]), 
        .Z(n2134) );
  XOR4D1 U53 ( .A1(DataRead[1]), .A2(DataRead[0]), .A3(DataRead[3]), .A4(
        DataRead[2]), .Z(n2136) );
  XOR4D1 U54 ( .A1(DataRead[5]), .A2(DataRead[4]), .A3(DataRead[7]), .A4(
        DataRead[6]), .Z(n2135) );
  XOR4D1 U57 ( .A1(n2137), .A2(n2138), .A3(DataRead[16]), .A4(DataRead[17]), 
        .Z(n2131) );
  XOR4D1 U58 ( .A1(DataRead[25]), .A2(DataRead[24]), .A3(DataRead[27]), .A4(
        DataRead[26]), .Z(n2138) );
  XOR4D1 U59 ( .A1(DataRead[29]), .A2(DataRead[28]), .A3(DataRead[31]), .A4(
        DataRead[30]), .Z(n2137) );
  Bit_0 \WordArray[0].Word[0].Cell  ( .Q(\WordArray[0].Word[0].QWire ), .D(
        n103), .Clk(_9_net_) );
  Bit_1055 \WordArray[0].Word[1].Cell  ( .Q(\WordArray[0].Word[1].QWire ), .D(
        n105), .Clk(_9_net_) );
  Bit_1054 \WordArray[0].Word[2].Cell  ( .Q(\WordArray[0].Word[2].QWire ), .D(
        n107), .Clk(_9_net_) );
  Bit_1053 \WordArray[0].Word[3].Cell  ( .Q(\WordArray[0].Word[3].QWire ), .D(
        n109), .Clk(_9_net_) );
  Bit_1052 \WordArray[0].Word[4].Cell  ( .Q(\WordArray[0].Word[4].QWire ), .D(
        n111), .Clk(_9_net_) );
  Bit_1051 \WordArray[0].Word[5].Cell  ( .Q(\WordArray[0].Word[5].QWire ), .D(
        n113), .Clk(_9_net_) );
  Bit_1050 \WordArray[0].Word[6].Cell  ( .Q(\WordArray[0].Word[6].QWire ), .D(
        n115), .Clk(_9_net_) );
  Bit_1049 \WordArray[0].Word[7].Cell  ( .Q(\WordArray[0].Word[7].QWire ), .D(
        n117), .Clk(_9_net_) );
  Bit_1048 \WordArray[0].Word[8].Cell  ( .Q(\WordArray[0].Word[8].QWire ), .D(
        n119), .Clk(_9_net_) );
  Bit_1047 \WordArray[0].Word[9].Cell  ( .Q(\WordArray[0].Word[9].QWire ), .D(
        n121), .Clk(_9_net_) );
  Bit_1046 \WordArray[0].Word[10].Cell  ( .Q(\WordArray[0].Word[10].QWire ), 
        .D(n123), .Clk(_9_net_) );
  Bit_1045 \WordArray[0].Word[11].Cell  ( .Q(\WordArray[0].Word[11].QWire ), 
        .D(n125), .Clk(_9_net_) );
  Bit_1044 \WordArray[0].Word[12].Cell  ( .Q(\WordArray[0].Word[12].QWire ), 
        .D(n127), .Clk(_9_net_) );
  Bit_1043 \WordArray[0].Word[13].Cell  ( .Q(\WordArray[0].Word[13].QWire ), 
        .D(n129), .Clk(_9_net_) );
  Bit_1042 \WordArray[0].Word[14].Cell  ( .Q(\WordArray[0].Word[14].QWire ), 
        .D(n131), .Clk(_9_net_) );
  Bit_1041 \WordArray[0].Word[15].Cell  ( .Q(\WordArray[0].Word[15].QWire ), 
        .D(n133), .Clk(_9_net_) );
  Bit_1040 \WordArray[0].Word[16].Cell  ( .Q(\WordArray[0].Word[16].QWire ), 
        .D(n135), .Clk(_9_net_) );
  Bit_1039 \WordArray[0].Word[17].Cell  ( .Q(\WordArray[0].Word[17].QWire ), 
        .D(n137), .Clk(_9_net_) );
  Bit_1038 \WordArray[0].Word[18].Cell  ( .Q(\WordArray[0].Word[18].QWire ), 
        .D(n139), .Clk(_9_net_) );
  Bit_1037 \WordArray[0].Word[19].Cell  ( .Q(\WordArray[0].Word[19].QWire ), 
        .D(n141), .Clk(_9_net_) );
  Bit_1036 \WordArray[0].Word[20].Cell  ( .Q(\WordArray[0].Word[20].QWire ), 
        .D(n143), .Clk(_9_net_) );
  Bit_1035 \WordArray[0].Word[21].Cell  ( .Q(\WordArray[0].Word[21].QWire ), 
        .D(n145), .Clk(_9_net_) );
  Bit_1034 \WordArray[0].Word[22].Cell  ( .Q(\WordArray[0].Word[22].QWire ), 
        .D(n147), .Clk(_9_net_) );
  Bit_1033 \WordArray[0].Word[23].Cell  ( .Q(\WordArray[0].Word[23].QWire ), 
        .D(n149), .Clk(_9_net_) );
  Bit_1032 \WordArray[0].Word[24].Cell  ( .Q(\WordArray[0].Word[24].QWire ), 
        .D(n151), .Clk(_9_net_) );
  Bit_1031 \WordArray[0].Word[25].Cell  ( .Q(\WordArray[0].Word[25].QWire ), 
        .D(n153), .Clk(_9_net_) );
  Bit_1030 \WordArray[0].Word[26].Cell  ( .Q(\WordArray[0].Word[26].QWire ), 
        .D(n155), .Clk(_9_net_) );
  Bit_1029 \WordArray[0].Word[27].Cell  ( .Q(\WordArray[0].Word[27].QWire ), 
        .D(n157), .Clk(_9_net_) );
  Bit_1028 \WordArray[0].Word[28].Cell  ( .Q(\WordArray[0].Word[28].QWire ), 
        .D(n159), .Clk(_9_net_) );
  Bit_1027 \WordArray[0].Word[29].Cell  ( .Q(\WordArray[0].Word[29].QWire ), 
        .D(n161), .Clk(_9_net_) );
  Bit_1026 \WordArray[0].Word[30].Cell  ( .Q(\WordArray[0].Word[30].QWire ), 
        .D(n163), .Clk(_9_net_) );
  Bit_1025 \WordArray[0].Word[31].Cell  ( .Q(\WordArray[0].Word[31].QWire ), 
        .D(n165), .Clk(_9_net_) );
  Bit_1024 \WordArray[0].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _9_net_) );
  Bit_1023 \WordArray[1].Word[0].Cell  ( .Q(\WordArray[1].Word[0].QWire ), .D(
        n103), .Clk(_65_net_) );
  Bit_1022 \WordArray[1].Word[1].Cell  ( .Q(\WordArray[1].Word[1].QWire ), .D(
        n105), .Clk(_65_net_) );
  Bit_1021 \WordArray[1].Word[2].Cell  ( .Q(\WordArray[1].Word[2].QWire ), .D(
        n107), .Clk(_65_net_) );
  Bit_1020 \WordArray[1].Word[3].Cell  ( .Q(\WordArray[1].Word[3].QWire ), .D(
        n109), .Clk(_65_net_) );
  Bit_1019 \WordArray[1].Word[4].Cell  ( .Q(\WordArray[1].Word[4].QWire ), .D(
        n111), .Clk(_65_net_) );
  Bit_1018 \WordArray[1].Word[5].Cell  ( .Q(\WordArray[1].Word[5].QWire ), .D(
        n113), .Clk(_65_net_) );
  Bit_1017 \WordArray[1].Word[6].Cell  ( .Q(\WordArray[1].Word[6].QWire ), .D(
        n115), .Clk(_65_net_) );
  Bit_1016 \WordArray[1].Word[7].Cell  ( .Q(\WordArray[1].Word[7].QWire ), .D(
        n117), .Clk(_65_net_) );
  Bit_1015 \WordArray[1].Word[8].Cell  ( .Q(\WordArray[1].Word[8].QWire ), .D(
        n119), .Clk(_65_net_) );
  Bit_1014 \WordArray[1].Word[9].Cell  ( .Q(\WordArray[1].Word[9].QWire ), .D(
        n121), .Clk(_65_net_) );
  Bit_1013 \WordArray[1].Word[10].Cell  ( .Q(\WordArray[1].Word[10].QWire ), 
        .D(n123), .Clk(_65_net_) );
  Bit_1012 \WordArray[1].Word[11].Cell  ( .Q(\WordArray[1].Word[11].QWire ), 
        .D(n125), .Clk(_65_net_) );
  Bit_1011 \WordArray[1].Word[12].Cell  ( .Q(\WordArray[1].Word[12].QWire ), 
        .D(n127), .Clk(_65_net_) );
  Bit_1010 \WordArray[1].Word[13].Cell  ( .Q(\WordArray[1].Word[13].QWire ), 
        .D(n129), .Clk(_65_net_) );
  Bit_1009 \WordArray[1].Word[14].Cell  ( .Q(\WordArray[1].Word[14].QWire ), 
        .D(n131), .Clk(_65_net_) );
  Bit_1008 \WordArray[1].Word[15].Cell  ( .Q(\WordArray[1].Word[15].QWire ), 
        .D(n133), .Clk(_65_net_) );
  Bit_1007 \WordArray[1].Word[16].Cell  ( .Q(\WordArray[1].Word[16].QWire ), 
        .D(n135), .Clk(_65_net_) );
  Bit_1006 \WordArray[1].Word[17].Cell  ( .Q(\WordArray[1].Word[17].QWire ), 
        .D(n137), .Clk(_65_net_) );
  Bit_1005 \WordArray[1].Word[18].Cell  ( .Q(\WordArray[1].Word[18].QWire ), 
        .D(n139), .Clk(_65_net_) );
  Bit_1004 \WordArray[1].Word[19].Cell  ( .Q(\WordArray[1].Word[19].QWire ), 
        .D(n141), .Clk(_65_net_) );
  Bit_1003 \WordArray[1].Word[20].Cell  ( .Q(\WordArray[1].Word[20].QWire ), 
        .D(n143), .Clk(_65_net_) );
  Bit_1002 \WordArray[1].Word[21].Cell  ( .Q(\WordArray[1].Word[21].QWire ), 
        .D(n145), .Clk(_65_net_) );
  Bit_1001 \WordArray[1].Word[22].Cell  ( .Q(\WordArray[1].Word[22].QWire ), 
        .D(n147), .Clk(_65_net_) );
  Bit_1000 \WordArray[1].Word[23].Cell  ( .Q(\WordArray[1].Word[23].QWire ), 
        .D(n149), .Clk(_65_net_) );
  Bit_999 \WordArray[1].Word[24].Cell  ( .Q(\WordArray[1].Word[24].QWire ), 
        .D(n151), .Clk(_65_net_) );
  Bit_998 \WordArray[1].Word[25].Cell  ( .Q(\WordArray[1].Word[25].QWire ), 
        .D(n153), .Clk(_65_net_) );
  Bit_997 \WordArray[1].Word[26].Cell  ( .Q(\WordArray[1].Word[26].QWire ), 
        .D(n155), .Clk(_65_net_) );
  Bit_996 \WordArray[1].Word[27].Cell  ( .Q(\WordArray[1].Word[27].QWire ), 
        .D(n157), .Clk(_65_net_) );
  Bit_995 \WordArray[1].Word[28].Cell  ( .Q(\WordArray[1].Word[28].QWire ), 
        .D(n159), .Clk(_65_net_) );
  Bit_994 \WordArray[1].Word[29].Cell  ( .Q(\WordArray[1].Word[29].QWire ), 
        .D(n161), .Clk(_65_net_) );
  Bit_993 \WordArray[1].Word[30].Cell  ( .Q(\WordArray[1].Word[30].QWire ), 
        .D(n163), .Clk(_65_net_) );
  Bit_992 \WordArray[1].Word[31].Cell  ( .Q(\WordArray[1].Word[31].QWire ), 
        .D(n165), .Clk(_65_net_) );
  Bit_991 \WordArray[1].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _65_net_) );
  Bit_990 \WordArray[2].Word[0].Cell  ( .Q(\WordArray[2].Word[0].QWire ), .D(
        n103), .Clk(_98_net_) );
  Bit_989 \WordArray[2].Word[1].Cell  ( .Q(\WordArray[2].Word[1].QWire ), .D(
        n105), .Clk(_98_net_) );
  Bit_988 \WordArray[2].Word[2].Cell  ( .Q(\WordArray[2].Word[2].QWire ), .D(
        n107), .Clk(_98_net_) );
  Bit_987 \WordArray[2].Word[3].Cell  ( .Q(\WordArray[2].Word[3].QWire ), .D(
        n109), .Clk(_98_net_) );
  Bit_986 \WordArray[2].Word[4].Cell  ( .Q(\WordArray[2].Word[4].QWire ), .D(
        n111), .Clk(_98_net_) );
  Bit_985 \WordArray[2].Word[5].Cell  ( .Q(\WordArray[2].Word[5].QWire ), .D(
        n113), .Clk(_98_net_) );
  Bit_984 \WordArray[2].Word[6].Cell  ( .Q(\WordArray[2].Word[6].QWire ), .D(
        n115), .Clk(_98_net_) );
  Bit_983 \WordArray[2].Word[7].Cell  ( .Q(\WordArray[2].Word[7].QWire ), .D(
        n117), .Clk(_98_net_) );
  Bit_982 \WordArray[2].Word[8].Cell  ( .Q(\WordArray[2].Word[8].QWire ), .D(
        n119), .Clk(_98_net_) );
  Bit_981 \WordArray[2].Word[9].Cell  ( .Q(\WordArray[2].Word[9].QWire ), .D(
        n121), .Clk(_98_net_) );
  Bit_980 \WordArray[2].Word[10].Cell  ( .Q(\WordArray[2].Word[10].QWire ), 
        .D(n123), .Clk(_98_net_) );
  Bit_979 \WordArray[2].Word[11].Cell  ( .Q(\WordArray[2].Word[11].QWire ), 
        .D(n125), .Clk(_98_net_) );
  Bit_978 \WordArray[2].Word[12].Cell  ( .Q(\WordArray[2].Word[12].QWire ), 
        .D(n127), .Clk(_98_net_) );
  Bit_977 \WordArray[2].Word[13].Cell  ( .Q(\WordArray[2].Word[13].QWire ), 
        .D(n129), .Clk(_98_net_) );
  Bit_976 \WordArray[2].Word[14].Cell  ( .Q(\WordArray[2].Word[14].QWire ), 
        .D(n131), .Clk(_98_net_) );
  Bit_975 \WordArray[2].Word[15].Cell  ( .Q(\WordArray[2].Word[15].QWire ), 
        .D(n133), .Clk(_98_net_) );
  Bit_974 \WordArray[2].Word[16].Cell  ( .Q(\WordArray[2].Word[16].QWire ), 
        .D(n135), .Clk(_98_net_) );
  Bit_973 \WordArray[2].Word[17].Cell  ( .Q(\WordArray[2].Word[17].QWire ), 
        .D(n137), .Clk(_98_net_) );
  Bit_972 \WordArray[2].Word[18].Cell  ( .Q(\WordArray[2].Word[18].QWire ), 
        .D(n139), .Clk(_98_net_) );
  Bit_971 \WordArray[2].Word[19].Cell  ( .Q(\WordArray[2].Word[19].QWire ), 
        .D(n141), .Clk(_98_net_) );
  Bit_970 \WordArray[2].Word[20].Cell  ( .Q(\WordArray[2].Word[20].QWire ), 
        .D(n143), .Clk(_98_net_) );
  Bit_969 \WordArray[2].Word[21].Cell  ( .Q(\WordArray[2].Word[21].QWire ), 
        .D(n145), .Clk(_98_net_) );
  Bit_968 \WordArray[2].Word[22].Cell  ( .Q(\WordArray[2].Word[22].QWire ), 
        .D(n147), .Clk(_98_net_) );
  Bit_967 \WordArray[2].Word[23].Cell  ( .Q(\WordArray[2].Word[23].QWire ), 
        .D(n149), .Clk(_98_net_) );
  Bit_966 \WordArray[2].Word[24].Cell  ( .Q(\WordArray[2].Word[24].QWire ), 
        .D(n151), .Clk(_98_net_) );
  Bit_965 \WordArray[2].Word[25].Cell  ( .Q(\WordArray[2].Word[25].QWire ), 
        .D(n153), .Clk(_98_net_) );
  Bit_964 \WordArray[2].Word[26].Cell  ( .Q(\WordArray[2].Word[26].QWire ), 
        .D(n155), .Clk(_98_net_) );
  Bit_963 \WordArray[2].Word[27].Cell  ( .Q(\WordArray[2].Word[27].QWire ), 
        .D(n157), .Clk(_98_net_) );
  Bit_962 \WordArray[2].Word[28].Cell  ( .Q(\WordArray[2].Word[28].QWire ), 
        .D(n159), .Clk(_98_net_) );
  Bit_961 \WordArray[2].Word[29].Cell  ( .Q(\WordArray[2].Word[29].QWire ), 
        .D(n161), .Clk(_98_net_) );
  Bit_960 \WordArray[2].Word[30].Cell  ( .Q(\WordArray[2].Word[30].QWire ), 
        .D(n163), .Clk(_98_net_) );
  Bit_959 \WordArray[2].Word[31].Cell  ( .Q(\WordArray[2].Word[31].QWire ), 
        .D(n165), .Clk(_98_net_) );
  Bit_958 \WordArray[2].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _98_net_) );
  Bit_957 \WordArray[3].Word[0].Cell  ( .Q(\WordArray[3].Word[0].QWire ), .D(
        n103), .Clk(_99_net_) );
  Bit_956 \WordArray[3].Word[1].Cell  ( .Q(\WordArray[3].Word[1].QWire ), .D(
        n105), .Clk(_99_net_) );
  Bit_955 \WordArray[3].Word[2].Cell  ( .Q(\WordArray[3].Word[2].QWire ), .D(
        n107), .Clk(_99_net_) );
  Bit_954 \WordArray[3].Word[3].Cell  ( .Q(\WordArray[3].Word[3].QWire ), .D(
        n109), .Clk(_99_net_) );
  Bit_953 \WordArray[3].Word[4].Cell  ( .Q(\WordArray[3].Word[4].QWire ), .D(
        n111), .Clk(_99_net_) );
  Bit_952 \WordArray[3].Word[5].Cell  ( .Q(\WordArray[3].Word[5].QWire ), .D(
        n113), .Clk(_99_net_) );
  Bit_951 \WordArray[3].Word[6].Cell  ( .Q(\WordArray[3].Word[6].QWire ), .D(
        n115), .Clk(_99_net_) );
  Bit_950 \WordArray[3].Word[7].Cell  ( .Q(\WordArray[3].Word[7].QWire ), .D(
        n117), .Clk(_99_net_) );
  Bit_949 \WordArray[3].Word[8].Cell  ( .Q(\WordArray[3].Word[8].QWire ), .D(
        n119), .Clk(_99_net_) );
  Bit_948 \WordArray[3].Word[9].Cell  ( .Q(\WordArray[3].Word[9].QWire ), .D(
        n121), .Clk(_99_net_) );
  Bit_947 \WordArray[3].Word[10].Cell  ( .Q(\WordArray[3].Word[10].QWire ), 
        .D(n123), .Clk(_99_net_) );
  Bit_946 \WordArray[3].Word[11].Cell  ( .Q(\WordArray[3].Word[11].QWire ), 
        .D(n125), .Clk(_99_net_) );
  Bit_945 \WordArray[3].Word[12].Cell  ( .Q(\WordArray[3].Word[12].QWire ), 
        .D(n127), .Clk(_99_net_) );
  Bit_944 \WordArray[3].Word[13].Cell  ( .Q(\WordArray[3].Word[13].QWire ), 
        .D(n129), .Clk(_99_net_) );
  Bit_943 \WordArray[3].Word[14].Cell  ( .Q(\WordArray[3].Word[14].QWire ), 
        .D(n131), .Clk(_99_net_) );
  Bit_942 \WordArray[3].Word[15].Cell  ( .Q(\WordArray[3].Word[15].QWire ), 
        .D(n133), .Clk(_99_net_) );
  Bit_941 \WordArray[3].Word[16].Cell  ( .Q(\WordArray[3].Word[16].QWire ), 
        .D(n135), .Clk(_99_net_) );
  Bit_940 \WordArray[3].Word[17].Cell  ( .Q(\WordArray[3].Word[17].QWire ), 
        .D(n137), .Clk(_99_net_) );
  Bit_939 \WordArray[3].Word[18].Cell  ( .Q(\WordArray[3].Word[18].QWire ), 
        .D(n139), .Clk(_99_net_) );
  Bit_938 \WordArray[3].Word[19].Cell  ( .Q(\WordArray[3].Word[19].QWire ), 
        .D(n141), .Clk(_99_net_) );
  Bit_937 \WordArray[3].Word[20].Cell  ( .Q(\WordArray[3].Word[20].QWire ), 
        .D(n143), .Clk(_99_net_) );
  Bit_936 \WordArray[3].Word[21].Cell  ( .Q(\WordArray[3].Word[21].QWire ), 
        .D(n145), .Clk(_99_net_) );
  Bit_935 \WordArray[3].Word[22].Cell  ( .Q(\WordArray[3].Word[22].QWire ), 
        .D(n147), .Clk(_99_net_) );
  Bit_934 \WordArray[3].Word[23].Cell  ( .Q(\WordArray[3].Word[23].QWire ), 
        .D(n149), .Clk(_99_net_) );
  Bit_933 \WordArray[3].Word[24].Cell  ( .Q(\WordArray[3].Word[24].QWire ), 
        .D(n151), .Clk(_99_net_) );
  Bit_932 \WordArray[3].Word[25].Cell  ( .Q(\WordArray[3].Word[25].QWire ), 
        .D(n153), .Clk(_99_net_) );
  Bit_931 \WordArray[3].Word[26].Cell  ( .Q(\WordArray[3].Word[26].QWire ), 
        .D(n155), .Clk(_99_net_) );
  Bit_930 \WordArray[3].Word[27].Cell  ( .Q(\WordArray[3].Word[27].QWire ), 
        .D(n157), .Clk(_99_net_) );
  Bit_929 \WordArray[3].Word[28].Cell  ( .Q(\WordArray[3].Word[28].QWire ), 
        .D(n159), .Clk(_99_net_) );
  Bit_928 \WordArray[3].Word[29].Cell  ( .Q(\WordArray[3].Word[29].QWire ), 
        .D(n161), .Clk(_99_net_) );
  Bit_927 \WordArray[3].Word[30].Cell  ( .Q(\WordArray[3].Word[30].QWire ), 
        .D(n163), .Clk(_99_net_) );
  Bit_926 \WordArray[3].Word[31].Cell  ( .Q(\WordArray[3].Word[31].QWire ), 
        .D(n165), .Clk(_99_net_) );
  Bit_925 \WordArray[3].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _99_net_) );
  Bit_924 \WordArray[4].Word[0].Cell  ( .Q(\WordArray[4].Word[0].QWire ), .D(
        n103), .Clk(_164_net_) );
  Bit_923 \WordArray[4].Word[1].Cell  ( .Q(\WordArray[4].Word[1].QWire ), .D(
        n105), .Clk(_164_net_) );
  Bit_922 \WordArray[4].Word[2].Cell  ( .Q(\WordArray[4].Word[2].QWire ), .D(
        n107), .Clk(_164_net_) );
  Bit_921 \WordArray[4].Word[3].Cell  ( .Q(\WordArray[4].Word[3].QWire ), .D(
        n109), .Clk(_164_net_) );
  Bit_920 \WordArray[4].Word[4].Cell  ( .Q(\WordArray[4].Word[4].QWire ), .D(
        n111), .Clk(_164_net_) );
  Bit_919 \WordArray[4].Word[5].Cell  ( .Q(\WordArray[4].Word[5].QWire ), .D(
        n113), .Clk(_164_net_) );
  Bit_918 \WordArray[4].Word[6].Cell  ( .Q(\WordArray[4].Word[6].QWire ), .D(
        n115), .Clk(_164_net_) );
  Bit_917 \WordArray[4].Word[7].Cell  ( .Q(\WordArray[4].Word[7].QWire ), .D(
        n117), .Clk(_164_net_) );
  Bit_916 \WordArray[4].Word[8].Cell  ( .Q(\WordArray[4].Word[8].QWire ), .D(
        n119), .Clk(_164_net_) );
  Bit_915 \WordArray[4].Word[9].Cell  ( .Q(\WordArray[4].Word[9].QWire ), .D(
        n121), .Clk(_164_net_) );
  Bit_914 \WordArray[4].Word[10].Cell  ( .Q(\WordArray[4].Word[10].QWire ), 
        .D(n123), .Clk(_164_net_) );
  Bit_913 \WordArray[4].Word[11].Cell  ( .Q(\WordArray[4].Word[11].QWire ), 
        .D(n125), .Clk(_164_net_) );
  Bit_912 \WordArray[4].Word[12].Cell  ( .Q(\WordArray[4].Word[12].QWire ), 
        .D(n127), .Clk(_164_net_) );
  Bit_911 \WordArray[4].Word[13].Cell  ( .Q(\WordArray[4].Word[13].QWire ), 
        .D(n129), .Clk(_164_net_) );
  Bit_910 \WordArray[4].Word[14].Cell  ( .Q(\WordArray[4].Word[14].QWire ), 
        .D(n131), .Clk(_164_net_) );
  Bit_909 \WordArray[4].Word[15].Cell  ( .Q(\WordArray[4].Word[15].QWire ), 
        .D(n133), .Clk(_164_net_) );
  Bit_908 \WordArray[4].Word[16].Cell  ( .Q(\WordArray[4].Word[16].QWire ), 
        .D(n135), .Clk(_164_net_) );
  Bit_907 \WordArray[4].Word[17].Cell  ( .Q(\WordArray[4].Word[17].QWire ), 
        .D(n137), .Clk(_164_net_) );
  Bit_906 \WordArray[4].Word[18].Cell  ( .Q(\WordArray[4].Word[18].QWire ), 
        .D(n139), .Clk(_164_net_) );
  Bit_905 \WordArray[4].Word[19].Cell  ( .Q(\WordArray[4].Word[19].QWire ), 
        .D(n141), .Clk(_164_net_) );
  Bit_904 \WordArray[4].Word[20].Cell  ( .Q(\WordArray[4].Word[20].QWire ), 
        .D(n143), .Clk(_164_net_) );
  Bit_903 \WordArray[4].Word[21].Cell  ( .Q(\WordArray[4].Word[21].QWire ), 
        .D(n145), .Clk(_164_net_) );
  Bit_902 \WordArray[4].Word[22].Cell  ( .Q(\WordArray[4].Word[22].QWire ), 
        .D(n147), .Clk(_164_net_) );
  Bit_901 \WordArray[4].Word[23].Cell  ( .Q(\WordArray[4].Word[23].QWire ), 
        .D(n149), .Clk(_164_net_) );
  Bit_900 \WordArray[4].Word[24].Cell  ( .Q(\WordArray[4].Word[24].QWire ), 
        .D(n151), .Clk(_164_net_) );
  Bit_899 \WordArray[4].Word[25].Cell  ( .Q(\WordArray[4].Word[25].QWire ), 
        .D(n153), .Clk(_164_net_) );
  Bit_898 \WordArray[4].Word[26].Cell  ( .Q(\WordArray[4].Word[26].QWire ), 
        .D(n155), .Clk(_164_net_) );
  Bit_897 \WordArray[4].Word[27].Cell  ( .Q(\WordArray[4].Word[27].QWire ), 
        .D(n157), .Clk(_164_net_) );
  Bit_896 \WordArray[4].Word[28].Cell  ( .Q(\WordArray[4].Word[28].QWire ), 
        .D(n159), .Clk(_164_net_) );
  Bit_895 \WordArray[4].Word[29].Cell  ( .Q(\WordArray[4].Word[29].QWire ), 
        .D(n161), .Clk(_164_net_) );
  Bit_894 \WordArray[4].Word[30].Cell  ( .Q(\WordArray[4].Word[30].QWire ), 
        .D(n163), .Clk(_164_net_) );
  Bit_893 \WordArray[4].Word[31].Cell  ( .Q(\WordArray[4].Word[31].QWire ), 
        .D(n165), .Clk(_164_net_) );
  Bit_892 \WordArray[4].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _164_net_) );
  Bit_891 \WordArray[5].Word[0].Cell  ( .Q(\WordArray[5].Word[0].QWire ), .D(
        n103), .Clk(_197_net_) );
  Bit_890 \WordArray[5].Word[1].Cell  ( .Q(\WordArray[5].Word[1].QWire ), .D(
        n105), .Clk(_197_net_) );
  Bit_889 \WordArray[5].Word[2].Cell  ( .Q(\WordArray[5].Word[2].QWire ), .D(
        n107), .Clk(_197_net_) );
  Bit_888 \WordArray[5].Word[3].Cell  ( .Q(\WordArray[5].Word[3].QWire ), .D(
        n109), .Clk(_197_net_) );
  Bit_887 \WordArray[5].Word[4].Cell  ( .Q(\WordArray[5].Word[4].QWire ), .D(
        n111), .Clk(_197_net_) );
  Bit_886 \WordArray[5].Word[5].Cell  ( .Q(\WordArray[5].Word[5].QWire ), .D(
        n113), .Clk(_197_net_) );
  Bit_885 \WordArray[5].Word[6].Cell  ( .Q(\WordArray[5].Word[6].QWire ), .D(
        n115), .Clk(_197_net_) );
  Bit_884 \WordArray[5].Word[7].Cell  ( .Q(\WordArray[5].Word[7].QWire ), .D(
        n117), .Clk(_197_net_) );
  Bit_883 \WordArray[5].Word[8].Cell  ( .Q(\WordArray[5].Word[8].QWire ), .D(
        n119), .Clk(_197_net_) );
  Bit_882 \WordArray[5].Word[9].Cell  ( .Q(\WordArray[5].Word[9].QWire ), .D(
        n121), .Clk(_197_net_) );
  Bit_881 \WordArray[5].Word[10].Cell  ( .Q(\WordArray[5].Word[10].QWire ), 
        .D(n123), .Clk(_197_net_) );
  Bit_880 \WordArray[5].Word[11].Cell  ( .Q(\WordArray[5].Word[11].QWire ), 
        .D(n125), .Clk(_197_net_) );
  Bit_879 \WordArray[5].Word[12].Cell  ( .Q(\WordArray[5].Word[12].QWire ), 
        .D(n127), .Clk(_197_net_) );
  Bit_878 \WordArray[5].Word[13].Cell  ( .Q(\WordArray[5].Word[13].QWire ), 
        .D(n129), .Clk(_197_net_) );
  Bit_877 \WordArray[5].Word[14].Cell  ( .Q(\WordArray[5].Word[14].QWire ), 
        .D(n131), .Clk(_197_net_) );
  Bit_876 \WordArray[5].Word[15].Cell  ( .Q(\WordArray[5].Word[15].QWire ), 
        .D(n133), .Clk(_197_net_) );
  Bit_875 \WordArray[5].Word[16].Cell  ( .Q(\WordArray[5].Word[16].QWire ), 
        .D(n135), .Clk(_197_net_) );
  Bit_874 \WordArray[5].Word[17].Cell  ( .Q(\WordArray[5].Word[17].QWire ), 
        .D(n137), .Clk(_197_net_) );
  Bit_873 \WordArray[5].Word[18].Cell  ( .Q(\WordArray[5].Word[18].QWire ), 
        .D(n139), .Clk(_197_net_) );
  Bit_872 \WordArray[5].Word[19].Cell  ( .Q(\WordArray[5].Word[19].QWire ), 
        .D(n141), .Clk(_197_net_) );
  Bit_871 \WordArray[5].Word[20].Cell  ( .Q(\WordArray[5].Word[20].QWire ), 
        .D(n143), .Clk(_197_net_) );
  Bit_870 \WordArray[5].Word[21].Cell  ( .Q(\WordArray[5].Word[21].QWire ), 
        .D(n145), .Clk(_197_net_) );
  Bit_869 \WordArray[5].Word[22].Cell  ( .Q(\WordArray[5].Word[22].QWire ), 
        .D(n147), .Clk(_197_net_) );
  Bit_868 \WordArray[5].Word[23].Cell  ( .Q(\WordArray[5].Word[23].QWire ), 
        .D(n149), .Clk(_197_net_) );
  Bit_867 \WordArray[5].Word[24].Cell  ( .Q(\WordArray[5].Word[24].QWire ), 
        .D(n151), .Clk(_197_net_) );
  Bit_866 \WordArray[5].Word[25].Cell  ( .Q(\WordArray[5].Word[25].QWire ), 
        .D(n153), .Clk(_197_net_) );
  Bit_865 \WordArray[5].Word[26].Cell  ( .Q(\WordArray[5].Word[26].QWire ), 
        .D(n155), .Clk(_197_net_) );
  Bit_864 \WordArray[5].Word[27].Cell  ( .Q(\WordArray[5].Word[27].QWire ), 
        .D(n157), .Clk(_197_net_) );
  Bit_863 \WordArray[5].Word[28].Cell  ( .Q(\WordArray[5].Word[28].QWire ), 
        .D(n159), .Clk(_197_net_) );
  Bit_862 \WordArray[5].Word[29].Cell  ( .Q(\WordArray[5].Word[29].QWire ), 
        .D(n161), .Clk(_197_net_) );
  Bit_861 \WordArray[5].Word[30].Cell  ( .Q(\WordArray[5].Word[30].QWire ), 
        .D(n163), .Clk(_197_net_) );
  Bit_860 \WordArray[5].Word[31].Cell  ( .Q(\WordArray[5].Word[31].QWire ), 
        .D(n165), .Clk(_197_net_) );
  Bit_859 \WordArray[5].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _197_net_) );
  Bit_858 \WordArray[6].Word[0].Cell  ( .Q(\WordArray[6].Word[0].QWire ), .D(
        n103), .Clk(_230_net_) );
  Bit_857 \WordArray[6].Word[1].Cell  ( .Q(\WordArray[6].Word[1].QWire ), .D(
        n105), .Clk(_230_net_) );
  Bit_856 \WordArray[6].Word[2].Cell  ( .Q(\WordArray[6].Word[2].QWire ), .D(
        n107), .Clk(_230_net_) );
  Bit_855 \WordArray[6].Word[3].Cell  ( .Q(\WordArray[6].Word[3].QWire ), .D(
        n109), .Clk(_230_net_) );
  Bit_854 \WordArray[6].Word[4].Cell  ( .Q(\WordArray[6].Word[4].QWire ), .D(
        n111), .Clk(_230_net_) );
  Bit_853 \WordArray[6].Word[5].Cell  ( .Q(\WordArray[6].Word[5].QWire ), .D(
        n113), .Clk(_230_net_) );
  Bit_852 \WordArray[6].Word[6].Cell  ( .Q(\WordArray[6].Word[6].QWire ), .D(
        n115), .Clk(_230_net_) );
  Bit_851 \WordArray[6].Word[7].Cell  ( .Q(\WordArray[6].Word[7].QWire ), .D(
        n117), .Clk(_230_net_) );
  Bit_850 \WordArray[6].Word[8].Cell  ( .Q(\WordArray[6].Word[8].QWire ), .D(
        n119), .Clk(_230_net_) );
  Bit_849 \WordArray[6].Word[9].Cell  ( .Q(\WordArray[6].Word[9].QWire ), .D(
        n121), .Clk(_230_net_) );
  Bit_848 \WordArray[6].Word[10].Cell  ( .Q(\WordArray[6].Word[10].QWire ), 
        .D(n123), .Clk(_230_net_) );
  Bit_847 \WordArray[6].Word[11].Cell  ( .Q(\WordArray[6].Word[11].QWire ), 
        .D(n125), .Clk(_230_net_) );
  Bit_846 \WordArray[6].Word[12].Cell  ( .Q(\WordArray[6].Word[12].QWire ), 
        .D(n127), .Clk(_230_net_) );
  Bit_845 \WordArray[6].Word[13].Cell  ( .Q(\WordArray[6].Word[13].QWire ), 
        .D(n129), .Clk(_230_net_) );
  Bit_844 \WordArray[6].Word[14].Cell  ( .Q(\WordArray[6].Word[14].QWire ), 
        .D(n131), .Clk(_230_net_) );
  Bit_843 \WordArray[6].Word[15].Cell  ( .Q(\WordArray[6].Word[15].QWire ), 
        .D(n133), .Clk(_230_net_) );
  Bit_842 \WordArray[6].Word[16].Cell  ( .Q(\WordArray[6].Word[16].QWire ), 
        .D(n135), .Clk(_230_net_) );
  Bit_841 \WordArray[6].Word[17].Cell  ( .Q(\WordArray[6].Word[17].QWire ), 
        .D(n137), .Clk(_230_net_) );
  Bit_840 \WordArray[6].Word[18].Cell  ( .Q(\WordArray[6].Word[18].QWire ), 
        .D(n139), .Clk(_230_net_) );
  Bit_839 \WordArray[6].Word[19].Cell  ( .Q(\WordArray[6].Word[19].QWire ), 
        .D(n141), .Clk(_230_net_) );
  Bit_838 \WordArray[6].Word[20].Cell  ( .Q(\WordArray[6].Word[20].QWire ), 
        .D(n143), .Clk(_230_net_) );
  Bit_837 \WordArray[6].Word[21].Cell  ( .Q(\WordArray[6].Word[21].QWire ), 
        .D(n145), .Clk(_230_net_) );
  Bit_836 \WordArray[6].Word[22].Cell  ( .Q(\WordArray[6].Word[22].QWire ), 
        .D(n147), .Clk(_230_net_) );
  Bit_835 \WordArray[6].Word[23].Cell  ( .Q(\WordArray[6].Word[23].QWire ), 
        .D(n149), .Clk(_230_net_) );
  Bit_834 \WordArray[6].Word[24].Cell  ( .Q(\WordArray[6].Word[24].QWire ), 
        .D(n151), .Clk(_230_net_) );
  Bit_833 \WordArray[6].Word[25].Cell  ( .Q(\WordArray[6].Word[25].QWire ), 
        .D(n153), .Clk(_230_net_) );
  Bit_832 \WordArray[6].Word[26].Cell  ( .Q(\WordArray[6].Word[26].QWire ), 
        .D(n155), .Clk(_230_net_) );
  Bit_831 \WordArray[6].Word[27].Cell  ( .Q(\WordArray[6].Word[27].QWire ), 
        .D(n157), .Clk(_230_net_) );
  Bit_830 \WordArray[6].Word[28].Cell  ( .Q(\WordArray[6].Word[28].QWire ), 
        .D(n159), .Clk(_230_net_) );
  Bit_829 \WordArray[6].Word[29].Cell  ( .Q(\WordArray[6].Word[29].QWire ), 
        .D(n161), .Clk(_230_net_) );
  Bit_828 \WordArray[6].Word[30].Cell  ( .Q(\WordArray[6].Word[30].QWire ), 
        .D(n163), .Clk(_230_net_) );
  Bit_827 \WordArray[6].Word[31].Cell  ( .Q(\WordArray[6].Word[31].QWire ), 
        .D(n165), .Clk(_230_net_) );
  Bit_826 \WordArray[6].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _230_net_) );
  Bit_825 \WordArray[7].Word[0].Cell  ( .Q(\WordArray[7].Word[0].QWire ), .D(
        n103), .Clk(_263_net_) );
  Bit_824 \WordArray[7].Word[1].Cell  ( .Q(\WordArray[7].Word[1].QWire ), .D(
        n105), .Clk(_263_net_) );
  Bit_823 \WordArray[7].Word[2].Cell  ( .Q(\WordArray[7].Word[2].QWire ), .D(
        n107), .Clk(_263_net_) );
  Bit_822 \WordArray[7].Word[3].Cell  ( .Q(\WordArray[7].Word[3].QWire ), .D(
        n109), .Clk(_263_net_) );
  Bit_821 \WordArray[7].Word[4].Cell  ( .Q(\WordArray[7].Word[4].QWire ), .D(
        n111), .Clk(_263_net_) );
  Bit_820 \WordArray[7].Word[5].Cell  ( .Q(\WordArray[7].Word[5].QWire ), .D(
        n113), .Clk(_263_net_) );
  Bit_819 \WordArray[7].Word[6].Cell  ( .Q(\WordArray[7].Word[6].QWire ), .D(
        n115), .Clk(_263_net_) );
  Bit_818 \WordArray[7].Word[7].Cell  ( .Q(\WordArray[7].Word[7].QWire ), .D(
        n117), .Clk(_263_net_) );
  Bit_817 \WordArray[7].Word[8].Cell  ( .Q(\WordArray[7].Word[8].QWire ), .D(
        n119), .Clk(_263_net_) );
  Bit_816 \WordArray[7].Word[9].Cell  ( .Q(\WordArray[7].Word[9].QWire ), .D(
        n121), .Clk(_263_net_) );
  Bit_815 \WordArray[7].Word[10].Cell  ( .Q(\WordArray[7].Word[10].QWire ), 
        .D(n123), .Clk(_263_net_) );
  Bit_814 \WordArray[7].Word[11].Cell  ( .Q(\WordArray[7].Word[11].QWire ), 
        .D(n125), .Clk(_263_net_) );
  Bit_813 \WordArray[7].Word[12].Cell  ( .Q(\WordArray[7].Word[12].QWire ), 
        .D(n127), .Clk(_263_net_) );
  Bit_812 \WordArray[7].Word[13].Cell  ( .Q(\WordArray[7].Word[13].QWire ), 
        .D(n129), .Clk(_263_net_) );
  Bit_811 \WordArray[7].Word[14].Cell  ( .Q(\WordArray[7].Word[14].QWire ), 
        .D(n131), .Clk(_263_net_) );
  Bit_810 \WordArray[7].Word[15].Cell  ( .Q(\WordArray[7].Word[15].QWire ), 
        .D(n133), .Clk(_263_net_) );
  Bit_809 \WordArray[7].Word[16].Cell  ( .Q(\WordArray[7].Word[16].QWire ), 
        .D(n135), .Clk(_263_net_) );
  Bit_808 \WordArray[7].Word[17].Cell  ( .Q(\WordArray[7].Word[17].QWire ), 
        .D(n137), .Clk(_263_net_) );
  Bit_807 \WordArray[7].Word[18].Cell  ( .Q(\WordArray[7].Word[18].QWire ), 
        .D(n139), .Clk(_263_net_) );
  Bit_806 \WordArray[7].Word[19].Cell  ( .Q(\WordArray[7].Word[19].QWire ), 
        .D(n141), .Clk(_263_net_) );
  Bit_805 \WordArray[7].Word[20].Cell  ( .Q(\WordArray[7].Word[20].QWire ), 
        .D(n143), .Clk(_263_net_) );
  Bit_804 \WordArray[7].Word[21].Cell  ( .Q(\WordArray[7].Word[21].QWire ), 
        .D(n145), .Clk(_263_net_) );
  Bit_803 \WordArray[7].Word[22].Cell  ( .Q(\WordArray[7].Word[22].QWire ), 
        .D(n147), .Clk(_263_net_) );
  Bit_802 \WordArray[7].Word[23].Cell  ( .Q(\WordArray[7].Word[23].QWire ), 
        .D(n149), .Clk(_263_net_) );
  Bit_801 \WordArray[7].Word[24].Cell  ( .Q(\WordArray[7].Word[24].QWire ), 
        .D(n151), .Clk(_263_net_) );
  Bit_800 \WordArray[7].Word[25].Cell  ( .Q(\WordArray[7].Word[25].QWire ), 
        .D(n153), .Clk(_263_net_) );
  Bit_799 \WordArray[7].Word[26].Cell  ( .Q(\WordArray[7].Word[26].QWire ), 
        .D(n155), .Clk(_263_net_) );
  Bit_798 \WordArray[7].Word[27].Cell  ( .Q(\WordArray[7].Word[27].QWire ), 
        .D(n157), .Clk(_263_net_) );
  Bit_797 \WordArray[7].Word[28].Cell  ( .Q(\WordArray[7].Word[28].QWire ), 
        .D(n159), .Clk(_263_net_) );
  Bit_796 \WordArray[7].Word[29].Cell  ( .Q(\WordArray[7].Word[29].QWire ), 
        .D(n161), .Clk(_263_net_) );
  Bit_795 \WordArray[7].Word[30].Cell  ( .Q(\WordArray[7].Word[30].QWire ), 
        .D(n163), .Clk(_263_net_) );
  Bit_794 \WordArray[7].Word[31].Cell  ( .Q(\WordArray[7].Word[31].QWire ), 
        .D(n165), .Clk(_263_net_) );
  Bit_793 \WordArray[7].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _263_net_) );
  Bit_792 \WordArray[8].Word[0].Cell  ( .Q(\WordArray[8].Word[0].QWire ), .D(
        n103), .Clk(_296_net_) );
  Bit_791 \WordArray[8].Word[1].Cell  ( .Q(\WordArray[8].Word[1].QWire ), .D(
        n105), .Clk(_296_net_) );
  Bit_790 \WordArray[8].Word[2].Cell  ( .Q(\WordArray[8].Word[2].QWire ), .D(
        n107), .Clk(_296_net_) );
  Bit_789 \WordArray[8].Word[3].Cell  ( .Q(\WordArray[8].Word[3].QWire ), .D(
        n109), .Clk(_296_net_) );
  Bit_788 \WordArray[8].Word[4].Cell  ( .Q(\WordArray[8].Word[4].QWire ), .D(
        n111), .Clk(_296_net_) );
  Bit_787 \WordArray[8].Word[5].Cell  ( .Q(\WordArray[8].Word[5].QWire ), .D(
        n113), .Clk(_296_net_) );
  Bit_786 \WordArray[8].Word[6].Cell  ( .Q(\WordArray[8].Word[6].QWire ), .D(
        n115), .Clk(_296_net_) );
  Bit_785 \WordArray[8].Word[7].Cell  ( .Q(\WordArray[8].Word[7].QWire ), .D(
        n117), .Clk(_296_net_) );
  Bit_784 \WordArray[8].Word[8].Cell  ( .Q(\WordArray[8].Word[8].QWire ), .D(
        n119), .Clk(_296_net_) );
  Bit_783 \WordArray[8].Word[9].Cell  ( .Q(\WordArray[8].Word[9].QWire ), .D(
        n121), .Clk(_296_net_) );
  Bit_782 \WordArray[8].Word[10].Cell  ( .Q(\WordArray[8].Word[10].QWire ), 
        .D(n123), .Clk(_296_net_) );
  Bit_781 \WordArray[8].Word[11].Cell  ( .Q(\WordArray[8].Word[11].QWire ), 
        .D(n125), .Clk(_296_net_) );
  Bit_780 \WordArray[8].Word[12].Cell  ( .Q(\WordArray[8].Word[12].QWire ), 
        .D(n127), .Clk(_296_net_) );
  Bit_779 \WordArray[8].Word[13].Cell  ( .Q(\WordArray[8].Word[13].QWire ), 
        .D(n129), .Clk(_296_net_) );
  Bit_778 \WordArray[8].Word[14].Cell  ( .Q(\WordArray[8].Word[14].QWire ), 
        .D(n131), .Clk(_296_net_) );
  Bit_777 \WordArray[8].Word[15].Cell  ( .Q(\WordArray[8].Word[15].QWire ), 
        .D(n133), .Clk(_296_net_) );
  Bit_776 \WordArray[8].Word[16].Cell  ( .Q(\WordArray[8].Word[16].QWire ), 
        .D(n135), .Clk(_296_net_) );
  Bit_775 \WordArray[8].Word[17].Cell  ( .Q(\WordArray[8].Word[17].QWire ), 
        .D(n137), .Clk(_296_net_) );
  Bit_774 \WordArray[8].Word[18].Cell  ( .Q(\WordArray[8].Word[18].QWire ), 
        .D(n139), .Clk(_296_net_) );
  Bit_773 \WordArray[8].Word[19].Cell  ( .Q(\WordArray[8].Word[19].QWire ), 
        .D(n141), .Clk(_296_net_) );
  Bit_772 \WordArray[8].Word[20].Cell  ( .Q(\WordArray[8].Word[20].QWire ), 
        .D(n143), .Clk(_296_net_) );
  Bit_771 \WordArray[8].Word[21].Cell  ( .Q(\WordArray[8].Word[21].QWire ), 
        .D(n145), .Clk(_296_net_) );
  Bit_770 \WordArray[8].Word[22].Cell  ( .Q(\WordArray[8].Word[22].QWire ), 
        .D(n147), .Clk(_296_net_) );
  Bit_769 \WordArray[8].Word[23].Cell  ( .Q(\WordArray[8].Word[23].QWire ), 
        .D(n149), .Clk(_296_net_) );
  Bit_768 \WordArray[8].Word[24].Cell  ( .Q(\WordArray[8].Word[24].QWire ), 
        .D(n151), .Clk(_296_net_) );
  Bit_767 \WordArray[8].Word[25].Cell  ( .Q(\WordArray[8].Word[25].QWire ), 
        .D(n153), .Clk(_296_net_) );
  Bit_766 \WordArray[8].Word[26].Cell  ( .Q(\WordArray[8].Word[26].QWire ), 
        .D(n155), .Clk(_296_net_) );
  Bit_765 \WordArray[8].Word[27].Cell  ( .Q(\WordArray[8].Word[27].QWire ), 
        .D(n157), .Clk(_296_net_) );
  Bit_764 \WordArray[8].Word[28].Cell  ( .Q(\WordArray[8].Word[28].QWire ), 
        .D(n159), .Clk(_296_net_) );
  Bit_763 \WordArray[8].Word[29].Cell  ( .Q(\WordArray[8].Word[29].QWire ), 
        .D(n161), .Clk(_296_net_) );
  Bit_762 \WordArray[8].Word[30].Cell  ( .Q(\WordArray[8].Word[30].QWire ), 
        .D(n163), .Clk(_296_net_) );
  Bit_761 \WordArray[8].Word[31].Cell  ( .Q(\WordArray[8].Word[31].QWire ), 
        .D(n165), .Clk(_296_net_) );
  Bit_760 \WordArray[8].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _296_net_) );
  Bit_759 \WordArray[9].Word[0].Cell  ( .Q(\WordArray[9].Word[0].QWire ), .D(
        n103), .Clk(_329_net_) );
  Bit_758 \WordArray[9].Word[1].Cell  ( .Q(\WordArray[9].Word[1].QWire ), .D(
        n105), .Clk(_329_net_) );
  Bit_757 \WordArray[9].Word[2].Cell  ( .Q(\WordArray[9].Word[2].QWire ), .D(
        n107), .Clk(_329_net_) );
  Bit_756 \WordArray[9].Word[3].Cell  ( .Q(\WordArray[9].Word[3].QWire ), .D(
        n109), .Clk(_329_net_) );
  Bit_755 \WordArray[9].Word[4].Cell  ( .Q(\WordArray[9].Word[4].QWire ), .D(
        n111), .Clk(_329_net_) );
  Bit_754 \WordArray[9].Word[5].Cell  ( .Q(\WordArray[9].Word[5].QWire ), .D(
        n113), .Clk(_329_net_) );
  Bit_753 \WordArray[9].Word[6].Cell  ( .Q(\WordArray[9].Word[6].QWire ), .D(
        n115), .Clk(_329_net_) );
  Bit_752 \WordArray[9].Word[7].Cell  ( .Q(\WordArray[9].Word[7].QWire ), .D(
        n117), .Clk(_329_net_) );
  Bit_751 \WordArray[9].Word[8].Cell  ( .Q(\WordArray[9].Word[8].QWire ), .D(
        n119), .Clk(_329_net_) );
  Bit_750 \WordArray[9].Word[9].Cell  ( .Q(\WordArray[9].Word[9].QWire ), .D(
        n121), .Clk(_329_net_) );
  Bit_749 \WordArray[9].Word[10].Cell  ( .Q(\WordArray[9].Word[10].QWire ), 
        .D(n123), .Clk(_329_net_) );
  Bit_748 \WordArray[9].Word[11].Cell  ( .Q(\WordArray[9].Word[11].QWire ), 
        .D(n125), .Clk(_329_net_) );
  Bit_747 \WordArray[9].Word[12].Cell  ( .Q(\WordArray[9].Word[12].QWire ), 
        .D(n127), .Clk(_329_net_) );
  Bit_746 \WordArray[9].Word[13].Cell  ( .Q(\WordArray[9].Word[13].QWire ), 
        .D(n129), .Clk(_329_net_) );
  Bit_745 \WordArray[9].Word[14].Cell  ( .Q(\WordArray[9].Word[14].QWire ), 
        .D(n131), .Clk(_329_net_) );
  Bit_744 \WordArray[9].Word[15].Cell  ( .Q(\WordArray[9].Word[15].QWire ), 
        .D(n133), .Clk(_329_net_) );
  Bit_743 \WordArray[9].Word[16].Cell  ( .Q(\WordArray[9].Word[16].QWire ), 
        .D(n135), .Clk(_329_net_) );
  Bit_742 \WordArray[9].Word[17].Cell  ( .Q(\WordArray[9].Word[17].QWire ), 
        .D(n137), .Clk(_329_net_) );
  Bit_741 \WordArray[9].Word[18].Cell  ( .Q(\WordArray[9].Word[18].QWire ), 
        .D(n139), .Clk(_329_net_) );
  Bit_740 \WordArray[9].Word[19].Cell  ( .Q(\WordArray[9].Word[19].QWire ), 
        .D(n141), .Clk(_329_net_) );
  Bit_739 \WordArray[9].Word[20].Cell  ( .Q(\WordArray[9].Word[20].QWire ), 
        .D(n143), .Clk(_329_net_) );
  Bit_738 \WordArray[9].Word[21].Cell  ( .Q(\WordArray[9].Word[21].QWire ), 
        .D(n145), .Clk(_329_net_) );
  Bit_737 \WordArray[9].Word[22].Cell  ( .Q(\WordArray[9].Word[22].QWire ), 
        .D(n147), .Clk(_329_net_) );
  Bit_736 \WordArray[9].Word[23].Cell  ( .Q(\WordArray[9].Word[23].QWire ), 
        .D(n149), .Clk(_329_net_) );
  Bit_735 \WordArray[9].Word[24].Cell  ( .Q(\WordArray[9].Word[24].QWire ), 
        .D(n151), .Clk(_329_net_) );
  Bit_734 \WordArray[9].Word[25].Cell  ( .Q(\WordArray[9].Word[25].QWire ), 
        .D(n153), .Clk(_329_net_) );
  Bit_733 \WordArray[9].Word[26].Cell  ( .Q(\WordArray[9].Word[26].QWire ), 
        .D(n155), .Clk(_329_net_) );
  Bit_732 \WordArray[9].Word[27].Cell  ( .Q(\WordArray[9].Word[27].QWire ), 
        .D(n157), .Clk(_329_net_) );
  Bit_731 \WordArray[9].Word[28].Cell  ( .Q(\WordArray[9].Word[28].QWire ), 
        .D(n159), .Clk(_329_net_) );
  Bit_730 \WordArray[9].Word[29].Cell  ( .Q(\WordArray[9].Word[29].QWire ), 
        .D(n161), .Clk(_329_net_) );
  Bit_729 \WordArray[9].Word[30].Cell  ( .Q(\WordArray[9].Word[30].QWire ), 
        .D(n163), .Clk(_329_net_) );
  Bit_728 \WordArray[9].Word[31].Cell  ( .Q(\WordArray[9].Word[31].QWire ), 
        .D(n165), .Clk(_329_net_) );
  Bit_727 \WordArray[9].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _329_net_) );
  Bit_726 \WordArray[10].Word[0].Cell  ( .Q(\WordArray[10].Word[0].QWire ), 
        .D(n103), .Clk(_362_net_) );
  Bit_725 \WordArray[10].Word[1].Cell  ( .Q(\WordArray[10].Word[1].QWire ), 
        .D(n105), .Clk(_362_net_) );
  Bit_724 \WordArray[10].Word[2].Cell  ( .Q(\WordArray[10].Word[2].QWire ), 
        .D(n107), .Clk(_362_net_) );
  Bit_723 \WordArray[10].Word[3].Cell  ( .Q(\WordArray[10].Word[3].QWire ), 
        .D(n109), .Clk(_362_net_) );
  Bit_722 \WordArray[10].Word[4].Cell  ( .Q(\WordArray[10].Word[4].QWire ), 
        .D(n111), .Clk(_362_net_) );
  Bit_721 \WordArray[10].Word[5].Cell  ( .Q(\WordArray[10].Word[5].QWire ), 
        .D(n113), .Clk(_362_net_) );
  Bit_720 \WordArray[10].Word[6].Cell  ( .Q(\WordArray[10].Word[6].QWire ), 
        .D(n115), .Clk(_362_net_) );
  Bit_719 \WordArray[10].Word[7].Cell  ( .Q(\WordArray[10].Word[7].QWire ), 
        .D(n117), .Clk(_362_net_) );
  Bit_718 \WordArray[10].Word[8].Cell  ( .Q(\WordArray[10].Word[8].QWire ), 
        .D(n119), .Clk(_362_net_) );
  Bit_717 \WordArray[10].Word[9].Cell  ( .Q(\WordArray[10].Word[9].QWire ), 
        .D(n121), .Clk(_362_net_) );
  Bit_716 \WordArray[10].Word[10].Cell  ( .Q(\WordArray[10].Word[10].QWire ), 
        .D(n123), .Clk(_362_net_) );
  Bit_715 \WordArray[10].Word[11].Cell  ( .Q(\WordArray[10].Word[11].QWire ), 
        .D(n125), .Clk(_362_net_) );
  Bit_714 \WordArray[10].Word[12].Cell  ( .Q(\WordArray[10].Word[12].QWire ), 
        .D(n127), .Clk(_362_net_) );
  Bit_713 \WordArray[10].Word[13].Cell  ( .Q(\WordArray[10].Word[13].QWire ), 
        .D(n129), .Clk(_362_net_) );
  Bit_712 \WordArray[10].Word[14].Cell  ( .Q(\WordArray[10].Word[14].QWire ), 
        .D(n131), .Clk(_362_net_) );
  Bit_711 \WordArray[10].Word[15].Cell  ( .Q(\WordArray[10].Word[15].QWire ), 
        .D(n133), .Clk(_362_net_) );
  Bit_710 \WordArray[10].Word[16].Cell  ( .Q(\WordArray[10].Word[16].QWire ), 
        .D(n135), .Clk(_362_net_) );
  Bit_709 \WordArray[10].Word[17].Cell  ( .Q(\WordArray[10].Word[17].QWire ), 
        .D(n137), .Clk(_362_net_) );
  Bit_708 \WordArray[10].Word[18].Cell  ( .Q(\WordArray[10].Word[18].QWire ), 
        .D(n139), .Clk(_362_net_) );
  Bit_707 \WordArray[10].Word[19].Cell  ( .Q(\WordArray[10].Word[19].QWire ), 
        .D(n141), .Clk(_362_net_) );
  Bit_706 \WordArray[10].Word[20].Cell  ( .Q(\WordArray[10].Word[20].QWire ), 
        .D(n143), .Clk(_362_net_) );
  Bit_705 \WordArray[10].Word[21].Cell  ( .Q(\WordArray[10].Word[21].QWire ), 
        .D(n145), .Clk(_362_net_) );
  Bit_704 \WordArray[10].Word[22].Cell  ( .Q(\WordArray[10].Word[22].QWire ), 
        .D(n147), .Clk(_362_net_) );
  Bit_703 \WordArray[10].Word[23].Cell  ( .Q(\WordArray[10].Word[23].QWire ), 
        .D(n149), .Clk(_362_net_) );
  Bit_702 \WordArray[10].Word[24].Cell  ( .Q(\WordArray[10].Word[24].QWire ), 
        .D(n151), .Clk(_362_net_) );
  Bit_701 \WordArray[10].Word[25].Cell  ( .Q(\WordArray[10].Word[25].QWire ), 
        .D(n153), .Clk(_362_net_) );
  Bit_700 \WordArray[10].Word[26].Cell  ( .Q(\WordArray[10].Word[26].QWire ), 
        .D(n155), .Clk(_362_net_) );
  Bit_699 \WordArray[10].Word[27].Cell  ( .Q(\WordArray[10].Word[27].QWire ), 
        .D(n157), .Clk(_362_net_) );
  Bit_698 \WordArray[10].Word[28].Cell  ( .Q(\WordArray[10].Word[28].QWire ), 
        .D(n159), .Clk(_362_net_) );
  Bit_697 \WordArray[10].Word[29].Cell  ( .Q(\WordArray[10].Word[29].QWire ), 
        .D(n161), .Clk(_362_net_) );
  Bit_696 \WordArray[10].Word[30].Cell  ( .Q(\WordArray[10].Word[30].QWire ), 
        .D(n163), .Clk(_362_net_) );
  Bit_695 \WordArray[10].Word[31].Cell  ( .Q(\WordArray[10].Word[31].QWire ), 
        .D(n165), .Clk(_362_net_) );
  Bit_694 \WordArray[10].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _362_net_) );
  Bit_693 \WordArray[11].Word[0].Cell  ( .Q(\WordArray[11].Word[0].QWire ), 
        .D(n103), .Clk(_395_net_) );
  Bit_692 \WordArray[11].Word[1].Cell  ( .Q(\WordArray[11].Word[1].QWire ), 
        .D(n105), .Clk(_395_net_) );
  Bit_691 \WordArray[11].Word[2].Cell  ( .Q(\WordArray[11].Word[2].QWire ), 
        .D(DataI[2]), .Clk(_395_net_) );
  Bit_690 \WordArray[11].Word[3].Cell  ( .Q(\WordArray[11].Word[3].QWire ), 
        .D(n109), .Clk(_395_net_) );
  Bit_689 \WordArray[11].Word[4].Cell  ( .Q(\WordArray[11].Word[4].QWire ), 
        .D(n111), .Clk(_395_net_) );
  Bit_688 \WordArray[11].Word[5].Cell  ( .Q(\WordArray[11].Word[5].QWire ), 
        .D(DataI[5]), .Clk(_395_net_) );
  Bit_687 \WordArray[11].Word[6].Cell  ( .Q(\WordArray[11].Word[6].QWire ), 
        .D(n115), .Clk(_395_net_) );
  Bit_686 \WordArray[11].Word[7].Cell  ( .Q(\WordArray[11].Word[7].QWire ), 
        .D(n117), .Clk(_395_net_) );
  Bit_685 \WordArray[11].Word[8].Cell  ( .Q(\WordArray[11].Word[8].QWire ), 
        .D(n119), .Clk(_395_net_) );
  Bit_684 \WordArray[11].Word[9].Cell  ( .Q(\WordArray[11].Word[9].QWire ), 
        .D(n121), .Clk(_395_net_) );
  Bit_683 \WordArray[11].Word[10].Cell  ( .Q(\WordArray[11].Word[10].QWire ), 
        .D(n123), .Clk(_395_net_) );
  Bit_682 \WordArray[11].Word[11].Cell  ( .Q(\WordArray[11].Word[11].QWire ), 
        .D(n125), .Clk(_395_net_) );
  Bit_681 \WordArray[11].Word[12].Cell  ( .Q(\WordArray[11].Word[12].QWire ), 
        .D(n127), .Clk(_395_net_) );
  Bit_680 \WordArray[11].Word[13].Cell  ( .Q(\WordArray[11].Word[13].QWire ), 
        .D(n129), .Clk(_395_net_) );
  Bit_679 \WordArray[11].Word[14].Cell  ( .Q(\WordArray[11].Word[14].QWire ), 
        .D(n131), .Clk(_395_net_) );
  Bit_678 \WordArray[11].Word[15].Cell  ( .Q(\WordArray[11].Word[15].QWire ), 
        .D(n133), .Clk(_395_net_) );
  Bit_677 \WordArray[11].Word[16].Cell  ( .Q(\WordArray[11].Word[16].QWire ), 
        .D(n135), .Clk(_395_net_) );
  Bit_676 \WordArray[11].Word[17].Cell  ( .Q(\WordArray[11].Word[17].QWire ), 
        .D(n137), .Clk(_395_net_) );
  Bit_675 \WordArray[11].Word[18].Cell  ( .Q(\WordArray[11].Word[18].QWire ), 
        .D(n139), .Clk(_395_net_) );
  Bit_674 \WordArray[11].Word[19].Cell  ( .Q(\WordArray[11].Word[19].QWire ), 
        .D(n141), .Clk(_395_net_) );
  Bit_673 \WordArray[11].Word[20].Cell  ( .Q(\WordArray[11].Word[20].QWire ), 
        .D(n143), .Clk(_395_net_) );
  Bit_672 \WordArray[11].Word[21].Cell  ( .Q(\WordArray[11].Word[21].QWire ), 
        .D(n145), .Clk(_395_net_) );
  Bit_671 \WordArray[11].Word[22].Cell  ( .Q(\WordArray[11].Word[22].QWire ), 
        .D(n147), .Clk(_395_net_) );
  Bit_670 \WordArray[11].Word[23].Cell  ( .Q(\WordArray[11].Word[23].QWire ), 
        .D(n149), .Clk(_395_net_) );
  Bit_669 \WordArray[11].Word[24].Cell  ( .Q(\WordArray[11].Word[24].QWire ), 
        .D(n151), .Clk(_395_net_) );
  Bit_668 \WordArray[11].Word[25].Cell  ( .Q(\WordArray[11].Word[25].QWire ), 
        .D(n153), .Clk(_395_net_) );
  Bit_667 \WordArray[11].Word[26].Cell  ( .Q(\WordArray[11].Word[26].QWire ), 
        .D(n155), .Clk(_395_net_) );
  Bit_666 \WordArray[11].Word[27].Cell  ( .Q(\WordArray[11].Word[27].QWire ), 
        .D(n157), .Clk(_395_net_) );
  Bit_665 \WordArray[11].Word[28].Cell  ( .Q(\WordArray[11].Word[28].QWire ), 
        .D(n159), .Clk(_395_net_) );
  Bit_664 \WordArray[11].Word[29].Cell  ( .Q(\WordArray[11].Word[29].QWire ), 
        .D(n161), .Clk(_395_net_) );
  Bit_663 \WordArray[11].Word[30].Cell  ( .Q(\WordArray[11].Word[30].QWire ), 
        .D(n163), .Clk(_395_net_) );
  Bit_662 \WordArray[11].Word[31].Cell  ( .Q(\WordArray[11].Word[31].QWire ), 
        .D(n165), .Clk(_395_net_) );
  Bit_661 \WordArray[11].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _395_net_) );
  Bit_660 \WordArray[12].Word[0].Cell  ( .Q(\WordArray[12].Word[0].QWire ), 
        .D(DataI[0]), .Clk(_428_net_) );
  Bit_659 \WordArray[12].Word[1].Cell  ( .Q(\WordArray[12].Word[1].QWire ), 
        .D(n105), .Clk(_428_net_) );
  Bit_658 \WordArray[12].Word[2].Cell  ( .Q(\WordArray[12].Word[2].QWire ), 
        .D(n107), .Clk(_428_net_) );
  Bit_657 \WordArray[12].Word[3].Cell  ( .Q(\WordArray[12].Word[3].QWire ), 
        .D(n109), .Clk(_428_net_) );
  Bit_656 \WordArray[12].Word[4].Cell  ( .Q(\WordArray[12].Word[4].QWire ), 
        .D(n111), .Clk(_428_net_) );
  Bit_655 \WordArray[12].Word[5].Cell  ( .Q(\WordArray[12].Word[5].QWire ), 
        .D(n113), .Clk(_428_net_) );
  Bit_654 \WordArray[12].Word[6].Cell  ( .Q(\WordArray[12].Word[6].QWire ), 
        .D(n115), .Clk(_428_net_) );
  Bit_653 \WordArray[12].Word[7].Cell  ( .Q(\WordArray[12].Word[7].QWire ), 
        .D(n117), .Clk(_428_net_) );
  Bit_652 \WordArray[12].Word[8].Cell  ( .Q(\WordArray[12].Word[8].QWire ), 
        .D(n119), .Clk(_428_net_) );
  Bit_651 \WordArray[12].Word[9].Cell  ( .Q(\WordArray[12].Word[9].QWire ), 
        .D(n121), .Clk(_428_net_) );
  Bit_650 \WordArray[12].Word[10].Cell  ( .Q(\WordArray[12].Word[10].QWire ), 
        .D(n123), .Clk(_428_net_) );
  Bit_649 \WordArray[12].Word[11].Cell  ( .Q(\WordArray[12].Word[11].QWire ), 
        .D(n125), .Clk(_428_net_) );
  Bit_648 \WordArray[12].Word[12].Cell  ( .Q(\WordArray[12].Word[12].QWire ), 
        .D(n127), .Clk(_428_net_) );
  Bit_647 \WordArray[12].Word[13].Cell  ( .Q(\WordArray[12].Word[13].QWire ), 
        .D(n129), .Clk(_428_net_) );
  Bit_646 \WordArray[12].Word[14].Cell  ( .Q(\WordArray[12].Word[14].QWire ), 
        .D(n131), .Clk(_428_net_) );
  Bit_645 \WordArray[12].Word[15].Cell  ( .Q(\WordArray[12].Word[15].QWire ), 
        .D(n133), .Clk(_428_net_) );
  Bit_644 \WordArray[12].Word[16].Cell  ( .Q(\WordArray[12].Word[16].QWire ), 
        .D(n135), .Clk(_428_net_) );
  Bit_643 \WordArray[12].Word[17].Cell  ( .Q(\WordArray[12].Word[17].QWire ), 
        .D(n137), .Clk(_428_net_) );
  Bit_642 \WordArray[12].Word[18].Cell  ( .Q(\WordArray[12].Word[18].QWire ), 
        .D(n139), .Clk(_428_net_) );
  Bit_641 \WordArray[12].Word[19].Cell  ( .Q(\WordArray[12].Word[19].QWire ), 
        .D(n141), .Clk(_428_net_) );
  Bit_640 \WordArray[12].Word[20].Cell  ( .Q(\WordArray[12].Word[20].QWire ), 
        .D(n143), .Clk(_428_net_) );
  Bit_639 \WordArray[12].Word[21].Cell  ( .Q(\WordArray[12].Word[21].QWire ), 
        .D(n145), .Clk(_428_net_) );
  Bit_638 \WordArray[12].Word[22].Cell  ( .Q(\WordArray[12].Word[22].QWire ), 
        .D(n147), .Clk(_428_net_) );
  Bit_637 \WordArray[12].Word[23].Cell  ( .Q(\WordArray[12].Word[23].QWire ), 
        .D(n149), .Clk(_428_net_) );
  Bit_636 \WordArray[12].Word[24].Cell  ( .Q(\WordArray[12].Word[24].QWire ), 
        .D(n151), .Clk(_428_net_) );
  Bit_635 \WordArray[12].Word[25].Cell  ( .Q(\WordArray[12].Word[25].QWire ), 
        .D(n153), .Clk(_428_net_) );
  Bit_634 \WordArray[12].Word[26].Cell  ( .Q(\WordArray[12].Word[26].QWire ), 
        .D(n155), .Clk(_428_net_) );
  Bit_633 \WordArray[12].Word[27].Cell  ( .Q(\WordArray[12].Word[27].QWire ), 
        .D(n157), .Clk(_428_net_) );
  Bit_632 \WordArray[12].Word[28].Cell  ( .Q(\WordArray[12].Word[28].QWire ), 
        .D(n159), .Clk(_428_net_) );
  Bit_631 \WordArray[12].Word[29].Cell  ( .Q(\WordArray[12].Word[29].QWire ), 
        .D(n161), .Clk(_428_net_) );
  Bit_630 \WordArray[12].Word[30].Cell  ( .Q(\WordArray[12].Word[30].QWire ), 
        .D(n163), .Clk(_428_net_) );
  Bit_629 \WordArray[12].Word[31].Cell  ( .Q(\WordArray[12].Word[31].QWire ), 
        .D(n165), .Clk(_428_net_) );
  Bit_628 \WordArray[12].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _428_net_) );
  Bit_627 \WordArray[13].Word[0].Cell  ( .Q(\WordArray[13].Word[0].QWire ), 
        .D(n103), .Clk(_461_net_) );
  Bit_626 \WordArray[13].Word[1].Cell  ( .Q(\WordArray[13].Word[1].QWire ), 
        .D(n105), .Clk(_461_net_) );
  Bit_625 \WordArray[13].Word[2].Cell  ( .Q(\WordArray[13].Word[2].QWire ), 
        .D(n107), .Clk(_461_net_) );
  Bit_624 \WordArray[13].Word[3].Cell  ( .Q(\WordArray[13].Word[3].QWire ), 
        .D(n109), .Clk(_461_net_) );
  Bit_623 \WordArray[13].Word[4].Cell  ( .Q(\WordArray[13].Word[4].QWire ), 
        .D(n111), .Clk(_461_net_) );
  Bit_622 \WordArray[13].Word[5].Cell  ( .Q(\WordArray[13].Word[5].QWire ), 
        .D(n113), .Clk(_461_net_) );
  Bit_621 \WordArray[13].Word[6].Cell  ( .Q(\WordArray[13].Word[6].QWire ), 
        .D(n115), .Clk(_461_net_) );
  Bit_620 \WordArray[13].Word[7].Cell  ( .Q(\WordArray[13].Word[7].QWire ), 
        .D(n117), .Clk(_461_net_) );
  Bit_619 \WordArray[13].Word[8].Cell  ( .Q(\WordArray[13].Word[8].QWire ), 
        .D(n119), .Clk(_461_net_) );
  Bit_618 \WordArray[13].Word[9].Cell  ( .Q(\WordArray[13].Word[9].QWire ), 
        .D(n121), .Clk(_461_net_) );
  Bit_617 \WordArray[13].Word[10].Cell  ( .Q(\WordArray[13].Word[10].QWire ), 
        .D(n123), .Clk(_461_net_) );
  Bit_616 \WordArray[13].Word[11].Cell  ( .Q(\WordArray[13].Word[11].QWire ), 
        .D(n125), .Clk(_461_net_) );
  Bit_615 \WordArray[13].Word[12].Cell  ( .Q(\WordArray[13].Word[12].QWire ), 
        .D(n127), .Clk(_461_net_) );
  Bit_614 \WordArray[13].Word[13].Cell  ( .Q(\WordArray[13].Word[13].QWire ), 
        .D(n129), .Clk(_461_net_) );
  Bit_613 \WordArray[13].Word[14].Cell  ( .Q(\WordArray[13].Word[14].QWire ), 
        .D(n131), .Clk(_461_net_) );
  Bit_612 \WordArray[13].Word[15].Cell  ( .Q(\WordArray[13].Word[15].QWire ), 
        .D(n133), .Clk(_461_net_) );
  Bit_611 \WordArray[13].Word[16].Cell  ( .Q(\WordArray[13].Word[16].QWire ), 
        .D(n135), .Clk(_461_net_) );
  Bit_610 \WordArray[13].Word[17].Cell  ( .Q(\WordArray[13].Word[17].QWire ), 
        .D(n137), .Clk(_461_net_) );
  Bit_609 \WordArray[13].Word[18].Cell  ( .Q(\WordArray[13].Word[18].QWire ), 
        .D(n139), .Clk(_461_net_) );
  Bit_608 \WordArray[13].Word[19].Cell  ( .Q(\WordArray[13].Word[19].QWire ), 
        .D(n141), .Clk(_461_net_) );
  Bit_607 \WordArray[13].Word[20].Cell  ( .Q(\WordArray[13].Word[20].QWire ), 
        .D(n143), .Clk(_461_net_) );
  Bit_606 \WordArray[13].Word[21].Cell  ( .Q(\WordArray[13].Word[21].QWire ), 
        .D(n145), .Clk(_461_net_) );
  Bit_605 \WordArray[13].Word[22].Cell  ( .Q(\WordArray[13].Word[22].QWire ), 
        .D(n147), .Clk(_461_net_) );
  Bit_604 \WordArray[13].Word[23].Cell  ( .Q(\WordArray[13].Word[23].QWire ), 
        .D(n149), .Clk(_461_net_) );
  Bit_603 \WordArray[13].Word[24].Cell  ( .Q(\WordArray[13].Word[24].QWire ), 
        .D(n151), .Clk(_461_net_) );
  Bit_602 \WordArray[13].Word[25].Cell  ( .Q(\WordArray[13].Word[25].QWire ), 
        .D(n153), .Clk(_461_net_) );
  Bit_601 \WordArray[13].Word[26].Cell  ( .Q(\WordArray[13].Word[26].QWire ), 
        .D(n155), .Clk(_461_net_) );
  Bit_600 \WordArray[13].Word[27].Cell  ( .Q(\WordArray[13].Word[27].QWire ), 
        .D(n157), .Clk(_461_net_) );
  Bit_599 \WordArray[13].Word[28].Cell  ( .Q(\WordArray[13].Word[28].QWire ), 
        .D(n159), .Clk(_461_net_) );
  Bit_598 \WordArray[13].Word[29].Cell  ( .Q(\WordArray[13].Word[29].QWire ), 
        .D(n161), .Clk(_461_net_) );
  Bit_597 \WordArray[13].Word[30].Cell  ( .Q(\WordArray[13].Word[30].QWire ), 
        .D(n163), .Clk(_461_net_) );
  Bit_596 \WordArray[13].Word[31].Cell  ( .Q(\WordArray[13].Word[31].QWire ), 
        .D(n165), .Clk(_461_net_) );
  Bit_595 \WordArray[13].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _461_net_) );
  Bit_594 \WordArray[14].Word[0].Cell  ( .Q(\WordArray[14].Word[0].QWire ), 
        .D(n103), .Clk(_494_net_) );
  Bit_593 \WordArray[14].Word[1].Cell  ( .Q(\WordArray[14].Word[1].QWire ), 
        .D(n105), .Clk(_494_net_) );
  Bit_592 \WordArray[14].Word[2].Cell  ( .Q(\WordArray[14].Word[2].QWire ), 
        .D(n107), .Clk(_494_net_) );
  Bit_591 \WordArray[14].Word[3].Cell  ( .Q(\WordArray[14].Word[3].QWire ), 
        .D(n109), .Clk(_494_net_) );
  Bit_590 \WordArray[14].Word[4].Cell  ( .Q(\WordArray[14].Word[4].QWire ), 
        .D(n111), .Clk(_494_net_) );
  Bit_589 \WordArray[14].Word[5].Cell  ( .Q(\WordArray[14].Word[5].QWire ), 
        .D(n113), .Clk(_494_net_) );
  Bit_588 \WordArray[14].Word[6].Cell  ( .Q(\WordArray[14].Word[6].QWire ), 
        .D(n115), .Clk(_494_net_) );
  Bit_587 \WordArray[14].Word[7].Cell  ( .Q(\WordArray[14].Word[7].QWire ), 
        .D(n117), .Clk(_494_net_) );
  Bit_586 \WordArray[14].Word[8].Cell  ( .Q(\WordArray[14].Word[8].QWire ), 
        .D(n119), .Clk(_494_net_) );
  Bit_585 \WordArray[14].Word[9].Cell  ( .Q(\WordArray[14].Word[9].QWire ), 
        .D(n121), .Clk(_494_net_) );
  Bit_584 \WordArray[14].Word[10].Cell  ( .Q(\WordArray[14].Word[10].QWire ), 
        .D(n123), .Clk(_494_net_) );
  Bit_583 \WordArray[14].Word[11].Cell  ( .Q(\WordArray[14].Word[11].QWire ), 
        .D(n125), .Clk(_494_net_) );
  Bit_582 \WordArray[14].Word[12].Cell  ( .Q(\WordArray[14].Word[12].QWire ), 
        .D(n127), .Clk(_494_net_) );
  Bit_581 \WordArray[14].Word[13].Cell  ( .Q(\WordArray[14].Word[13].QWire ), 
        .D(n129), .Clk(_494_net_) );
  Bit_580 \WordArray[14].Word[14].Cell  ( .Q(\WordArray[14].Word[14].QWire ), 
        .D(n131), .Clk(_494_net_) );
  Bit_579 \WordArray[14].Word[15].Cell  ( .Q(\WordArray[14].Word[15].QWire ), 
        .D(n133), .Clk(_494_net_) );
  Bit_578 \WordArray[14].Word[16].Cell  ( .Q(\WordArray[14].Word[16].QWire ), 
        .D(n135), .Clk(_494_net_) );
  Bit_577 \WordArray[14].Word[17].Cell  ( .Q(\WordArray[14].Word[17].QWire ), 
        .D(n137), .Clk(_494_net_) );
  Bit_576 \WordArray[14].Word[18].Cell  ( .Q(\WordArray[14].Word[18].QWire ), 
        .D(n139), .Clk(_494_net_) );
  Bit_575 \WordArray[14].Word[19].Cell  ( .Q(\WordArray[14].Word[19].QWire ), 
        .D(n141), .Clk(_494_net_) );
  Bit_574 \WordArray[14].Word[20].Cell  ( .Q(\WordArray[14].Word[20].QWire ), 
        .D(n143), .Clk(_494_net_) );
  Bit_573 \WordArray[14].Word[21].Cell  ( .Q(\WordArray[14].Word[21].QWire ), 
        .D(n145), .Clk(_494_net_) );
  Bit_572 \WordArray[14].Word[22].Cell  ( .Q(\WordArray[14].Word[22].QWire ), 
        .D(n147), .Clk(_494_net_) );
  Bit_571 \WordArray[14].Word[23].Cell  ( .Q(\WordArray[14].Word[23].QWire ), 
        .D(n149), .Clk(_494_net_) );
  Bit_570 \WordArray[14].Word[24].Cell  ( .Q(\WordArray[14].Word[24].QWire ), 
        .D(n151), .Clk(_494_net_) );
  Bit_569 \WordArray[14].Word[25].Cell  ( .Q(\WordArray[14].Word[25].QWire ), 
        .D(n153), .Clk(_494_net_) );
  Bit_568 \WordArray[14].Word[26].Cell  ( .Q(\WordArray[14].Word[26].QWire ), 
        .D(n155), .Clk(_494_net_) );
  Bit_567 \WordArray[14].Word[27].Cell  ( .Q(\WordArray[14].Word[27].QWire ), 
        .D(n157), .Clk(_494_net_) );
  Bit_566 \WordArray[14].Word[28].Cell  ( .Q(\WordArray[14].Word[28].QWire ), 
        .D(n159), .Clk(_494_net_) );
  Bit_565 \WordArray[14].Word[29].Cell  ( .Q(\WordArray[14].Word[29].QWire ), 
        .D(n161), .Clk(_494_net_) );
  Bit_564 \WordArray[14].Word[30].Cell  ( .Q(\WordArray[14].Word[30].QWire ), 
        .D(n163), .Clk(_494_net_) );
  Bit_563 \WordArray[14].Word[31].Cell  ( .Q(\WordArray[14].Word[31].QWire ), 
        .D(n165), .Clk(_494_net_) );
  Bit_562 \WordArray[14].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _494_net_) );
  Bit_561 \WordArray[15].Word[0].Cell  ( .Q(\WordArray[15].Word[0].QWire ), 
        .D(n103), .Clk(_527_net_) );
  Bit_560 \WordArray[15].Word[1].Cell  ( .Q(\WordArray[15].Word[1].QWire ), 
        .D(n105), .Clk(_527_net_) );
  Bit_559 \WordArray[15].Word[2].Cell  ( .Q(\WordArray[15].Word[2].QWire ), 
        .D(n107), .Clk(_527_net_) );
  Bit_558 \WordArray[15].Word[3].Cell  ( .Q(\WordArray[15].Word[3].QWire ), 
        .D(n109), .Clk(_527_net_) );
  Bit_557 \WordArray[15].Word[4].Cell  ( .Q(\WordArray[15].Word[4].QWire ), 
        .D(n111), .Clk(_527_net_) );
  Bit_556 \WordArray[15].Word[5].Cell  ( .Q(\WordArray[15].Word[5].QWire ), 
        .D(n113), .Clk(_527_net_) );
  Bit_555 \WordArray[15].Word[6].Cell  ( .Q(\WordArray[15].Word[6].QWire ), 
        .D(n115), .Clk(_527_net_) );
  Bit_554 \WordArray[15].Word[7].Cell  ( .Q(\WordArray[15].Word[7].QWire ), 
        .D(n117), .Clk(_527_net_) );
  Bit_553 \WordArray[15].Word[8].Cell  ( .Q(\WordArray[15].Word[8].QWire ), 
        .D(n119), .Clk(_527_net_) );
  Bit_552 \WordArray[15].Word[9].Cell  ( .Q(\WordArray[15].Word[9].QWire ), 
        .D(n121), .Clk(_527_net_) );
  Bit_551 \WordArray[15].Word[10].Cell  ( .Q(\WordArray[15].Word[10].QWire ), 
        .D(n123), .Clk(_527_net_) );
  Bit_550 \WordArray[15].Word[11].Cell  ( .Q(\WordArray[15].Word[11].QWire ), 
        .D(n125), .Clk(_527_net_) );
  Bit_549 \WordArray[15].Word[12].Cell  ( .Q(\WordArray[15].Word[12].QWire ), 
        .D(n127), .Clk(_527_net_) );
  Bit_548 \WordArray[15].Word[13].Cell  ( .Q(\WordArray[15].Word[13].QWire ), 
        .D(n129), .Clk(_527_net_) );
  Bit_547 \WordArray[15].Word[14].Cell  ( .Q(\WordArray[15].Word[14].QWire ), 
        .D(n131), .Clk(_527_net_) );
  Bit_546 \WordArray[15].Word[15].Cell  ( .Q(\WordArray[15].Word[15].QWire ), 
        .D(n133), .Clk(_527_net_) );
  Bit_545 \WordArray[15].Word[16].Cell  ( .Q(\WordArray[15].Word[16].QWire ), 
        .D(n135), .Clk(_527_net_) );
  Bit_544 \WordArray[15].Word[17].Cell  ( .Q(\WordArray[15].Word[17].QWire ), 
        .D(n137), .Clk(_527_net_) );
  Bit_543 \WordArray[15].Word[18].Cell  ( .Q(\WordArray[15].Word[18].QWire ), 
        .D(n139), .Clk(_527_net_) );
  Bit_542 \WordArray[15].Word[19].Cell  ( .Q(\WordArray[15].Word[19].QWire ), 
        .D(n141), .Clk(_527_net_) );
  Bit_541 \WordArray[15].Word[20].Cell  ( .Q(\WordArray[15].Word[20].QWire ), 
        .D(n143), .Clk(_527_net_) );
  Bit_540 \WordArray[15].Word[21].Cell  ( .Q(\WordArray[15].Word[21].QWire ), 
        .D(n145), .Clk(_527_net_) );
  Bit_539 \WordArray[15].Word[22].Cell  ( .Q(\WordArray[15].Word[22].QWire ), 
        .D(n147), .Clk(_527_net_) );
  Bit_538 \WordArray[15].Word[23].Cell  ( .Q(\WordArray[15].Word[23].QWire ), 
        .D(n149), .Clk(_527_net_) );
  Bit_537 \WordArray[15].Word[24].Cell  ( .Q(\WordArray[15].Word[24].QWire ), 
        .D(n151), .Clk(_527_net_) );
  Bit_536 \WordArray[15].Word[25].Cell  ( .Q(\WordArray[15].Word[25].QWire ), 
        .D(n153), .Clk(_527_net_) );
  Bit_535 \WordArray[15].Word[26].Cell  ( .Q(\WordArray[15].Word[26].QWire ), 
        .D(n155), .Clk(_527_net_) );
  Bit_534 \WordArray[15].Word[27].Cell  ( .Q(\WordArray[15].Word[27].QWire ), 
        .D(n157), .Clk(_527_net_) );
  Bit_533 \WordArray[15].Word[28].Cell  ( .Q(\WordArray[15].Word[28].QWire ), 
        .D(n159), .Clk(_527_net_) );
  Bit_532 \WordArray[15].Word[29].Cell  ( .Q(\WordArray[15].Word[29].QWire ), 
        .D(n161), .Clk(_527_net_) );
  Bit_531 \WordArray[15].Word[30].Cell  ( .Q(\WordArray[15].Word[30].QWire ), 
        .D(n163), .Clk(_527_net_) );
  Bit_530 \WordArray[15].Word[31].Cell  ( .Q(\WordArray[15].Word[31].QWire ), 
        .D(n165), .Clk(_527_net_) );
  Bit_529 \WordArray[15].Word[32].Cell  ( .D(n34), .Clk(_527_net_) );
  Bit_528 \WordArray[16].Word[0].Cell  ( .Q(\WordArray[16].Word[0].QWire ), 
        .D(n103), .Clk(_560_net_) );
  Bit_527 \WordArray[16].Word[1].Cell  ( .Q(\WordArray[16].Word[1].QWire ), 
        .D(n105), .Clk(_560_net_) );
  Bit_526 \WordArray[16].Word[2].Cell  ( .Q(\WordArray[16].Word[2].QWire ), 
        .D(n107), .Clk(_560_net_) );
  Bit_525 \WordArray[16].Word[3].Cell  ( .Q(\WordArray[16].Word[3].QWire ), 
        .D(n109), .Clk(_560_net_) );
  Bit_524 \WordArray[16].Word[4].Cell  ( .Q(\WordArray[16].Word[4].QWire ), 
        .D(n111), .Clk(_560_net_) );
  Bit_523 \WordArray[16].Word[5].Cell  ( .Q(\WordArray[16].Word[5].QWire ), 
        .D(n113), .Clk(_560_net_) );
  Bit_522 \WordArray[16].Word[6].Cell  ( .Q(\WordArray[16].Word[6].QWire ), 
        .D(n115), .Clk(_560_net_) );
  Bit_521 \WordArray[16].Word[7].Cell  ( .Q(\WordArray[16].Word[7].QWire ), 
        .D(n117), .Clk(_560_net_) );
  Bit_520 \WordArray[16].Word[8].Cell  ( .Q(\WordArray[16].Word[8].QWire ), 
        .D(n119), .Clk(_560_net_) );
  Bit_519 \WordArray[16].Word[9].Cell  ( .Q(\WordArray[16].Word[9].QWire ), 
        .D(n121), .Clk(_560_net_) );
  Bit_518 \WordArray[16].Word[10].Cell  ( .Q(\WordArray[16].Word[10].QWire ), 
        .D(n123), .Clk(_560_net_) );
  Bit_517 \WordArray[16].Word[11].Cell  ( .Q(\WordArray[16].Word[11].QWire ), 
        .D(n125), .Clk(_560_net_) );
  Bit_516 \WordArray[16].Word[12].Cell  ( .Q(\WordArray[16].Word[12].QWire ), 
        .D(n127), .Clk(_560_net_) );
  Bit_515 \WordArray[16].Word[13].Cell  ( .Q(\WordArray[16].Word[13].QWire ), 
        .D(n129), .Clk(_560_net_) );
  Bit_514 \WordArray[16].Word[14].Cell  ( .Q(\WordArray[16].Word[14].QWire ), 
        .D(n131), .Clk(_560_net_) );
  Bit_513 \WordArray[16].Word[15].Cell  ( .Q(\WordArray[16].Word[15].QWire ), 
        .D(n133), .Clk(_560_net_) );
  Bit_512 \WordArray[16].Word[16].Cell  ( .Q(\WordArray[16].Word[16].QWire ), 
        .D(n135), .Clk(_560_net_) );
  Bit_511 \WordArray[16].Word[17].Cell  ( .Q(\WordArray[16].Word[17].QWire ), 
        .D(n137), .Clk(_560_net_) );
  Bit_510 \WordArray[16].Word[18].Cell  ( .Q(\WordArray[16].Word[18].QWire ), 
        .D(n139), .Clk(_560_net_) );
  Bit_509 \WordArray[16].Word[19].Cell  ( .Q(\WordArray[16].Word[19].QWire ), 
        .D(n141), .Clk(_560_net_) );
  Bit_508 \WordArray[16].Word[20].Cell  ( .Q(\WordArray[16].Word[20].QWire ), 
        .D(n143), .Clk(_560_net_) );
  Bit_507 \WordArray[16].Word[21].Cell  ( .Q(\WordArray[16].Word[21].QWire ), 
        .D(n145), .Clk(_560_net_) );
  Bit_506 \WordArray[16].Word[22].Cell  ( .Q(\WordArray[16].Word[22].QWire ), 
        .D(n147), .Clk(_560_net_) );
  Bit_505 \WordArray[16].Word[23].Cell  ( .Q(\WordArray[16].Word[23].QWire ), 
        .D(n149), .Clk(_560_net_) );
  Bit_504 \WordArray[16].Word[24].Cell  ( .Q(\WordArray[16].Word[24].QWire ), 
        .D(n151), .Clk(_560_net_) );
  Bit_503 \WordArray[16].Word[25].Cell  ( .Q(\WordArray[16].Word[25].QWire ), 
        .D(n153), .Clk(_560_net_) );
  Bit_502 \WordArray[16].Word[26].Cell  ( .Q(\WordArray[16].Word[26].QWire ), 
        .D(n155), .Clk(_560_net_) );
  Bit_501 \WordArray[16].Word[27].Cell  ( .Q(\WordArray[16].Word[27].QWire ), 
        .D(n157), .Clk(_560_net_) );
  Bit_500 \WordArray[16].Word[28].Cell  ( .Q(\WordArray[16].Word[28].QWire ), 
        .D(n159), .Clk(_560_net_) );
  Bit_499 \WordArray[16].Word[29].Cell  ( .Q(\WordArray[16].Word[29].QWire ), 
        .D(n161), .Clk(_560_net_) );
  Bit_498 \WordArray[16].Word[30].Cell  ( .Q(\WordArray[16].Word[30].QWire ), 
        .D(n163), .Clk(_560_net_) );
  Bit_497 \WordArray[16].Word[31].Cell  ( .Q(\WordArray[16].Word[31].QWire ), 
        .D(n165), .Clk(_560_net_) );
  Bit_496 \WordArray[16].Word[32].Cell  ( .D(n34), .Clk(_560_net_) );
  Bit_495 \WordArray[17].Word[0].Cell  ( .Q(\WordArray[17].Word[0].QWire ), 
        .D(n103), .Clk(_593_net_) );
  Bit_494 \WordArray[17].Word[1].Cell  ( .Q(\WordArray[17].Word[1].QWire ), 
        .D(n105), .Clk(_593_net_) );
  Bit_493 \WordArray[17].Word[2].Cell  ( .Q(\WordArray[17].Word[2].QWire ), 
        .D(n107), .Clk(_593_net_) );
  Bit_492 \WordArray[17].Word[3].Cell  ( .Q(\WordArray[17].Word[3].QWire ), 
        .D(n109), .Clk(_593_net_) );
  Bit_491 \WordArray[17].Word[4].Cell  ( .Q(\WordArray[17].Word[4].QWire ), 
        .D(n111), .Clk(_593_net_) );
  Bit_490 \WordArray[17].Word[5].Cell  ( .Q(\WordArray[17].Word[5].QWire ), 
        .D(n113), .Clk(_593_net_) );
  Bit_489 \WordArray[17].Word[6].Cell  ( .Q(\WordArray[17].Word[6].QWire ), 
        .D(n115), .Clk(_593_net_) );
  Bit_488 \WordArray[17].Word[7].Cell  ( .Q(\WordArray[17].Word[7].QWire ), 
        .D(n117), .Clk(_593_net_) );
  Bit_487 \WordArray[17].Word[8].Cell  ( .Q(\WordArray[17].Word[8].QWire ), 
        .D(n119), .Clk(_593_net_) );
  Bit_486 \WordArray[17].Word[9].Cell  ( .Q(\WordArray[17].Word[9].QWire ), 
        .D(n121), .Clk(_593_net_) );
  Bit_485 \WordArray[17].Word[10].Cell  ( .Q(\WordArray[17].Word[10].QWire ), 
        .D(n123), .Clk(_593_net_) );
  Bit_484 \WordArray[17].Word[11].Cell  ( .Q(\WordArray[17].Word[11].QWire ), 
        .D(n125), .Clk(_593_net_) );
  Bit_483 \WordArray[17].Word[12].Cell  ( .Q(\WordArray[17].Word[12].QWire ), 
        .D(n127), .Clk(_593_net_) );
  Bit_482 \WordArray[17].Word[13].Cell  ( .Q(\WordArray[17].Word[13].QWire ), 
        .D(n129), .Clk(_593_net_) );
  Bit_481 \WordArray[17].Word[14].Cell  ( .Q(\WordArray[17].Word[14].QWire ), 
        .D(n131), .Clk(_593_net_) );
  Bit_480 \WordArray[17].Word[15].Cell  ( .Q(\WordArray[17].Word[15].QWire ), 
        .D(n133), .Clk(_593_net_) );
  Bit_479 \WordArray[17].Word[16].Cell  ( .Q(\WordArray[17].Word[16].QWire ), 
        .D(n135), .Clk(_593_net_) );
  Bit_478 \WordArray[17].Word[17].Cell  ( .Q(\WordArray[17].Word[17].QWire ), 
        .D(n137), .Clk(_593_net_) );
  Bit_477 \WordArray[17].Word[18].Cell  ( .Q(\WordArray[17].Word[18].QWire ), 
        .D(n139), .Clk(_593_net_) );
  Bit_476 \WordArray[17].Word[19].Cell  ( .Q(\WordArray[17].Word[19].QWire ), 
        .D(n141), .Clk(_593_net_) );
  Bit_475 \WordArray[17].Word[20].Cell  ( .Q(\WordArray[17].Word[20].QWire ), 
        .D(n143), .Clk(_593_net_) );
  Bit_474 \WordArray[17].Word[21].Cell  ( .Q(\WordArray[17].Word[21].QWire ), 
        .D(n145), .Clk(_593_net_) );
  Bit_473 \WordArray[17].Word[22].Cell  ( .Q(\WordArray[17].Word[22].QWire ), 
        .D(n147), .Clk(_593_net_) );
  Bit_472 \WordArray[17].Word[23].Cell  ( .Q(\WordArray[17].Word[23].QWire ), 
        .D(n149), .Clk(_593_net_) );
  Bit_471 \WordArray[17].Word[24].Cell  ( .Q(\WordArray[17].Word[24].QWire ), 
        .D(n151), .Clk(_593_net_) );
  Bit_470 \WordArray[17].Word[25].Cell  ( .Q(\WordArray[17].Word[25].QWire ), 
        .D(n153), .Clk(_593_net_) );
  Bit_469 \WordArray[17].Word[26].Cell  ( .Q(\WordArray[17].Word[26].QWire ), 
        .D(n155), .Clk(_593_net_) );
  Bit_468 \WordArray[17].Word[27].Cell  ( .Q(\WordArray[17].Word[27].QWire ), 
        .D(n157), .Clk(_593_net_) );
  Bit_467 \WordArray[17].Word[28].Cell  ( .Q(\WordArray[17].Word[28].QWire ), 
        .D(n159), .Clk(_593_net_) );
  Bit_466 \WordArray[17].Word[29].Cell  ( .Q(\WordArray[17].Word[29].QWire ), 
        .D(n161), .Clk(_593_net_) );
  Bit_465 \WordArray[17].Word[30].Cell  ( .Q(\WordArray[17].Word[30].QWire ), 
        .D(n163), .Clk(_593_net_) );
  Bit_464 \WordArray[17].Word[31].Cell  ( .Q(\WordArray[17].Word[31].QWire ), 
        .D(n165), .Clk(_593_net_) );
  Bit_463 \WordArray[17].Word[32].Cell  ( .D(n34), .Clk(_593_net_) );
  Bit_462 \WordArray[18].Word[0].Cell  ( .Q(\WordArray[18].Word[0].QWire ), 
        .D(n103), .Clk(_626_net_) );
  Bit_461 \WordArray[18].Word[1].Cell  ( .Q(\WordArray[18].Word[1].QWire ), 
        .D(n105), .Clk(_626_net_) );
  Bit_460 \WordArray[18].Word[2].Cell  ( .Q(\WordArray[18].Word[2].QWire ), 
        .D(n107), .Clk(_626_net_) );
  Bit_459 \WordArray[18].Word[3].Cell  ( .Q(\WordArray[18].Word[3].QWire ), 
        .D(n109), .Clk(_626_net_) );
  Bit_458 \WordArray[18].Word[4].Cell  ( .Q(\WordArray[18].Word[4].QWire ), 
        .D(n111), .Clk(_626_net_) );
  Bit_457 \WordArray[18].Word[5].Cell  ( .Q(\WordArray[18].Word[5].QWire ), 
        .D(n113), .Clk(_626_net_) );
  Bit_456 \WordArray[18].Word[6].Cell  ( .Q(\WordArray[18].Word[6].QWire ), 
        .D(n115), .Clk(_626_net_) );
  Bit_455 \WordArray[18].Word[7].Cell  ( .Q(\WordArray[18].Word[7].QWire ), 
        .D(n117), .Clk(_626_net_) );
  Bit_454 \WordArray[18].Word[8].Cell  ( .Q(\WordArray[18].Word[8].QWire ), 
        .D(n119), .Clk(_626_net_) );
  Bit_453 \WordArray[18].Word[9].Cell  ( .Q(\WordArray[18].Word[9].QWire ), 
        .D(n121), .Clk(_626_net_) );
  Bit_452 \WordArray[18].Word[10].Cell  ( .Q(\WordArray[18].Word[10].QWire ), 
        .D(n123), .Clk(_626_net_) );
  Bit_451 \WordArray[18].Word[11].Cell  ( .Q(\WordArray[18].Word[11].QWire ), 
        .D(n125), .Clk(_626_net_) );
  Bit_450 \WordArray[18].Word[12].Cell  ( .Q(\WordArray[18].Word[12].QWire ), 
        .D(n127), .Clk(_626_net_) );
  Bit_449 \WordArray[18].Word[13].Cell  ( .Q(\WordArray[18].Word[13].QWire ), 
        .D(n129), .Clk(_626_net_) );
  Bit_448 \WordArray[18].Word[14].Cell  ( .Q(\WordArray[18].Word[14].QWire ), 
        .D(n131), .Clk(_626_net_) );
  Bit_447 \WordArray[18].Word[15].Cell  ( .Q(\WordArray[18].Word[15].QWire ), 
        .D(n133), .Clk(_626_net_) );
  Bit_446 \WordArray[18].Word[16].Cell  ( .Q(\WordArray[18].Word[16].QWire ), 
        .D(n135), .Clk(_626_net_) );
  Bit_445 \WordArray[18].Word[17].Cell  ( .Q(\WordArray[18].Word[17].QWire ), 
        .D(n137), .Clk(_626_net_) );
  Bit_444 \WordArray[18].Word[18].Cell  ( .Q(\WordArray[18].Word[18].QWire ), 
        .D(n139), .Clk(_626_net_) );
  Bit_443 \WordArray[18].Word[19].Cell  ( .Q(\WordArray[18].Word[19].QWire ), 
        .D(n141), .Clk(_626_net_) );
  Bit_442 \WordArray[18].Word[20].Cell  ( .Q(\WordArray[18].Word[20].QWire ), 
        .D(n143), .Clk(_626_net_) );
  Bit_441 \WordArray[18].Word[21].Cell  ( .Q(\WordArray[18].Word[21].QWire ), 
        .D(n145), .Clk(_626_net_) );
  Bit_440 \WordArray[18].Word[22].Cell  ( .Q(\WordArray[18].Word[22].QWire ), 
        .D(n147), .Clk(_626_net_) );
  Bit_439 \WordArray[18].Word[23].Cell  ( .Q(\WordArray[18].Word[23].QWire ), 
        .D(n149), .Clk(_626_net_) );
  Bit_438 \WordArray[18].Word[24].Cell  ( .Q(\WordArray[18].Word[24].QWire ), 
        .D(n151), .Clk(_626_net_) );
  Bit_437 \WordArray[18].Word[25].Cell  ( .Q(\WordArray[18].Word[25].QWire ), 
        .D(n153), .Clk(_626_net_) );
  Bit_436 \WordArray[18].Word[26].Cell  ( .Q(\WordArray[18].Word[26].QWire ), 
        .D(n155), .Clk(_626_net_) );
  Bit_435 \WordArray[18].Word[27].Cell  ( .Q(\WordArray[18].Word[27].QWire ), 
        .D(n157), .Clk(_626_net_) );
  Bit_434 \WordArray[18].Word[28].Cell  ( .Q(\WordArray[18].Word[28].QWire ), 
        .D(n159), .Clk(_626_net_) );
  Bit_433 \WordArray[18].Word[29].Cell  ( .Q(\WordArray[18].Word[29].QWire ), 
        .D(n161), .Clk(_626_net_) );
  Bit_432 \WordArray[18].Word[30].Cell  ( .Q(\WordArray[18].Word[30].QWire ), 
        .D(n163), .Clk(_626_net_) );
  Bit_431 \WordArray[18].Word[31].Cell  ( .Q(\WordArray[18].Word[31].QWire ), 
        .D(n165), .Clk(_626_net_) );
  Bit_430 \WordArray[18].Word[32].Cell  ( .D(n34), .Clk(_626_net_) );
  Bit_429 \WordArray[19].Word[0].Cell  ( .Q(\WordArray[19].Word[0].QWire ), 
        .D(n103), .Clk(_659_net_) );
  Bit_428 \WordArray[19].Word[1].Cell  ( .Q(\WordArray[19].Word[1].QWire ), 
        .D(n105), .Clk(_659_net_) );
  Bit_427 \WordArray[19].Word[2].Cell  ( .Q(\WordArray[19].Word[2].QWire ), 
        .D(n107), .Clk(_659_net_) );
  Bit_426 \WordArray[19].Word[3].Cell  ( .Q(\WordArray[19].Word[3].QWire ), 
        .D(n109), .Clk(_659_net_) );
  Bit_425 \WordArray[19].Word[4].Cell  ( .Q(\WordArray[19].Word[4].QWire ), 
        .D(n111), .Clk(_659_net_) );
  Bit_424 \WordArray[19].Word[5].Cell  ( .Q(\WordArray[19].Word[5].QWire ), 
        .D(n113), .Clk(_659_net_) );
  Bit_423 \WordArray[19].Word[6].Cell  ( .Q(\WordArray[19].Word[6].QWire ), 
        .D(n115), .Clk(_659_net_) );
  Bit_422 \WordArray[19].Word[7].Cell  ( .Q(\WordArray[19].Word[7].QWire ), 
        .D(n117), .Clk(_659_net_) );
  Bit_421 \WordArray[19].Word[8].Cell  ( .Q(\WordArray[19].Word[8].QWire ), 
        .D(n119), .Clk(_659_net_) );
  Bit_420 \WordArray[19].Word[9].Cell  ( .Q(\WordArray[19].Word[9].QWire ), 
        .D(n121), .Clk(_659_net_) );
  Bit_419 \WordArray[19].Word[10].Cell  ( .Q(\WordArray[19].Word[10].QWire ), 
        .D(n123), .Clk(_659_net_) );
  Bit_418 \WordArray[19].Word[11].Cell  ( .Q(\WordArray[19].Word[11].QWire ), 
        .D(n125), .Clk(_659_net_) );
  Bit_417 \WordArray[19].Word[12].Cell  ( .Q(\WordArray[19].Word[12].QWire ), 
        .D(n127), .Clk(_659_net_) );
  Bit_416 \WordArray[19].Word[13].Cell  ( .Q(\WordArray[19].Word[13].QWire ), 
        .D(n129), .Clk(_659_net_) );
  Bit_415 \WordArray[19].Word[14].Cell  ( .Q(\WordArray[19].Word[14].QWire ), 
        .D(n131), .Clk(_659_net_) );
  Bit_414 \WordArray[19].Word[15].Cell  ( .Q(\WordArray[19].Word[15].QWire ), 
        .D(n133), .Clk(_659_net_) );
  Bit_413 \WordArray[19].Word[16].Cell  ( .Q(\WordArray[19].Word[16].QWire ), 
        .D(n135), .Clk(_659_net_) );
  Bit_412 \WordArray[19].Word[17].Cell  ( .Q(\WordArray[19].Word[17].QWire ), 
        .D(n137), .Clk(_659_net_) );
  Bit_411 \WordArray[19].Word[18].Cell  ( .Q(\WordArray[19].Word[18].QWire ), 
        .D(n139), .Clk(_659_net_) );
  Bit_410 \WordArray[19].Word[19].Cell  ( .Q(\WordArray[19].Word[19].QWire ), 
        .D(n141), .Clk(_659_net_) );
  Bit_409 \WordArray[19].Word[20].Cell  ( .Q(\WordArray[19].Word[20].QWire ), 
        .D(n143), .Clk(_659_net_) );
  Bit_408 \WordArray[19].Word[21].Cell  ( .Q(\WordArray[19].Word[21].QWire ), 
        .D(n145), .Clk(_659_net_) );
  Bit_407 \WordArray[19].Word[22].Cell  ( .Q(\WordArray[19].Word[22].QWire ), 
        .D(n147), .Clk(_659_net_) );
  Bit_406 \WordArray[19].Word[23].Cell  ( .Q(\WordArray[19].Word[23].QWire ), 
        .D(n149), .Clk(_659_net_) );
  Bit_405 \WordArray[19].Word[24].Cell  ( .Q(\WordArray[19].Word[24].QWire ), 
        .D(n151), .Clk(_659_net_) );
  Bit_404 \WordArray[19].Word[25].Cell  ( .Q(\WordArray[19].Word[25].QWire ), 
        .D(n153), .Clk(_659_net_) );
  Bit_403 \WordArray[19].Word[26].Cell  ( .Q(\WordArray[19].Word[26].QWire ), 
        .D(n155), .Clk(_659_net_) );
  Bit_402 \WordArray[19].Word[27].Cell  ( .Q(\WordArray[19].Word[27].QWire ), 
        .D(n157), .Clk(_659_net_) );
  Bit_401 \WordArray[19].Word[28].Cell  ( .Q(\WordArray[19].Word[28].QWire ), 
        .D(n159), .Clk(_659_net_) );
  Bit_400 \WordArray[19].Word[29].Cell  ( .Q(\WordArray[19].Word[29].QWire ), 
        .D(n161), .Clk(_659_net_) );
  Bit_399 \WordArray[19].Word[30].Cell  ( .Q(\WordArray[19].Word[30].QWire ), 
        .D(n163), .Clk(_659_net_) );
  Bit_398 \WordArray[19].Word[31].Cell  ( .Q(\WordArray[19].Word[31].QWire ), 
        .D(n165), .Clk(_659_net_) );
  Bit_397 \WordArray[19].Word[32].Cell  ( .D(n34), .Clk(_659_net_) );
  Bit_396 \WordArray[20].Word[0].Cell  ( .Q(\WordArray[20].Word[0].QWire ), 
        .D(n103), .Clk(_692_net_) );
  Bit_395 \WordArray[20].Word[1].Cell  ( .Q(\WordArray[20].Word[1].QWire ), 
        .D(n105), .Clk(_692_net_) );
  Bit_394 \WordArray[20].Word[2].Cell  ( .Q(\WordArray[20].Word[2].QWire ), 
        .D(n107), .Clk(_692_net_) );
  Bit_393 \WordArray[20].Word[3].Cell  ( .Q(\WordArray[20].Word[3].QWire ), 
        .D(n109), .Clk(_692_net_) );
  Bit_392 \WordArray[20].Word[4].Cell  ( .Q(\WordArray[20].Word[4].QWire ), 
        .D(n111), .Clk(_692_net_) );
  Bit_391 \WordArray[20].Word[5].Cell  ( .Q(\WordArray[20].Word[5].QWire ), 
        .D(n113), .Clk(_692_net_) );
  Bit_390 \WordArray[20].Word[6].Cell  ( .Q(\WordArray[20].Word[6].QWire ), 
        .D(n115), .Clk(_692_net_) );
  Bit_389 \WordArray[20].Word[7].Cell  ( .Q(\WordArray[20].Word[7].QWire ), 
        .D(n117), .Clk(_692_net_) );
  Bit_388 \WordArray[20].Word[8].Cell  ( .Q(\WordArray[20].Word[8].QWire ), 
        .D(n119), .Clk(_692_net_) );
  Bit_387 \WordArray[20].Word[9].Cell  ( .Q(\WordArray[20].Word[9].QWire ), 
        .D(n121), .Clk(_692_net_) );
  Bit_386 \WordArray[20].Word[10].Cell  ( .Q(\WordArray[20].Word[10].QWire ), 
        .D(n123), .Clk(_692_net_) );
  Bit_385 \WordArray[20].Word[11].Cell  ( .Q(\WordArray[20].Word[11].QWire ), 
        .D(n125), .Clk(_692_net_) );
  Bit_384 \WordArray[20].Word[12].Cell  ( .Q(\WordArray[20].Word[12].QWire ), 
        .D(n127), .Clk(_692_net_) );
  Bit_383 \WordArray[20].Word[13].Cell  ( .Q(\WordArray[20].Word[13].QWire ), 
        .D(n129), .Clk(_692_net_) );
  Bit_382 \WordArray[20].Word[14].Cell  ( .Q(\WordArray[20].Word[14].QWire ), 
        .D(n131), .Clk(_692_net_) );
  Bit_381 \WordArray[20].Word[15].Cell  ( .Q(\WordArray[20].Word[15].QWire ), 
        .D(n133), .Clk(_692_net_) );
  Bit_380 \WordArray[20].Word[16].Cell  ( .Q(\WordArray[20].Word[16].QWire ), 
        .D(n135), .Clk(_692_net_) );
  Bit_379 \WordArray[20].Word[17].Cell  ( .Q(\WordArray[20].Word[17].QWire ), 
        .D(n137), .Clk(_692_net_) );
  Bit_378 \WordArray[20].Word[18].Cell  ( .Q(\WordArray[20].Word[18].QWire ), 
        .D(n139), .Clk(_692_net_) );
  Bit_377 \WordArray[20].Word[19].Cell  ( .Q(\WordArray[20].Word[19].QWire ), 
        .D(n141), .Clk(_692_net_) );
  Bit_376 \WordArray[20].Word[20].Cell  ( .Q(\WordArray[20].Word[20].QWire ), 
        .D(n143), .Clk(_692_net_) );
  Bit_375 \WordArray[20].Word[21].Cell  ( .Q(\WordArray[20].Word[21].QWire ), 
        .D(n145), .Clk(_692_net_) );
  Bit_374 \WordArray[20].Word[22].Cell  ( .Q(\WordArray[20].Word[22].QWire ), 
        .D(n147), .Clk(_692_net_) );
  Bit_373 \WordArray[20].Word[23].Cell  ( .Q(\WordArray[20].Word[23].QWire ), 
        .D(n149), .Clk(_692_net_) );
  Bit_372 \WordArray[20].Word[24].Cell  ( .Q(\WordArray[20].Word[24].QWire ), 
        .D(n151), .Clk(_692_net_) );
  Bit_371 \WordArray[20].Word[25].Cell  ( .Q(\WordArray[20].Word[25].QWire ), 
        .D(n153), .Clk(_692_net_) );
  Bit_370 \WordArray[20].Word[26].Cell  ( .Q(\WordArray[20].Word[26].QWire ), 
        .D(n155), .Clk(_692_net_) );
  Bit_369 \WordArray[20].Word[27].Cell  ( .Q(\WordArray[20].Word[27].QWire ), 
        .D(n157), .Clk(_692_net_) );
  Bit_368 \WordArray[20].Word[28].Cell  ( .Q(\WordArray[20].Word[28].QWire ), 
        .D(n159), .Clk(_692_net_) );
  Bit_367 \WordArray[20].Word[29].Cell  ( .Q(\WordArray[20].Word[29].QWire ), 
        .D(n161), .Clk(_692_net_) );
  Bit_366 \WordArray[20].Word[30].Cell  ( .Q(\WordArray[20].Word[30].QWire ), 
        .D(n163), .Clk(_692_net_) );
  Bit_365 \WordArray[20].Word[31].Cell  ( .Q(\WordArray[20].Word[31].QWire ), 
        .D(n165), .Clk(_692_net_) );
  Bit_364 \WordArray[20].Word[32].Cell  ( .D(n34), .Clk(_692_net_) );
  Bit_363 \WordArray[21].Word[0].Cell  ( .Q(\WordArray[21].Word[0].QWire ), 
        .D(n103), .Clk(_725_net_) );
  Bit_362 \WordArray[21].Word[1].Cell  ( .Q(\WordArray[21].Word[1].QWire ), 
        .D(n105), .Clk(_725_net_) );
  Bit_361 \WordArray[21].Word[2].Cell  ( .Q(\WordArray[21].Word[2].QWire ), 
        .D(n107), .Clk(_725_net_) );
  Bit_360 \WordArray[21].Word[3].Cell  ( .Q(\WordArray[21].Word[3].QWire ), 
        .D(n109), .Clk(_725_net_) );
  Bit_359 \WordArray[21].Word[4].Cell  ( .Q(\WordArray[21].Word[4].QWire ), 
        .D(n111), .Clk(_725_net_) );
  Bit_358 \WordArray[21].Word[5].Cell  ( .Q(\WordArray[21].Word[5].QWire ), 
        .D(n113), .Clk(_725_net_) );
  Bit_357 \WordArray[21].Word[6].Cell  ( .Q(\WordArray[21].Word[6].QWire ), 
        .D(n115), .Clk(_725_net_) );
  Bit_356 \WordArray[21].Word[7].Cell  ( .Q(\WordArray[21].Word[7].QWire ), 
        .D(n117), .Clk(_725_net_) );
  Bit_355 \WordArray[21].Word[8].Cell  ( .Q(\WordArray[21].Word[8].QWire ), 
        .D(n119), .Clk(_725_net_) );
  Bit_354 \WordArray[21].Word[9].Cell  ( .Q(\WordArray[21].Word[9].QWire ), 
        .D(n121), .Clk(_725_net_) );
  Bit_353 \WordArray[21].Word[10].Cell  ( .Q(\WordArray[21].Word[10].QWire ), 
        .D(n123), .Clk(_725_net_) );
  Bit_352 \WordArray[21].Word[11].Cell  ( .Q(\WordArray[21].Word[11].QWire ), 
        .D(n125), .Clk(_725_net_) );
  Bit_351 \WordArray[21].Word[12].Cell  ( .Q(\WordArray[21].Word[12].QWire ), 
        .D(n127), .Clk(_725_net_) );
  Bit_350 \WordArray[21].Word[13].Cell  ( .Q(\WordArray[21].Word[13].QWire ), 
        .D(n129), .Clk(_725_net_) );
  Bit_349 \WordArray[21].Word[14].Cell  ( .Q(\WordArray[21].Word[14].QWire ), 
        .D(n131), .Clk(_725_net_) );
  Bit_348 \WordArray[21].Word[15].Cell  ( .Q(\WordArray[21].Word[15].QWire ), 
        .D(n133), .Clk(_725_net_) );
  Bit_347 \WordArray[21].Word[16].Cell  ( .Q(\WordArray[21].Word[16].QWire ), 
        .D(n135), .Clk(_725_net_) );
  Bit_346 \WordArray[21].Word[17].Cell  ( .Q(\WordArray[21].Word[17].QWire ), 
        .D(n137), .Clk(_725_net_) );
  Bit_345 \WordArray[21].Word[18].Cell  ( .Q(\WordArray[21].Word[18].QWire ), 
        .D(n139), .Clk(_725_net_) );
  Bit_344 \WordArray[21].Word[19].Cell  ( .Q(\WordArray[21].Word[19].QWire ), 
        .D(n141), .Clk(_725_net_) );
  Bit_343 \WordArray[21].Word[20].Cell  ( .Q(\WordArray[21].Word[20].QWire ), 
        .D(n143), .Clk(_725_net_) );
  Bit_342 \WordArray[21].Word[21].Cell  ( .Q(\WordArray[21].Word[21].QWire ), 
        .D(n145), .Clk(_725_net_) );
  Bit_341 \WordArray[21].Word[22].Cell  ( .Q(\WordArray[21].Word[22].QWire ), 
        .D(n147), .Clk(_725_net_) );
  Bit_340 \WordArray[21].Word[23].Cell  ( .Q(\WordArray[21].Word[23].QWire ), 
        .D(n149), .Clk(_725_net_) );
  Bit_339 \WordArray[21].Word[24].Cell  ( .Q(\WordArray[21].Word[24].QWire ), 
        .D(n151), .Clk(_725_net_) );
  Bit_338 \WordArray[21].Word[25].Cell  ( .Q(\WordArray[21].Word[25].QWire ), 
        .D(n153), .Clk(_725_net_) );
  Bit_337 \WordArray[21].Word[26].Cell  ( .Q(\WordArray[21].Word[26].QWire ), 
        .D(n155), .Clk(_725_net_) );
  Bit_336 \WordArray[21].Word[27].Cell  ( .Q(\WordArray[21].Word[27].QWire ), 
        .D(n157), .Clk(_725_net_) );
  Bit_335 \WordArray[21].Word[28].Cell  ( .Q(\WordArray[21].Word[28].QWire ), 
        .D(n159), .Clk(_725_net_) );
  Bit_334 \WordArray[21].Word[29].Cell  ( .Q(\WordArray[21].Word[29].QWire ), 
        .D(n161), .Clk(_725_net_) );
  Bit_333 \WordArray[21].Word[30].Cell  ( .Q(\WordArray[21].Word[30].QWire ), 
        .D(n163), .Clk(_725_net_) );
  Bit_332 \WordArray[21].Word[31].Cell  ( .Q(\WordArray[21].Word[31].QWire ), 
        .D(n165), .Clk(_725_net_) );
  Bit_331 \WordArray[21].Word[32].Cell  ( .D(n34), .Clk(_725_net_) );
  Bit_330 \WordArray[22].Word[0].Cell  ( .Q(\WordArray[22].Word[0].QWire ), 
        .D(n103), .Clk(_758_net_) );
  Bit_329 \WordArray[22].Word[1].Cell  ( .Q(\WordArray[22].Word[1].QWire ), 
        .D(DataI[1]), .Clk(_758_net_) );
  Bit_328 \WordArray[22].Word[2].Cell  ( .Q(\WordArray[22].Word[2].QWire ), 
        .D(n107), .Clk(_758_net_) );
  Bit_327 \WordArray[22].Word[3].Cell  ( .Q(\WordArray[22].Word[3].QWire ), 
        .D(DataI[3]), .Clk(_758_net_) );
  Bit_326 \WordArray[22].Word[4].Cell  ( .Q(\WordArray[22].Word[4].QWire ), 
        .D(DataI[4]), .Clk(_758_net_) );
  Bit_325 \WordArray[22].Word[5].Cell  ( .Q(\WordArray[22].Word[5].QWire ), 
        .D(n113), .Clk(_758_net_) );
  Bit_324 \WordArray[22].Word[6].Cell  ( .Q(\WordArray[22].Word[6].QWire ), 
        .D(DataI[6]), .Clk(_758_net_) );
  Bit_323 \WordArray[22].Word[7].Cell  ( .Q(\WordArray[22].Word[7].QWire ), 
        .D(DataI[7]), .Clk(_758_net_) );
  Bit_322 \WordArray[22].Word[8].Cell  ( .Q(\WordArray[22].Word[8].QWire ), 
        .D(DataI[8]), .Clk(_758_net_) );
  Bit_321 \WordArray[22].Word[9].Cell  ( .Q(\WordArray[22].Word[9].QWire ), 
        .D(DataI[9]), .Clk(_758_net_) );
  Bit_320 \WordArray[22].Word[10].Cell  ( .Q(\WordArray[22].Word[10].QWire ), 
        .D(DataI[10]), .Clk(_758_net_) );
  Bit_319 \WordArray[22].Word[11].Cell  ( .Q(\WordArray[22].Word[11].QWire ), 
        .D(DataI[11]), .Clk(_758_net_) );
  Bit_318 \WordArray[22].Word[12].Cell  ( .Q(\WordArray[22].Word[12].QWire ), 
        .D(DataI[12]), .Clk(_758_net_) );
  Bit_317 \WordArray[22].Word[13].Cell  ( .Q(\WordArray[22].Word[13].QWire ), 
        .D(DataI[13]), .Clk(_758_net_) );
  Bit_316 \WordArray[22].Word[14].Cell  ( .Q(\WordArray[22].Word[14].QWire ), 
        .D(DataI[14]), .Clk(_758_net_) );
  Bit_315 \WordArray[22].Word[15].Cell  ( .Q(\WordArray[22].Word[15].QWire ), 
        .D(DataI[15]), .Clk(_758_net_) );
  Bit_314 \WordArray[22].Word[16].Cell  ( .Q(\WordArray[22].Word[16].QWire ), 
        .D(DataI[16]), .Clk(_758_net_) );
  Bit_313 \WordArray[22].Word[17].Cell  ( .Q(\WordArray[22].Word[17].QWire ), 
        .D(DataI[17]), .Clk(_758_net_) );
  Bit_312 \WordArray[22].Word[18].Cell  ( .Q(\WordArray[22].Word[18].QWire ), 
        .D(DataI[18]), .Clk(_758_net_) );
  Bit_311 \WordArray[22].Word[19].Cell  ( .Q(\WordArray[22].Word[19].QWire ), 
        .D(DataI[19]), .Clk(_758_net_) );
  Bit_310 \WordArray[22].Word[20].Cell  ( .Q(\WordArray[22].Word[20].QWire ), 
        .D(DataI[20]), .Clk(_758_net_) );
  Bit_309 \WordArray[22].Word[21].Cell  ( .Q(\WordArray[22].Word[21].QWire ), 
        .D(DataI[21]), .Clk(_758_net_) );
  Bit_308 \WordArray[22].Word[22].Cell  ( .Q(\WordArray[22].Word[22].QWire ), 
        .D(DataI[22]), .Clk(_758_net_) );
  Bit_307 \WordArray[22].Word[23].Cell  ( .Q(\WordArray[22].Word[23].QWire ), 
        .D(DataI[23]), .Clk(_758_net_) );
  Bit_306 \WordArray[22].Word[24].Cell  ( .Q(\WordArray[22].Word[24].QWire ), 
        .D(DataI[24]), .Clk(_758_net_) );
  Bit_305 \WordArray[22].Word[25].Cell  ( .Q(\WordArray[22].Word[25].QWire ), 
        .D(DataI[25]), .Clk(_758_net_) );
  Bit_304 \WordArray[22].Word[26].Cell  ( .Q(\WordArray[22].Word[26].QWire ), 
        .D(DataI[26]), .Clk(_758_net_) );
  Bit_303 \WordArray[22].Word[27].Cell  ( .Q(\WordArray[22].Word[27].QWire ), 
        .D(DataI[27]), .Clk(_758_net_) );
  Bit_302 \WordArray[22].Word[28].Cell  ( .Q(\WordArray[22].Word[28].QWire ), 
        .D(DataI[28]), .Clk(_758_net_) );
  Bit_301 \WordArray[22].Word[29].Cell  ( .Q(\WordArray[22].Word[29].QWire ), 
        .D(DataI[29]), .Clk(_758_net_) );
  Bit_300 \WordArray[22].Word[30].Cell  ( .Q(\WordArray[22].Word[30].QWire ), 
        .D(DataI[30]), .Clk(_758_net_) );
  Bit_299 \WordArray[22].Word[31].Cell  ( .Q(\WordArray[22].Word[31].QWire ), 
        .D(DataI[31]), .Clk(_758_net_) );
  Bit_298 \WordArray[22].Word[32].Cell  ( .D(n34), .Clk(_758_net_) );
  Bit_297 \WordArray[23].Word[0].Cell  ( .Q(\WordArray[23].Word[0].QWire ), 
        .D(n103), .Clk(_791_net_) );
  Bit_296 \WordArray[23].Word[1].Cell  ( .Q(\WordArray[23].Word[1].QWire ), 
        .D(n105), .Clk(_791_net_) );
  Bit_295 \WordArray[23].Word[2].Cell  ( .Q(\WordArray[23].Word[2].QWire ), 
        .D(n107), .Clk(_791_net_) );
  Bit_294 \WordArray[23].Word[3].Cell  ( .Q(\WordArray[23].Word[3].QWire ), 
        .D(n109), .Clk(_791_net_) );
  Bit_293 \WordArray[23].Word[4].Cell  ( .Q(\WordArray[23].Word[4].QWire ), 
        .D(n111), .Clk(_791_net_) );
  Bit_292 \WordArray[23].Word[5].Cell  ( .Q(\WordArray[23].Word[5].QWire ), 
        .D(n113), .Clk(_791_net_) );
  Bit_291 \WordArray[23].Word[6].Cell  ( .Q(\WordArray[23].Word[6].QWire ), 
        .D(n115), .Clk(_791_net_) );
  Bit_290 \WordArray[23].Word[7].Cell  ( .Q(\WordArray[23].Word[7].QWire ), 
        .D(DataI[7]), .Clk(_791_net_) );
  Bit_289 \WordArray[23].Word[8].Cell  ( .Q(\WordArray[23].Word[8].QWire ), 
        .D(DataI[8]), .Clk(_791_net_) );
  Bit_288 \WordArray[23].Word[9].Cell  ( .Q(\WordArray[23].Word[9].QWire ), 
        .D(n121), .Clk(_791_net_) );
  Bit_287 \WordArray[23].Word[10].Cell  ( .Q(\WordArray[23].Word[10].QWire ), 
        .D(n123), .Clk(_791_net_) );
  Bit_286 \WordArray[23].Word[11].Cell  ( .Q(\WordArray[23].Word[11].QWire ), 
        .D(n125), .Clk(_791_net_) );
  Bit_285 \WordArray[23].Word[12].Cell  ( .Q(\WordArray[23].Word[12].QWire ), 
        .D(n127), .Clk(_791_net_) );
  Bit_284 \WordArray[23].Word[13].Cell  ( .Q(\WordArray[23].Word[13].QWire ), 
        .D(n129), .Clk(_791_net_) );
  Bit_283 \WordArray[23].Word[14].Cell  ( .Q(\WordArray[23].Word[14].QWire ), 
        .D(DataI[14]), .Clk(_791_net_) );
  Bit_282 \WordArray[23].Word[15].Cell  ( .Q(\WordArray[23].Word[15].QWire ), 
        .D(DataI[15]), .Clk(_791_net_) );
  Bit_281 \WordArray[23].Word[16].Cell  ( .Q(\WordArray[23].Word[16].QWire ), 
        .D(n135), .Clk(_791_net_) );
  Bit_280 \WordArray[23].Word[17].Cell  ( .Q(\WordArray[23].Word[17].QWire ), 
        .D(n137), .Clk(_791_net_) );
  Bit_279 \WordArray[23].Word[18].Cell  ( .Q(\WordArray[23].Word[18].QWire ), 
        .D(n139), .Clk(_791_net_) );
  Bit_278 \WordArray[23].Word[19].Cell  ( .Q(\WordArray[23].Word[19].QWire ), 
        .D(n141), .Clk(_791_net_) );
  Bit_277 \WordArray[23].Word[20].Cell  ( .Q(\WordArray[23].Word[20].QWire ), 
        .D(n143), .Clk(_791_net_) );
  Bit_276 \WordArray[23].Word[21].Cell  ( .Q(\WordArray[23].Word[21].QWire ), 
        .D(DataI[21]), .Clk(_791_net_) );
  Bit_275 \WordArray[23].Word[22].Cell  ( .Q(\WordArray[23].Word[22].QWire ), 
        .D(DataI[22]), .Clk(_791_net_) );
  Bit_274 \WordArray[23].Word[23].Cell  ( .Q(\WordArray[23].Word[23].QWire ), 
        .D(n149), .Clk(_791_net_) );
  Bit_273 \WordArray[23].Word[24].Cell  ( .Q(\WordArray[23].Word[24].QWire ), 
        .D(n151), .Clk(_791_net_) );
  Bit_272 \WordArray[23].Word[25].Cell  ( .Q(\WordArray[23].Word[25].QWire ), 
        .D(DataI[25]), .Clk(_791_net_) );
  Bit_271 \WordArray[23].Word[26].Cell  ( .Q(\WordArray[23].Word[26].QWire ), 
        .D(DataI[26]), .Clk(_791_net_) );
  Bit_270 \WordArray[23].Word[27].Cell  ( .Q(\WordArray[23].Word[27].QWire ), 
        .D(n157), .Clk(_791_net_) );
  Bit_269 \WordArray[23].Word[28].Cell  ( .Q(\WordArray[23].Word[28].QWire ), 
        .D(n159), .Clk(_791_net_) );
  Bit_268 \WordArray[23].Word[29].Cell  ( .Q(\WordArray[23].Word[29].QWire ), 
        .D(DataI[29]), .Clk(_791_net_) );
  Bit_267 \WordArray[23].Word[30].Cell  ( .Q(\WordArray[23].Word[30].QWire ), 
        .D(DataI[30]), .Clk(_791_net_) );
  Bit_266 \WordArray[23].Word[31].Cell  ( .Q(\WordArray[23].Word[31].QWire ), 
        .D(n165), .Clk(_791_net_) );
  Bit_265 \WordArray[23].Word[32].Cell  ( .D(n34), .Clk(_791_net_) );
  Bit_264 \WordArray[24].Word[0].Cell  ( .Q(\WordArray[24].Word[0].QWire ), 
        .D(n103), .Clk(_824_net_) );
  Bit_263 \WordArray[24].Word[1].Cell  ( .Q(\WordArray[24].Word[1].QWire ), 
        .D(DataI[1]), .Clk(_824_net_) );
  Bit_262 \WordArray[24].Word[2].Cell  ( .Q(\WordArray[24].Word[2].QWire ), 
        .D(DataI[2]), .Clk(_824_net_) );
  Bit_261 \WordArray[24].Word[3].Cell  ( .Q(\WordArray[24].Word[3].QWire ), 
        .D(DataI[3]), .Clk(_824_net_) );
  Bit_260 \WordArray[24].Word[4].Cell  ( .Q(\WordArray[24].Word[4].QWire ), 
        .D(DataI[4]), .Clk(_824_net_) );
  Bit_259 \WordArray[24].Word[5].Cell  ( .Q(\WordArray[24].Word[5].QWire ), 
        .D(DataI[5]), .Clk(_824_net_) );
  Bit_258 \WordArray[24].Word[6].Cell  ( .Q(\WordArray[24].Word[6].QWire ), 
        .D(DataI[6]), .Clk(_824_net_) );
  Bit_257 \WordArray[24].Word[7].Cell  ( .Q(\WordArray[24].Word[7].QWire ), 
        .D(DataI[7]), .Clk(_824_net_) );
  Bit_256 \WordArray[24].Word[8].Cell  ( .Q(\WordArray[24].Word[8].QWire ), 
        .D(DataI[8]), .Clk(_824_net_) );
  Bit_255 \WordArray[24].Word[9].Cell  ( .Q(\WordArray[24].Word[9].QWire ), 
        .D(DataI[9]), .Clk(_824_net_) );
  Bit_254 \WordArray[24].Word[10].Cell  ( .Q(\WordArray[24].Word[10].QWire ), 
        .D(DataI[10]), .Clk(_824_net_) );
  Bit_253 \WordArray[24].Word[11].Cell  ( .Q(\WordArray[24].Word[11].QWire ), 
        .D(DataI[11]), .Clk(_824_net_) );
  Bit_252 \WordArray[24].Word[12].Cell  ( .Q(\WordArray[24].Word[12].QWire ), 
        .D(DataI[12]), .Clk(_824_net_) );
  Bit_251 \WordArray[24].Word[13].Cell  ( .Q(\WordArray[24].Word[13].QWire ), 
        .D(DataI[13]), .Clk(_824_net_) );
  Bit_250 \WordArray[24].Word[14].Cell  ( .Q(\WordArray[24].Word[14].QWire ), 
        .D(DataI[14]), .Clk(_824_net_) );
  Bit_249 \WordArray[24].Word[15].Cell  ( .Q(\WordArray[24].Word[15].QWire ), 
        .D(DataI[15]), .Clk(_824_net_) );
  Bit_248 \WordArray[24].Word[16].Cell  ( .Q(\WordArray[24].Word[16].QWire ), 
        .D(DataI[16]), .Clk(_824_net_) );
  Bit_247 \WordArray[24].Word[17].Cell  ( .Q(\WordArray[24].Word[17].QWire ), 
        .D(DataI[17]), .Clk(_824_net_) );
  Bit_246 \WordArray[24].Word[18].Cell  ( .Q(\WordArray[24].Word[18].QWire ), 
        .D(DataI[18]), .Clk(_824_net_) );
  Bit_245 \WordArray[24].Word[19].Cell  ( .Q(\WordArray[24].Word[19].QWire ), 
        .D(DataI[19]), .Clk(_824_net_) );
  Bit_244 \WordArray[24].Word[20].Cell  ( .Q(\WordArray[24].Word[20].QWire ), 
        .D(DataI[20]), .Clk(_824_net_) );
  Bit_243 \WordArray[24].Word[21].Cell  ( .Q(\WordArray[24].Word[21].QWire ), 
        .D(DataI[21]), .Clk(_824_net_) );
  Bit_242 \WordArray[24].Word[22].Cell  ( .Q(\WordArray[24].Word[22].QWire ), 
        .D(DataI[22]), .Clk(_824_net_) );
  Bit_241 \WordArray[24].Word[23].Cell  ( .Q(\WordArray[24].Word[23].QWire ), 
        .D(DataI[23]), .Clk(_824_net_) );
  Bit_240 \WordArray[24].Word[24].Cell  ( .Q(\WordArray[24].Word[24].QWire ), 
        .D(DataI[24]), .Clk(_824_net_) );
  Bit_239 \WordArray[24].Word[25].Cell  ( .Q(\WordArray[24].Word[25].QWire ), 
        .D(DataI[25]), .Clk(_824_net_) );
  Bit_238 \WordArray[24].Word[26].Cell  ( .Q(\WordArray[24].Word[26].QWire ), 
        .D(DataI[26]), .Clk(_824_net_) );
  Bit_237 \WordArray[24].Word[27].Cell  ( .Q(\WordArray[24].Word[27].QWire ), 
        .D(DataI[27]), .Clk(_824_net_) );
  Bit_236 \WordArray[24].Word[28].Cell  ( .Q(\WordArray[24].Word[28].QWire ), 
        .D(DataI[28]), .Clk(_824_net_) );
  Bit_235 \WordArray[24].Word[29].Cell  ( .Q(\WordArray[24].Word[29].QWire ), 
        .D(DataI[29]), .Clk(_824_net_) );
  Bit_234 \WordArray[24].Word[30].Cell  ( .Q(\WordArray[24].Word[30].QWire ), 
        .D(DataI[30]), .Clk(_824_net_) );
  Bit_233 \WordArray[24].Word[31].Cell  ( .Q(\WordArray[24].Word[31].QWire ), 
        .D(DataI[31]), .Clk(_824_net_) );
  Bit_232 \WordArray[24].Word[32].Cell  ( .D(n34), .Clk(_824_net_) );
  Bit_231 \WordArray[25].Word[0].Cell  ( .Q(\WordArray[25].Word[0].QWire ), 
        .D(DataI[0]), .Clk(_857_net_) );
  Bit_230 \WordArray[25].Word[1].Cell  ( .Q(\WordArray[25].Word[1].QWire ), 
        .D(n105), .Clk(_857_net_) );
  Bit_229 \WordArray[25].Word[2].Cell  ( .Q(\WordArray[25].Word[2].QWire ), 
        .D(n107), .Clk(_857_net_) );
  Bit_228 \WordArray[25].Word[3].Cell  ( .Q(\WordArray[25].Word[3].QWire ), 
        .D(n109), .Clk(_857_net_) );
  Bit_227 \WordArray[25].Word[4].Cell  ( .Q(\WordArray[25].Word[4].QWire ), 
        .D(n111), .Clk(_857_net_) );
  Bit_226 \WordArray[25].Word[5].Cell  ( .Q(\WordArray[25].Word[5].QWire ), 
        .D(n113), .Clk(_857_net_) );
  Bit_225 \WordArray[25].Word[6].Cell  ( .Q(\WordArray[25].Word[6].QWire ), 
        .D(n115), .Clk(_857_net_) );
  Bit_224 \WordArray[25].Word[7].Cell  ( .Q(\WordArray[25].Word[7].QWire ), 
        .D(n117), .Clk(_857_net_) );
  Bit_223 \WordArray[25].Word[8].Cell  ( .Q(\WordArray[25].Word[8].QWire ), 
        .D(n119), .Clk(_857_net_) );
  Bit_222 \WordArray[25].Word[9].Cell  ( .Q(\WordArray[25].Word[9].QWire ), 
        .D(n121), .Clk(_857_net_) );
  Bit_221 \WordArray[25].Word[10].Cell  ( .Q(\WordArray[25].Word[10].QWire ), 
        .D(n123), .Clk(_857_net_) );
  Bit_220 \WordArray[25].Word[11].Cell  ( .Q(\WordArray[25].Word[11].QWire ), 
        .D(n125), .Clk(_857_net_) );
  Bit_219 \WordArray[25].Word[12].Cell  ( .Q(\WordArray[25].Word[12].QWire ), 
        .D(n127), .Clk(_857_net_) );
  Bit_218 \WordArray[25].Word[13].Cell  ( .Q(\WordArray[25].Word[13].QWire ), 
        .D(n129), .Clk(_857_net_) );
  Bit_217 \WordArray[25].Word[14].Cell  ( .Q(\WordArray[25].Word[14].QWire ), 
        .D(n131), .Clk(_857_net_) );
  Bit_216 \WordArray[25].Word[15].Cell  ( .Q(\WordArray[25].Word[15].QWire ), 
        .D(n133), .Clk(_857_net_) );
  Bit_215 \WordArray[25].Word[16].Cell  ( .Q(\WordArray[25].Word[16].QWire ), 
        .D(n135), .Clk(_857_net_) );
  Bit_214 \WordArray[25].Word[17].Cell  ( .Q(\WordArray[25].Word[17].QWire ), 
        .D(n137), .Clk(_857_net_) );
  Bit_213 \WordArray[25].Word[18].Cell  ( .Q(\WordArray[25].Word[18].QWire ), 
        .D(n139), .Clk(_857_net_) );
  Bit_212 \WordArray[25].Word[19].Cell  ( .Q(\WordArray[25].Word[19].QWire ), 
        .D(n141), .Clk(_857_net_) );
  Bit_211 \WordArray[25].Word[20].Cell  ( .Q(\WordArray[25].Word[20].QWire ), 
        .D(n143), .Clk(_857_net_) );
  Bit_210 \WordArray[25].Word[21].Cell  ( .Q(\WordArray[25].Word[21].QWire ), 
        .D(n145), .Clk(_857_net_) );
  Bit_209 \WordArray[25].Word[22].Cell  ( .Q(\WordArray[25].Word[22].QWire ), 
        .D(n147), .Clk(_857_net_) );
  Bit_208 \WordArray[25].Word[23].Cell  ( .Q(\WordArray[25].Word[23].QWire ), 
        .D(n149), .Clk(_857_net_) );
  Bit_207 \WordArray[25].Word[24].Cell  ( .Q(\WordArray[25].Word[24].QWire ), 
        .D(n151), .Clk(_857_net_) );
  Bit_206 \WordArray[25].Word[25].Cell  ( .Q(\WordArray[25].Word[25].QWire ), 
        .D(n153), .Clk(_857_net_) );
  Bit_205 \WordArray[25].Word[26].Cell  ( .Q(\WordArray[25].Word[26].QWire ), 
        .D(n155), .Clk(_857_net_) );
  Bit_204 \WordArray[25].Word[27].Cell  ( .Q(\WordArray[25].Word[27].QWire ), 
        .D(n157), .Clk(_857_net_) );
  Bit_203 \WordArray[25].Word[28].Cell  ( .Q(\WordArray[25].Word[28].QWire ), 
        .D(n159), .Clk(_857_net_) );
  Bit_202 \WordArray[25].Word[29].Cell  ( .Q(\WordArray[25].Word[29].QWire ), 
        .D(n161), .Clk(_857_net_) );
  Bit_201 \WordArray[25].Word[30].Cell  ( .Q(\WordArray[25].Word[30].QWire ), 
        .D(n163), .Clk(_857_net_) );
  Bit_200 \WordArray[25].Word[31].Cell  ( .Q(\WordArray[25].Word[31].QWire ), 
        .D(n165), .Clk(_857_net_) );
  Bit_199 \WordArray[25].Word[32].Cell  ( .D(n34), .Clk(_857_net_) );
  Bit_198 \WordArray[26].Word[0].Cell  ( .Q(\WordArray[26].Word[0].QWire ), 
        .D(n103), .Clk(_890_net_) );
  Bit_197 \WordArray[26].Word[1].Cell  ( .Q(\WordArray[26].Word[1].QWire ), 
        .D(n105), .Clk(_890_net_) );
  Bit_196 \WordArray[26].Word[2].Cell  ( .Q(\WordArray[26].Word[2].QWire ), 
        .D(DataI[2]), .Clk(_890_net_) );
  Bit_195 \WordArray[26].Word[3].Cell  ( .Q(\WordArray[26].Word[3].QWire ), 
        .D(n109), .Clk(_890_net_) );
  Bit_194 \WordArray[26].Word[4].Cell  ( .Q(\WordArray[26].Word[4].QWire ), 
        .D(n111), .Clk(_890_net_) );
  Bit_193 \WordArray[26].Word[5].Cell  ( .Q(\WordArray[26].Word[5].QWire ), 
        .D(DataI[5]), .Clk(_890_net_) );
  Bit_192 \WordArray[26].Word[6].Cell  ( .Q(\WordArray[26].Word[6].QWire ), 
        .D(n115), .Clk(_890_net_) );
  Bit_191 \WordArray[26].Word[7].Cell  ( .Q(\WordArray[26].Word[7].QWire ), 
        .D(n117), .Clk(_890_net_) );
  Bit_190 \WordArray[26].Word[8].Cell  ( .Q(\WordArray[26].Word[8].QWire ), 
        .D(n119), .Clk(_890_net_) );
  Bit_189 \WordArray[26].Word[9].Cell  ( .Q(\WordArray[26].Word[9].QWire ), 
        .D(n121), .Clk(_890_net_) );
  Bit_188 \WordArray[26].Word[10].Cell  ( .Q(\WordArray[26].Word[10].QWire ), 
        .D(n123), .Clk(_890_net_) );
  Bit_187 \WordArray[26].Word[11].Cell  ( .Q(\WordArray[26].Word[11].QWire ), 
        .D(n125), .Clk(_890_net_) );
  Bit_186 \WordArray[26].Word[12].Cell  ( .Q(\WordArray[26].Word[12].QWire ), 
        .D(n127), .Clk(_890_net_) );
  Bit_185 \WordArray[26].Word[13].Cell  ( .Q(\WordArray[26].Word[13].QWire ), 
        .D(n129), .Clk(_890_net_) );
  Bit_184 \WordArray[26].Word[14].Cell  ( .Q(\WordArray[26].Word[14].QWire ), 
        .D(n131), .Clk(_890_net_) );
  Bit_183 \WordArray[26].Word[15].Cell  ( .Q(\WordArray[26].Word[15].QWire ), 
        .D(n133), .Clk(_890_net_) );
  Bit_182 \WordArray[26].Word[16].Cell  ( .Q(\WordArray[26].Word[16].QWire ), 
        .D(n135), .Clk(_890_net_) );
  Bit_181 \WordArray[26].Word[17].Cell  ( .Q(\WordArray[26].Word[17].QWire ), 
        .D(n137), .Clk(_890_net_) );
  Bit_180 \WordArray[26].Word[18].Cell  ( .Q(\WordArray[26].Word[18].QWire ), 
        .D(n139), .Clk(_890_net_) );
  Bit_179 \WordArray[26].Word[19].Cell  ( .Q(\WordArray[26].Word[19].QWire ), 
        .D(n141), .Clk(_890_net_) );
  Bit_178 \WordArray[26].Word[20].Cell  ( .Q(\WordArray[26].Word[20].QWire ), 
        .D(n143), .Clk(_890_net_) );
  Bit_177 \WordArray[26].Word[21].Cell  ( .Q(\WordArray[26].Word[21].QWire ), 
        .D(n145), .Clk(_890_net_) );
  Bit_176 \WordArray[26].Word[22].Cell  ( .Q(\WordArray[26].Word[22].QWire ), 
        .D(n147), .Clk(_890_net_) );
  Bit_175 \WordArray[26].Word[23].Cell  ( .Q(\WordArray[26].Word[23].QWire ), 
        .D(n149), .Clk(_890_net_) );
  Bit_174 \WordArray[26].Word[24].Cell  ( .Q(\WordArray[26].Word[24].QWire ), 
        .D(n151), .Clk(_890_net_) );
  Bit_173 \WordArray[26].Word[25].Cell  ( .Q(\WordArray[26].Word[25].QWire ), 
        .D(n153), .Clk(_890_net_) );
  Bit_172 \WordArray[26].Word[26].Cell  ( .Q(\WordArray[26].Word[26].QWire ), 
        .D(n155), .Clk(_890_net_) );
  Bit_171 \WordArray[26].Word[27].Cell  ( .Q(\WordArray[26].Word[27].QWire ), 
        .D(n157), .Clk(_890_net_) );
  Bit_170 \WordArray[26].Word[28].Cell  ( .Q(\WordArray[26].Word[28].QWire ), 
        .D(n159), .Clk(_890_net_) );
  Bit_169 \WordArray[26].Word[29].Cell  ( .Q(\WordArray[26].Word[29].QWire ), 
        .D(n161), .Clk(_890_net_) );
  Bit_168 \WordArray[26].Word[30].Cell  ( .Q(\WordArray[26].Word[30].QWire ), 
        .D(n163), .Clk(_890_net_) );
  Bit_167 \WordArray[26].Word[31].Cell  ( .Q(\WordArray[26].Word[31].QWire ), 
        .D(n165), .Clk(_890_net_) );
  Bit_166 \WordArray[26].Word[32].Cell  ( .D(n34), .Clk(_890_net_) );
  Bit_165 \WordArray[27].Word[0].Cell  ( .Q(\WordArray[27].Word[0].QWire ), 
        .D(DataI[0]), .Clk(_923_net_) );
  Bit_164 \WordArray[27].Word[1].Cell  ( .Q(\WordArray[27].Word[1].QWire ), 
        .D(n105), .Clk(_923_net_) );
  Bit_163 \WordArray[27].Word[2].Cell  ( .Q(\WordArray[27].Word[2].QWire ), 
        .D(n107), .Clk(_923_net_) );
  Bit_162 \WordArray[27].Word[3].Cell  ( .Q(\WordArray[27].Word[3].QWire ), 
        .D(n109), .Clk(_923_net_) );
  Bit_161 \WordArray[27].Word[4].Cell  ( .Q(\WordArray[27].Word[4].QWire ), 
        .D(n111), .Clk(_923_net_) );
  Bit_160 \WordArray[27].Word[5].Cell  ( .Q(\WordArray[27].Word[5].QWire ), 
        .D(n113), .Clk(_923_net_) );
  Bit_159 \WordArray[27].Word[6].Cell  ( .Q(\WordArray[27].Word[6].QWire ), 
        .D(n115), .Clk(_923_net_) );
  Bit_158 \WordArray[27].Word[7].Cell  ( .Q(\WordArray[27].Word[7].QWire ), 
        .D(n117), .Clk(_923_net_) );
  Bit_157 \WordArray[27].Word[8].Cell  ( .Q(\WordArray[27].Word[8].QWire ), 
        .D(n119), .Clk(_923_net_) );
  Bit_156 \WordArray[27].Word[9].Cell  ( .Q(\WordArray[27].Word[9].QWire ), 
        .D(n121), .Clk(_923_net_) );
  Bit_155 \WordArray[27].Word[10].Cell  ( .Q(\WordArray[27].Word[10].QWire ), 
        .D(n123), .Clk(_923_net_) );
  Bit_154 \WordArray[27].Word[11].Cell  ( .Q(\WordArray[27].Word[11].QWire ), 
        .D(n125), .Clk(_923_net_) );
  Bit_153 \WordArray[27].Word[12].Cell  ( .Q(\WordArray[27].Word[12].QWire ), 
        .D(n127), .Clk(_923_net_) );
  Bit_152 \WordArray[27].Word[13].Cell  ( .Q(\WordArray[27].Word[13].QWire ), 
        .D(n129), .Clk(_923_net_) );
  Bit_151 \WordArray[27].Word[14].Cell  ( .Q(\WordArray[27].Word[14].QWire ), 
        .D(n131), .Clk(_923_net_) );
  Bit_150 \WordArray[27].Word[15].Cell  ( .Q(\WordArray[27].Word[15].QWire ), 
        .D(n133), .Clk(_923_net_) );
  Bit_149 \WordArray[27].Word[16].Cell  ( .Q(\WordArray[27].Word[16].QWire ), 
        .D(n135), .Clk(_923_net_) );
  Bit_148 \WordArray[27].Word[17].Cell  ( .Q(\WordArray[27].Word[17].QWire ), 
        .D(n137), .Clk(_923_net_) );
  Bit_147 \WordArray[27].Word[18].Cell  ( .Q(\WordArray[27].Word[18].QWire ), 
        .D(n139), .Clk(_923_net_) );
  Bit_146 \WordArray[27].Word[19].Cell  ( .Q(\WordArray[27].Word[19].QWire ), 
        .D(n141), .Clk(_923_net_) );
  Bit_145 \WordArray[27].Word[20].Cell  ( .Q(\WordArray[27].Word[20].QWire ), 
        .D(n143), .Clk(_923_net_) );
  Bit_144 \WordArray[27].Word[21].Cell  ( .Q(\WordArray[27].Word[21].QWire ), 
        .D(n145), .Clk(_923_net_) );
  Bit_143 \WordArray[27].Word[22].Cell  ( .Q(\WordArray[27].Word[22].QWire ), 
        .D(n147), .Clk(_923_net_) );
  Bit_142 \WordArray[27].Word[23].Cell  ( .Q(\WordArray[27].Word[23].QWire ), 
        .D(n149), .Clk(_923_net_) );
  Bit_141 \WordArray[27].Word[24].Cell  ( .Q(\WordArray[27].Word[24].QWire ), 
        .D(n151), .Clk(_923_net_) );
  Bit_140 \WordArray[27].Word[25].Cell  ( .Q(\WordArray[27].Word[25].QWire ), 
        .D(n153), .Clk(_923_net_) );
  Bit_139 \WordArray[27].Word[26].Cell  ( .Q(\WordArray[27].Word[26].QWire ), 
        .D(n155), .Clk(_923_net_) );
  Bit_138 \WordArray[27].Word[27].Cell  ( .Q(\WordArray[27].Word[27].QWire ), 
        .D(n157), .Clk(_923_net_) );
  Bit_137 \WordArray[27].Word[28].Cell  ( .Q(\WordArray[27].Word[28].QWire ), 
        .D(n159), .Clk(_923_net_) );
  Bit_136 \WordArray[27].Word[29].Cell  ( .Q(\WordArray[27].Word[29].QWire ), 
        .D(n161), .Clk(_923_net_) );
  Bit_135 \WordArray[27].Word[30].Cell  ( .Q(\WordArray[27].Word[30].QWire ), 
        .D(n163), .Clk(_923_net_) );
  Bit_134 \WordArray[27].Word[31].Cell  ( .Q(\WordArray[27].Word[31].QWire ), 
        .D(n165), .Clk(_923_net_) );
  Bit_133 \WordArray[27].Word[32].Cell  ( .D(n34), .Clk(_923_net_) );
  Bit_132 \WordArray[28].Word[0].Cell  ( .Q(\WordArray[28].Word[0].QWire ), 
        .D(n103), .Clk(_956_net_) );
  Bit_131 \WordArray[28].Word[1].Cell  ( .Q(\WordArray[28].Word[1].QWire ), 
        .D(n105), .Clk(_956_net_) );
  Bit_130 \WordArray[28].Word[2].Cell  ( .Q(\WordArray[28].Word[2].QWire ), 
        .D(DataI[2]), .Clk(_956_net_) );
  Bit_129 \WordArray[28].Word[3].Cell  ( .Q(\WordArray[28].Word[3].QWire ), 
        .D(n109), .Clk(_956_net_) );
  Bit_128 \WordArray[28].Word[4].Cell  ( .Q(\WordArray[28].Word[4].QWire ), 
        .D(n111), .Clk(_956_net_) );
  Bit_127 \WordArray[28].Word[5].Cell  ( .Q(\WordArray[28].Word[5].QWire ), 
        .D(DataI[5]), .Clk(_956_net_) );
  Bit_126 \WordArray[28].Word[6].Cell  ( .Q(\WordArray[28].Word[6].QWire ), 
        .D(n115), .Clk(_956_net_) );
  Bit_125 \WordArray[28].Word[7].Cell  ( .Q(\WordArray[28].Word[7].QWire ), 
        .D(n117), .Clk(_956_net_) );
  Bit_124 \WordArray[28].Word[8].Cell  ( .Q(\WordArray[28].Word[8].QWire ), 
        .D(n119), .Clk(_956_net_) );
  Bit_123 \WordArray[28].Word[9].Cell  ( .Q(\WordArray[28].Word[9].QWire ), 
        .D(n121), .Clk(_956_net_) );
  Bit_122 \WordArray[28].Word[10].Cell  ( .Q(\WordArray[28].Word[10].QWire ), 
        .D(n123), .Clk(_956_net_) );
  Bit_121 \WordArray[28].Word[11].Cell  ( .Q(\WordArray[28].Word[11].QWire ), 
        .D(n125), .Clk(_956_net_) );
  Bit_120 \WordArray[28].Word[12].Cell  ( .Q(\WordArray[28].Word[12].QWire ), 
        .D(n127), .Clk(_956_net_) );
  Bit_119 \WordArray[28].Word[13].Cell  ( .Q(\WordArray[28].Word[13].QWire ), 
        .D(n129), .Clk(_956_net_) );
  Bit_118 \WordArray[28].Word[14].Cell  ( .Q(\WordArray[28].Word[14].QWire ), 
        .D(n131), .Clk(_956_net_) );
  Bit_117 \WordArray[28].Word[15].Cell  ( .Q(\WordArray[28].Word[15].QWire ), 
        .D(n133), .Clk(_956_net_) );
  Bit_116 \WordArray[28].Word[16].Cell  ( .Q(\WordArray[28].Word[16].QWire ), 
        .D(n135), .Clk(_956_net_) );
  Bit_115 \WordArray[28].Word[17].Cell  ( .Q(\WordArray[28].Word[17].QWire ), 
        .D(n137), .Clk(_956_net_) );
  Bit_114 \WordArray[28].Word[18].Cell  ( .Q(\WordArray[28].Word[18].QWire ), 
        .D(n139), .Clk(_956_net_) );
  Bit_113 \WordArray[28].Word[19].Cell  ( .Q(\WordArray[28].Word[19].QWire ), 
        .D(n141), .Clk(_956_net_) );
  Bit_112 \WordArray[28].Word[20].Cell  ( .Q(\WordArray[28].Word[20].QWire ), 
        .D(n143), .Clk(_956_net_) );
  Bit_111 \WordArray[28].Word[21].Cell  ( .Q(\WordArray[28].Word[21].QWire ), 
        .D(n145), .Clk(_956_net_) );
  Bit_110 \WordArray[28].Word[22].Cell  ( .Q(\WordArray[28].Word[22].QWire ), 
        .D(n147), .Clk(_956_net_) );
  Bit_109 \WordArray[28].Word[23].Cell  ( .Q(\WordArray[28].Word[23].QWire ), 
        .D(n149), .Clk(_956_net_) );
  Bit_108 \WordArray[28].Word[24].Cell  ( .Q(\WordArray[28].Word[24].QWire ), 
        .D(n151), .Clk(_956_net_) );
  Bit_107 \WordArray[28].Word[25].Cell  ( .Q(\WordArray[28].Word[25].QWire ), 
        .D(n153), .Clk(_956_net_) );
  Bit_106 \WordArray[28].Word[26].Cell  ( .Q(\WordArray[28].Word[26].QWire ), 
        .D(n155), .Clk(_956_net_) );
  Bit_105 \WordArray[28].Word[27].Cell  ( .Q(\WordArray[28].Word[27].QWire ), 
        .D(n157), .Clk(_956_net_) );
  Bit_104 \WordArray[28].Word[28].Cell  ( .Q(\WordArray[28].Word[28].QWire ), 
        .D(n159), .Clk(_956_net_) );
  Bit_103 \WordArray[28].Word[29].Cell  ( .Q(\WordArray[28].Word[29].QWire ), 
        .D(n161), .Clk(_956_net_) );
  Bit_102 \WordArray[28].Word[30].Cell  ( .Q(\WordArray[28].Word[30].QWire ), 
        .D(n163), .Clk(_956_net_) );
  Bit_101 \WordArray[28].Word[31].Cell  ( .Q(\WordArray[28].Word[31].QWire ), 
        .D(n165), .Clk(_956_net_) );
  Bit_100 \WordArray[28].Word[32].Cell  ( .D(n34), .Clk(_956_net_) );
  Bit_99 \WordArray[29].Word[0].Cell  ( .Q(\WordArray[29].Word[0].QWire ), .D(
        DataI[0]), .Clk(_989_net_) );
  Bit_98 \WordArray[29].Word[1].Cell  ( .Q(\WordArray[29].Word[1].QWire ), .D(
        DataI[1]), .Clk(_989_net_) );
  Bit_97 \WordArray[29].Word[2].Cell  ( .Q(\WordArray[29].Word[2].QWire ), .D(
        n107), .Clk(_989_net_) );
  Bit_96 \WordArray[29].Word[3].Cell  ( .Q(\WordArray[29].Word[3].QWire ), .D(
        DataI[3]), .Clk(_989_net_) );
  Bit_95 \WordArray[29].Word[4].Cell  ( .Q(\WordArray[29].Word[4].QWire ), .D(
        DataI[4]), .Clk(_989_net_) );
  Bit_94 \WordArray[29].Word[5].Cell  ( .Q(\WordArray[29].Word[5].QWire ), .D(
        n113), .Clk(_989_net_) );
  Bit_93 \WordArray[29].Word[6].Cell  ( .Q(\WordArray[29].Word[6].QWire ), .D(
        DataI[6]), .Clk(_989_net_) );
  Bit_92 \WordArray[29].Word[7].Cell  ( .Q(\WordArray[29].Word[7].QWire ), .D(
        DataI[7]), .Clk(_989_net_) );
  Bit_91 \WordArray[29].Word[8].Cell  ( .Q(\WordArray[29].Word[8].QWire ), .D(
        DataI[8]), .Clk(_989_net_) );
  Bit_90 \WordArray[29].Word[9].Cell  ( .Q(\WordArray[29].Word[9].QWire ), .D(
        DataI[9]), .Clk(_989_net_) );
  Bit_89 \WordArray[29].Word[10].Cell  ( .Q(\WordArray[29].Word[10].QWire ), 
        .D(DataI[10]), .Clk(_989_net_) );
  Bit_88 \WordArray[29].Word[11].Cell  ( .Q(\WordArray[29].Word[11].QWire ), 
        .D(DataI[11]), .Clk(_989_net_) );
  Bit_87 \WordArray[29].Word[12].Cell  ( .Q(\WordArray[29].Word[12].QWire ), 
        .D(DataI[12]), .Clk(_989_net_) );
  Bit_86 \WordArray[29].Word[13].Cell  ( .Q(\WordArray[29].Word[13].QWire ), 
        .D(DataI[13]), .Clk(_989_net_) );
  Bit_85 \WordArray[29].Word[14].Cell  ( .Q(\WordArray[29].Word[14].QWire ), 
        .D(DataI[14]), .Clk(_989_net_) );
  Bit_84 \WordArray[29].Word[15].Cell  ( .Q(\WordArray[29].Word[15].QWire ), 
        .D(DataI[15]), .Clk(_989_net_) );
  Bit_83 \WordArray[29].Word[16].Cell  ( .Q(\WordArray[29].Word[16].QWire ), 
        .D(DataI[16]), .Clk(_989_net_) );
  Bit_82 \WordArray[29].Word[17].Cell  ( .Q(\WordArray[29].Word[17].QWire ), 
        .D(DataI[17]), .Clk(_989_net_) );
  Bit_81 \WordArray[29].Word[18].Cell  ( .Q(\WordArray[29].Word[18].QWire ), 
        .D(DataI[18]), .Clk(_989_net_) );
  Bit_80 \WordArray[29].Word[19].Cell  ( .Q(\WordArray[29].Word[19].QWire ), 
        .D(DataI[19]), .Clk(_989_net_) );
  Bit_79 \WordArray[29].Word[20].Cell  ( .Q(\WordArray[29].Word[20].QWire ), 
        .D(DataI[20]), .Clk(_989_net_) );
  Bit_78 \WordArray[29].Word[21].Cell  ( .Q(\WordArray[29].Word[21].QWire ), 
        .D(DataI[21]), .Clk(_989_net_) );
  Bit_77 \WordArray[29].Word[22].Cell  ( .Q(\WordArray[29].Word[22].QWire ), 
        .D(DataI[22]), .Clk(_989_net_) );
  Bit_76 \WordArray[29].Word[23].Cell  ( .Q(\WordArray[29].Word[23].QWire ), 
        .D(DataI[23]), .Clk(_989_net_) );
  Bit_75 \WordArray[29].Word[24].Cell  ( .Q(\WordArray[29].Word[24].QWire ), 
        .D(DataI[24]), .Clk(_989_net_) );
  Bit_74 \WordArray[29].Word[25].Cell  ( .Q(\WordArray[29].Word[25].QWire ), 
        .D(DataI[25]), .Clk(_989_net_) );
  Bit_73 \WordArray[29].Word[26].Cell  ( .Q(\WordArray[29].Word[26].QWire ), 
        .D(DataI[26]), .Clk(_989_net_) );
  Bit_72 \WordArray[29].Word[27].Cell  ( .Q(\WordArray[29].Word[27].QWire ), 
        .D(DataI[27]), .Clk(_989_net_) );
  Bit_71 \WordArray[29].Word[28].Cell  ( .Q(\WordArray[29].Word[28].QWire ), 
        .D(DataI[28]), .Clk(_989_net_) );
  Bit_70 \WordArray[29].Word[29].Cell  ( .Q(\WordArray[29].Word[29].QWire ), 
        .D(DataI[29]), .Clk(_989_net_) );
  Bit_69 \WordArray[29].Word[30].Cell  ( .Q(\WordArray[29].Word[30].QWire ), 
        .D(DataI[30]), .Clk(_989_net_) );
  Bit_68 \WordArray[29].Word[31].Cell  ( .Q(\WordArray[29].Word[31].QWire ), 
        .D(DataI[31]), .Clk(_989_net_) );
  Bit_67 \WordArray[29].Word[32].Cell  ( .D(n34), .Clk(_989_net_) );
  Bit_66 \WordArray[30].Word[0].Cell  ( .Q(\WordArray[30].Word[0].QWire ), .D(
        n103), .Clk(_999_net_) );
  Bit_65 \WordArray[30].Word[1].Cell  ( .Q(\WordArray[30].Word[1].QWire ), .D(
        DataI[1]), .Clk(_999_net_) );
  Bit_64 \WordArray[30].Word[2].Cell  ( .Q(\WordArray[30].Word[2].QWire ), .D(
        DataI[2]), .Clk(_999_net_) );
  Bit_63 \WordArray[30].Word[3].Cell  ( .Q(\WordArray[30].Word[3].QWire ), .D(
        DataI[3]), .Clk(_999_net_) );
  Bit_62 \WordArray[30].Word[4].Cell  ( .Q(\WordArray[30].Word[4].QWire ), .D(
        DataI[4]), .Clk(_999_net_) );
  Bit_61 \WordArray[30].Word[5].Cell  ( .Q(\WordArray[30].Word[5].QWire ), .D(
        DataI[5]), .Clk(_999_net_) );
  Bit_60 \WordArray[30].Word[6].Cell  ( .Q(\WordArray[30].Word[6].QWire ), .D(
        DataI[6]), .Clk(_999_net_) );
  Bit_59 \WordArray[30].Word[7].Cell  ( .Q(\WordArray[30].Word[7].QWire ), .D(
        n117), .Clk(_999_net_) );
  Bit_58 \WordArray[30].Word[8].Cell  ( .Q(\WordArray[30].Word[8].QWire ), .D(
        n119), .Clk(_999_net_) );
  Bit_57 \WordArray[30].Word[9].Cell  ( .Q(\WordArray[30].Word[9].QWire ), .D(
        DataI[9]), .Clk(_999_net_) );
  Bit_56 \WordArray[30].Word[10].Cell  ( .Q(\WordArray[30].Word[10].QWire ), 
        .D(DataI[10]), .Clk(_999_net_) );
  Bit_55 \WordArray[30].Word[11].Cell  ( .Q(\WordArray[30].Word[11].QWire ), 
        .D(DataI[11]), .Clk(_999_net_) );
  Bit_54 \WordArray[30].Word[12].Cell  ( .Q(\WordArray[30].Word[12].QWire ), 
        .D(DataI[12]), .Clk(_999_net_) );
  Bit_53 \WordArray[30].Word[13].Cell  ( .Q(\WordArray[30].Word[13].QWire ), 
        .D(DataI[13]), .Clk(_999_net_) );
  Bit_52 \WordArray[30].Word[14].Cell  ( .Q(\WordArray[30].Word[14].QWire ), 
        .D(n131), .Clk(_999_net_) );
  Bit_51 \WordArray[30].Word[15].Cell  ( .Q(\WordArray[30].Word[15].QWire ), 
        .D(n133), .Clk(_999_net_) );
  Bit_50 \WordArray[30].Word[16].Cell  ( .Q(\WordArray[30].Word[16].QWire ), 
        .D(DataI[16]), .Clk(_999_net_) );
  Bit_49 \WordArray[30].Word[17].Cell  ( .Q(\WordArray[30].Word[17].QWire ), 
        .D(DataI[17]), .Clk(_999_net_) );
  Bit_48 \WordArray[30].Word[18].Cell  ( .Q(\WordArray[30].Word[18].QWire ), 
        .D(DataI[18]), .Clk(_999_net_) );
  Bit_47 \WordArray[30].Word[19].Cell  ( .Q(\WordArray[30].Word[19].QWire ), 
        .D(DataI[19]), .Clk(_999_net_) );
  Bit_46 \WordArray[30].Word[20].Cell  ( .Q(\WordArray[30].Word[20].QWire ), 
        .D(DataI[20]), .Clk(_999_net_) );
  Bit_45 \WordArray[30].Word[21].Cell  ( .Q(\WordArray[30].Word[21].QWire ), 
        .D(n145), .Clk(_999_net_) );
  Bit_44 \WordArray[30].Word[22].Cell  ( .Q(\WordArray[30].Word[22].QWire ), 
        .D(n147), .Clk(_999_net_) );
  Bit_43 \WordArray[30].Word[23].Cell  ( .Q(\WordArray[30].Word[23].QWire ), 
        .D(DataI[23]), .Clk(_999_net_) );
  Bit_42 \WordArray[30].Word[24].Cell  ( .Q(\WordArray[30].Word[24].QWire ), 
        .D(DataI[24]), .Clk(_999_net_) );
  Bit_41 \WordArray[30].Word[25].Cell  ( .Q(\WordArray[30].Word[25].QWire ), 
        .D(n153), .Clk(_999_net_) );
  Bit_40 \WordArray[30].Word[26].Cell  ( .Q(\WordArray[30].Word[26].QWire ), 
        .D(n155), .Clk(_999_net_) );
  Bit_39 \WordArray[30].Word[27].Cell  ( .Q(\WordArray[30].Word[27].QWire ), 
        .D(DataI[27]), .Clk(_999_net_) );
  Bit_38 \WordArray[30].Word[28].Cell  ( .Q(\WordArray[30].Word[28].QWire ), 
        .D(DataI[28]), .Clk(_999_net_) );
  Bit_37 \WordArray[30].Word[29].Cell  ( .Q(\WordArray[30].Word[29].QWire ), 
        .D(n161), .Clk(_999_net_) );
  Bit_36 \WordArray[30].Word[30].Cell  ( .Q(\WordArray[30].Word[30].QWire ), 
        .D(n163), .Clk(_999_net_) );
  Bit_35 \WordArray[30].Word[31].Cell  ( .Q(\WordArray[30].Word[31].QWire ), 
        .D(DataI[31]), .Clk(_999_net_) );
  Bit_34 \WordArray[30].Word[32].Cell  ( .D(n34), .Clk(_999_net_) );
  Bit_33 \WordArray[31].Word[0].Cell  ( .Q(\WordArray[31].Word[0].QWire ), .D(
        DataI[0]), .Clk(_1055_net_) );
  Bit_32 \WordArray[31].Word[1].Cell  ( .Q(\WordArray[31].Word[1].QWire ), .D(
        DataI[1]), .Clk(_1055_net_) );
  Bit_31 \WordArray[31].Word[2].Cell  ( .Q(\WordArray[31].Word[2].QWire ), .D(
        n107), .Clk(_1055_net_) );
  Bit_30 \WordArray[31].Word[3].Cell  ( .Q(\WordArray[31].Word[3].QWire ), .D(
        DataI[3]), .Clk(_1055_net_) );
  Bit_29 \WordArray[31].Word[4].Cell  ( .Q(\WordArray[31].Word[4].QWire ), .D(
        DataI[4]), .Clk(_1055_net_) );
  Bit_28 \WordArray[31].Word[5].Cell  ( .Q(\WordArray[31].Word[5].QWire ), .D(
        n113), .Clk(_1055_net_) );
  Bit_27 \WordArray[31].Word[6].Cell  ( .Q(\WordArray[31].Word[6].QWire ), .D(
        DataI[6]), .Clk(_1055_net_) );
  Bit_26 \WordArray[31].Word[7].Cell  ( .Q(\WordArray[31].Word[7].QWire ), .D(
        DataI[7]), .Clk(_1055_net_) );
  Bit_25 \WordArray[31].Word[8].Cell  ( .Q(\WordArray[31].Word[8].QWire ), .D(
        DataI[8]), .Clk(_1055_net_) );
  Bit_24 \WordArray[31].Word[9].Cell  ( .Q(\WordArray[31].Word[9].QWire ), .D(
        DataI[9]), .Clk(_1055_net_) );
  Bit_23 \WordArray[31].Word[10].Cell  ( .Q(\WordArray[31].Word[10].QWire ), 
        .D(DataI[10]), .Clk(_1055_net_) );
  Bit_22 \WordArray[31].Word[11].Cell  ( .Q(\WordArray[31].Word[11].QWire ), 
        .D(DataI[11]), .Clk(_1055_net_) );
  Bit_21 \WordArray[31].Word[12].Cell  ( .Q(\WordArray[31].Word[12].QWire ), 
        .D(DataI[12]), .Clk(_1055_net_) );
  Bit_20 \WordArray[31].Word[13].Cell  ( .Q(\WordArray[31].Word[13].QWire ), 
        .D(DataI[13]), .Clk(_1055_net_) );
  Bit_19 \WordArray[31].Word[14].Cell  ( .Q(\WordArray[31].Word[14].QWire ), 
        .D(DataI[14]), .Clk(_1055_net_) );
  Bit_18 \WordArray[31].Word[15].Cell  ( .Q(\WordArray[31].Word[15].QWire ), 
        .D(DataI[15]), .Clk(_1055_net_) );
  Bit_17 \WordArray[31].Word[16].Cell  ( .Q(\WordArray[31].Word[16].QWire ), 
        .D(DataI[16]), .Clk(_1055_net_) );
  Bit_16 \WordArray[31].Word[17].Cell  ( .Q(\WordArray[31].Word[17].QWire ), 
        .D(DataI[17]), .Clk(_1055_net_) );
  Bit_15 \WordArray[31].Word[18].Cell  ( .Q(\WordArray[31].Word[18].QWire ), 
        .D(DataI[18]), .Clk(_1055_net_) );
  Bit_14 \WordArray[31].Word[19].Cell  ( .Q(\WordArray[31].Word[19].QWire ), 
        .D(DataI[19]), .Clk(_1055_net_) );
  Bit_13 \WordArray[31].Word[20].Cell  ( .Q(\WordArray[31].Word[20].QWire ), 
        .D(DataI[20]), .Clk(_1055_net_) );
  Bit_12 \WordArray[31].Word[21].Cell  ( .Q(\WordArray[31].Word[21].QWire ), 
        .D(DataI[21]), .Clk(_1055_net_) );
  Bit_11 \WordArray[31].Word[22].Cell  ( .Q(\WordArray[31].Word[22].QWire ), 
        .D(DataI[22]), .Clk(_1055_net_) );
  Bit_10 \WordArray[31].Word[23].Cell  ( .Q(\WordArray[31].Word[23].QWire ), 
        .D(DataI[23]), .Clk(_1055_net_) );
  Bit_9 \WordArray[31].Word[24].Cell  ( .Q(\WordArray[31].Word[24].QWire ), 
        .D(DataI[24]), .Clk(_1055_net_) );
  Bit_8 \WordArray[31].Word[25].Cell  ( .Q(\WordArray[31].Word[25].QWire ), 
        .D(DataI[25]), .Clk(_1055_net_) );
  Bit_7 \WordArray[31].Word[26].Cell  ( .Q(\WordArray[31].Word[26].QWire ), 
        .D(DataI[26]), .Clk(_1055_net_) );
  Bit_6 \WordArray[31].Word[27].Cell  ( .Q(\WordArray[31].Word[27].QWire ), 
        .D(DataI[27]), .Clk(_1055_net_) );
  Bit_5 \WordArray[31].Word[28].Cell  ( .Q(\WordArray[31].Word[28].QWire ), 
        .D(DataI[28]), .Clk(_1055_net_) );
  Bit_4 \WordArray[31].Word[29].Cell  ( .Q(\WordArray[31].Word[29].QWire ), 
        .D(DataI[29]), .Clk(_1055_net_) );
  Bit_3 \WordArray[31].Word[30].Cell  ( .Q(\WordArray[31].Word[30].QWire ), 
        .D(DataI[30]), .Clk(_1055_net_) );
  Bit_2 \WordArray[31].Word[31].Cell  ( .Q(\WordArray[31].Word[31].QWire ), 
        .D(DataI[31]), .Clk(_1055_net_) );
  Bit_1 \WordArray[31].Word[32].Cell  ( .D(\WordArray[9].CoreIn[32] ), .Clk(
        _1055_net_) );
  DFQD1 ParityErrReg_reg ( .D(N1127), .CP(ChipClock), .Q(ParityErr) );
  AN2D1 U3 ( .A1(ClockIn), .A2(n102), .Z(ChipClock) );
  OA21D1 U4 ( .A1(n2140), .A2(n2141), .B(n100), .Z(n1) );
  INVD0 U5 ( .I(Write), .ZN(n2083) );
  INVD1 U6 ( .I(DataI[3]), .ZN(n110) );
  INVD1 U7 ( .I(DataI[10]), .ZN(n124) );
  INVD1 U8 ( .I(DataI[11]), .ZN(n126) );
  INVD1 U9 ( .I(DataI[12]), .ZN(n128) );
  INVD1 U10 ( .I(DataI[13]), .ZN(n130) );
  INVD1 U11 ( .I(DataI[14]), .ZN(n132) );
  INVD1 U12 ( .I(DataI[15]), .ZN(n134) );
  INVD1 U13 ( .I(DataI[16]), .ZN(n136) );
  INVD1 U14 ( .I(DataI[17]), .ZN(n138) );
  INVD1 U15 ( .I(DataI[18]), .ZN(n140) );
  INVD1 U16 ( .I(DataI[19]), .ZN(n142) );
  INVD1 U17 ( .I(DataI[20]), .ZN(n144) );
  INVD1 U18 ( .I(DataI[21]), .ZN(n146) );
  INVD1 U19 ( .I(DataI[22]), .ZN(n148) );
  INVD1 U20 ( .I(DataI[23]), .ZN(n150) );
  INVD1 U21 ( .I(DataI[24]), .ZN(n152) );
  INVD1 U22 ( .I(DataI[25]), .ZN(n154) );
  INVD1 U23 ( .I(DataI[26]), .ZN(n156) );
  INVD1 U24 ( .I(DataI[27]), .ZN(n158) );
  INVD1 U25 ( .I(DataI[28]), .ZN(n160) );
  INVD1 U26 ( .I(DataI[29]), .ZN(n162) );
  INVD1 U27 ( .I(DataI[30]), .ZN(n164) );
  INVD1 U28 ( .I(DataI[31]), .ZN(n166) );
  INVD1 U29 ( .I(DataI[1]), .ZN(n106) );
  INVD1 U30 ( .I(DataI[2]), .ZN(n108) );
  INVD1 U31 ( .I(DataI[4]), .ZN(n112) );
  INVD1 U32 ( .I(DataI[5]), .ZN(n114) );
  INVD1 U33 ( .I(DataI[6]), .ZN(n116) );
  INVD1 U34 ( .I(DataI[7]), .ZN(n118) );
  INVD1 U35 ( .I(DataI[8]), .ZN(n120) );
  INVD1 U36 ( .I(DataI[9]), .ZN(n122) );
  INVD1 U37 ( .I(DataI[0]), .ZN(n104) );
  INVD1 U38 ( .I(n2), .ZN(n97) );
  INVD1 U39 ( .I(n2), .ZN(n98) );
  INVD1 U40 ( .I(n3), .ZN(n93) );
  INVD1 U41 ( .I(n3), .ZN(n94) );
  INVD1 U42 ( .I(n4), .ZN(n91) );
  INVD1 U48 ( .I(n4), .ZN(n92) );
  INVD1 U55 ( .I(n5), .ZN(n89) );
  INVD1 U56 ( .I(n5), .ZN(n90) );
  INVD1 U60 ( .I(n6), .ZN(n87) );
  INVD1 U61 ( .I(n6), .ZN(n88) );
  INVD1 U62 ( .I(n7), .ZN(n85) );
  INVD1 U63 ( .I(n7), .ZN(n86) );
  INVD1 U64 ( .I(n8), .ZN(n83) );
  INVD1 U65 ( .I(n8), .ZN(n84) );
  INVD1 U66 ( .I(n9), .ZN(n41) );
  INVD1 U67 ( .I(n9), .ZN(n42) );
  INVD1 U68 ( .I(n10), .ZN(n39) );
  INVD1 U69 ( .I(n10), .ZN(n40) );
  INVD1 U70 ( .I(n11), .ZN(n37) );
  INVD1 U71 ( .I(n11), .ZN(n38) );
  INVD1 U72 ( .I(n12), .ZN(n95) );
  INVD1 U73 ( .I(n12), .ZN(n96) );
  INVD1 U74 ( .I(n13), .ZN(n81) );
  INVD1 U75 ( .I(n13), .ZN(n82) );
  INVD1 U76 ( .I(n14), .ZN(n79) );
  INVD1 U77 ( .I(n14), .ZN(n80) );
  INVD1 U78 ( .I(n15), .ZN(n77) );
  INVD1 U79 ( .I(n15), .ZN(n78) );
  INVD1 U80 ( .I(n16), .ZN(n75) );
  INVD1 U81 ( .I(n16), .ZN(n76) );
  INVD1 U82 ( .I(n17), .ZN(n65) );
  INVD1 U83 ( .I(n17), .ZN(n66) );
  INVD1 U84 ( .I(n18), .ZN(n63) );
  INVD1 U85 ( .I(n18), .ZN(n64) );
  INVD1 U86 ( .I(n19), .ZN(n61) );
  INVD1 U87 ( .I(n19), .ZN(n62) );
  INVD1 U88 ( .I(n20), .ZN(n59) );
  INVD1 U89 ( .I(n20), .ZN(n60) );
  INVD1 U90 ( .I(n21), .ZN(n49) );
  INVD1 U91 ( .I(n21), .ZN(n50) );
  INVD1 U92 ( .I(n22), .ZN(n47) );
  INVD1 U93 ( .I(n22), .ZN(n48) );
  INVD1 U94 ( .I(n23), .ZN(n45) );
  INVD1 U95 ( .I(n23), .ZN(n46) );
  INVD1 U96 ( .I(n24), .ZN(n43) );
  INVD1 U97 ( .I(n24), .ZN(n44) );
  INVD1 U98 ( .I(n25), .ZN(n73) );
  INVD1 U99 ( .I(n25), .ZN(n74) );
  INVD1 U100 ( .I(n26), .ZN(n71) );
  INVD1 U101 ( .I(n26), .ZN(n72) );
  INVD1 U102 ( .I(n27), .ZN(n69) );
  INVD1 U103 ( .I(n27), .ZN(n70) );
  INVD1 U104 ( .I(n28), .ZN(n67) );
  INVD1 U105 ( .I(n28), .ZN(n68) );
  INVD1 U106 ( .I(n29), .ZN(n57) );
  INVD1 U107 ( .I(n29), .ZN(n58) );
  INVD1 U108 ( .I(n30), .ZN(n55) );
  INVD1 U109 ( .I(n30), .ZN(n56) );
  INVD1 U110 ( .I(n31), .ZN(n53) );
  INVD1 U111 ( .I(n31), .ZN(n54) );
  INVD1 U112 ( .I(n32), .ZN(n51) );
  INVD1 U113 ( .I(n32), .ZN(n52) );
  INVD1 U114 ( .I(n33), .ZN(n35) );
  INVD1 U115 ( .I(n33), .ZN(n36) );
  BUFFD1 U116 ( .I(\WordArray[9].CoreIn[32] ), .Z(n34) );
  AN2D1 U117 ( .A1(n102), .A2(Read), .Z(Dready) );
  ND2D1 U118 ( .A1(n2151), .A2(n2166), .ZN(n2) );
  ND2D1 U119 ( .A1(n2150), .A2(n2166), .ZN(n3) );
  ND2D1 U120 ( .A1(n2150), .A2(n2167), .ZN(n4) );
  ND2D1 U121 ( .A1(n2149), .A2(n2166), .ZN(n5) );
  ND2D1 U122 ( .A1(n2149), .A2(n2167), .ZN(n6) );
  ND2D1 U123 ( .A1(n2146), .A2(n2166), .ZN(n7) );
  ND2D1 U124 ( .A1(n2146), .A2(n2167), .ZN(n8) );
  ND2D1 U125 ( .A1(n2149), .A2(n2147), .ZN(n9) );
  ND2D1 U126 ( .A1(n2149), .A2(n2148), .ZN(n10) );
  ND2D1 U127 ( .A1(n2146), .A2(n2147), .ZN(n11) );
  ND2D1 U128 ( .A1(n2167), .A2(n2151), .ZN(n12) );
  ND2D1 U129 ( .A1(n2163), .A2(n2151), .ZN(n13) );
  ND2D1 U130 ( .A1(n2164), .A2(n2151), .ZN(n14) );
  ND2D1 U131 ( .A1(n2163), .A2(n2150), .ZN(n15) );
  ND2D1 U132 ( .A1(n2164), .A2(n2150), .ZN(n16) );
  ND2D1 U133 ( .A1(n2156), .A2(n2151), .ZN(n17) );
  ND2D1 U134 ( .A1(n2157), .A2(n2151), .ZN(n18) );
  ND2D1 U135 ( .A1(n2156), .A2(n2150), .ZN(n19) );
  ND2D1 U136 ( .A1(n2157), .A2(n2150), .ZN(n20) );
  ND2D1 U137 ( .A1(n2147), .A2(n2151), .ZN(n21) );
  ND2D1 U138 ( .A1(n2148), .A2(n2151), .ZN(n22) );
  ND2D1 U139 ( .A1(n2147), .A2(n2150), .ZN(n23) );
  ND2D1 U140 ( .A1(n2148), .A2(n2150), .ZN(n24) );
  ND2D1 U141 ( .A1(n2163), .A2(n2149), .ZN(n25) );
  ND2D1 U142 ( .A1(n2164), .A2(n2149), .ZN(n26) );
  ND2D1 U143 ( .A1(n2163), .A2(n2146), .ZN(n27) );
  ND2D1 U144 ( .A1(n2164), .A2(n2146), .ZN(n28) );
  ND2D1 U145 ( .A1(n2156), .A2(n2149), .ZN(n29) );
  ND2D1 U146 ( .A1(n2157), .A2(n2149), .ZN(n30) );
  ND2D1 U147 ( .A1(n2156), .A2(n2146), .ZN(n31) );
  ND2D1 U148 ( .A1(n2157), .A2(n2146), .ZN(n32) );
  ND2D1 U149 ( .A1(n2148), .A2(n2146), .ZN(n33) );
  AN2D1 U150 ( .A1(n2169), .A2(n2153), .Z(n2166) );
  AN2D1 U151 ( .A1(n2152), .A2(n2153), .Z(n2147) );
  AN2D1 U152 ( .A1(n2165), .A2(n2153), .Z(n2163) );
  AN2D1 U153 ( .A1(n2158), .A2(n2153), .Z(n2156) );
  NR2D1 U154 ( .A1(n2154), .A2(n2155), .ZN(n2152) );
  BUFFD1 U155 ( .I(n101), .Z(n102) );
  ND4D1 U156 ( .A1(n2142), .A2(n2143), .A3(n2144), .A4(n2145), .ZN(n2141) );
  ND4D1 U157 ( .A1(n2159), .A2(n2160), .A3(n2161), .A4(n2162), .ZN(n2140) );
  AN4D1 U158 ( .A1(n2100), .A2(n2101), .A3(n2098), .A4(n2099), .Z(n2142) );
  AN4D1 U159 ( .A1(n2097), .A2(n2082), .A3(n2084), .A4(n2086), .Z(n2159) );
  AN4D1 U160 ( .A1(n2112), .A2(n2113), .A3(n2110), .A4(n2111), .Z(n2160) );
  AN4D1 U161 ( .A1(n2095), .A2(n2096), .A3(n2093), .A4(n2094), .Z(n2143) );
  AN4D1 U162 ( .A1(n2108), .A2(n2109), .A3(n2106), .A4(n2107), .Z(n2161) );
  AN4D1 U163 ( .A1(n2091), .A2(n2092), .A3(n2089), .A4(n2090), .Z(n2144) );
  AN4D1 U164 ( .A1(n2104), .A2(n2105), .A3(n2102), .A4(n2103), .Z(n2162) );
  AN4D1 U165 ( .A1(n2087), .A2(n2088), .A3(n2114), .A4(n2085), .Z(n2145) );
  XOR3D1 U166 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n2124), .Z(n2123) );
  XOR3D1 U167 ( .A1(n2125), .A2(DataI[17]), .A3(n2126), .Z(n2124) );
  XOR3D1 U168 ( .A1(n2119), .A2(DataI[3]), .A3(n2120), .Z(n2118) );
  XOR3D1 U169 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n2121), .Z(n2120) );
  XOR3D1 U170 ( .A1(n2122), .A2(DataI[10]), .A3(n2123), .Z(n2121) );
  XOR3D1 U171 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n2115), .Z(
        \WordArray[9].CoreIn[32] ) );
  XOR3D1 U172 ( .A1(DataI[0]), .A2(n2116), .A3(n2117), .Z(n2115) );
  XOR3D1 U173 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n2118), .Z(n2117) );
  NR2D3 U174 ( .A1(n99), .A2(n2097), .ZN(_65_net_) );
  NR2D3 U175 ( .A1(n2083), .A2(n2086), .ZN(_98_net_) );
  NR2D3 U176 ( .A1(n2083), .A2(n2084), .ZN(_99_net_) );
  NR2D3 U177 ( .A1(n100), .A2(n2113), .ZN(_164_net_) );
  NR2D3 U178 ( .A1(n100), .A2(n2112), .ZN(_197_net_) );
  NR2D3 U179 ( .A1(n100), .A2(n2111), .ZN(_230_net_) );
  NR2D3 U180 ( .A1(n100), .A2(n2110), .ZN(_263_net_) );
  NR2D3 U181 ( .A1(n100), .A2(n2109), .ZN(_296_net_) );
  NR2D3 U182 ( .A1(n100), .A2(n2108), .ZN(_329_net_) );
  NR2D3 U183 ( .A1(n100), .A2(n2107), .ZN(_362_net_) );
  NR2D3 U184 ( .A1(n100), .A2(n2106), .ZN(_395_net_) );
  NR2D3 U185 ( .A1(n100), .A2(n2105), .ZN(_428_net_) );
  NR2D3 U186 ( .A1(n99), .A2(n2104), .ZN(_461_net_) );
  NR2D3 U187 ( .A1(n99), .A2(n2103), .ZN(_494_net_) );
  NR2D3 U188 ( .A1(n99), .A2(n2102), .ZN(_527_net_) );
  NR2D3 U189 ( .A1(n99), .A2(n2101), .ZN(_560_net_) );
  NR2D3 U190 ( .A1(n99), .A2(n2100), .ZN(_593_net_) );
  NR2D3 U191 ( .A1(n99), .A2(n2099), .ZN(_626_net_) );
  NR2D3 U192 ( .A1(n99), .A2(n2098), .ZN(_659_net_) );
  NR2D3 U193 ( .A1(n99), .A2(n2096), .ZN(_692_net_) );
  NR2D3 U194 ( .A1(n99), .A2(n2095), .ZN(_725_net_) );
  NR2D3 U195 ( .A1(n99), .A2(n2094), .ZN(_758_net_) );
  NR2D3 U196 ( .A1(n2083), .A2(n2093), .ZN(_791_net_) );
  NR2D3 U197 ( .A1(n2083), .A2(n2092), .ZN(_824_net_) );
  NR2D3 U198 ( .A1(n2083), .A2(n2091), .ZN(_857_net_) );
  NR2D3 U199 ( .A1(n2083), .A2(n2090), .ZN(_890_net_) );
  NR2D3 U200 ( .A1(n99), .A2(n2089), .ZN(_923_net_) );
  NR2D3 U201 ( .A1(n99), .A2(n2088), .ZN(_956_net_) );
  NR2D3 U202 ( .A1(n99), .A2(n2087), .ZN(_989_net_) );
  NR2D3 U203 ( .A1(n99), .A2(n2085), .ZN(_999_net_) );
  NR2D3 U204 ( .A1(n100), .A2(n2114), .ZN(_1055_net_) );
  NR2D3 U205 ( .A1(n2082), .A2(n99), .ZN(_9_net_) );
  NR2D1 U206 ( .A1(Addr[1]), .A2(Addr[2]), .ZN(n2151) );
  NR2D1 U207 ( .A1(n2168), .A2(Addr[2]), .ZN(n2150) );
  AN2D1 U208 ( .A1(Addr[2]), .A2(Addr[1]), .Z(n2146) );
  AN2D1 U209 ( .A1(Addr[2]), .A2(n2168), .Z(n2149) );
  INVD1 U210 ( .I(Addr[0]), .ZN(n2153) );
  INVD1 U211 ( .I(Addr[3]), .ZN(n2155) );
  INVD1 U212 ( .I(Addr[4]), .ZN(n2154) );
  AN2D1 U213 ( .A1(n2169), .A2(Addr[0]), .Z(n2167) );
  AN2D1 U214 ( .A1(n2152), .A2(Addr[0]), .Z(n2148) );
  AN2D1 U215 ( .A1(n2165), .A2(Addr[0]), .Z(n2164) );
  AN2D1 U216 ( .A1(n2158), .A2(Addr[0]), .Z(n2157) );
  INVD1 U217 ( .I(Addr[1]), .ZN(n2168) );
  NR2D1 U218 ( .A1(Addr[3]), .A2(Addr[4]), .ZN(n2169) );
  NR2D1 U219 ( .A1(n2155), .A2(Addr[4]), .ZN(n2165) );
  NR2D1 U220 ( .A1(n2154), .A2(Addr[3]), .ZN(n2158) );
  BUFFD1 U221 ( .I(ChipEna), .Z(n101) );
  ND2D1 U222 ( .A1(n69), .A2(ChipClock), .ZN(n2103) );
  ND2D1 U223 ( .A1(n85), .A2(ChipClock), .ZN(n2111) );
  ND2D1 U224 ( .A1(n77), .A2(ChipClock), .ZN(n2107) );
  ND2D1 U225 ( .A1(n93), .A2(ChipClock), .ZN(n2086) );
  ND2D1 U226 ( .A1(n37), .A2(ChipClock), .ZN(n2085) );
  ND2D1 U227 ( .A1(n53), .A2(ChipClock), .ZN(n2094) );
  ND2D1 U228 ( .A1(n45), .A2(ChipClock), .ZN(n2090) );
  ND2D1 U229 ( .A1(n61), .A2(ChipClock), .ZN(n2099) );
  ND2D1 U230 ( .A1(n67), .A2(ChipClock), .ZN(n2102) );
  ND2D1 U231 ( .A1(n83), .A2(ChipClock), .ZN(n2110) );
  ND2D1 U232 ( .A1(n75), .A2(ChipClock), .ZN(n2106) );
  ND2D1 U233 ( .A1(n91), .A2(ChipClock), .ZN(n2084) );
  ND2D1 U234 ( .A1(n35), .A2(ChipClock), .ZN(n2114) );
  ND2D1 U235 ( .A1(n51), .A2(ChipClock), .ZN(n2093) );
  ND2D1 U236 ( .A1(n43), .A2(ChipClock), .ZN(n2089) );
  ND2D1 U237 ( .A1(n59), .A2(ChipClock), .ZN(n2098) );
  ND2D1 U238 ( .A1(n73), .A2(ChipClock), .ZN(n2105) );
  ND2D1 U239 ( .A1(n89), .A2(ChipClock), .ZN(n2113) );
  ND2D1 U240 ( .A1(n81), .A2(ChipClock), .ZN(n2109) );
  ND2D1 U241 ( .A1(n41), .A2(ChipClock), .ZN(n2088) );
  ND2D1 U242 ( .A1(n57), .A2(ChipClock), .ZN(n2096) );
  ND2D1 U243 ( .A1(n49), .A2(ChipClock), .ZN(n2092) );
  ND2D1 U244 ( .A1(n65), .A2(ChipClock), .ZN(n2101) );
  ND2D1 U245 ( .A1(ChipClock), .A2(n97), .ZN(n2082) );
  ND2D1 U246 ( .A1(n71), .A2(ChipClock), .ZN(n2104) );
  ND2D1 U247 ( .A1(n87), .A2(ChipClock), .ZN(n2112) );
  ND2D1 U248 ( .A1(n79), .A2(ChipClock), .ZN(n2108) );
  ND2D1 U249 ( .A1(n95), .A2(ChipClock), .ZN(n2097) );
  ND2D1 U250 ( .A1(n39), .A2(ChipClock), .ZN(n2087) );
  ND2D1 U251 ( .A1(n55), .A2(ChipClock), .ZN(n2095) );
  ND2D1 U252 ( .A1(n47), .A2(ChipClock), .ZN(n2091) );
  ND2D1 U253 ( .A1(n63), .A2(ChipClock), .ZN(n2100) );
  INVD1 U254 ( .I(Write), .ZN(n100) );
  INVD1 U255 ( .I(n106), .ZN(n105) );
  INVD1 U256 ( .I(n108), .ZN(n107) );
  INVD1 U257 ( .I(n110), .ZN(n109) );
  INVD1 U258 ( .I(n112), .ZN(n111) );
  INVD1 U259 ( .I(n114), .ZN(n113) );
  INVD1 U260 ( .I(n116), .ZN(n115) );
  INVD1 U261 ( .I(n118), .ZN(n117) );
  INVD1 U262 ( .I(n120), .ZN(n119) );
  INVD1 U263 ( .I(n122), .ZN(n121) );
  INVD1 U264 ( .I(n124), .ZN(n123) );
  INVD1 U265 ( .I(n126), .ZN(n125) );
  INVD1 U266 ( .I(n128), .ZN(n127) );
  INVD1 U267 ( .I(n130), .ZN(n129) );
  INVD1 U268 ( .I(n132), .ZN(n131) );
  INVD1 U269 ( .I(n134), .ZN(n133) );
  INVD1 U270 ( .I(n136), .ZN(n135) );
  INVD1 U271 ( .I(n138), .ZN(n137) );
  INVD1 U272 ( .I(n140), .ZN(n139) );
  INVD1 U273 ( .I(n142), .ZN(n141) );
  INVD1 U274 ( .I(n144), .ZN(n143) );
  INVD1 U275 ( .I(n146), .ZN(n145) );
  INVD1 U276 ( .I(n148), .ZN(n147) );
  INVD1 U277 ( .I(n150), .ZN(n149) );
  INVD1 U278 ( .I(n152), .ZN(n151) );
  INVD1 U279 ( .I(n154), .ZN(n153) );
  INVD1 U280 ( .I(n156), .ZN(n155) );
  INVD1 U281 ( .I(n158), .ZN(n157) );
  INVD1 U282 ( .I(n160), .ZN(n159) );
  INVD1 U283 ( .I(n162), .ZN(n161) );
  INVD1 U284 ( .I(n164), .ZN(n163) );
  INVD1 U285 ( .I(n166), .ZN(n165) );
  INVD1 U286 ( .I(n104), .ZN(n103) );
  INVD1 U287 ( .I(Write), .ZN(n99) );
  AN3D1 U288 ( .A1(n1), .A2(n2128), .A3(Read), .Z(N1127) );
  XNR3D1 U289 ( .A1(DataRead[9]), .A2(DataRead[8]), .A3(DataRead[15]), .ZN(
        n2133) );
  XNR3D1 U290 ( .A1(DataRead[20]), .A2(DataRead[19]), .A3(DataRead[18]), .ZN(
        n2132) );
endmodule


module Bit_0 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_2 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_3 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_4 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_5 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_6 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_7 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_8 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_9 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_10 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_11 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_12 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_13 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_14 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_15 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_16 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_17 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_18 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_19 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_20 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_21 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_22 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_23 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_24 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_25 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_26 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_27 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_28 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_29 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_30 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_31 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_32 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_33 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_34 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_35 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_36 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_37 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_38 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_39 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_40 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_41 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_42 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_43 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_44 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_45 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_46 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_47 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_48 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_49 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_50 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_51 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_52 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_53 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_54 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_55 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_56 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_57 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_58 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_59 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_60 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_61 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_62 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_63 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_64 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_65 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_66 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_67 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_68 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_69 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_70 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_71 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_72 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_73 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_74 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_75 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_76 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_77 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_78 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_79 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_80 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_81 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_82 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_83 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_84 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_85 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_86 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_87 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_88 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_89 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_90 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_91 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_92 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_93 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_94 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_95 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_96 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_97 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_98 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_99 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_100 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_101 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_102 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_103 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_104 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_105 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_106 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_107 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_108 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_109 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_110 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_111 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_112 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_113 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_114 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_115 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_116 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_117 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_118 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_119 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_120 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_121 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_122 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_123 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_124 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_125 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_126 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_127 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_128 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_129 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_130 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_131 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_132 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_133 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_134 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_135 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_136 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_137 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_138 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_139 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_140 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_141 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_142 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_143 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_144 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_145 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_146 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_147 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_148 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_149 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_150 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_151 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_152 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_153 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_154 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_155 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_156 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_157 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_158 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_159 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_160 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_161 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_162 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_163 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_164 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_165 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_166 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_167 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_168 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_169 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_170 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_171 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_172 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_173 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_174 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_175 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_176 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_177 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_178 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_179 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_180 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_181 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_182 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_183 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_184 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_185 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_186 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_187 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_188 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_189 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_190 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_191 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_192 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_193 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_194 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_195 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_196 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_197 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_198 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_199 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_200 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_201 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_202 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_203 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_204 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_205 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_206 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_207 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_208 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_209 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_210 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_211 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_212 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_213 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_214 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_215 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_216 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_217 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_218 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_219 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_220 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_221 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_222 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_223 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_224 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_225 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_226 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_227 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_228 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_229 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_230 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_231 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_232 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_233 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_234 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_235 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_236 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_237 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_238 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_239 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_240 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_241 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_242 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_243 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_244 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_245 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_246 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_247 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_248 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_249 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_250 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_251 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_252 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_253 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_254 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_255 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_256 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_257 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_258 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_259 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_260 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_261 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_262 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_263 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_264 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_265 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_266 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_267 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_268 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_269 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_270 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_271 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_272 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_273 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_274 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_275 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_276 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_277 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_278 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_279 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_280 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_281 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_282 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_283 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_284 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_285 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_286 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_287 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_288 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_289 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_290 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_291 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_292 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_293 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_294 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_295 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_296 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_297 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_298 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_299 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_300 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_301 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_302 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_303 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_304 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_305 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_306 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_307 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_308 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_309 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_310 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_311 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_312 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_313 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_314 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_315 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_316 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_317 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_318 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_319 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_320 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_321 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_322 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_323 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_324 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_325 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_326 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_327 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_328 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_329 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_330 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_331 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_332 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_333 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_334 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_335 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_336 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_337 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_338 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_339 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_340 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_341 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_342 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_343 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_344 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_345 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_346 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_347 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_348 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_349 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_350 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_351 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_352 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_353 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_354 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_355 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_356 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_357 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_358 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_359 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_360 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_361 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_362 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_363 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_364 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_365 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_366 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_367 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_368 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_369 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_370 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_371 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_372 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_373 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_374 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_375 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_376 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_377 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_378 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_379 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_380 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_381 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_382 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_383 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_384 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_385 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_386 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_387 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_388 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_389 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_390 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_391 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_392 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_393 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_394 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_395 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_396 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_397 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_398 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_399 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_400 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_401 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_402 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_403 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_404 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_405 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_406 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_407 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_408 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_409 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_410 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_411 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_412 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_413 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_414 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_415 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_416 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_417 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_418 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_419 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_420 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_421 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_422 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_423 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_424 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_425 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_426 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_427 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_428 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_429 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_430 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_431 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_432 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_433 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_434 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_435 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_436 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_437 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_438 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_439 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_440 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_441 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_442 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_443 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_444 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_445 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_446 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_447 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_448 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_449 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_450 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_451 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_452 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_453 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_454 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_455 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_456 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_457 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_458 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_459 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_460 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_461 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_462 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_463 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_464 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_465 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_466 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_467 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_468 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_469 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_470 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_471 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_472 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_473 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_474 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_475 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_476 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_477 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_478 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_479 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_480 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_481 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_482 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_483 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_484 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_485 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_486 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_487 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_488 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_489 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_490 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_491 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_492 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_493 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_494 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_495 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_496 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_497 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_498 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_499 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_500 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_501 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_502 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_503 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_504 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_505 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_506 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_507 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_508 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_509 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_510 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_511 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_512 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_513 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_514 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_515 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_516 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_517 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_518 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_519 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_520 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_521 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_522 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_523 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_524 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_525 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_526 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_527 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_528 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_529 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_530 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_531 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_532 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_533 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_534 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_535 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_536 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_537 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_538 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_539 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_540 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_541 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_542 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_543 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_544 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_545 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_546 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_547 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_548 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_549 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_550 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_551 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_552 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_553 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_554 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_555 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_556 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_557 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_558 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_559 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_560 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_561 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_562 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_563 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_564 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_565 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_566 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_567 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_568 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_569 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_570 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_571 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_572 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_573 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_574 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_575 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_576 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_577 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_578 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_579 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_580 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_581 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_582 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_583 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_584 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_585 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_586 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_587 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_588 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_589 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_590 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_591 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_592 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_593 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_594 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_595 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_596 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_597 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_598 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_599 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_600 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_601 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_602 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_603 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_604 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_605 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_606 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_607 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_608 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_609 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_610 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_611 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_612 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_613 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_614 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_615 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_616 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_617 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_618 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_619 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_620 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_621 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_622 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_623 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_624 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_625 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_626 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_627 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_628 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_629 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_630 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_631 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_632 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_633 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_634 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_635 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_636 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_637 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_638 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_639 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_640 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_641 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_642 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_643 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_644 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_645 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_646 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_647 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_648 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_649 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_650 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_651 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_652 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_653 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_654 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_655 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_656 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_657 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_658 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_659 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_660 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_661 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_662 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_663 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_664 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_665 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_666 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_667 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_668 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_669 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_670 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_671 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_672 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_673 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_674 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_675 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_676 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_677 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_678 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_679 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_680 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_681 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_682 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_683 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_684 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_685 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_686 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_687 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_688 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_689 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_690 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_691 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_692 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_693 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_694 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_695 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_696 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_697 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_698 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_699 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_700 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_701 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_702 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_703 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_704 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_705 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_706 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_707 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_708 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_709 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_710 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_711 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_712 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_713 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_714 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_715 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_716 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_717 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_718 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_719 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_720 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_721 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_722 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_723 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_724 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_725 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_726 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_727 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_728 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_729 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_730 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_731 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_732 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_733 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_734 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_735 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_736 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_737 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_738 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_739 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_740 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_741 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_742 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_743 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_744 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_745 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_746 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_747 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_748 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_749 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_750 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_751 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_752 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_753 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_754 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_755 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_756 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_757 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_758 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_759 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_760 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_761 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_762 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_763 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_764 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_765 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_766 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_767 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_768 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_769 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_770 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_771 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_772 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_773 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_774 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_775 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_776 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_777 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_778 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_779 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_780 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_781 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_782 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_783 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_784 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_785 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_786 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_787 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_788 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_789 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_790 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_791 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_792 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_793 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_794 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_795 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_796 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_797 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_798 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_799 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_800 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_801 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_802 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_803 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_804 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_805 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_806 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_807 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_808 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_809 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_810 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_811 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_812 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_813 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_814 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_815 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_816 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_817 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_818 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_819 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_820 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_821 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_822 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_823 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_824 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_825 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_826 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_827 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_828 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_829 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_830 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_831 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_832 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_833 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_834 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_835 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_836 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_837 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_838 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_839 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_840 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_841 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_842 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_843 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_844 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_845 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_846 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_847 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_848 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_849 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_850 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_851 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_852 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_853 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_854 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_855 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_856 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_857 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_858 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_859 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_860 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_861 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_862 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_863 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_864 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_865 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_866 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_867 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_868 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_869 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_870 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_871 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_872 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_873 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_874 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_875 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_876 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_877 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_878 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_879 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_880 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_881 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_882 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_883 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_884 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_885 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_886 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_887 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_888 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_889 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_890 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_891 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_892 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_893 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_894 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_895 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_896 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_897 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_898 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_899 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_900 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_901 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_902 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_903 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_904 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_905 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_906 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_907 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_908 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_909 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_910 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_911 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_912 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_913 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_914 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_915 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_916 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_917 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_918 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_919 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_920 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_921 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_922 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_923 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_924 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_925 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_926 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_927 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_928 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_929 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_930 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_931 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_932 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_933 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_934 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_935 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_936 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_937 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_938 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_939 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_940 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_941 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_942 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_943 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_944 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_945 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_946 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_947 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_948 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_949 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_950 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_951 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_952 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_953 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_954 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_955 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_956 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_957 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_958 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_959 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_960 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_961 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_962 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_963 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_964 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_965 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_966 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_967 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_968 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_969 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_970 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_971 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_972 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_973 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_974 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_975 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_976 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_977 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_978 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_979 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_980 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_981 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_982 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_983 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_984 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_985 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_986 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_987 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_988 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_989 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_990 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_991 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_992 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_993 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_994 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_995 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_996 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_997 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_998 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_999 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1000 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1001 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1002 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1003 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1004 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1005 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1006 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1007 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1008 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1009 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1010 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1011 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1012 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1013 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1014 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1015 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1016 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1017 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1018 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1019 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1020 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1021 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1022 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1023 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1024 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1025 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1026 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1027 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1028 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1029 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1030 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1031 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1032 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1033 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1034 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1035 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1036 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1037 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1038 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1039 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1040 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1041 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1042 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1043 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1044 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1045 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1046 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1047 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1048 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1049 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1050 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1051 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1052 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1053 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1054 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module Bit_1055 ( Q, D, Clk );
  input D, Clk;
  output Q;


  DFQD1 QReg_reg ( .D(D), .CP(Clk), .Q(Q) );
endmodule


module FIFOStateM_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_4 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

