library verilog;
use verilog.vl_types.all;
entity uart_eeprom_tb is
end uart_eeprom_tb;
