
`ifndef RKV_I2C_TESTS_SVH
`define RKV_I2C_TESTS_SVH

`include "rkv_i2c_base_test.sv"
`include "rkv_i2c_quick_reg_access_test.sv"
`include "rkv_i2c_master_directed_interrupt_test.sv"
`include "rkv_i2c_master_directed_write_packet_test.sv"
`include "rkv_i2c_master_directed_read_packet_test.sv"

`endif // RKV_I2C_TESTS_SVH
