
module FIFO_Top ( Dout, Din, ReadIn, WriteIn, Clocker, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, Clocker, Reseter;
  wire   E_FIFO, F_FIFO, Mem_Enable, ReadWire, WriteWire, _0_net_, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40;
  wire   [4:0] SM_MemAddr;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(E_FIFO), .FullFIFO(F_FIFO), .ReadCmd(ReadWire), .WriteCmd(
        WriteWire), .ReadReq(ReadIn), .WriteReq(WriteIn), .Clk(Clocker), 
        .Reset(Reseter) );
  Mem1kx32 RegFile1 ( .DataO(Dout), .DataI({n23, n39, n36, n10, n14, n35, n32, 
        n19, n20, n31, n30, n16, n12, n27, n24, n8, n33, n34, n11, n13, n26, 
        n29, n17, n37, n38, n21, n9, n25, n28, n18, n22, n15}), .Addr({
        SM_MemAddr[4], n7, SM_MemAddr[2:0]}), .ClockIn(_0_net_), .ChipEna(
        Mem_Enable), .Read(ReadWire), .Write(WriteWire) );
  AO211D1 U10 ( .A1(WriteWire), .A2(ReadWire), .B(F_FIFO), .C(E_FIFO), .Z(n6)
         );
  INVD1 U11 ( .I(n6), .ZN(Mem_Enable) );
  MUX2D0 U12 ( .I0(SM_WriteAddr[3]), .I1(SM_ReadAddr[3]), .S(n40), .Z(n7) );
  MUX2D0 U13 ( .I0(SM_WriteAddr[4]), .I1(SM_ReadAddr[4]), .S(n40), .Z(
        SM_MemAddr[4]) );
  BUFFD1 U14 ( .I(Din[16]), .Z(n8) );
  BUFFD1 U15 ( .I(Din[5]), .Z(n9) );
  BUFFD1 U16 ( .I(Din[28]), .Z(n10) );
  BUFFD1 U17 ( .I(Din[13]), .Z(n11) );
  BUFFD1 U18 ( .I(Din[19]), .Z(n12) );
  BUFFD1 U19 ( .I(Din[12]), .Z(n13) );
  BUFFD1 U20 ( .I(Din[27]), .Z(n14) );
  BUFFD1 U21 ( .I(Din[0]), .Z(n15) );
  BUFFD1 U22 ( .I(Din[20]), .Z(n16) );
  BUFFD1 U23 ( .I(Din[9]), .Z(n17) );
  BUFFD1 U24 ( .I(Din[2]), .Z(n18) );
  BUFFD1 U25 ( .I(Din[24]), .Z(n19) );
  BUFFD1 U26 ( .I(Din[23]), .Z(n20) );
  BUFFD1 U27 ( .I(Din[6]), .Z(n21) );
  BUFFD1 U28 ( .I(Din[1]), .Z(n22) );
  BUFFD1 U29 ( .I(Din[31]), .Z(n23) );
  BUFFD1 U30 ( .I(Din[17]), .Z(n24) );
  BUFFD1 U31 ( .I(Din[4]), .Z(n25) );
  BUFFD1 U32 ( .I(Din[11]), .Z(n26) );
  BUFFD1 U33 ( .I(Din[18]), .Z(n27) );
  BUFFD1 U34 ( .I(Din[3]), .Z(n28) );
  BUFFD1 U35 ( .I(Din[10]), .Z(n29) );
  BUFFD1 U36 ( .I(Din[21]), .Z(n30) );
  BUFFD1 U37 ( .I(Din[22]), .Z(n31) );
  BUFFD1 U38 ( .I(Din[25]), .Z(n32) );
  BUFFD1 U39 ( .I(Din[15]), .Z(n33) );
  BUFFD1 U40 ( .I(Din[14]), .Z(n34) );
  BUFFD1 U41 ( .I(Din[26]), .Z(n35) );
  BUFFD1 U42 ( .I(Din[29]), .Z(n36) );
  BUFFD1 U43 ( .I(Din[8]), .Z(n37) );
  BUFFD1 U44 ( .I(Din[7]), .Z(n38) );
  BUFFD1 U45 ( .I(Din[30]), .Z(n39) );
  CKND0 U46 ( .CLK(Clocker), .CN(_0_net_) );
  MUX2D0 U47 ( .I0(SM_WriteAddr[2]), .I1(SM_ReadAddr[2]), .S(n40), .Z(
        SM_MemAddr[2]) );
  MUX2D0 U48 ( .I0(SM_WriteAddr[1]), .I1(SM_ReadAddr[1]), .S(n40), .Z(
        SM_MemAddr[1]) );
  MUX2D0 U49 ( .I0(SM_WriteAddr[0]), .I1(SM_ReadAddr[0]), .S(n40), .Z(
        SM_MemAddr[0]) );
  INR2D0 U50 ( .A1(ReadWire), .B1(WriteWire), .ZN(n40) );
endmodule


module FIFOStateM ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, Clk, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, Clk, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, \CurState[1] , N72, N73, N74,
         N75, N76, N88, N89, N90, N91, N92, N93, N106, N107, N108, N109, N110,
         N111, N124, N125, N126, N127, N128, N144, N146, N148, N150, N152,
         N155, N158, N161, N164, N167, N169, N172, N175, N178, N181, N184,
         N186, N187, N190, N191, N200, N201, N202, N211, N212, N213, N214,
         N217, N220, N223, N226, N229, N232, N235, N238, N241, n2, \U3/U1/Z_0 ,
         \U3/U1/Z_1 , \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n1, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71;
  wire   [2:0] NextState;

  LHQD1 \WriteCount_tri_enable_reg[0]  ( .E(N200), .D(N201), .Q(N9) );
  LHQD1 \NextState_reg[0]  ( .E(N190), .D(N144), .Q(NextState[0]) );
  LHQD1 \WriteCount_reg[1]  ( .E(N200), .D(N155), .Q(N238) );
  LHQD1 \ReadCount_reg[1]  ( .E(N211), .D(N172), .Q(N223) );
  LHQD1 \WriteCount_reg[4]  ( .E(N200), .D(N164), .Q(N229) );
  LHQD1 \ReadCount_reg[4]  ( .E(N211), .D(N181), .Q(N214) );
  LHQD1 \NextState_reg[1]  ( .E(N190), .D(N146), .Q(NextState[1]) );
  LHQD1 \NextState_reg[2]  ( .E(N190), .D(N148), .Q(NextState[2]) );
  LHQD1 EmptyFIFOReg_reg ( .E(N213), .D(N184), .Q(EmptyFIFO) );
  LHQD1 \ReadCount_tri_enable_reg[4]  ( .E(N211), .D(N212), .Q(N0) );
  LHQD1 \ReadCount_tri_enable_reg[2]  ( .E(N211), .D(N212), .Q(N2) );
  LHQD1 \ReadCount_tri_enable_reg[0]  ( .E(N211), .D(N212), .Q(N4) );
  LHQD1 \ReadCount_tri_enable_reg[1]  ( .E(N211), .D(N212), .Q(N3) );
  LHQD1 \ReadCount_tri_enable_reg[3]  ( .E(N211), .D(N212), .Q(N1) );
  LHQD1 \WriteCount_tri_enable_reg[4]  ( .E(N200), .D(N201), .Q(N5) );
  LHQD1 \WriteCount_tri_enable_reg[2]  ( .E(N200), .D(N201), .Q(N7) );
  LHQD1 \WriteCount_tri_enable_reg[1]  ( .E(N200), .D(N201), .Q(N8) );
  LHQD1 \WriteCount_tri_enable_reg[3]  ( .E(N200), .D(N201), .Q(N6) );
  LHQD1 FullFIFOReg_reg ( .E(N191), .D(N150), .Q(FullFIFO) );
  LHQD1 ReadCmdReg_reg ( .E(N187), .D(N186), .Q(ReadCmd) );
  LHQD1 WriteCmdReg_reg ( .E(N202), .D(N167), .Q(WriteCmd) );
  LHQD1 \ReadCount_reg[2]  ( .E(N211), .D(N175), .Q(N220) );
  LHQD1 \WriteCount_reg[2]  ( .E(N200), .D(N158), .Q(N235) );
  LHQD1 \WriteCount_reg[3]  ( .E(N200), .D(N161), .Q(N232) );
  LHQD1 \ReadCount_reg[3]  ( .E(N211), .D(N178), .Q(N217) );
  LHQD1 \ReadCount_reg[0]  ( .E(N211), .D(N169), .Q(N226) );
  LHQD1 \WriteCount_reg[0]  ( .E(N200), .D(N152), .Q(N241) );
  BUFTD1 \WriteCount_tri[0]  ( .I(N241), .OE(n96), .Z(WriteAddr[0]) );
  BUFTD1 \WriteCount_tri[1]  ( .I(N238), .OE(n95), .Z(WriteAddr[1]) );
  BUFTD1 \WriteCount_tri[2]  ( .I(N235), .OE(n94), .Z(WriteAddr[2]) );
  BUFTD1 \WriteCount_tri[3]  ( .I(N232), .OE(n93), .Z(WriteAddr[3]) );
  BUFTD1 \WriteCount_tri[4]  ( .I(N229), .OE(n92), .Z(WriteAddr[4]) );
  BUFTD1 \ReadCount_tri[0]  ( .I(N226), .OE(n91), .Z(ReadAddr[0]) );
  BUFTD1 \ReadCount_tri[1]  ( .I(N223), .OE(n90), .Z(ReadAddr[1]) );
  BUFTD1 \ReadCount_tri[2]  ( .I(N220), .OE(n89), .Z(ReadAddr[2]) );
  BUFTD1 \ReadCount_tri[3]  ( .I(N217), .OE(n88), .Z(ReadAddr[3]) );
  BUFTD1 \ReadCount_tri[4]  ( .I(N214), .OE(n87), .Z(ReadAddr[4]) );
  FIFOStateM_DW01_inc_0 add_199 ( .A({n2, N76, N75, N74, N73, N72}), .SUM({N93, 
        N92, N91, N90, N89, N88}) );
  FIFOStateM_DW01_inc_1 r147 ( .A(WriteAddr), .SUM({N76, N75, N74, N73, N72})
         );
  FIFOStateM_DW01_inc_2 add_211 ( .A({n2, N128, N127, N126, N125, N124}), 
        .SUM({N111, N110, N109, N108, N107, N106}) );
  FIFOStateM_DW01_inc_3 r133 ( .A({\U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , 
        \U3/U1/Z_1 , \U3/U1/Z_0 }), .SUM({N128, N127, N126, N125, N124}) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(Clk), .CDN(n97), .Q(
        \CurState[1] ) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(Clk), .CDN(n97), .Q(n70), 
        .QN(n1) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(Clk), .CDN(n97), .Q(n71) );
  AOI31D0 U3 ( .A1(n34), .A2(n53), .A3(n19), .B(n32), .ZN(n6) );
  ND3D1 U4 ( .A1(n1), .A2(n71), .A3(\CurState[1] ), .ZN(n53) );
  OAI21D1 U5 ( .A1(n55), .A2(n17), .B(n38), .ZN(n37) );
  AOI21D1 U6 ( .A1(n13), .A2(n22), .B(Clk), .ZN(N211) );
  TIEL U7 ( .ZN(n2) );
  CKND0 U8 ( .CLK(N9), .CN(n96) );
  CKND0 U9 ( .CLK(N8), .CN(n95) );
  CKND0 U10 ( .CLK(N7), .CN(n94) );
  CKND0 U11 ( .CLK(N6), .CN(n93) );
  CKND0 U12 ( .CLK(N5), .CN(n92) );
  CKND0 U13 ( .CLK(N4), .CN(n91) );
  CKND0 U14 ( .CLK(N3), .CN(n90) );
  CKND0 U15 ( .CLK(N2), .CN(n89) );
  CKND0 U16 ( .CLK(N1), .CN(n88) );
  CKND0 U17 ( .CLK(N0), .CN(n87) );
  IOA22D0 U18 ( .B1(n4), .B2(n5), .A1(n6), .A2(ReadAddr[4]), .ZN(\U3/U1/Z_4 )
         );
  IOA22D0 U19 ( .B1(n4), .B2(n7), .A1(n6), .A2(ReadAddr[3]), .ZN(\U3/U1/Z_3 )
         );
  IOA22D0 U20 ( .B1(n4), .B2(n8), .A1(n6), .A2(ReadAddr[2]), .ZN(\U3/U1/Z_2 )
         );
  IOA22D0 U21 ( .B1(n4), .B2(n9), .A1(n6), .A2(ReadAddr[1]), .ZN(\U3/U1/Z_1 )
         );
  IOA22D0 U22 ( .B1(n4), .B2(n10), .A1(n6), .A2(ReadAddr[0]), .ZN(\U3/U1/Z_0 )
         );
  CKND2D0 U23 ( .A1(n11), .A2(n97), .ZN(n4) );
  AOI21D0 U24 ( .A1(n12), .A2(n13), .B(Clk), .ZN(N213) );
  INR2D0 U25 ( .A1(N184), .B1(Clk), .ZN(N212) );
  AOI31D0 U26 ( .A1(n14), .A2(n15), .A3(n16), .B(Clk), .ZN(N202) );
  CKND0 U27 ( .CLK(N186), .CN(n15) );
  CKND2D0 U28 ( .A1(n17), .A2(n18), .ZN(n14) );
  INR2D0 U29 ( .A1(N150), .B1(Clk), .ZN(N201) );
  AOI21D0 U30 ( .A1(n16), .A2(n19), .B(Clk), .ZN(N200) );
  AOI21D0 U31 ( .A1(n20), .A2(n21), .B(Clk), .ZN(N191) );
  AOI31D0 U32 ( .A1(n16), .A2(n22), .A3(n23), .B(Clk), .ZN(N190) );
  NR2D0 U33 ( .A1(n24), .A2(n25), .ZN(n23) );
  MUX2ND0 U34 ( .I0(n26), .I1(n71), .S(n70), .ZN(n25) );
  CKND2D0 U35 ( .A1(n71), .A2(n27), .ZN(n26) );
  INR3D0 U36 ( .A1(n21), .B1(n28), .B2(n11), .ZN(n16) );
  CKND2D0 U37 ( .A1(n29), .A2(Reset), .ZN(n21) );
  IND2D0 U38 ( .A1(N211), .B1(n30), .ZN(N187) );
  OAI21D0 U39 ( .A1(n28), .A2(n24), .B(n31), .ZN(n30) );
  CKND0 U40 ( .CLK(Clk), .CN(n31) );
  OAI22D0 U41 ( .A1(n32), .A2(n12), .B1(n33), .B2(n34), .ZN(n24) );
  NR2D0 U42 ( .A1(n33), .A2(n35), .ZN(n28) );
  CKND0 U43 ( .CLK(n6), .CN(n22) );
  ND3D0 U44 ( .A1(n36), .A2(n19), .A3(n37), .ZN(N186) );
  NR2D0 U45 ( .A1(n13), .A2(n18), .ZN(N184) );
  CKND0 U46 ( .CLK(n29), .CN(n13) );
  OAI22D0 U47 ( .A1(n39), .A2(n40), .B1(n5), .B2(n41), .ZN(N181) );
  CKND0 U48 ( .CLK(N128), .CN(n40) );
  OAI22D0 U49 ( .A1(n39), .A2(n42), .B1(n7), .B2(n41), .ZN(N178) );
  CKND0 U50 ( .CLK(N127), .CN(n42) );
  OAI22D0 U51 ( .A1(n39), .A2(n43), .B1(n8), .B2(n41), .ZN(N175) );
  CKND0 U52 ( .CLK(WriteAddr[2]), .CN(n8) );
  CKND0 U53 ( .CLK(N126), .CN(n43) );
  OAI22D0 U54 ( .A1(n39), .A2(n44), .B1(n9), .B2(n41), .ZN(N172) );
  CKND0 U55 ( .CLK(N125), .CN(n44) );
  OAI22D0 U56 ( .A1(n39), .A2(n45), .B1(n10), .B2(n41), .ZN(N169) );
  CKND2D0 U57 ( .A1(n29), .A2(n97), .ZN(n41) );
  CKND0 U58 ( .CLK(Reset), .CN(n97) );
  CKND0 U59 ( .CLK(WriteAddr[0]), .CN(n10) );
  CKND0 U60 ( .CLK(N124), .CN(n45) );
  INR2D0 U61 ( .A1(n20), .B1(n46), .ZN(n39) );
  OAI21D0 U62 ( .A1(n38), .A2(n47), .B(n48), .ZN(N167) );
  NR2D0 U63 ( .A1(n17), .A2(n49), .ZN(n47) );
  AO222D0 U64 ( .A1(ReadAddr[4]), .A2(n50), .B1(N128), .B2(n11), .C1(N76), 
        .C2(n49), .Z(N164) );
  AO222D0 U65 ( .A1(ReadAddr[3]), .A2(n50), .B1(N127), .B2(n11), .C1(N75), 
        .C2(n49), .Z(N161) );
  AO222D0 U66 ( .A1(ReadAddr[2]), .A2(n50), .B1(N126), .B2(n11), .C1(N74), 
        .C2(n49), .Z(N158) );
  AO222D0 U67 ( .A1(ReadAddr[1]), .A2(n50), .B1(N125), .B2(n11), .C1(N73), 
        .C2(n49), .Z(N155) );
  AO222D0 U68 ( .A1(ReadAddr[0]), .A2(n50), .B1(N124), .B2(n11), .C1(N72), 
        .C2(n49), .Z(N152) );
  CKND0 U69 ( .CLK(n48), .CN(n11) );
  NR2D0 U70 ( .A1(n19), .A2(n38), .ZN(N150) );
  OAI21D0 U71 ( .A1(n38), .A2(n51), .B(n19), .ZN(N148) );
  IAO21D0 U72 ( .A1(n52), .A2(n53), .B(n17), .ZN(n51) );
  ND4D0 U73 ( .A1(n36), .A2(n34), .A3(n48), .A4(n54), .ZN(N146) );
  AOI22D0 U74 ( .A1(n46), .A2(n52), .B1(n55), .B2(n32), .ZN(n54) );
  CKND0 U75 ( .CLK(n38), .CN(n32) );
  ND4D0 U76 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(n52) );
  NR3D0 U77 ( .A1(n60), .A2(N93), .A3(n61), .ZN(n59) );
  CKXOR2D0 U78 ( .A1(ReadAddr[0]), .A2(N88), .Z(n61) );
  CKXOR2D0 U79 ( .A1(ReadAddr[4]), .A2(N92), .Z(n60) );
  XNR2D0 U80 ( .A1(N90), .A2(ReadAddr[2]), .ZN(n58) );
  XNR2D0 U81 ( .A1(N91), .A2(ReadAddr[3]), .ZN(n57) );
  XNR2D0 U82 ( .A1(N89), .A2(ReadAddr[1]), .ZN(n56) );
  CKND2D0 U83 ( .A1(n18), .A2(n29), .ZN(n48) );
  NR3D0 U84 ( .A1(n71), .A2(n70), .A3(\CurState[1] ), .ZN(n29) );
  CKND0 U85 ( .CLK(n33), .CN(n18) );
  CKND2D0 U86 ( .A1(WriteReq), .A2(n62), .ZN(n33) );
  CKND2D0 U87 ( .A1(n38), .A2(n46), .ZN(n36) );
  CKND0 U88 ( .CLK(n53), .CN(n46) );
  OAI221D0 U89 ( .A1(n63), .A2(n53), .B1(n38), .B2(n35), .C(n20), .ZN(N144) );
  NR2D0 U90 ( .A1(n50), .A2(n17), .ZN(n20) );
  CKND0 U91 ( .CLK(n34), .CN(n17) );
  ND3D0 U92 ( .A1(n71), .A2(n27), .A3(n70), .ZN(n34) );
  CKND0 U93 ( .CLK(n19), .CN(n50) );
  ND3D0 U94 ( .A1(n71), .A2(\CurState[1] ), .A3(n70), .ZN(n19) );
  CKND0 U95 ( .CLK(n49), .CN(n35) );
  CKND2D0 U96 ( .A1(n12), .A2(n53), .ZN(n49) );
  CKND0 U97 ( .CLK(n55), .CN(n12) );
  NR3D0 U98 ( .A1(n71), .A2(n70), .A3(n27), .ZN(n55) );
  CKND0 U99 ( .CLK(\CurState[1] ), .CN(n27) );
  NR2D0 U100 ( .A1(n62), .A2(WriteReq), .ZN(n38) );
  CKND0 U101 ( .CLK(ReadReq), .CN(n62) );
  NR4D0 U102 ( .A1(n64), .A2(n65), .A3(N111), .A4(n66), .ZN(n63) );
  CKXOR2D0 U103 ( .A1(WriteAddr[2]), .A2(N108), .Z(n66) );
  CKXOR2D0 U104 ( .A1(WriteAddr[0]), .A2(N106), .Z(n65) );
  ND3D0 U105 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n64) );
  CKXOR2D0 U106 ( .A1(N110), .A2(n5), .Z(n69) );
  CKND0 U107 ( .CLK(WriteAddr[4]), .CN(n5) );
  CKXOR2D0 U108 ( .A1(N107), .A2(n9), .Z(n68) );
  CKND0 U109 ( .CLK(WriteAddr[1]), .CN(n9) );
  CKXOR2D0 U110 ( .A1(N109), .A2(n7), .Z(n67) );
  CKND0 U111 ( .CLK(WriteAddr[3]), .CN(n7) );
endmodule


module Mem1kx32 ( Dready, ParityErr, DataO, DataI, Addr, ClockIn, ChipEna, 
        Read, Write );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] Addr;
  input ClockIn, ChipEna, Read, Write;
  output Dready, ParityErr;
  wire   N43, N44, N45, N46, N47, ChipClock, DreadyReg, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N84, N2262, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799;
  wire   [31:0] DataOreg;
  assign N43 = Addr[0];
  assign N44 = Addr[1];
  assign N45 = Addr[2];
  assign N46 = Addr[3];
  assign N47 = Addr[4];

  EDFQD1 \Storage_reg[26][32]  ( .D(n202), .E(n153), .CP(n239), .Q(
        \Storage[26][32] ) );
  EDFQD1 \Storage_reg[26][31]  ( .D(n63), .E(n153), .CP(n238), .Q(
        \Storage[26][31] ) );
  EDFQD1 \Storage_reg[26][30]  ( .D(n62), .E(n154), .CP(n238), .Q(
        \Storage[26][30] ) );
  EDFQD1 \Storage_reg[26][29]  ( .D(n58), .E(n154), .CP(n238), .Q(
        \Storage[26][29] ) );
  EDFQD1 \Storage_reg[26][28]  ( .D(n53), .E(n153), .CP(n238), .Q(
        \Storage[26][28] ) );
  EDFQD1 \Storage_reg[26][27]  ( .D(n49), .E(n152), .CP(n238), .Q(
        \Storage[26][27] ) );
  EDFQD1 \Storage_reg[26][26]  ( .D(n46), .E(n152), .CP(n238), .Q(
        \Storage[26][26] ) );
  EDFQD1 \Storage_reg[26][25]  ( .D(n42), .E(n153), .CP(n238), .Q(
        \Storage[26][25] ) );
  EDFQD1 \Storage_reg[26][24]  ( .D(n37), .E(n152), .CP(n238), .Q(
        \Storage[26][24] ) );
  EDFQD1 \Storage_reg[26][23]  ( .D(n33), .E(n154), .CP(n238), .Q(
        \Storage[26][23] ) );
  EDFQD1 \Storage_reg[26][22]  ( .D(n30), .E(n153), .CP(n238), .Q(
        \Storage[26][22] ) );
  EDFQD1 \Storage_reg[26][21]  ( .D(n26), .E(n152), .CP(n238), .Q(
        \Storage[26][21] ) );
  EDFQD1 \Storage_reg[26][20]  ( .D(n21), .E(n154), .CP(n237), .Q(
        \Storage[26][20] ) );
  EDFQD1 \Storage_reg[26][19]  ( .D(n17), .E(n152), .CP(n237), .Q(
        \Storage[26][19] ) );
  EDFQD1 \Storage_reg[26][18]  ( .D(n14), .E(n152), .CP(n237), .Q(
        \Storage[26][18] ) );
  EDFQD1 \Storage_reg[26][17]  ( .D(n10), .E(n153), .CP(n237), .Q(
        \Storage[26][17] ) );
  EDFQD1 \Storage_reg[26][16]  ( .D(n5), .E(n154), .CP(n237), .Q(
        \Storage[26][16] ) );
  EDFQD1 \Storage_reg[26][15]  ( .D(n2), .E(n154), .CP(n237), .Q(
        \Storage[26][15] ) );
  EDFQD1 \Storage_reg[26][14]  ( .D(n4), .E(n153), .CP(n237), .Q(
        \Storage[26][14] ) );
  EDFQD1 \Storage_reg[26][13]  ( .D(n7), .E(n152), .CP(n237), .Q(
        \Storage[26][13] ) );
  EDFQD1 \Storage_reg[26][12]  ( .D(n11), .E(n152), .CP(n237), .Q(
        \Storage[26][12] ) );
  EDFQD1 \Storage_reg[26][11]  ( .D(n16), .E(n153), .CP(n237), .Q(
        \Storage[26][11] ) );
  EDFQD1 \Storage_reg[26][10]  ( .D(n20), .E(n154), .CP(n237), .Q(
        \Storage[26][10] ) );
  EDFQD1 \Storage_reg[26][9]  ( .D(n23), .E(n154), .CP(n236), .Q(
        \Storage[26][9] ) );
  EDFQD1 \Storage_reg[26][8]  ( .D(n28), .E(n153), .CP(n236), .Q(
        \Storage[26][8] ) );
  EDFQD1 \Storage_reg[26][7]  ( .D(n32), .E(n152), .CP(n236), .Q(
        \Storage[26][7] ) );
  EDFQD1 \Storage_reg[26][6]  ( .D(n35), .E(n152), .CP(n236), .Q(
        \Storage[26][6] ) );
  EDFQD1 \Storage_reg[26][5]  ( .D(n39), .E(n153), .CP(n236), .Q(
        \Storage[26][5] ) );
  EDFQD1 \Storage_reg[26][4]  ( .D(n44), .E(n154), .CP(n236), .Q(
        \Storage[26][4] ) );
  EDFQD1 \Storage_reg[26][3]  ( .D(n48), .E(n154), .CP(n236), .Q(
        \Storage[26][3] ) );
  EDFQD1 \Storage_reg[26][2]  ( .D(n51), .E(n153), .CP(n236), .Q(
        \Storage[26][2] ) );
  EDFQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(n154), .CP(n236), .Q(
        \Storage[26][1] ) );
  EDFQD1 \Storage_reg[26][0]  ( .D(n59), .E(n152), .CP(n236), .Q(
        \Storage[26][0] ) );
  EDFQD1 \Storage_reg[24][32]  ( .D(n202), .E(n137), .CP(n233), .Q(
        \Storage[24][32] ) );
  EDFQD1 \Storage_reg[24][31]  ( .D(n64), .E(n137), .CP(n232), .Q(
        \Storage[24][31] ) );
  EDFQD1 \Storage_reg[24][30]  ( .D(n62), .E(n138), .CP(n232), .Q(
        \Storage[24][30] ) );
  EDFQD1 \Storage_reg[24][29]  ( .D(n58), .E(n138), .CP(n232), .Q(
        \Storage[24][29] ) );
  EDFQD1 \Storage_reg[24][28]  ( .D(n54), .E(n137), .CP(n232), .Q(
        \Storage[24][28] ) );
  EDFQD1 \Storage_reg[24][27]  ( .D(n50), .E(n136), .CP(n232), .Q(
        \Storage[24][27] ) );
  EDFQD1 \Storage_reg[24][26]  ( .D(n46), .E(n136), .CP(n232), .Q(
        \Storage[24][26] ) );
  EDFQD1 \Storage_reg[24][25]  ( .D(n42), .E(n137), .CP(n232), .Q(
        \Storage[24][25] ) );
  EDFQD1 \Storage_reg[24][24]  ( .D(n38), .E(n136), .CP(n232), .Q(
        \Storage[24][24] ) );
  EDFQD1 \Storage_reg[24][23]  ( .D(n34), .E(n138), .CP(n232), .Q(
        \Storage[24][23] ) );
  EDFQD1 \Storage_reg[24][22]  ( .D(n30), .E(n137), .CP(n232), .Q(
        \Storage[24][22] ) );
  EDFQD1 \Storage_reg[24][21]  ( .D(n26), .E(n136), .CP(n232), .Q(
        \Storage[24][21] ) );
  EDFQD1 \Storage_reg[24][20]  ( .D(n22), .E(n138), .CP(n231), .Q(
        \Storage[24][20] ) );
  EDFQD1 \Storage_reg[24][19]  ( .D(n18), .E(n136), .CP(n231), .Q(
        \Storage[24][19] ) );
  EDFQD1 \Storage_reg[24][18]  ( .D(n14), .E(n136), .CP(n231), .Q(
        \Storage[24][18] ) );
  EDFQD1 \Storage_reg[24][17]  ( .D(n10), .E(n137), .CP(n231), .Q(
        \Storage[24][17] ) );
  EDFQD1 \Storage_reg[24][16]  ( .D(n6), .E(n138), .CP(n231), .Q(
        \Storage[24][16] ) );
  EDFQD1 \Storage_reg[24][15]  ( .D(n2), .E(n138), .CP(n231), .Q(
        \Storage[24][15] ) );
  EDFQD1 \Storage_reg[24][14]  ( .D(n4), .E(n137), .CP(n231), .Q(
        \Storage[24][14] ) );
  EDFQD1 \Storage_reg[24][13]  ( .D(n8), .E(n136), .CP(n231), .Q(
        \Storage[24][13] ) );
  EDFQD1 \Storage_reg[24][12]  ( .D(n12), .E(n136), .CP(n231), .Q(
        \Storage[24][12] ) );
  EDFQD1 \Storage_reg[24][11]  ( .D(n16), .E(n137), .CP(n231), .Q(
        \Storage[24][11] ) );
  EDFQD1 \Storage_reg[24][10]  ( .D(n20), .E(n138), .CP(n231), .Q(
        \Storage[24][10] ) );
  EDFQD1 \Storage_reg[24][9]  ( .D(n24), .E(n138), .CP(n230), .Q(
        \Storage[24][9] ) );
  EDFQD1 \Storage_reg[24][8]  ( .D(n28), .E(n137), .CP(n230), .Q(
        \Storage[24][8] ) );
  EDFQD1 \Storage_reg[24][7]  ( .D(n32), .E(n136), .CP(n230), .Q(
        \Storage[24][7] ) );
  EDFQD1 \Storage_reg[24][6]  ( .D(n36), .E(n136), .CP(n230), .Q(
        \Storage[24][6] ) );
  EDFQD1 \Storage_reg[24][5]  ( .D(n40), .E(n137), .CP(n230), .Q(
        \Storage[24][5] ) );
  EDFQD1 \Storage_reg[24][4]  ( .D(n44), .E(n138), .CP(n230), .Q(
        \Storage[24][4] ) );
  EDFQD1 \Storage_reg[24][3]  ( .D(n48), .E(n138), .CP(n230), .Q(
        \Storage[24][3] ) );
  EDFQD1 \Storage_reg[24][2]  ( .D(n51), .E(n137), .CP(n230), .Q(
        \Storage[24][2] ) );
  EDFQD1 \Storage_reg[24][1]  ( .D(n56), .E(n138), .CP(n230), .Q(
        \Storage[24][1] ) );
  EDFQD1 \Storage_reg[24][0]  ( .D(n60), .E(n136), .CP(n230), .Q(
        \Storage[24][0] ) );
  EDFQD1 \Storage_reg[30][32]  ( .D(n201), .E(n185), .CP(n251), .Q(
        \Storage[30][32] ) );
  EDFQD1 \Storage_reg[30][31]  ( .D(n63), .E(n185), .CP(n250), .Q(
        \Storage[30][31] ) );
  EDFQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n186), .CP(n250), .Q(
        \Storage[30][30] ) );
  EDFQD1 \Storage_reg[30][29]  ( .D(n57), .E(n186), .CP(n250), .Q(
        \Storage[30][29] ) );
  EDFQD1 \Storage_reg[30][28]  ( .D(n53), .E(n185), .CP(n250), .Q(
        \Storage[30][28] ) );
  EDFQD1 \Storage_reg[30][27]  ( .D(n49), .E(n184), .CP(n250), .Q(
        \Storage[30][27] ) );
  EDFQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n184), .CP(n250), .Q(
        \Storage[30][26] ) );
  EDFQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n185), .CP(n250), .Q(
        \Storage[30][25] ) );
  EDFQD1 \Storage_reg[30][24]  ( .D(n37), .E(n184), .CP(n250), .Q(
        \Storage[30][24] ) );
  EDFQD1 \Storage_reg[30][23]  ( .D(n33), .E(n186), .CP(n250), .Q(
        \Storage[30][23] ) );
  EDFQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(n185), .CP(n250), .Q(
        \Storage[30][22] ) );
  EDFQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n184), .CP(n250), .Q(
        \Storage[30][21] ) );
  EDFQD1 \Storage_reg[30][20]  ( .D(n21), .E(n186), .CP(n249), .Q(
        \Storage[30][20] ) );
  EDFQD1 \Storage_reg[30][19]  ( .D(n17), .E(n184), .CP(n249), .Q(
        \Storage[30][19] ) );
  EDFQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n184), .CP(n249), .Q(
        \Storage[30][18] ) );
  EDFQD1 \Storage_reg[30][17]  ( .D(n9), .E(n185), .CP(n249), .Q(
        \Storage[30][17] ) );
  EDFQD1 \Storage_reg[30][16]  ( .D(n5), .E(n186), .CP(n249), .Q(
        \Storage[30][16] ) );
  EDFQD1 \Storage_reg[30][15]  ( .D(n1), .E(n186), .CP(n249), .Q(
        \Storage[30][15] ) );
  EDFQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n185), .CP(n249), .Q(
        \Storage[30][14] ) );
  EDFQD1 \Storage_reg[30][13]  ( .D(n7), .E(n184), .CP(n249), .Q(
        \Storage[30][13] ) );
  EDFQD1 \Storage_reg[30][12]  ( .D(n11), .E(n184), .CP(n249), .Q(
        \Storage[30][12] ) );
  EDFQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n185), .CP(n249), .Q(
        \Storage[30][11] ) );
  EDFQD1 \Storage_reg[30][10]  ( .D(n19), .E(n186), .CP(n249), .Q(
        \Storage[30][10] ) );
  EDFQD1 \Storage_reg[30][9]  ( .D(n23), .E(n186), .CP(n248), .Q(
        \Storage[30][9] ) );
  EDFQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n185), .CP(n248), .Q(
        \Storage[30][8] ) );
  EDFQD1 \Storage_reg[30][7]  ( .D(n31), .E(n184), .CP(n248), .Q(
        \Storage[30][7] ) );
  EDFQD1 \Storage_reg[30][6]  ( .D(n35), .E(n184), .CP(n248), .Q(
        \Storage[30][6] ) );
  EDFQD1 \Storage_reg[30][5]  ( .D(n39), .E(n185), .CP(n248), .Q(
        \Storage[30][5] ) );
  EDFQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(n186), .CP(n248), .Q(
        \Storage[30][4] ) );
  EDFQD1 \Storage_reg[30][3]  ( .D(n47), .E(n186), .CP(n248), .Q(
        \Storage[30][3] ) );
  EDFQD1 \Storage_reg[30][2]  ( .D(n52), .E(n185), .CP(n248), .Q(
        \Storage[30][2] ) );
  EDFQD1 \Storage_reg[30][1]  ( .D(n56), .E(n186), .CP(n248), .Q(
        \Storage[30][1] ) );
  EDFQD1 \Storage_reg[30][0]  ( .D(n59), .E(n184), .CP(n248), .Q(
        \Storage[30][0] ) );
  EDFQD1 \Storage_reg[29][32]  ( .D(n200), .E(n177), .CP(n248), .Q(
        \Storage[29][32] ) );
  EDFQD1 \Storage_reg[29][31]  ( .D(n63), .E(n177), .CP(n247), .Q(
        \Storage[29][31] ) );
  EDFQD1 \Storage_reg[29][30]  ( .D(n61), .E(n178), .CP(n247), .Q(
        \Storage[29][30] ) );
  EDFQD1 \Storage_reg[29][29]  ( .D(n58), .E(n178), .CP(n247), .Q(
        \Storage[29][29] ) );
  EDFQD1 \Storage_reg[29][28]  ( .D(n53), .E(n177), .CP(n247), .Q(
        \Storage[29][28] ) );
  EDFQD1 \Storage_reg[29][27]  ( .D(n49), .E(n176), .CP(n247), .Q(
        \Storage[29][27] ) );
  EDFQD1 \Storage_reg[29][26]  ( .D(n45), .E(n176), .CP(n247), .Q(
        \Storage[29][26] ) );
  EDFQD1 \Storage_reg[29][25]  ( .D(n41), .E(n177), .CP(n247), .Q(
        \Storage[29][25] ) );
  EDFQD1 \Storage_reg[29][24]  ( .D(n37), .E(n176), .CP(n247), .Q(
        \Storage[29][24] ) );
  EDFQD1 \Storage_reg[29][23]  ( .D(n33), .E(n178), .CP(n247), .Q(
        \Storage[29][23] ) );
  EDFQD1 \Storage_reg[29][22]  ( .D(n29), .E(n177), .CP(n247), .Q(
        \Storage[29][22] ) );
  EDFQD1 \Storage_reg[29][21]  ( .D(n25), .E(n176), .CP(n247), .Q(
        \Storage[29][21] ) );
  EDFQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(n178), .CP(n246), .Q(
        \Storage[29][20] ) );
  EDFQD1 \Storage_reg[29][19]  ( .D(n17), .E(n176), .CP(n246), .Q(
        \Storage[29][19] ) );
  EDFQD1 \Storage_reg[29][18]  ( .D(n13), .E(n176), .CP(n246), .Q(
        \Storage[29][18] ) );
  EDFQD1 \Storage_reg[29][17]  ( .D(n10), .E(n177), .CP(n246), .Q(
        \Storage[29][17] ) );
  EDFQD1 \Storage_reg[29][16]  ( .D(n5), .E(n178), .CP(n246), .Q(
        \Storage[29][16] ) );
  EDFQD1 \Storage_reg[29][15]  ( .D(n2), .E(n178), .CP(n246), .Q(
        \Storage[29][15] ) );
  EDFQD1 \Storage_reg[29][14]  ( .D(n3), .E(n177), .CP(n246), .Q(
        \Storage[29][14] ) );
  EDFQD1 \Storage_reg[29][13]  ( .D(n7), .E(n176), .CP(n246), .Q(
        \Storage[29][13] ) );
  EDFQD1 \Storage_reg[29][12]  ( .D(n11), .E(n176), .CP(n246), .Q(
        \Storage[29][12] ) );
  EDFQD1 \Storage_reg[29][11]  ( .D(n15), .E(n177), .CP(n246), .Q(
        \Storage[29][11] ) );
  EDFQD1 \Storage_reg[29][10]  ( .D(n20), .E(n178), .CP(n246), .Q(
        \Storage[29][10] ) );
  EDFQD1 \Storage_reg[29][9]  ( .D(n23), .E(n178), .CP(n245), .Q(
        \Storage[29][9] ) );
  EDFQD1 \Storage_reg[29][8]  ( .D(n27), .E(n177), .CP(n245), .Q(
        \Storage[29][8] ) );
  EDFQD1 \Storage_reg[29][7]  ( .D(n32), .E(n176), .CP(n245), .Q(
        \Storage[29][7] ) );
  EDFQD1 \Storage_reg[29][6]  ( .D(n35), .E(n176), .CP(n245), .Q(
        \Storage[29][6] ) );
  EDFQD1 \Storage_reg[29][5]  ( .D(n39), .E(n177), .CP(n245), .Q(
        \Storage[29][5] ) );
  EDFQD1 \Storage_reg[29][4]  ( .D(n43), .E(n178), .CP(n245), .Q(
        \Storage[29][4] ) );
  EDFQD1 \Storage_reg[29][3]  ( .D(n48), .E(n178), .CP(n245), .Q(
        \Storage[29][3] ) );
  EDFQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(n177), .CP(n245), .Q(
        \Storage[29][2] ) );
  EDFQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(n178), .CP(n245), .Q(
        \Storage[29][1] ) );
  EDFQD1 \Storage_reg[29][0]  ( .D(n59), .E(n176), .CP(n245), .Q(
        \Storage[29][0] ) );
  EDFQD1 \Storage_reg[28][32]  ( .D(n201), .E(n169), .CP(n245), .Q(
        \Storage[28][32] ) );
  EDFQD1 \Storage_reg[28][31]  ( .D(n64), .E(n169), .CP(n244), .Q(
        \Storage[28][31] ) );
  EDFQD1 \Storage_reg[28][30]  ( .D(n62), .E(n170), .CP(n244), .Q(
        \Storage[28][30] ) );
  EDFQD1 \Storage_reg[28][29]  ( .D(n58), .E(n170), .CP(n244), .Q(
        \Storage[28][29] ) );
  EDFQD1 \Storage_reg[28][28]  ( .D(n54), .E(n169), .CP(n244), .Q(
        \Storage[28][28] ) );
  EDFQD1 \Storage_reg[28][27]  ( .D(n50), .E(n168), .CP(n244), .Q(
        \Storage[28][27] ) );
  EDFQD1 \Storage_reg[28][26]  ( .D(n46), .E(n168), .CP(n244), .Q(
        \Storage[28][26] ) );
  EDFQD1 \Storage_reg[28][25]  ( .D(n42), .E(n169), .CP(n244), .Q(
        \Storage[28][25] ) );
  EDFQD1 \Storage_reg[28][24]  ( .D(n38), .E(n168), .CP(n244), .Q(
        \Storage[28][24] ) );
  EDFQD1 \Storage_reg[28][23]  ( .D(n34), .E(n170), .CP(n244), .Q(
        \Storage[28][23] ) );
  EDFQD1 \Storage_reg[28][22]  ( .D(n30), .E(n169), .CP(n244), .Q(
        \Storage[28][22] ) );
  EDFQD1 \Storage_reg[28][21]  ( .D(n26), .E(n168), .CP(n244), .Q(
        \Storage[28][21] ) );
  EDFQD1 \Storage_reg[28][20]  ( .D(n22), .E(n170), .CP(n243), .Q(
        \Storage[28][20] ) );
  EDFQD1 \Storage_reg[28][19]  ( .D(n18), .E(n168), .CP(n243), .Q(
        \Storage[28][19] ) );
  EDFQD1 \Storage_reg[28][18]  ( .D(n14), .E(n168), .CP(n243), .Q(
        \Storage[28][18] ) );
  EDFQD1 \Storage_reg[28][17]  ( .D(n10), .E(n169), .CP(n243), .Q(
        \Storage[28][17] ) );
  EDFQD1 \Storage_reg[28][16]  ( .D(n6), .E(n170), .CP(n243), .Q(
        \Storage[28][16] ) );
  EDFQD1 \Storage_reg[28][15]  ( .D(n2), .E(n170), .CP(n243), .Q(
        \Storage[28][15] ) );
  EDFQD1 \Storage_reg[28][14]  ( .D(n4), .E(n169), .CP(n243), .Q(
        \Storage[28][14] ) );
  EDFQD1 \Storage_reg[28][13]  ( .D(n8), .E(n168), .CP(n243), .Q(
        \Storage[28][13] ) );
  EDFQD1 \Storage_reg[28][12]  ( .D(n12), .E(n168), .CP(n243), .Q(
        \Storage[28][12] ) );
  EDFQD1 \Storage_reg[28][11]  ( .D(n16), .E(n169), .CP(n243), .Q(
        \Storage[28][11] ) );
  EDFQD1 \Storage_reg[28][10]  ( .D(n20), .E(n170), .CP(n243), .Q(
        \Storage[28][10] ) );
  EDFQD1 \Storage_reg[28][9]  ( .D(n24), .E(n170), .CP(n242), .Q(
        \Storage[28][9] ) );
  EDFQD1 \Storage_reg[28][8]  ( .D(n28), .E(n169), .CP(n242), .Q(
        \Storage[28][8] ) );
  EDFQD1 \Storage_reg[28][7]  ( .D(n32), .E(n168), .CP(n242), .Q(
        \Storage[28][7] ) );
  EDFQD1 \Storage_reg[28][6]  ( .D(n36), .E(n168), .CP(n242), .Q(
        \Storage[28][6] ) );
  EDFQD1 \Storage_reg[28][5]  ( .D(n40), .E(n169), .CP(n242), .Q(
        \Storage[28][5] ) );
  EDFQD1 \Storage_reg[28][4]  ( .D(n44), .E(n170), .CP(n242), .Q(
        \Storage[28][4] ) );
  EDFQD1 \Storage_reg[28][3]  ( .D(n48), .E(n170), .CP(n242), .Q(
        \Storage[28][3] ) );
  EDFQD1 \Storage_reg[28][2]  ( .D(n51), .E(n169), .CP(n242), .Q(
        \Storage[28][2] ) );
  EDFQD1 \Storage_reg[28][1]  ( .D(n55), .E(n170), .CP(n242), .Q(
        \Storage[28][1] ) );
  EDFQD1 \Storage_reg[28][0]  ( .D(n60), .E(n168), .CP(n242), .Q(
        \Storage[28][0] ) );
  EDFQD1 \Storage_reg[27][32]  ( .D(n202), .E(n161), .CP(n242), .Q(
        \Storage[27][32] ) );
  EDFQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(n161), .CP(n241), .Q(
        \Storage[27][31] ) );
  EDFQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(n162), .CP(n241), .Q(
        \Storage[27][30] ) );
  EDFQD1 \Storage_reg[27][29]  ( .D(n57), .E(n162), .CP(n241), .Q(
        \Storage[27][29] ) );
  EDFQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(n161), .CP(n241), .Q(
        \Storage[27][28] ) );
  EDFQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(n160), .CP(n241), .Q(
        \Storage[27][27] ) );
  EDFQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(n160), .CP(n241), .Q(
        \Storage[27][26] ) );
  EDFQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(n161), .CP(n241), .Q(
        \Storage[27][25] ) );
  EDFQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(n160), .CP(n241), .Q(
        \Storage[27][24] ) );
  EDFQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(n162), .CP(n241), .Q(
        \Storage[27][23] ) );
  EDFQD1 \Storage_reg[27][22]  ( .D(DataI[22]), .E(n161), .CP(n241), .Q(
        \Storage[27][22] ) );
  EDFQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(n160), .CP(n241), .Q(
        \Storage[27][21] ) );
  EDFQD1 \Storage_reg[27][20]  ( .D(n21), .E(n162), .CP(n240), .Q(
        \Storage[27][20] ) );
  EDFQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(n160), .CP(n240), .Q(
        \Storage[27][19] ) );
  EDFQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(n160), .CP(n240), .Q(
        \Storage[27][18] ) );
  EDFQD1 \Storage_reg[27][17]  ( .D(n9), .E(n161), .CP(n240), .Q(
        \Storage[27][17] ) );
  EDFQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(n162), .CP(n240), .Q(
        \Storage[27][16] ) );
  EDFQD1 \Storage_reg[27][15]  ( .D(n1), .E(n162), .CP(n240), .Q(
        \Storage[27][15] ) );
  EDFQD1 \Storage_reg[27][14]  ( .D(DataI[14]), .E(n161), .CP(n240), .Q(
        \Storage[27][14] ) );
  EDFQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(n160), .CP(n240), .Q(
        \Storage[27][13] ) );
  EDFQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(n160), .CP(n240), .Q(
        \Storage[27][12] ) );
  EDFQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(n161), .CP(n240), .Q(
        \Storage[27][11] ) );
  EDFQD1 \Storage_reg[27][10]  ( .D(n19), .E(n162), .CP(n240), .Q(
        \Storage[27][10] ) );
  EDFQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(n162), .CP(n239), .Q(
        \Storage[27][9] ) );
  EDFQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(n161), .CP(n239), .Q(
        \Storage[27][8] ) );
  EDFQD1 \Storage_reg[27][7]  ( .D(n31), .E(n160), .CP(n239), .Q(
        \Storage[27][7] ) );
  EDFQD1 \Storage_reg[27][6]  ( .D(DataI[6]), .E(n160), .CP(n239), .Q(
        \Storage[27][6] ) );
  EDFQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(n161), .CP(n239), .Q(
        \Storage[27][5] ) );
  EDFQD1 \Storage_reg[27][4]  ( .D(DataI[4]), .E(n162), .CP(n239), .Q(
        \Storage[27][4] ) );
  EDFQD1 \Storage_reg[27][3]  ( .D(n47), .E(n162), .CP(n239), .Q(
        \Storage[27][3] ) );
  EDFQD1 \Storage_reg[27][2]  ( .D(n52), .E(n161), .CP(n239), .Q(
        \Storage[27][2] ) );
  EDFQD1 \Storage_reg[27][1]  ( .D(n56), .E(n162), .CP(n239), .Q(
        \Storage[27][1] ) );
  EDFQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(n160), .CP(n239), .Q(
        \Storage[27][0] ) );
  EDFQD1 \Storage_reg[25][32]  ( .D(n201), .E(n145), .CP(n236), .Q(
        \Storage[25][32] ) );
  EDFQD1 \Storage_reg[25][31]  ( .D(n63), .E(n145), .CP(n235), .Q(
        \Storage[25][31] ) );
  EDFQD1 \Storage_reg[25][30]  ( .D(n61), .E(n146), .CP(n235), .Q(
        \Storage[25][30] ) );
  EDFQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(n146), .CP(n235), .Q(
        \Storage[25][29] ) );
  EDFQD1 \Storage_reg[25][28]  ( .D(n53), .E(n145), .CP(n235), .Q(
        \Storage[25][28] ) );
  EDFQD1 \Storage_reg[25][27]  ( .D(n49), .E(n144), .CP(n235), .Q(
        \Storage[25][27] ) );
  EDFQD1 \Storage_reg[25][26]  ( .D(n45), .E(n144), .CP(n235), .Q(
        \Storage[25][26] ) );
  EDFQD1 \Storage_reg[25][25]  ( .D(n41), .E(n145), .CP(n235), .Q(
        \Storage[25][25] ) );
  EDFQD1 \Storage_reg[25][24]  ( .D(n37), .E(n144), .CP(n235), .Q(
        \Storage[25][24] ) );
  EDFQD1 \Storage_reg[25][23]  ( .D(n33), .E(n146), .CP(n235), .Q(
        \Storage[25][23] ) );
  EDFQD1 \Storage_reg[25][22]  ( .D(n29), .E(n145), .CP(n235), .Q(
        \Storage[25][22] ) );
  EDFQD1 \Storage_reg[25][21]  ( .D(n25), .E(n144), .CP(n235), .Q(
        \Storage[25][21] ) );
  EDFQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(n146), .CP(n234), .Q(
        \Storage[25][20] ) );
  EDFQD1 \Storage_reg[25][19]  ( .D(n17), .E(n144), .CP(n234), .Q(
        \Storage[25][19] ) );
  EDFQD1 \Storage_reg[25][18]  ( .D(n13), .E(n144), .CP(n234), .Q(
        \Storage[25][18] ) );
  EDFQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(n145), .CP(n234), .Q(
        \Storage[25][17] ) );
  EDFQD1 \Storage_reg[25][16]  ( .D(n5), .E(n146), .CP(n234), .Q(
        \Storage[25][16] ) );
  EDFQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(n146), .CP(n234), .Q(
        \Storage[25][15] ) );
  EDFQD1 \Storage_reg[25][14]  ( .D(n3), .E(n145), .CP(n234), .Q(
        \Storage[25][14] ) );
  EDFQD1 \Storage_reg[25][13]  ( .D(n7), .E(n144), .CP(n234), .Q(
        \Storage[25][13] ) );
  EDFQD1 \Storage_reg[25][12]  ( .D(n11), .E(n144), .CP(n234), .Q(
        \Storage[25][12] ) );
  EDFQD1 \Storage_reg[25][11]  ( .D(n15), .E(n145), .CP(n234), .Q(
        \Storage[25][11] ) );
  EDFQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(n146), .CP(n234), .Q(
        \Storage[25][10] ) );
  EDFQD1 \Storage_reg[25][9]  ( .D(n23), .E(n146), .CP(n233), .Q(
        \Storage[25][9] ) );
  EDFQD1 \Storage_reg[25][8]  ( .D(n27), .E(n145), .CP(n233), .Q(
        \Storage[25][8] ) );
  EDFQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(n144), .CP(n233), .Q(
        \Storage[25][7] ) );
  EDFQD1 \Storage_reg[25][6]  ( .D(n35), .E(n144), .CP(n233), .Q(
        \Storage[25][6] ) );
  EDFQD1 \Storage_reg[25][5]  ( .D(n39), .E(n145), .CP(n233), .Q(
        \Storage[25][5] ) );
  EDFQD1 \Storage_reg[25][4]  ( .D(n43), .E(n146), .CP(n233), .Q(
        \Storage[25][4] ) );
  EDFQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(n146), .CP(n233), .Q(
        \Storage[25][3] ) );
  EDFQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(n145), .CP(n233), .Q(
        \Storage[25][2] ) );
  EDFQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(n146), .CP(n233), .Q(
        \Storage[25][1] ) );
  EDFQD1 \Storage_reg[25][0]  ( .D(n59), .E(n144), .CP(n233), .Q(
        \Storage[25][0] ) );
  EDFQD1 \Storage_reg[22][32]  ( .D(n200), .E(n121), .CP(n227), .Q(
        \Storage[22][32] ) );
  EDFQD1 \Storage_reg[22][31]  ( .D(n64), .E(n121), .CP(n226), .Q(
        \Storage[22][31] ) );
  EDFQD1 \Storage_reg[22][30]  ( .D(n62), .E(n122), .CP(n226), .Q(
        \Storage[22][30] ) );
  EDFQD1 \Storage_reg[22][29]  ( .D(n58), .E(n122), .CP(n226), .Q(
        \Storage[22][29] ) );
  EDFQD1 \Storage_reg[22][28]  ( .D(n54), .E(n121), .CP(n226), .Q(
        \Storage[22][28] ) );
  EDFQD1 \Storage_reg[22][27]  ( .D(n50), .E(n120), .CP(n226), .Q(
        \Storage[22][27] ) );
  EDFQD1 \Storage_reg[22][26]  ( .D(n46), .E(n120), .CP(n226), .Q(
        \Storage[22][26] ) );
  EDFQD1 \Storage_reg[22][25]  ( .D(n42), .E(n121), .CP(n226), .Q(
        \Storage[22][25] ) );
  EDFQD1 \Storage_reg[22][24]  ( .D(n38), .E(n120), .CP(n226), .Q(
        \Storage[22][24] ) );
  EDFQD1 \Storage_reg[22][23]  ( .D(n34), .E(n122), .CP(n226), .Q(
        \Storage[22][23] ) );
  EDFQD1 \Storage_reg[22][22]  ( .D(n30), .E(n121), .CP(n226), .Q(
        \Storage[22][22] ) );
  EDFQD1 \Storage_reg[22][21]  ( .D(n26), .E(n120), .CP(n226), .Q(
        \Storage[22][21] ) );
  EDFQD1 \Storage_reg[22][20]  ( .D(n22), .E(n122), .CP(n225), .Q(
        \Storage[22][20] ) );
  EDFQD1 \Storage_reg[22][19]  ( .D(n18), .E(n120), .CP(n225), .Q(
        \Storage[22][19] ) );
  EDFQD1 \Storage_reg[22][18]  ( .D(n14), .E(n120), .CP(n225), .Q(
        \Storage[22][18] ) );
  EDFQD1 \Storage_reg[22][17]  ( .D(n10), .E(n121), .CP(n225), .Q(
        \Storage[22][17] ) );
  EDFQD1 \Storage_reg[22][16]  ( .D(n6), .E(n122), .CP(n225), .Q(
        \Storage[22][16] ) );
  EDFQD1 \Storage_reg[22][15]  ( .D(n2), .E(n122), .CP(n225), .Q(
        \Storage[22][15] ) );
  EDFQD1 \Storage_reg[22][14]  ( .D(n4), .E(n121), .CP(n225), .Q(
        \Storage[22][14] ) );
  EDFQD1 \Storage_reg[22][13]  ( .D(n8), .E(n120), .CP(n225), .Q(
        \Storage[22][13] ) );
  EDFQD1 \Storage_reg[22][12]  ( .D(n12), .E(n120), .CP(n225), .Q(
        \Storage[22][12] ) );
  EDFQD1 \Storage_reg[22][11]  ( .D(n16), .E(n121), .CP(n225), .Q(
        \Storage[22][11] ) );
  EDFQD1 \Storage_reg[22][10]  ( .D(n20), .E(n122), .CP(n225), .Q(
        \Storage[22][10] ) );
  EDFQD1 \Storage_reg[22][9]  ( .D(n24), .E(n122), .CP(n224), .Q(
        \Storage[22][9] ) );
  EDFQD1 \Storage_reg[22][8]  ( .D(n28), .E(n121), .CP(n224), .Q(
        \Storage[22][8] ) );
  EDFQD1 \Storage_reg[22][7]  ( .D(n32), .E(n120), .CP(n224), .Q(
        \Storage[22][7] ) );
  EDFQD1 \Storage_reg[22][6]  ( .D(n36), .E(n120), .CP(n224), .Q(
        \Storage[22][6] ) );
  EDFQD1 \Storage_reg[22][5]  ( .D(n40), .E(n121), .CP(n224), .Q(
        \Storage[22][5] ) );
  EDFQD1 \Storage_reg[22][4]  ( .D(n44), .E(n122), .CP(n224), .Q(
        \Storage[22][4] ) );
  EDFQD1 \Storage_reg[22][3]  ( .D(n48), .E(n122), .CP(n224), .Q(
        \Storage[22][3] ) );
  EDFQD1 \Storage_reg[22][2]  ( .D(n51), .E(n121), .CP(n224), .Q(
        \Storage[22][2] ) );
  EDFQD1 \Storage_reg[22][1]  ( .D(n55), .E(n122), .CP(n224), .Q(
        \Storage[22][1] ) );
  EDFQD1 \Storage_reg[22][0]  ( .D(n60), .E(n120), .CP(n224), .Q(
        \Storage[22][0] ) );
  EDFQD1 \Storage_reg[21][32]  ( .D(n201), .E(n113), .CP(n224), .Q(
        \Storage[21][32] ) );
  EDFQD1 \Storage_reg[21][31]  ( .D(DataI[31]), .E(n113), .CP(n223), .Q(
        \Storage[21][31] ) );
  EDFQD1 \Storage_reg[21][30]  ( .D(DataI[30]), .E(n114), .CP(n223), .Q(
        \Storage[21][30] ) );
  EDFQD1 \Storage_reg[21][29]  ( .D(n57), .E(n114), .CP(n223), .Q(
        \Storage[21][29] ) );
  EDFQD1 \Storage_reg[21][28]  ( .D(DataI[28]), .E(n113), .CP(n223), .Q(
        \Storage[21][28] ) );
  EDFQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(n112), .CP(n223), .Q(
        \Storage[21][27] ) );
  EDFQD1 \Storage_reg[21][26]  ( .D(DataI[26]), .E(n112), .CP(n223), .Q(
        \Storage[21][26] ) );
  EDFQD1 \Storage_reg[21][25]  ( .D(DataI[25]), .E(n113), .CP(n223), .Q(
        \Storage[21][25] ) );
  EDFQD1 \Storage_reg[21][24]  ( .D(DataI[24]), .E(n112), .CP(n223), .Q(
        \Storage[21][24] ) );
  EDFQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(n114), .CP(n223), .Q(
        \Storage[21][23] ) );
  EDFQD1 \Storage_reg[21][22]  ( .D(DataI[22]), .E(n113), .CP(n223), .Q(
        \Storage[21][22] ) );
  EDFQD1 \Storage_reg[21][21]  ( .D(DataI[21]), .E(n112), .CP(n223), .Q(
        \Storage[21][21] ) );
  EDFQD1 \Storage_reg[21][20]  ( .D(n21), .E(n114), .CP(n222), .Q(
        \Storage[21][20] ) );
  EDFQD1 \Storage_reg[21][19]  ( .D(DataI[19]), .E(n112), .CP(n222), .Q(
        \Storage[21][19] ) );
  EDFQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(n112), .CP(n222), .Q(
        \Storage[21][18] ) );
  EDFQD1 \Storage_reg[21][17]  ( .D(n9), .E(n113), .CP(n222), .Q(
        \Storage[21][17] ) );
  EDFQD1 \Storage_reg[21][16]  ( .D(DataI[16]), .E(n114), .CP(n222), .Q(
        \Storage[21][16] ) );
  EDFQD1 \Storage_reg[21][15]  ( .D(n1), .E(n114), .CP(n222), .Q(
        \Storage[21][15] ) );
  EDFQD1 \Storage_reg[21][14]  ( .D(DataI[14]), .E(n113), .CP(n222), .Q(
        \Storage[21][14] ) );
  EDFQD1 \Storage_reg[21][13]  ( .D(DataI[13]), .E(n112), .CP(n222), .Q(
        \Storage[21][13] ) );
  EDFQD1 \Storage_reg[21][12]  ( .D(DataI[12]), .E(n112), .CP(n222), .Q(
        \Storage[21][12] ) );
  EDFQD1 \Storage_reg[21][11]  ( .D(DataI[11]), .E(n113), .CP(n222), .Q(
        \Storage[21][11] ) );
  EDFQD1 \Storage_reg[21][10]  ( .D(n19), .E(n114), .CP(n222), .Q(
        \Storage[21][10] ) );
  EDFQD1 \Storage_reg[21][9]  ( .D(DataI[9]), .E(n114), .CP(n221), .Q(
        \Storage[21][9] ) );
  EDFQD1 \Storage_reg[21][8]  ( .D(DataI[8]), .E(n113), .CP(n221), .Q(
        \Storage[21][8] ) );
  EDFQD1 \Storage_reg[21][7]  ( .D(n31), .E(n112), .CP(n221), .Q(
        \Storage[21][7] ) );
  EDFQD1 \Storage_reg[21][6]  ( .D(DataI[6]), .E(n112), .CP(n221), .Q(
        \Storage[21][6] ) );
  EDFQD1 \Storage_reg[21][5]  ( .D(DataI[5]), .E(n113), .CP(n221), .Q(
        \Storage[21][5] ) );
  EDFQD1 \Storage_reg[21][4]  ( .D(DataI[4]), .E(n114), .CP(n221), .Q(
        \Storage[21][4] ) );
  EDFQD1 \Storage_reg[21][3]  ( .D(n47), .E(n114), .CP(n221), .Q(
        \Storage[21][3] ) );
  EDFQD1 \Storage_reg[21][2]  ( .D(n52), .E(n113), .CP(n221), .Q(
        \Storage[21][2] ) );
  EDFQD1 \Storage_reg[21][1]  ( .D(n56), .E(n114), .CP(n221), .Q(
        \Storage[21][1] ) );
  EDFQD1 \Storage_reg[21][0]  ( .D(DataI[0]), .E(n112), .CP(n221), .Q(
        \Storage[21][0] ) );
  EDFQD1 \Storage_reg[18][32]  ( .D(n202), .E(n89), .CP(n215), .Q(
        \Storage[18][32] ) );
  EDFQD1 \Storage_reg[18][31]  ( .D(n63), .E(n89), .CP(n214), .Q(
        \Storage[18][31] ) );
  EDFQD1 \Storage_reg[18][30]  ( .D(n61), .E(n90), .CP(n214), .Q(
        \Storage[18][30] ) );
  EDFQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(n90), .CP(n214), .Q(
        \Storage[18][29] ) );
  EDFQD1 \Storage_reg[18][28]  ( .D(n53), .E(n89), .CP(n214), .Q(
        \Storage[18][28] ) );
  EDFQD1 \Storage_reg[18][27]  ( .D(n49), .E(n88), .CP(n214), .Q(
        \Storage[18][27] ) );
  EDFQD1 \Storage_reg[18][26]  ( .D(n45), .E(n88), .CP(n214), .Q(
        \Storage[18][26] ) );
  EDFQD1 \Storage_reg[18][25]  ( .D(n41), .E(n89), .CP(n214), .Q(
        \Storage[18][25] ) );
  EDFQD1 \Storage_reg[18][24]  ( .D(n37), .E(n88), .CP(n214), .Q(
        \Storage[18][24] ) );
  EDFQD1 \Storage_reg[18][23]  ( .D(n33), .E(n90), .CP(n214), .Q(
        \Storage[18][23] ) );
  EDFQD1 \Storage_reg[18][22]  ( .D(n29), .E(n89), .CP(n214), .Q(
        \Storage[18][22] ) );
  EDFQD1 \Storage_reg[18][21]  ( .D(n25), .E(n88), .CP(n214), .Q(
        \Storage[18][21] ) );
  EDFQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(n90), .CP(n213), .Q(
        \Storage[18][20] ) );
  EDFQD1 \Storage_reg[18][19]  ( .D(n17), .E(n88), .CP(n213), .Q(
        \Storage[18][19] ) );
  EDFQD1 \Storage_reg[18][18]  ( .D(n13), .E(n88), .CP(n213), .Q(
        \Storage[18][18] ) );
  EDFQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(n89), .CP(n213), .Q(
        \Storage[18][17] ) );
  EDFQD1 \Storage_reg[18][16]  ( .D(n5), .E(n90), .CP(n213), .Q(
        \Storage[18][16] ) );
  EDFQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(n90), .CP(n213), .Q(
        \Storage[18][15] ) );
  EDFQD1 \Storage_reg[18][14]  ( .D(n3), .E(n89), .CP(n213), .Q(
        \Storage[18][14] ) );
  EDFQD1 \Storage_reg[18][13]  ( .D(n7), .E(n88), .CP(n213), .Q(
        \Storage[18][13] ) );
  EDFQD1 \Storage_reg[18][12]  ( .D(n11), .E(n88), .CP(n213), .Q(
        \Storage[18][12] ) );
  EDFQD1 \Storage_reg[18][11]  ( .D(n15), .E(n89), .CP(n213), .Q(
        \Storage[18][11] ) );
  EDFQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(n90), .CP(n213), .Q(
        \Storage[18][10] ) );
  EDFQD1 \Storage_reg[18][9]  ( .D(n23), .E(n90), .CP(n212), .Q(
        \Storage[18][9] ) );
  EDFQD1 \Storage_reg[18][8]  ( .D(n27), .E(n89), .CP(n212), .Q(
        \Storage[18][8] ) );
  EDFQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(n88), .CP(n212), .Q(
        \Storage[18][7] ) );
  EDFQD1 \Storage_reg[18][6]  ( .D(n35), .E(n88), .CP(n212), .Q(
        \Storage[18][6] ) );
  EDFQD1 \Storage_reg[18][5]  ( .D(n39), .E(n89), .CP(n212), .Q(
        \Storage[18][5] ) );
  EDFQD1 \Storage_reg[18][4]  ( .D(n43), .E(n90), .CP(n212), .Q(
        \Storage[18][4] ) );
  EDFQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(n90), .CP(n212), .Q(
        \Storage[18][3] ) );
  EDFQD1 \Storage_reg[18][2]  ( .D(DataI[2]), .E(n89), .CP(n212), .Q(
        \Storage[18][2] ) );
  EDFQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(n90), .CP(n212), .Q(
        \Storage[18][1] ) );
  EDFQD1 \Storage_reg[18][0]  ( .D(n59), .E(n88), .CP(n212), .Q(
        \Storage[18][0] ) );
  EDFQD1 \Storage_reg[17][32]  ( .D(n200), .E(n81), .CP(n212), .Q(
        \Storage[17][32] ) );
  EDFQD1 \Storage_reg[17][31]  ( .D(n64), .E(n81), .CP(n211), .Q(
        \Storage[17][31] ) );
  EDFQD1 \Storage_reg[17][30]  ( .D(n62), .E(n82), .CP(n211), .Q(
        \Storage[17][30] ) );
  EDFQD1 \Storage_reg[17][29]  ( .D(n58), .E(n82), .CP(n211), .Q(
        \Storage[17][29] ) );
  EDFQD1 \Storage_reg[17][28]  ( .D(n54), .E(n81), .CP(n211), .Q(
        \Storage[17][28] ) );
  EDFQD1 \Storage_reg[17][27]  ( .D(n50), .E(n80), .CP(n211), .Q(
        \Storage[17][27] ) );
  EDFQD1 \Storage_reg[17][26]  ( .D(n46), .E(n80), .CP(n211), .Q(
        \Storage[17][26] ) );
  EDFQD1 \Storage_reg[17][25]  ( .D(n42), .E(n81), .CP(n211), .Q(
        \Storage[17][25] ) );
  EDFQD1 \Storage_reg[17][24]  ( .D(n38), .E(n80), .CP(n211), .Q(
        \Storage[17][24] ) );
  EDFQD1 \Storage_reg[17][23]  ( .D(n34), .E(n82), .CP(n211), .Q(
        \Storage[17][23] ) );
  EDFQD1 \Storage_reg[17][22]  ( .D(n30), .E(n81), .CP(n211), .Q(
        \Storage[17][22] ) );
  EDFQD1 \Storage_reg[17][21]  ( .D(n26), .E(n80), .CP(n211), .Q(
        \Storage[17][21] ) );
  EDFQD1 \Storage_reg[17][20]  ( .D(n22), .E(n82), .CP(n210), .Q(
        \Storage[17][20] ) );
  EDFQD1 \Storage_reg[17][19]  ( .D(n18), .E(n80), .CP(n210), .Q(
        \Storage[17][19] ) );
  EDFQD1 \Storage_reg[17][18]  ( .D(n14), .E(n80), .CP(n210), .Q(
        \Storage[17][18] ) );
  EDFQD1 \Storage_reg[17][17]  ( .D(n10), .E(n81), .CP(n210), .Q(
        \Storage[17][17] ) );
  EDFQD1 \Storage_reg[17][16]  ( .D(n6), .E(n82), .CP(n210), .Q(
        \Storage[17][16] ) );
  EDFQD1 \Storage_reg[17][15]  ( .D(n2), .E(n82), .CP(n210), .Q(
        \Storage[17][15] ) );
  EDFQD1 \Storage_reg[17][14]  ( .D(n4), .E(n81), .CP(n210), .Q(
        \Storage[17][14] ) );
  EDFQD1 \Storage_reg[17][13]  ( .D(n8), .E(n80), .CP(n210), .Q(
        \Storage[17][13] ) );
  EDFQD1 \Storage_reg[17][12]  ( .D(n12), .E(n80), .CP(n210), .Q(
        \Storage[17][12] ) );
  EDFQD1 \Storage_reg[17][11]  ( .D(n16), .E(n81), .CP(n210), .Q(
        \Storage[17][11] ) );
  EDFQD1 \Storage_reg[17][10]  ( .D(n20), .E(n82), .CP(n210), .Q(
        \Storage[17][10] ) );
  EDFQD1 \Storage_reg[17][9]  ( .D(n24), .E(n82), .CP(n209), .Q(
        \Storage[17][9] ) );
  EDFQD1 \Storage_reg[17][8]  ( .D(n28), .E(n81), .CP(n209), .Q(
        \Storage[17][8] ) );
  EDFQD1 \Storage_reg[17][7]  ( .D(n32), .E(n80), .CP(n209), .Q(
        \Storage[17][7] ) );
  EDFQD1 \Storage_reg[17][6]  ( .D(n36), .E(n80), .CP(n209), .Q(
        \Storage[17][6] ) );
  EDFQD1 \Storage_reg[17][5]  ( .D(n40), .E(n81), .CP(n209), .Q(
        \Storage[17][5] ) );
  EDFQD1 \Storage_reg[17][4]  ( .D(n44), .E(n82), .CP(n209), .Q(
        \Storage[17][4] ) );
  EDFQD1 \Storage_reg[17][3]  ( .D(n48), .E(n82), .CP(n209), .Q(
        \Storage[17][3] ) );
  EDFQD1 \Storage_reg[17][2]  ( .D(n51), .E(n81), .CP(n209), .Q(
        \Storage[17][2] ) );
  EDFQD1 \Storage_reg[17][1]  ( .D(n55), .E(n82), .CP(n209), .Q(
        \Storage[17][1] ) );
  EDFQD1 \Storage_reg[17][0]  ( .D(n60), .E(n80), .CP(n209), .Q(
        \Storage[17][0] ) );
  EDFQD1 \Storage_reg[14][32]  ( .D(n200), .E(n85), .CP(n205), .Q(
        \Storage[14][32] ) );
  EDFQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(n85), .CP(n204), .Q(
        \Storage[14][31] ) );
  EDFQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(n86), .CP(n204), .Q(
        \Storage[14][30] ) );
  EDFQD1 \Storage_reg[14][29]  ( .D(n57), .E(n86), .CP(n204), .Q(
        \Storage[14][29] ) );
  EDFQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n85), .CP(n204), .Q(
        \Storage[14][28] ) );
  EDFQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n84), .CP(n204), .Q(
        \Storage[14][27] ) );
  EDFQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n84), .CP(n204), .Q(
        \Storage[14][26] ) );
  EDFQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(n85), .CP(n204), .Q(
        \Storage[14][25] ) );
  EDFQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n84), .CP(n204), .Q(
        \Storage[14][24] ) );
  EDFQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n86), .CP(n204), .Q(
        \Storage[14][23] ) );
  EDFQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(n85), .CP(n204), .Q(
        \Storage[14][22] ) );
  EDFQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n84), .CP(n204), .Q(
        \Storage[14][21] ) );
  EDFQD1 \Storage_reg[14][20]  ( .D(n21), .E(n86), .CP(n203), .Q(
        \Storage[14][20] ) );
  EDFQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n84), .CP(n203), .Q(
        \Storage[14][19] ) );
  EDFQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(n84), .CP(n203), .Q(
        \Storage[14][18] ) );
  EDFQD1 \Storage_reg[14][17]  ( .D(n9), .E(n85), .CP(n203), .Q(
        \Storage[14][17] ) );
  EDFQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(n86), .CP(n203), .Q(
        \Storage[14][16] ) );
  EDFQD1 \Storage_reg[14][15]  ( .D(n1), .E(n86), .CP(n203), .Q(
        \Storage[14][15] ) );
  EDFQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(n85), .CP(n203), .Q(
        \Storage[14][14] ) );
  EDFQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(n84), .CP(n203), .Q(
        \Storage[14][13] ) );
  EDFQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(n84), .CP(n203), .Q(
        \Storage[14][12] ) );
  EDFQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n85), .CP(n203), .Q(
        \Storage[14][11] ) );
  EDFQD1 \Storage_reg[14][10]  ( .D(n19), .E(n86), .CP(n203), .Q(
        \Storage[14][10] ) );
  EDFQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(n86), .CP(n240), .Q(
        \Storage[14][9] ) );
  EDFQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n85), .CP(n266), .Q(
        \Storage[14][8] ) );
  EDFQD1 \Storage_reg[14][7]  ( .D(n31), .E(n84), .CP(n251), .Q(
        \Storage[14][7] ) );
  EDFQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(n84), .CP(n250), .Q(
        \Storage[14][6] ) );
  EDFQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(n85), .CP(n249), .Q(
        \Storage[14][5] ) );
  EDFQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(n86), .CP(n248), .Q(
        \Storage[14][4] ) );
  EDFQD1 \Storage_reg[14][3]  ( .D(n47), .E(n86), .CP(n247), .Q(
        \Storage[14][3] ) );
  EDFQD1 \Storage_reg[14][2]  ( .D(n52), .E(n85), .CP(n246), .Q(
        \Storage[14][2] ) );
  EDFQD1 \Storage_reg[14][1]  ( .D(n56), .E(n86), .CP(n245), .Q(
        \Storage[14][1] ) );
  EDFQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(n84), .CP(n244), .Q(
        \Storage[14][0] ) );
  EDFQD1 \Storage_reg[13][32]  ( .D(n201), .E(n93), .CP(n243), .Q(
        \Storage[13][32] ) );
  EDFQD1 \Storage_reg[13][31]  ( .D(n63), .E(n93), .CP(n203), .Q(
        \Storage[13][31] ) );
  EDFQD1 \Storage_reg[13][30]  ( .D(n61), .E(n94), .CP(n265), .Q(
        \Storage[13][30] ) );
  EDFQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n94), .CP(n241), .Q(
        \Storage[13][29] ) );
  EDFQD1 \Storage_reg[13][28]  ( .D(n53), .E(n93), .CP(n242), .Q(
        \Storage[13][28] ) );
  EDFQD1 \Storage_reg[13][27]  ( .D(n49), .E(n92), .CP(n239), .Q(
        \Storage[13][27] ) );
  EDFQD1 \Storage_reg[13][26]  ( .D(n45), .E(n92), .CP(n238), .Q(
        \Storage[13][26] ) );
  EDFQD1 \Storage_reg[13][25]  ( .D(n41), .E(n93), .CP(n237), .Q(
        \Storage[13][25] ) );
  EDFQD1 \Storage_reg[13][24]  ( .D(n37), .E(n92), .CP(n236), .Q(
        \Storage[13][24] ) );
  EDFQD1 \Storage_reg[13][23]  ( .D(n33), .E(n94), .CP(n235), .Q(
        \Storage[13][23] ) );
  EDFQD1 \Storage_reg[13][22]  ( .D(n29), .E(n93), .CP(n234), .Q(
        \Storage[13][22] ) );
  EDFQD1 \Storage_reg[13][21]  ( .D(n25), .E(n92), .CP(n206), .Q(
        \Storage[13][21] ) );
  EDFQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n94), .CP(n264), .Q(
        \Storage[13][20] ) );
  EDFQD1 \Storage_reg[13][19]  ( .D(n17), .E(n92), .CP(n204), .Q(
        \Storage[13][19] ) );
  EDFQD1 \Storage_reg[13][18]  ( .D(n13), .E(n92), .CP(n205), .Q(
        \Storage[13][18] ) );
  EDFQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n93), .CP(n270), .Q(
        \Storage[13][17] ) );
  EDFQD1 \Storage_reg[13][16]  ( .D(n5), .E(n94), .CP(n275), .Q(
        \Storage[13][16] ) );
  EDFQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n94), .CP(n275), .Q(
        \Storage[13][15] ) );
  EDFQD1 \Storage_reg[13][14]  ( .D(n3), .E(n93), .CP(n278), .Q(
        \Storage[13][14] ) );
  EDFQD1 \Storage_reg[13][13]  ( .D(n7), .E(n92), .CP(n279), .Q(
        \Storage[13][13] ) );
  EDFQD1 \Storage_reg[13][12]  ( .D(n11), .E(n92), .CP(n272), .Q(
        \Storage[13][12] ) );
  EDFQD1 \Storage_reg[13][11]  ( .D(n15), .E(n93), .CP(n267), .Q(
        \Storage[13][11] ) );
  EDFQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n94), .CP(n268), .Q(
        \Storage[13][10] ) );
  EDFQD1 \Storage_reg[13][9]  ( .D(n23), .E(n94), .CP(n259), .Q(
        \Storage[13][9] ) );
  EDFQD1 \Storage_reg[13][8]  ( .D(n27), .E(n93), .CP(n218), .Q(
        \Storage[13][8] ) );
  EDFQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(n92), .CP(n258), .Q(
        \Storage[13][7] ) );
  EDFQD1 \Storage_reg[13][6]  ( .D(n35), .E(n92), .CP(n278), .Q(
        \Storage[13][6] ) );
  EDFQD1 \Storage_reg[13][5]  ( .D(n39), .E(n93), .CP(n274), .Q(
        \Storage[13][5] ) );
  EDFQD1 \Storage_reg[13][4]  ( .D(n43), .E(n94), .CP(n263), .Q(
        \Storage[13][4] ) );
  EDFQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(n94), .CP(n267), .Q(
        \Storage[13][3] ) );
  EDFQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(n93), .CP(n268), .Q(
        \Storage[13][2] ) );
  EDFQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n94), .CP(n269), .Q(
        \Storage[13][1] ) );
  EDFQD1 \Storage_reg[13][0]  ( .D(n59), .E(n92), .CP(n276), .Q(
        \Storage[13][0] ) );
  EDFQD1 \Storage_reg[10][32]  ( .D(n200), .E(n117), .CP(n232), .Q(
        \Storage[10][32] ) );
  EDFQD1 \Storage_reg[10][31]  ( .D(n64), .E(n117), .CP(n212), .Q(
        \Storage[10][31] ) );
  EDFQD1 \Storage_reg[10][30]  ( .D(n62), .E(n118), .CP(n206), .Q(
        \Storage[10][30] ) );
  EDFQD1 \Storage_reg[10][29]  ( .D(n58), .E(n118), .CP(n231), .Q(
        \Storage[10][29] ) );
  EDFQD1 \Storage_reg[10][28]  ( .D(n54), .E(n117), .CP(n230), .Q(
        \Storage[10][28] ) );
  EDFQD1 \Storage_reg[10][27]  ( .D(n50), .E(n116), .CP(n229), .Q(
        \Storage[10][27] ) );
  EDFQD1 \Storage_reg[10][26]  ( .D(n46), .E(n116), .CP(n228), .Q(
        \Storage[10][26] ) );
  EDFQD1 \Storage_reg[10][25]  ( .D(n42), .E(n117), .CP(n227), .Q(
        \Storage[10][25] ) );
  EDFQD1 \Storage_reg[10][24]  ( .D(n38), .E(n116), .CP(n226), .Q(
        \Storage[10][24] ) );
  EDFQD1 \Storage_reg[10][23]  ( .D(n34), .E(n118), .CP(n225), .Q(
        \Storage[10][23] ) );
  EDFQD1 \Storage_reg[10][22]  ( .D(n30), .E(n117), .CP(n209), .Q(
        \Storage[10][22] ) );
  EDFQD1 \Storage_reg[10][21]  ( .D(n26), .E(n116), .CP(n208), .Q(
        \Storage[10][21] ) );
  EDFQD1 \Storage_reg[10][20]  ( .D(n22), .E(n118), .CP(n246), .Q(
        \Storage[10][20] ) );
  EDFQD1 \Storage_reg[10][19]  ( .D(n18), .E(n116), .CP(n211), .Q(
        \Storage[10][19] ) );
  EDFQD1 \Storage_reg[10][18]  ( .D(n14), .E(n116), .CP(n210), .Q(
        \Storage[10][18] ) );
  EDFQD1 \Storage_reg[10][17]  ( .D(n10), .E(n117), .CP(n213), .Q(
        \Storage[10][17] ) );
  EDFQD1 \Storage_reg[10][16]  ( .D(n6), .E(n118), .CP(n214), .Q(
        \Storage[10][16] ) );
  EDFQD1 \Storage_reg[10][15]  ( .D(n2), .E(n118), .CP(n215), .Q(
        \Storage[10][15] ) );
  EDFQD1 \Storage_reg[10][14]  ( .D(n4), .E(n117), .CP(n272), .Q(
        \Storage[10][14] ) );
  EDFQD1 \Storage_reg[10][13]  ( .D(n8), .E(n116), .CP(n251), .Q(
        \Storage[10][13] ) );
  EDFQD1 \Storage_reg[10][12]  ( .D(n12), .E(n116), .CP(n250), .Q(
        \Storage[10][12] ) );
  EDFQD1 \Storage_reg[10][11]  ( .D(n16), .E(n117), .CP(n249), .Q(
        \Storage[10][11] ) );
  EDFQD1 \Storage_reg[10][10]  ( .D(n20), .E(n118), .CP(n248), .Q(
        \Storage[10][10] ) );
  EDFQD1 \Storage_reg[10][9]  ( .D(n24), .E(n118), .CP(n269), .Q(
        \Storage[10][9] ) );
  EDFQD1 \Storage_reg[10][8]  ( .D(n28), .E(n117), .CP(n255), .Q(
        \Storage[10][8] ) );
  EDFQD1 \Storage_reg[10][7]  ( .D(n32), .E(n116), .CP(n236), .Q(
        \Storage[10][7] ) );
  EDFQD1 \Storage_reg[10][6]  ( .D(n36), .E(n116), .CP(n235), .Q(
        \Storage[10][6] ) );
  EDFQD1 \Storage_reg[10][5]  ( .D(n40), .E(n117), .CP(n234), .Q(
        \Storage[10][5] ) );
  EDFQD1 \Storage_reg[10][4]  ( .D(n44), .E(n118), .CP(n230), .Q(
        \Storage[10][4] ) );
  EDFQD1 \Storage_reg[10][3]  ( .D(n48), .E(n118), .CP(n208), .Q(
        \Storage[10][3] ) );
  EDFQD1 \Storage_reg[10][2]  ( .D(n51), .E(n117), .CP(n206), .Q(
        \Storage[10][2] ) );
  EDFQD1 \Storage_reg[10][1]  ( .D(n55), .E(n118), .CP(n205), .Q(
        \Storage[10][1] ) );
  EDFQD1 \Storage_reg[10][0]  ( .D(n60), .E(n116), .CP(n204), .Q(
        \Storage[10][0] ) );
  EDFQD1 \Storage_reg[9][32]  ( .D(n201), .E(n125), .CP(n203), .Q(
        \Storage[9][32] ) );
  EDFQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(n125), .CP(n278), .Q(
        \Storage[9][31] ) );
  EDFQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(n126), .CP(n257), .Q(
        \Storage[9][30] ) );
  EDFQD1 \Storage_reg[9][29]  ( .D(n57), .E(n126), .CP(n227), .Q(
        \Storage[9][29] ) );
  EDFQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(n125), .CP(n221), .Q(
        \Storage[9][28] ) );
  EDFQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(n124), .CP(n275), .Q(
        \Storage[9][27] ) );
  EDFQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(n124), .CP(n279), .Q(
        \Storage[9][26] ) );
  EDFQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(n125), .CP(n273), .Q(
        \Storage[9][25] ) );
  EDFQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(n124), .CP(n264), .Q(
        \Storage[9][24] ) );
  EDFQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(n126), .CP(n265), .Q(
        \Storage[9][23] ) );
  EDFQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n125), .CP(n266), .Q(
        \Storage[9][22] ) );
  EDFQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(n124), .CP(n261), .Q(
        \Storage[9][21] ) );
  EDFQD1 \Storage_reg[9][20]  ( .D(n21), .E(n126), .CP(n274), .Q(
        \Storage[9][20] ) );
  EDFQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(n124), .CP(n278), .Q(
        \Storage[9][19] ) );
  EDFQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(n124), .CP(n276), .Q(
        \Storage[9][18] ) );
  EDFQD1 \Storage_reg[9][17]  ( .D(n9), .E(n125), .CP(n259), .Q(
        \Storage[9][17] ) );
  EDFQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(n126), .CP(n237), .Q(
        \Storage[9][16] ) );
  EDFQD1 \Storage_reg[9][15]  ( .D(n1), .E(n126), .CP(n219), .Q(
        \Storage[9][15] ) );
  EDFQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(n125), .CP(n270), .Q(
        \Storage[9][14] ) );
  EDFQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(n124), .CP(n271), .Q(
        \Storage[9][13] ) );
  EDFQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n124), .CP(n263), .Q(
        \Storage[9][12] ) );
  EDFQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(n125), .CP(ChipClock), .Q(
        \Storage[9][11] ) );
  EDFQD1 \Storage_reg[9][10]  ( .D(n19), .E(n126), .CP(n254), .Q(
        \Storage[9][10] ) );
  EDFQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(n126), .CP(n207), .Q(
        \Storage[9][9] ) );
  EDFQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(n125), .CP(n256), .Q(
        \Storage[9][8] ) );
  EDFQD1 \Storage_reg[9][7]  ( .D(n31), .E(n124), .CP(n250), .Q(
        \Storage[9][7] ) );
  EDFQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(n124), .CP(n259), .Q(
        \Storage[9][6] ) );
  EDFQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(n125), .CP(n221), .Q(
        \Storage[9][5] ) );
  EDFQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n126), .CP(n270), .Q(
        \Storage[9][4] ) );
  EDFQD1 \Storage_reg[9][3]  ( .D(n47), .E(n126), .CP(n271), .Q(
        \Storage[9][3] ) );
  EDFQD1 \Storage_reg[9][2]  ( .D(n52), .E(n125), .CP(n261), .Q(
        \Storage[9][2] ) );
  EDFQD1 \Storage_reg[9][1]  ( .D(n56), .E(n126), .CP(n204), .Q(
        \Storage[9][1] ) );
  EDFQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n124), .CP(n225), .Q(
        \Storage[9][0] ) );
  EDFQD1 \Storage_reg[6][32]  ( .D(n202), .E(n149), .CP(n267), .Q(
        \Storage[6][32] ) );
  EDFQD1 \Storage_reg[6][31]  ( .D(n63), .E(n149), .CP(n277), .Q(
        \Storage[6][31] ) );
  EDFQD1 \Storage_reg[6][30]  ( .D(n61), .E(n150), .CP(n264), .Q(
        \Storage[6][30] ) );
  EDFQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n150), .CP(n268), .Q(
        \Storage[6][29] ) );
  EDFQD1 \Storage_reg[6][28]  ( .D(n53), .E(n149), .CP(n269), .Q(
        \Storage[6][28] ) );
  EDFQD1 \Storage_reg[6][27]  ( .D(n49), .E(n148), .CP(n270), .Q(
        \Storage[6][27] ) );
  EDFQD1 \Storage_reg[6][26]  ( .D(n45), .E(n148), .CP(n257), .Q(
        \Storage[6][26] ) );
  EDFQD1 \Storage_reg[6][25]  ( .D(n41), .E(n149), .CP(n255), .Q(
        \Storage[6][25] ) );
  EDFQD1 \Storage_reg[6][24]  ( .D(n37), .E(n148), .CP(n228), .Q(
        \Storage[6][24] ) );
  EDFQD1 \Storage_reg[6][23]  ( .D(n33), .E(n150), .CP(n233), .Q(
        \Storage[6][23] ) );
  EDFQD1 \Storage_reg[6][22]  ( .D(n29), .E(n149), .CP(n258), .Q(
        \Storage[6][22] ) );
  EDFQD1 \Storage_reg[6][21]  ( .D(n25), .E(n148), .CP(n239), .Q(
        \Storage[6][21] ) );
  EDFQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n150), .CP(n273), .Q(
        \Storage[6][20] ) );
  EDFQD1 \Storage_reg[6][19]  ( .D(n17), .E(n148), .CP(n277), .Q(
        \Storage[6][19] ) );
  EDFQD1 \Storage_reg[6][18]  ( .D(n13), .E(n148), .CP(n238), .Q(
        \Storage[6][18] ) );
  EDFQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n149), .CP(n254), .Q(
        \Storage[6][17] ) );
  EDFQD1 \Storage_reg[6][16]  ( .D(n5), .E(n150), .CP(n237), .Q(
        \Storage[6][16] ) );
  EDFQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n150), .CP(n279), .Q(
        \Storage[6][15] ) );
  EDFQD1 \Storage_reg[6][14]  ( .D(n3), .E(n149), .CP(n274), .Q(
        \Storage[6][14] ) );
  EDFQD1 \Storage_reg[6][13]  ( .D(n7), .E(n148), .CP(n271), .Q(
        \Storage[6][13] ) );
  EDFQD1 \Storage_reg[6][12]  ( .D(n11), .E(n148), .CP(n260), .Q(
        \Storage[6][12] ) );
  EDFQD1 \Storage_reg[6][11]  ( .D(n15), .E(n149), .CP(ChipClock), .Q(
        \Storage[6][11] ) );
  EDFQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n150), .CP(n267), .Q(
        \Storage[6][10] ) );
  EDFQD1 \Storage_reg[6][9]  ( .D(n23), .E(n150), .CP(n270), .Q(
        \Storage[6][9] ) );
  EDFQD1 \Storage_reg[6][8]  ( .D(n27), .E(n149), .CP(n267), .Q(
        \Storage[6][8] ) );
  EDFQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n148), .CP(n276), .Q(
        \Storage[6][7] ) );
  EDFQD1 \Storage_reg[6][6]  ( .D(n35), .E(n148), .CP(n222), .Q(
        \Storage[6][6] ) );
  EDFQD1 \Storage_reg[6][5]  ( .D(n39), .E(n149), .CP(n207), .Q(
        \Storage[6][5] ) );
  EDFQD1 \Storage_reg[6][4]  ( .D(n43), .E(n150), .CP(n272), .Q(
        \Storage[6][4] ) );
  EDFQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n150), .CP(n268), .Q(
        \Storage[6][3] ) );
  EDFQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n149), .CP(n269), .Q(
        \Storage[6][2] ) );
  EDFQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n150), .CP(n256), .Q(
        \Storage[6][1] ) );
  EDFQD1 \Storage_reg[6][0]  ( .D(n59), .E(n148), .CP(n261), .Q(
        \Storage[6][0] ) );
  EDFQD1 \Storage_reg[5][32]  ( .D(n201), .E(n157), .CP(n262), .Q(
        \Storage[5][32] ) );
  EDFQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n157), .CP(n279), .Q(
        \Storage[5][31] ) );
  EDFQD1 \Storage_reg[5][30]  ( .D(n61), .E(n158), .CP(n268), .Q(
        \Storage[5][30] ) );
  EDFQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n158), .CP(n254), .Q(
        \Storage[5][29] ) );
  EDFQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n157), .CP(ChipClock), .Q(
        \Storage[5][28] ) );
  EDFQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n156), .CP(n277), .Q(
        \Storage[5][27] ) );
  EDFQD1 \Storage_reg[5][26]  ( .D(n45), .E(n156), .CP(n269), .Q(
        \Storage[5][26] ) );
  EDFQD1 \Storage_reg[5][25]  ( .D(n41), .E(n157), .CP(n271), .Q(
        \Storage[5][25] ) );
  EDFQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n156), .CP(n258), .Q(
        \Storage[5][24] ) );
  EDFQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n158), .CP(n274), .Q(
        \Storage[5][23] ) );
  EDFQD1 \Storage_reg[5][22]  ( .D(n29), .E(n157), .CP(n260), .Q(
        \Storage[5][22] ) );
  EDFQD1 \Storage_reg[5][21]  ( .D(n25), .E(n156), .CP(n275), .Q(
        \Storage[5][21] ) );
  EDFQD1 \Storage_reg[5][20]  ( .D(n21), .E(n158), .CP(n272), .Q(
        \Storage[5][20] ) );
  EDFQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n156), .CP(n229), .Q(
        \Storage[5][19] ) );
  EDFQD1 \Storage_reg[5][18]  ( .D(n13), .E(n156), .CP(n277), .Q(
        \Storage[5][18] ) );
  EDFQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n157), .CP(n261), .Q(
        \Storage[5][17] ) );
  EDFQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n158), .CP(n262), .Q(
        \Storage[5][16] ) );
  EDFQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n158), .CP(n263), .Q(
        \Storage[5][15] ) );
  EDFQD1 \Storage_reg[5][14]  ( .D(n3), .E(n157), .CP(n273), .Q(
        \Storage[5][14] ) );
  EDFQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n156), .CP(n264), .Q(
        \Storage[5][13] ) );
  EDFQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n156), .CP(n265), .Q(
        \Storage[5][12] ) );
  EDFQD1 \Storage_reg[5][11]  ( .D(n15), .E(n157), .CP(n266), .Q(
        \Storage[5][11] ) );
  EDFQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n158), .CP(n247), .Q(
        \Storage[5][10] ) );
  EDFQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n158), .CP(n258), .Q(
        \Storage[5][9] ) );
  EDFQD1 \Storage_reg[5][8]  ( .D(n27), .E(n157), .CP(n279), .Q(
        \Storage[5][8] ) );
  EDFQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n156), .CP(n234), .Q(
        \Storage[5][7] ) );
  EDFQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n156), .CP(n257), .Q(
        \Storage[5][6] ) );
  EDFQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n157), .CP(ChipClock), .Q(
        \Storage[5][5] ) );
  EDFQD1 \Storage_reg[5][4]  ( .D(n43), .E(n158), .CP(n278), .Q(
        \Storage[5][4] ) );
  EDFQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n158), .CP(n276), .Q(
        \Storage[5][3] ) );
  EDFQD1 \Storage_reg[5][2]  ( .D(n51), .E(n157), .CP(n255), .Q(
        \Storage[5][2] ) );
  EDFQD1 \Storage_reg[5][1]  ( .D(n55), .E(n158), .CP(n256), .Q(
        \Storage[5][1] ) );
  EDFQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n156), .CP(n257), .Q(
        \Storage[5][0] ) );
  EDFQD1 \Storage_reg[2][32]  ( .D(n200), .E(n181), .CP(n256), .Q(
        \Storage[2][32] ) );
  EDFQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n181), .CP(n272), .Q(
        \Storage[2][31] ) );
  EDFQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n182), .CP(n232), .Q(
        \Storage[2][30] ) );
  EDFQD1 \Storage_reg[2][29]  ( .D(n57), .E(n182), .CP(n259), .Q(
        \Storage[2][29] ) );
  EDFQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n181), .CP(ChipClock), .Q(
        \Storage[2][28] ) );
  EDFQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n180), .CP(n274), .Q(
        \Storage[2][27] ) );
  EDFQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n180), .CP(n261), .Q(
        \Storage[2][26] ) );
  EDFQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n181), .CP(n262), .Q(
        \Storage[2][25] ) );
  EDFQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n180), .CP(n263), .Q(
        \Storage[2][24] ) );
  EDFQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n182), .CP(n264), .Q(
        \Storage[2][23] ) );
  EDFQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n181), .CP(n265), .Q(
        \Storage[2][22] ) );
  EDFQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n180), .CP(n266), .Q(
        \Storage[2][21] ) );
  EDFQD1 \Storage_reg[2][20]  ( .D(n21), .E(n182), .CP(n272), .Q(
        \Storage[2][20] ) );
  EDFQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n180), .CP(n231), .Q(
        \Storage[2][19] ) );
  EDFQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n180), .CP(n267), .Q(
        \Storage[2][18] ) );
  EDFQD1 \Storage_reg[2][17]  ( .D(n9), .E(n181), .CP(n268), .Q(
        \Storage[2][17] ) );
  EDFQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n182), .CP(n269), .Q(
        \Storage[2][16] ) );
  EDFQD1 \Storage_reg[2][15]  ( .D(n1), .E(n182), .CP(n222), .Q(
        \Storage[2][15] ) );
  EDFQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n181), .CP(n252), .Q(
        \Storage[2][14] ) );
  EDFQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n180), .CP(n254), .Q(
        \Storage[2][13] ) );
  EDFQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n180), .CP(n270), .Q(
        \Storage[2][12] ) );
  EDFQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n181), .CP(n271), .Q(
        \Storage[2][11] ) );
  EDFQD1 \Storage_reg[2][10]  ( .D(n19), .E(n182), .CP(n260), .Q(
        \Storage[2][10] ) );
  EDFQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n182), .CP(n259), .Q(
        \Storage[2][9] ) );
  EDFQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n181), .CP(ChipClock), .Q(
        \Storage[2][8] ) );
  EDFQD1 \Storage_reg[2][7]  ( .D(n31), .E(n180), .CP(n249), .Q(
        \Storage[2][7] ) );
  EDFQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n180), .CP(n205), .Q(
        \Storage[2][6] ) );
  EDFQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n181), .CP(n254), .Q(
        \Storage[2][5] ) );
  EDFQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n182), .CP(n277), .Q(
        \Storage[2][4] ) );
  EDFQD1 \Storage_reg[2][3]  ( .D(n47), .E(n182), .CP(n273), .Q(
        \Storage[2][3] ) );
  EDFQD1 \Storage_reg[2][2]  ( .D(n52), .E(n181), .CP(n260), .Q(
        \Storage[2][2] ) );
  EDFQD1 \Storage_reg[2][1]  ( .D(n55), .E(n182), .CP(n273), .Q(
        \Storage[2][1] ) );
  EDFQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n180), .CP(n243), .Q(
        \Storage[2][0] ) );
  EDFQD1 \Storage_reg[1][32]  ( .D(n201), .E(n189), .CP(n235), .Q(
        \Storage[1][32] ) );
  EDFQD1 \Storage_reg[1][31]  ( .D(n63), .E(n189), .CP(n267), .Q(
        \Storage[1][31] ) );
  EDFQD1 \Storage_reg[1][30]  ( .D(n61), .E(n190), .CP(n277), .Q(
        \Storage[1][30] ) );
  EDFQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n190), .CP(ChipClock), .Q(
        \Storage[1][29] ) );
  EDFQD1 \Storage_reg[1][28]  ( .D(n53), .E(n189), .CP(n275), .Q(
        \Storage[1][28] ) );
  EDFQD1 \Storage_reg[1][27]  ( .D(n49), .E(n188), .CP(n258), .Q(
        \Storage[1][27] ) );
  EDFQD1 \Storage_reg[1][26]  ( .D(n45), .E(n188), .CP(n259), .Q(
        \Storage[1][26] ) );
  EDFQD1 \Storage_reg[1][25]  ( .D(n41), .E(n189), .CP(n260), .Q(
        \Storage[1][25] ) );
  EDFQD1 \Storage_reg[1][24]  ( .D(n37), .E(n188), .CP(n276), .Q(
        \Storage[1][24] ) );
  EDFQD1 \Storage_reg[1][23]  ( .D(n33), .E(n190), .CP(n255), .Q(
        \Storage[1][23] ) );
  EDFQD1 \Storage_reg[1][22]  ( .D(n29), .E(n189), .CP(n256), .Q(
        \Storage[1][22] ) );
  EDFQD1 \Storage_reg[1][21]  ( .D(n25), .E(n188), .CP(n257), .Q(
        \Storage[1][21] ) );
  EDFQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n190), .CP(n258), .Q(
        \Storage[1][20] ) );
  EDFQD1 \Storage_reg[1][19]  ( .D(n17), .E(n188), .CP(n259), .Q(
        \Storage[1][19] ) );
  EDFQD1 \Storage_reg[1][18]  ( .D(n13), .E(n188), .CP(n268), .Q(
        \Storage[1][18] ) );
  EDFQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n189), .CP(n269), .Q(
        \Storage[1][17] ) );
  EDFQD1 \Storage_reg[1][16]  ( .D(n5), .E(n190), .CP(n264), .Q(
        \Storage[1][16] ) );
  EDFQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n190), .CP(n265), .Q(
        \Storage[1][15] ) );
  EDFQD1 \Storage_reg[1][14]  ( .D(n3), .E(n189), .CP(n266), .Q(
        \Storage[1][14] ) );
  EDFQD1 \Storage_reg[1][13]  ( .D(n7), .E(n188), .CP(n263), .Q(
        \Storage[1][13] ) );
  EDFQD1 \Storage_reg[1][12]  ( .D(n11), .E(n188), .CP(n262), .Q(
        \Storage[1][12] ) );
  EDFQD1 \Storage_reg[1][11]  ( .D(n15), .E(n189), .CP(n261), .Q(
        \Storage[1][11] ) );
  EDFQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n190), .CP(n253), .Q(
        \Storage[1][10] ) );
  EDFQD1 \Storage_reg[1][9]  ( .D(n23), .E(n190), .CP(n256), .Q(
        \Storage[1][9] ) );
  EDFQD1 \Storage_reg[1][8]  ( .D(n27), .E(n189), .CP(n253), .Q(
        \Storage[1][8] ) );
  EDFQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n188), .CP(n254), .Q(
        \Storage[1][7] ) );
  EDFQD1 \Storage_reg[1][6]  ( .D(n35), .E(n188), .CP(n271), .Q(
        \Storage[1][6] ) );
  EDFQD1 \Storage_reg[1][5]  ( .D(n39), .E(n189), .CP(n277), .Q(
        \Storage[1][5] ) );
  EDFQD1 \Storage_reg[1][4]  ( .D(n43), .E(n190), .CP(n242), .Q(
        \Storage[1][4] ) );
  EDFQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n190), .CP(n259), .Q(
        \Storage[1][3] ) );
  EDFQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n189), .CP(n240), .Q(
        \Storage[1][2] ) );
  EDFQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n190), .CP(n278), .Q(
        \Storage[1][1] ) );
  EDFQD1 \Storage_reg[1][0]  ( .D(n59), .E(n188), .CP(n276), .Q(
        \Storage[1][0] ) );
  EDFQD1 \Storage_reg[23][32]  ( .D(n202), .E(n129), .CP(n230), .Q(
        \Storage[23][32] ) );
  EDFQD1 \Storage_reg[23][31]  ( .D(n64), .E(n129), .CP(n229), .Q(
        \Storage[23][31] ) );
  EDFQD1 \Storage_reg[23][30]  ( .D(n62), .E(n130), .CP(n229), .Q(
        \Storage[23][30] ) );
  EDFQD1 \Storage_reg[23][29]  ( .D(n58), .E(n130), .CP(n229), .Q(
        \Storage[23][29] ) );
  EDFQD1 \Storage_reg[23][28]  ( .D(n54), .E(n129), .CP(n229), .Q(
        \Storage[23][28] ) );
  EDFQD1 \Storage_reg[23][27]  ( .D(n50), .E(n128), .CP(n229), .Q(
        \Storage[23][27] ) );
  EDFQD1 \Storage_reg[23][26]  ( .D(n46), .E(n128), .CP(n229), .Q(
        \Storage[23][26] ) );
  EDFQD1 \Storage_reg[23][25]  ( .D(n42), .E(n129), .CP(n229), .Q(
        \Storage[23][25] ) );
  EDFQD1 \Storage_reg[23][24]  ( .D(n38), .E(n128), .CP(n229), .Q(
        \Storage[23][24] ) );
  EDFQD1 \Storage_reg[23][23]  ( .D(n34), .E(n130), .CP(n229), .Q(
        \Storage[23][23] ) );
  EDFQD1 \Storage_reg[23][22]  ( .D(n30), .E(n129), .CP(n229), .Q(
        \Storage[23][22] ) );
  EDFQD1 \Storage_reg[23][21]  ( .D(n26), .E(n128), .CP(n229), .Q(
        \Storage[23][21] ) );
  EDFQD1 \Storage_reg[23][20]  ( .D(n22), .E(n130), .CP(n228), .Q(
        \Storage[23][20] ) );
  EDFQD1 \Storage_reg[23][19]  ( .D(n18), .E(n128), .CP(n228), .Q(
        \Storage[23][19] ) );
  EDFQD1 \Storage_reg[23][18]  ( .D(n14), .E(n128), .CP(n228), .Q(
        \Storage[23][18] ) );
  EDFQD1 \Storage_reg[23][17]  ( .D(n10), .E(n129), .CP(n228), .Q(
        \Storage[23][17] ) );
  EDFQD1 \Storage_reg[23][16]  ( .D(n6), .E(n130), .CP(n228), .Q(
        \Storage[23][16] ) );
  EDFQD1 \Storage_reg[23][15]  ( .D(n2), .E(n130), .CP(n228), .Q(
        \Storage[23][15] ) );
  EDFQD1 \Storage_reg[23][14]  ( .D(n4), .E(n129), .CP(n228), .Q(
        \Storage[23][14] ) );
  EDFQD1 \Storage_reg[23][13]  ( .D(n8), .E(n128), .CP(n228), .Q(
        \Storage[23][13] ) );
  EDFQD1 \Storage_reg[23][12]  ( .D(n12), .E(n128), .CP(n228), .Q(
        \Storage[23][12] ) );
  EDFQD1 \Storage_reg[23][11]  ( .D(n16), .E(n129), .CP(n228), .Q(
        \Storage[23][11] ) );
  EDFQD1 \Storage_reg[23][10]  ( .D(n20), .E(n130), .CP(n228), .Q(
        \Storage[23][10] ) );
  EDFQD1 \Storage_reg[23][9]  ( .D(n24), .E(n130), .CP(n227), .Q(
        \Storage[23][9] ) );
  EDFQD1 \Storage_reg[23][8]  ( .D(n28), .E(n129), .CP(n227), .Q(
        \Storage[23][8] ) );
  EDFQD1 \Storage_reg[23][7]  ( .D(n32), .E(n128), .CP(n227), .Q(
        \Storage[23][7] ) );
  EDFQD1 \Storage_reg[23][6]  ( .D(n36), .E(n128), .CP(n227), .Q(
        \Storage[23][6] ) );
  EDFQD1 \Storage_reg[23][5]  ( .D(n40), .E(n129), .CP(n227), .Q(
        \Storage[23][5] ) );
  EDFQD1 \Storage_reg[23][4]  ( .D(n44), .E(n130), .CP(n227), .Q(
        \Storage[23][4] ) );
  EDFQD1 \Storage_reg[23][3]  ( .D(n48), .E(n130), .CP(n227), .Q(
        \Storage[23][3] ) );
  EDFQD1 \Storage_reg[23][2]  ( .D(n51), .E(n129), .CP(n227), .Q(
        \Storage[23][2] ) );
  EDFQD1 \Storage_reg[23][1]  ( .D(n55), .E(n130), .CP(n227), .Q(
        \Storage[23][1] ) );
  EDFQD1 \Storage_reg[23][0]  ( .D(n60), .E(n128), .CP(n227), .Q(
        \Storage[23][0] ) );
  EDFQD1 \Storage_reg[20][32]  ( .D(n201), .E(n105), .CP(n221), .Q(
        \Storage[20][32] ) );
  EDFQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(n105), .CP(n220), .Q(
        \Storage[20][31] ) );
  EDFQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(n106), .CP(n220), .Q(
        \Storage[20][30] ) );
  EDFQD1 \Storage_reg[20][29]  ( .D(n57), .E(n106), .CP(n220), .Q(
        \Storage[20][29] ) );
  EDFQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(n105), .CP(n220), .Q(
        \Storage[20][28] ) );
  EDFQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(n104), .CP(n220), .Q(
        \Storage[20][27] ) );
  EDFQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(n104), .CP(n220), .Q(
        \Storage[20][26] ) );
  EDFQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(n105), .CP(n220), .Q(
        \Storage[20][25] ) );
  EDFQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(n104), .CP(n220), .Q(
        \Storage[20][24] ) );
  EDFQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(n106), .CP(n220), .Q(
        \Storage[20][23] ) );
  EDFQD1 \Storage_reg[20][22]  ( .D(DataI[22]), .E(n105), .CP(n220), .Q(
        \Storage[20][22] ) );
  EDFQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(n104), .CP(n220), .Q(
        \Storage[20][21] ) );
  EDFQD1 \Storage_reg[20][20]  ( .D(n21), .E(n106), .CP(n219), .Q(
        \Storage[20][20] ) );
  EDFQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(n104), .CP(n219), .Q(
        \Storage[20][19] ) );
  EDFQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(n104), .CP(n219), .Q(
        \Storage[20][18] ) );
  EDFQD1 \Storage_reg[20][17]  ( .D(n9), .E(n105), .CP(n219), .Q(
        \Storage[20][17] ) );
  EDFQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(n106), .CP(n219), .Q(
        \Storage[20][16] ) );
  EDFQD1 \Storage_reg[20][15]  ( .D(n1), .E(n106), .CP(n219), .Q(
        \Storage[20][15] ) );
  EDFQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(n105), .CP(n219), .Q(
        \Storage[20][14] ) );
  EDFQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(n104), .CP(n219), .Q(
        \Storage[20][13] ) );
  EDFQD1 \Storage_reg[20][12]  ( .D(DataI[12]), .E(n104), .CP(n219), .Q(
        \Storage[20][12] ) );
  EDFQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(n105), .CP(n219), .Q(
        \Storage[20][11] ) );
  EDFQD1 \Storage_reg[20][10]  ( .D(n19), .E(n106), .CP(n219), .Q(
        \Storage[20][10] ) );
  EDFQD1 \Storage_reg[20][9]  ( .D(DataI[9]), .E(n106), .CP(n218), .Q(
        \Storage[20][9] ) );
  EDFQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(n105), .CP(n218), .Q(
        \Storage[20][8] ) );
  EDFQD1 \Storage_reg[20][7]  ( .D(n31), .E(n104), .CP(n218), .Q(
        \Storage[20][7] ) );
  EDFQD1 \Storage_reg[20][6]  ( .D(DataI[6]), .E(n104), .CP(n218), .Q(
        \Storage[20][6] ) );
  EDFQD1 \Storage_reg[20][5]  ( .D(DataI[5]), .E(n105), .CP(n218), .Q(
        \Storage[20][5] ) );
  EDFQD1 \Storage_reg[20][4]  ( .D(DataI[4]), .E(n106), .CP(n218), .Q(
        \Storage[20][4] ) );
  EDFQD1 \Storage_reg[20][3]  ( .D(n47), .E(n106), .CP(n218), .Q(
        \Storage[20][3] ) );
  EDFQD1 \Storage_reg[20][2]  ( .D(n52), .E(n105), .CP(n218), .Q(
        \Storage[20][2] ) );
  EDFQD1 \Storage_reg[20][1]  ( .D(n56), .E(n106), .CP(n218), .Q(
        \Storage[20][1] ) );
  EDFQD1 \Storage_reg[20][0]  ( .D(DataI[0]), .E(n104), .CP(n218), .Q(
        \Storage[20][0] ) );
  EDFQD1 \Storage_reg[19][32]  ( .D(n202), .E(n97), .CP(n218), .Q(
        \Storage[19][32] ) );
  EDFQD1 \Storage_reg[19][31]  ( .D(n63), .E(n97), .CP(n217), .Q(
        \Storage[19][31] ) );
  EDFQD1 \Storage_reg[19][30]  ( .D(n61), .E(n98), .CP(n217), .Q(
        \Storage[19][30] ) );
  EDFQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(n98), .CP(n217), .Q(
        \Storage[19][29] ) );
  EDFQD1 \Storage_reg[19][28]  ( .D(n53), .E(n97), .CP(n217), .Q(
        \Storage[19][28] ) );
  EDFQD1 \Storage_reg[19][27]  ( .D(n49), .E(n96), .CP(n217), .Q(
        \Storage[19][27] ) );
  EDFQD1 \Storage_reg[19][26]  ( .D(n45), .E(n96), .CP(n217), .Q(
        \Storage[19][26] ) );
  EDFQD1 \Storage_reg[19][25]  ( .D(n41), .E(n97), .CP(n217), .Q(
        \Storage[19][25] ) );
  EDFQD1 \Storage_reg[19][24]  ( .D(n37), .E(n96), .CP(n217), .Q(
        \Storage[19][24] ) );
  EDFQD1 \Storage_reg[19][23]  ( .D(n33), .E(n98), .CP(n217), .Q(
        \Storage[19][23] ) );
  EDFQD1 \Storage_reg[19][22]  ( .D(n29), .E(n97), .CP(n217), .Q(
        \Storage[19][22] ) );
  EDFQD1 \Storage_reg[19][21]  ( .D(n25), .E(n96), .CP(n217), .Q(
        \Storage[19][21] ) );
  EDFQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(n98), .CP(n216), .Q(
        \Storage[19][20] ) );
  EDFQD1 \Storage_reg[19][19]  ( .D(n17), .E(n96), .CP(n216), .Q(
        \Storage[19][19] ) );
  EDFQD1 \Storage_reg[19][18]  ( .D(n13), .E(n96), .CP(n216), .Q(
        \Storage[19][18] ) );
  EDFQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(n97), .CP(n216), .Q(
        \Storage[19][17] ) );
  EDFQD1 \Storage_reg[19][16]  ( .D(n5), .E(n98), .CP(n216), .Q(
        \Storage[19][16] ) );
  EDFQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(n98), .CP(n216), .Q(
        \Storage[19][15] ) );
  EDFQD1 \Storage_reg[19][14]  ( .D(n3), .E(n97), .CP(n216), .Q(
        \Storage[19][14] ) );
  EDFQD1 \Storage_reg[19][13]  ( .D(n7), .E(n96), .CP(n216), .Q(
        \Storage[19][13] ) );
  EDFQD1 \Storage_reg[19][12]  ( .D(n11), .E(n96), .CP(n216), .Q(
        \Storage[19][12] ) );
  EDFQD1 \Storage_reg[19][11]  ( .D(n15), .E(n97), .CP(n216), .Q(
        \Storage[19][11] ) );
  EDFQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(n98), .CP(n216), .Q(
        \Storage[19][10] ) );
  EDFQD1 \Storage_reg[19][9]  ( .D(n23), .E(n98), .CP(n215), .Q(
        \Storage[19][9] ) );
  EDFQD1 \Storage_reg[19][8]  ( .D(n27), .E(n97), .CP(n215), .Q(
        \Storage[19][8] ) );
  EDFQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(n96), .CP(n215), .Q(
        \Storage[19][7] ) );
  EDFQD1 \Storage_reg[19][6]  ( .D(n35), .E(n96), .CP(n215), .Q(
        \Storage[19][6] ) );
  EDFQD1 \Storage_reg[19][5]  ( .D(n39), .E(n97), .CP(n215), .Q(
        \Storage[19][5] ) );
  EDFQD1 \Storage_reg[19][4]  ( .D(n43), .E(n98), .CP(n215), .Q(
        \Storage[19][4] ) );
  EDFQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(n98), .CP(n215), .Q(
        \Storage[19][3] ) );
  EDFQD1 \Storage_reg[19][2]  ( .D(DataI[2]), .E(n97), .CP(n215), .Q(
        \Storage[19][2] ) );
  EDFQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(n98), .CP(n215), .Q(
        \Storage[19][1] ) );
  EDFQD1 \Storage_reg[19][0]  ( .D(n59), .E(n96), .CP(n215), .Q(
        \Storage[19][0] ) );
  EDFQD1 \Storage_reg[16][32]  ( .D(n200), .E(n73), .CP(n209), .Q(
        \Storage[16][32] ) );
  EDFQD1 \Storage_reg[16][31]  ( .D(n64), .E(n73), .CP(n208), .Q(
        \Storage[16][31] ) );
  EDFQD1 \Storage_reg[16][30]  ( .D(n62), .E(n74), .CP(n208), .Q(
        \Storage[16][30] ) );
  EDFQD1 \Storage_reg[16][29]  ( .D(n58), .E(n74), .CP(n208), .Q(
        \Storage[16][29] ) );
  EDFQD1 \Storage_reg[16][28]  ( .D(n54), .E(n73), .CP(n208), .Q(
        \Storage[16][28] ) );
  EDFQD1 \Storage_reg[16][27]  ( .D(n50), .E(n72), .CP(n208), .Q(
        \Storage[16][27] ) );
  EDFQD1 \Storage_reg[16][26]  ( .D(n46), .E(n72), .CP(n208), .Q(
        \Storage[16][26] ) );
  EDFQD1 \Storage_reg[16][25]  ( .D(n42), .E(n73), .CP(n208), .Q(
        \Storage[16][25] ) );
  EDFQD1 \Storage_reg[16][24]  ( .D(n38), .E(n72), .CP(n208), .Q(
        \Storage[16][24] ) );
  EDFQD1 \Storage_reg[16][23]  ( .D(n34), .E(n74), .CP(n208), .Q(
        \Storage[16][23] ) );
  EDFQD1 \Storage_reg[16][22]  ( .D(n30), .E(n73), .CP(n208), .Q(
        \Storage[16][22] ) );
  EDFQD1 \Storage_reg[16][21]  ( .D(n26), .E(n72), .CP(n208), .Q(
        \Storage[16][21] ) );
  EDFQD1 \Storage_reg[16][20]  ( .D(n22), .E(n74), .CP(n207), .Q(
        \Storage[16][20] ) );
  EDFQD1 \Storage_reg[16][19]  ( .D(n18), .E(n72), .CP(n207), .Q(
        \Storage[16][19] ) );
  EDFQD1 \Storage_reg[16][18]  ( .D(n14), .E(n72), .CP(n207), .Q(
        \Storage[16][18] ) );
  EDFQD1 \Storage_reg[16][17]  ( .D(n10), .E(n73), .CP(n207), .Q(
        \Storage[16][17] ) );
  EDFQD1 \Storage_reg[16][16]  ( .D(n6), .E(n74), .CP(n207), .Q(
        \Storage[16][16] ) );
  EDFQD1 \Storage_reg[16][15]  ( .D(n2), .E(n74), .CP(n207), .Q(
        \Storage[16][15] ) );
  EDFQD1 \Storage_reg[16][14]  ( .D(n4), .E(n73), .CP(n207), .Q(
        \Storage[16][14] ) );
  EDFQD1 \Storage_reg[16][13]  ( .D(n8), .E(n72), .CP(n207), .Q(
        \Storage[16][13] ) );
  EDFQD1 \Storage_reg[16][12]  ( .D(n12), .E(n72), .CP(n207), .Q(
        \Storage[16][12] ) );
  EDFQD1 \Storage_reg[16][11]  ( .D(n16), .E(n73), .CP(n207), .Q(
        \Storage[16][11] ) );
  EDFQD1 \Storage_reg[16][10]  ( .D(n20), .E(n74), .CP(n207), .Q(
        \Storage[16][10] ) );
  EDFQD1 \Storage_reg[16][9]  ( .D(n24), .E(n74), .CP(n227), .Q(
        \Storage[16][9] ) );
  EDFQD1 \Storage_reg[16][8]  ( .D(n28), .E(n73), .CP(n270), .Q(
        \Storage[16][8] ) );
  EDFQD1 \Storage_reg[16][7]  ( .D(n32), .E(n72), .CP(n253), .Q(
        \Storage[16][7] ) );
  EDFQD1 \Storage_reg[16][6]  ( .D(n36), .E(n72), .CP(n252), .Q(
        \Storage[16][6] ) );
  EDFQD1 \Storage_reg[16][5]  ( .D(n40), .E(n73), .CP(n248), .Q(
        \Storage[16][5] ) );
  EDFQD1 \Storage_reg[16][4]  ( .D(n44), .E(n74), .CP(n245), .Q(
        \Storage[16][4] ) );
  EDFQD1 \Storage_reg[16][3]  ( .D(n48), .E(n74), .CP(n244), .Q(
        \Storage[16][3] ) );
  EDFQD1 \Storage_reg[16][2]  ( .D(n51), .E(n73), .CP(n243), .Q(
        \Storage[16][2] ) );
  EDFQD1 \Storage_reg[16][1]  ( .D(n55), .E(n74), .CP(n233), .Q(
        \Storage[16][1] ) );
  EDFQD1 \Storage_reg[16][0]  ( .D(n60), .E(n72), .CP(n232), .Q(
        \Storage[16][0] ) );
  EDFQD1 \Storage_reg[15][32]  ( .D(n200), .E(n77), .CP(n231), .Q(
        \Storage[15][32] ) );
  EDFQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n77), .CP(n205), .Q(
        \Storage[15][31] ) );
  EDFQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(n78), .CP(n270), .Q(
        \Storage[15][30] ) );
  EDFQD1 \Storage_reg[15][29]  ( .D(n57), .E(n78), .CP(n226), .Q(
        \Storage[15][29] ) );
  EDFQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(n77), .CP(n225), .Q(
        \Storage[15][28] ) );
  EDFQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(n76), .CP(n215), .Q(
        \Storage[15][27] ) );
  EDFQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(n76), .CP(n214), .Q(
        \Storage[15][26] ) );
  EDFQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(n77), .CP(n213), .Q(
        \Storage[15][25] ) );
  EDFQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(n76), .CP(n212), .Q(
        \Storage[15][24] ) );
  EDFQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(n78), .CP(n211), .Q(
        \Storage[15][23] ) );
  EDFQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(n77), .CP(n210), .Q(
        \Storage[15][22] ) );
  EDFQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n76), .CP(n209), .Q(
        \Storage[15][21] ) );
  EDFQD1 \Storage_reg[15][20]  ( .D(n21), .E(n78), .CP(n206), .Q(
        \Storage[15][20] ) );
  EDFQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n76), .CP(n206), .Q(
        \Storage[15][19] ) );
  EDFQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n76), .CP(n206), .Q(
        \Storage[15][18] ) );
  EDFQD1 \Storage_reg[15][17]  ( .D(n9), .E(n77), .CP(n206), .Q(
        \Storage[15][17] ) );
  EDFQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n78), .CP(n206), .Q(
        \Storage[15][16] ) );
  EDFQD1 \Storage_reg[15][15]  ( .D(n1), .E(n78), .CP(n206), .Q(
        \Storage[15][15] ) );
  EDFQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n77), .CP(n206), .Q(
        \Storage[15][14] ) );
  EDFQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n76), .CP(n206), .Q(
        \Storage[15][13] ) );
  EDFQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(n76), .CP(n206), .Q(
        \Storage[15][12] ) );
  EDFQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n77), .CP(n206), .Q(
        \Storage[15][11] ) );
  EDFQD1 \Storage_reg[15][10]  ( .D(n19), .E(n78), .CP(n206), .Q(
        \Storage[15][10] ) );
  EDFQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(n78), .CP(n205), .Q(
        \Storage[15][9] ) );
  EDFQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(n77), .CP(n205), .Q(
        \Storage[15][8] ) );
  EDFQD1 \Storage_reg[15][7]  ( .D(n31), .E(n76), .CP(n205), .Q(
        \Storage[15][7] ) );
  EDFQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(n76), .CP(n205), .Q(
        \Storage[15][6] ) );
  EDFQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(n77), .CP(n205), .Q(
        \Storage[15][5] ) );
  EDFQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(n78), .CP(n205), .Q(
        \Storage[15][4] ) );
  EDFQD1 \Storage_reg[15][3]  ( .D(n47), .E(n78), .CP(n205), .Q(
        \Storage[15][3] ) );
  EDFQD1 \Storage_reg[15][2]  ( .D(n52), .E(n77), .CP(n205), .Q(
        \Storage[15][2] ) );
  EDFQD1 \Storage_reg[15][1]  ( .D(n56), .E(n78), .CP(n205), .Q(
        \Storage[15][1] ) );
  EDFQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(n76), .CP(n205), .Q(
        \Storage[15][0] ) );
  EDFQD1 \Storage_reg[12][32]  ( .D(n202), .E(n101), .CP(n255), .Q(
        \Storage[12][32] ) );
  EDFQD1 \Storage_reg[12][31]  ( .D(n64), .E(n101), .CP(n215), .Q(
        \Storage[12][31] ) );
  EDFQD1 \Storage_reg[12][30]  ( .D(n62), .E(n102), .CP(n219), .Q(
        \Storage[12][30] ) );
  EDFQD1 \Storage_reg[12][29]  ( .D(n58), .E(n102), .CP(n216), .Q(
        \Storage[12][29] ) );
  EDFQD1 \Storage_reg[12][28]  ( .D(n54), .E(n101), .CP(n270), .Q(
        \Storage[12][28] ) );
  EDFQD1 \Storage_reg[12][27]  ( .D(n50), .E(n100), .CP(n271), .Q(
        \Storage[12][27] ) );
  EDFQD1 \Storage_reg[12][26]  ( .D(n46), .E(n100), .CP(n274), .Q(
        \Storage[12][26] ) );
  EDFQD1 \Storage_reg[12][25]  ( .D(n42), .E(n101), .CP(n260), .Q(
        \Storage[12][25] ) );
  EDFQD1 \Storage_reg[12][24]  ( .D(n38), .E(n100), .CP(ChipClock), .Q(
        \Storage[12][24] ) );
  EDFQD1 \Storage_reg[12][23]  ( .D(n34), .E(n102), .CP(n254), .Q(
        \Storage[12][23] ) );
  EDFQD1 \Storage_reg[12][22]  ( .D(n30), .E(n101), .CP(n242), .Q(
        \Storage[12][22] ) );
  EDFQD1 \Storage_reg[12][21]  ( .D(n26), .E(n100), .CP(n224), .Q(
        \Storage[12][21] ) );
  EDFQD1 \Storage_reg[12][20]  ( .D(n22), .E(n102), .CP(n220), .Q(
        \Storage[12][20] ) );
  EDFQD1 \Storage_reg[12][19]  ( .D(n18), .E(n100), .CP(n214), .Q(
        \Storage[12][19] ) );
  EDFQD1 \Storage_reg[12][18]  ( .D(n14), .E(n100), .CP(n213), .Q(
        \Storage[12][18] ) );
  EDFQD1 \Storage_reg[12][17]  ( .D(n10), .E(n101), .CP(n212), .Q(
        \Storage[12][17] ) );
  EDFQD1 \Storage_reg[12][16]  ( .D(n6), .E(n102), .CP(n211), .Q(
        \Storage[12][16] ) );
  EDFQD1 \Storage_reg[12][15]  ( .D(n2), .E(n102), .CP(n210), .Q(
        \Storage[12][15] ) );
  EDFQD1 \Storage_reg[12][14]  ( .D(n4), .E(n101), .CP(n209), .Q(
        \Storage[12][14] ) );
  EDFQD1 \Storage_reg[12][13]  ( .D(n8), .E(n100), .CP(n208), .Q(
        \Storage[12][13] ) );
  EDFQD1 \Storage_reg[12][12]  ( .D(n12), .E(n100), .CP(n207), .Q(
        \Storage[12][12] ) );
  EDFQD1 \Storage_reg[12][11]  ( .D(n16), .E(n101), .CP(n271), .Q(
        \Storage[12][11] ) );
  EDFQD1 \Storage_reg[12][10]  ( .D(n20), .E(n102), .CP(n223), .Q(
        \Storage[12][10] ) );
  EDFQD1 \Storage_reg[12][9]  ( .D(n24), .E(n102), .CP(n236), .Q(
        \Storage[12][9] ) );
  EDFQD1 \Storage_reg[12][8]  ( .D(n28), .E(n101), .CP(n235), .Q(
        \Storage[12][8] ) );
  EDFQD1 \Storage_reg[12][7]  ( .D(n32), .E(n100), .CP(n234), .Q(
        \Storage[12][7] ) );
  EDFQD1 \Storage_reg[12][6]  ( .D(n36), .E(n100), .CP(n237), .Q(
        \Storage[12][6] ) );
  EDFQD1 \Storage_reg[12][5]  ( .D(n40), .E(n101), .CP(n239), .Q(
        \Storage[12][5] ) );
  EDFQD1 \Storage_reg[12][4]  ( .D(n44), .E(n102), .CP(n238), .Q(
        \Storage[12][4] ) );
  EDFQD1 \Storage_reg[12][3]  ( .D(n48), .E(n102), .CP(n240), .Q(
        \Storage[12][3] ) );
  EDFQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(n101), .CP(n241), .Q(
        \Storage[12][2] ) );
  EDFQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(n102), .CP(n242), .Q(
        \Storage[12][1] ) );
  EDFQD1 \Storage_reg[12][0]  ( .D(n60), .E(n100), .CP(n251), .Q(
        \Storage[12][0] ) );
  EDFQD1 \Storage_reg[11][32]  ( .D(n202), .E(n109), .CP(n250), .Q(
        \Storage[11][32] ) );
  EDFQD1 \Storage_reg[11][31]  ( .D(n64), .E(n109), .CP(n264), .Q(
        \Storage[11][31] ) );
  EDFQD1 \Storage_reg[11][30]  ( .D(n62), .E(n110), .CP(n270), .Q(
        \Storage[11][30] ) );
  EDFQD1 \Storage_reg[11][29]  ( .D(n58), .E(n110), .CP(n258), .Q(
        \Storage[11][29] ) );
  EDFQD1 \Storage_reg[11][28]  ( .D(n54), .E(n109), .CP(n275), .Q(
        \Storage[11][28] ) );
  EDFQD1 \Storage_reg[11][27]  ( .D(n50), .E(n108), .CP(n278), .Q(
        \Storage[11][27] ) );
  EDFQD1 \Storage_reg[11][26]  ( .D(n46), .E(n108), .CP(n273), .Q(
        \Storage[11][26] ) );
  EDFQD1 \Storage_reg[11][25]  ( .D(n42), .E(n109), .CP(n279), .Q(
        \Storage[11][25] ) );
  EDFQD1 \Storage_reg[11][24]  ( .D(n38), .E(n108), .CP(n274), .Q(
        \Storage[11][24] ) );
  EDFQD1 \Storage_reg[11][23]  ( .D(n34), .E(n110), .CP(n261), .Q(
        \Storage[11][23] ) );
  EDFQD1 \Storage_reg[11][22]  ( .D(n30), .E(n109), .CP(n262), .Q(
        \Storage[11][22] ) );
  EDFQD1 \Storage_reg[11][21]  ( .D(n26), .E(n108), .CP(n263), .Q(
        \Storage[11][21] ) );
  EDFQD1 \Storage_reg[11][20]  ( .D(n22), .E(n110), .CP(n220), .Q(
        \Storage[11][20] ) );
  EDFQD1 \Storage_reg[11][19]  ( .D(n18), .E(n108), .CP(n271), .Q(
        \Storage[11][19] ) );
  EDFQD1 \Storage_reg[11][18]  ( .D(n14), .E(n108), .CP(n265), .Q(
        \Storage[11][18] ) );
  EDFQD1 \Storage_reg[11][17]  ( .D(n10), .E(n109), .CP(n266), .Q(
        \Storage[11][17] ) );
  EDFQD1 \Storage_reg[11][16]  ( .D(n6), .E(n110), .CP(n272), .Q(
        \Storage[11][16] ) );
  EDFQD1 \Storage_reg[11][15]  ( .D(n2), .E(n110), .CP(n267), .Q(
        \Storage[11][15] ) );
  EDFQD1 \Storage_reg[11][14]  ( .D(n4), .E(n109), .CP(n268), .Q(
        \Storage[11][14] ) );
  EDFQD1 \Storage_reg[11][13]  ( .D(n8), .E(n108), .CP(n269), .Q(
        \Storage[11][13] ) );
  EDFQD1 \Storage_reg[11][12]  ( .D(n12), .E(n108), .CP(n276), .Q(
        \Storage[11][12] ) );
  EDFQD1 \Storage_reg[11][11]  ( .D(n16), .E(n109), .CP(n255), .Q(
        \Storage[11][11] ) );
  EDFQD1 \Storage_reg[11][10]  ( .D(n20), .E(n110), .CP(n256), .Q(
        \Storage[11][10] ) );
  EDFQD1 \Storage_reg[11][9]  ( .D(n24), .E(n110), .CP(n203), .Q(
        \Storage[11][9] ) );
  EDFQD1 \Storage_reg[11][8]  ( .D(n28), .E(n109), .CP(n246), .Q(
        \Storage[11][8] ) );
  EDFQD1 \Storage_reg[11][7]  ( .D(n32), .E(n108), .CP(n223), .Q(
        \Storage[11][7] ) );
  EDFQD1 \Storage_reg[11][6]  ( .D(n36), .E(n108), .CP(n222), .Q(
        \Storage[11][6] ) );
  EDFQD1 \Storage_reg[11][5]  ( .D(n40), .E(n109), .CP(n219), .Q(
        \Storage[11][5] ) );
  EDFQD1 \Storage_reg[11][4]  ( .D(n44), .E(n110), .CP(n220), .Q(
        \Storage[11][4] ) );
  EDFQD1 \Storage_reg[11][3]  ( .D(n48), .E(n110), .CP(n221), .Q(
        \Storage[11][3] ) );
  EDFQD1 \Storage_reg[11][2]  ( .D(n51), .E(n109), .CP(n216), .Q(
        \Storage[11][2] ) );
  EDFQD1 \Storage_reg[11][1]  ( .D(n56), .E(n110), .CP(n217), .Q(
        \Storage[11][1] ) );
  EDFQD1 \Storage_reg[11][0]  ( .D(n60), .E(n108), .CP(n218), .Q(
        \Storage[11][0] ) );
  EDFQD1 \Storage_reg[8][32]  ( .D(n200), .E(n133), .CP(n277), .Q(
        \Storage[8][32] ) );
  EDFQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(n133), .CP(n262), .Q(
        \Storage[8][31] ) );
  EDFQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(n134), .CP(n279), .Q(
        \Storage[8][30] ) );
  EDFQD1 \Storage_reg[8][29]  ( .D(n57), .E(n134), .CP(n272), .Q(
        \Storage[8][29] ) );
  EDFQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(n133), .CP(n267), .Q(
        \Storage[8][28] ) );
  EDFQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(n132), .CP(n268), .Q(
        \Storage[8][27] ) );
  EDFQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(n132), .CP(n269), .Q(
        \Storage[8][26] ) );
  EDFQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(n133), .CP(n273), .Q(
        \Storage[8][25] ) );
  EDFQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(n132), .CP(n264), .Q(
        \Storage[8][24] ) );
  EDFQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(n134), .CP(n265), .Q(
        \Storage[8][23] ) );
  EDFQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(n133), .CP(n266), .Q(
        \Storage[8][22] ) );
  EDFQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(n132), .CP(n261), .Q(
        \Storage[8][21] ) );
  EDFQD1 \Storage_reg[8][20]  ( .D(n21), .E(n134), .CP(n248), .Q(
        \Storage[8][20] ) );
  EDFQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(n132), .CP(n240), .Q(
        \Storage[8][19] ) );
  EDFQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(n132), .CP(n263), .Q(
        \Storage[8][18] ) );
  EDFQD1 \Storage_reg[8][17]  ( .D(n9), .E(n133), .CP(n274), .Q(
        \Storage[8][17] ) );
  EDFQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(n134), .CP(n254), .Q(
        \Storage[8][16] ) );
  EDFQD1 \Storage_reg[8][15]  ( .D(n1), .E(n134), .CP(ChipClock), .Q(
        \Storage[8][15] ) );
  EDFQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(n133), .CP(n277), .Q(
        \Storage[8][14] ) );
  EDFQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(n132), .CP(n262), .Q(
        \Storage[8][13] ) );
  EDFQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n132), .CP(n245), .Q(
        \Storage[8][12] ) );
  EDFQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(n133), .CP(n244), .Q(
        \Storage[8][11] ) );
  EDFQD1 \Storage_reg[8][10]  ( .D(n19), .E(n134), .CP(n243), .Q(
        \Storage[8][10] ) );
  EDFQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(n134), .CP(n224), .Q(
        \Storage[8][9] ) );
  EDFQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(n133), .CP(n260), .Q(
        \Storage[8][8] ) );
  EDFQD1 \Storage_reg[8][7]  ( .D(n31), .E(n132), .CP(n213), .Q(
        \Storage[8][7] ) );
  EDFQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(n132), .CP(n214), .Q(
        \Storage[8][6] ) );
  EDFQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(n133), .CP(n215), .Q(
        \Storage[8][5] ) );
  EDFQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(n134), .CP(n210), .Q(
        \Storage[8][4] ) );
  EDFQD1 \Storage_reg[8][3]  ( .D(n47), .E(n134), .CP(n211), .Q(
        \Storage[8][3] ) );
  EDFQD1 \Storage_reg[8][2]  ( .D(n52), .E(n133), .CP(n212), .Q(
        \Storage[8][2] ) );
  EDFQD1 \Storage_reg[8][1]  ( .D(n56), .E(n134), .CP(n207), .Q(
        \Storage[8][1] ) );
  EDFQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n132), .CP(n208), .Q(
        \Storage[8][0] ) );
  EDFQD1 \Storage_reg[7][32]  ( .D(n200), .E(n141), .CP(n209), .Q(
        \Storage[7][32] ) );
  EDFQD1 \Storage_reg[7][31]  ( .D(n63), .E(n141), .CP(n229), .Q(
        \Storage[7][31] ) );
  EDFQD1 \Storage_reg[7][30]  ( .D(n61), .E(n142), .CP(n253), .Q(
        \Storage[7][30] ) );
  EDFQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n142), .CP(n223), .Q(
        \Storage[7][29] ) );
  EDFQD1 \Storage_reg[7][28]  ( .D(n53), .E(n141), .CP(n222), .Q(
        \Storage[7][28] ) );
  EDFQD1 \Storage_reg[7][27]  ( .D(n49), .E(n140), .CP(n221), .Q(
        \Storage[7][27] ) );
  EDFQD1 \Storage_reg[7][26]  ( .D(n45), .E(n140), .CP(n220), .Q(
        \Storage[7][26] ) );
  EDFQD1 \Storage_reg[7][25]  ( .D(n41), .E(n141), .CP(n219), .Q(
        \Storage[7][25] ) );
  EDFQD1 \Storage_reg[7][24]  ( .D(n37), .E(n140), .CP(n218), .Q(
        \Storage[7][24] ) );
  EDFQD1 \Storage_reg[7][23]  ( .D(n33), .E(n142), .CP(n217), .Q(
        \Storage[7][23] ) );
  EDFQD1 \Storage_reg[7][22]  ( .D(n29), .E(n141), .CP(n216), .Q(
        \Storage[7][22] ) );
  EDFQD1 \Storage_reg[7][21]  ( .D(n25), .E(n140), .CP(n230), .Q(
        \Storage[7][21] ) );
  EDFQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n142), .CP(n251), .Q(
        \Storage[7][20] ) );
  EDFQD1 \Storage_reg[7][19]  ( .D(n17), .E(n140), .CP(n228), .Q(
        \Storage[7][19] ) );
  EDFQD1 \Storage_reg[7][18]  ( .D(n13), .E(n140), .CP(n233), .Q(
        \Storage[7][18] ) );
  EDFQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n141), .CP(n232), .Q(
        \Storage[7][17] ) );
  EDFQD1 \Storage_reg[7][16]  ( .D(n5), .E(n142), .CP(n231), .Q(
        \Storage[7][16] ) );
  EDFQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n142), .CP(n225), .Q(
        \Storage[7][15] ) );
  EDFQD1 \Storage_reg[7][14]  ( .D(n3), .E(n141), .CP(n226), .Q(
        \Storage[7][14] ) );
  EDFQD1 \Storage_reg[7][13]  ( .D(n7), .E(n140), .CP(n227), .Q(
        \Storage[7][13] ) );
  EDFQD1 \Storage_reg[7][12]  ( .D(n11), .E(n140), .CP(n247), .Q(
        \Storage[7][12] ) );
  EDFQD1 \Storage_reg[7][11]  ( .D(n15), .E(n141), .CP(n246), .Q(
        \Storage[7][11] ) );
  EDFQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n142), .CP(n224), .Q(
        \Storage[7][10] ) );
  EDFQD1 \Storage_reg[7][9]  ( .D(n23), .E(n142), .CP(n233), .Q(
        \Storage[7][9] ) );
  EDFQD1 \Storage_reg[7][8]  ( .D(n27), .E(n141), .CP(n257), .Q(
        \Storage[7][8] ) );
  EDFQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n140), .CP(n261), .Q(
        \Storage[7][7] ) );
  EDFQD1 \Storage_reg[7][6]  ( .D(n35), .E(n140), .CP(n262), .Q(
        \Storage[7][6] ) );
  EDFQD1 \Storage_reg[7][5]  ( .D(n39), .E(n141), .CP(n263), .Q(
        \Storage[7][5] ) );
  EDFQD1 \Storage_reg[7][4]  ( .D(n43), .E(n142), .CP(n273), .Q(
        \Storage[7][4] ) );
  EDFQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n142), .CP(n264), .Q(
        \Storage[7][3] ) );
  EDFQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n141), .CP(n265), .Q(
        \Storage[7][2] ) );
  EDFQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n142), .CP(n266), .Q(
        \Storage[7][1] ) );
  EDFQD1 \Storage_reg[7][0]  ( .D(n59), .E(n140), .CP(n272), .Q(
        \Storage[7][0] ) );
  EDFQD1 \Storage_reg[4][32]  ( .D(n201), .E(n165), .CP(n275), .Q(
        \Storage[4][32] ) );
  EDFQD1 \Storage_reg[4][31]  ( .D(n63), .E(n165), .CP(n267), .Q(
        \Storage[4][31] ) );
  EDFQD1 \Storage_reg[4][30]  ( .D(n61), .E(n166), .CP(n257), .Q(
        \Storage[4][30] ) );
  EDFQD1 \Storage_reg[4][29]  ( .D(n57), .E(n166), .CP(n279), .Q(
        \Storage[4][29] ) );
  EDFQD1 \Storage_reg[4][28]  ( .D(n53), .E(n165), .CP(n274), .Q(
        \Storage[4][28] ) );
  EDFQD1 \Storage_reg[4][27]  ( .D(n49), .E(n164), .CP(n261), .Q(
        \Storage[4][27] ) );
  EDFQD1 \Storage_reg[4][26]  ( .D(n45), .E(n164), .CP(n262), .Q(
        \Storage[4][26] ) );
  EDFQD1 \Storage_reg[4][25]  ( .D(n41), .E(n165), .CP(n263), .Q(
        \Storage[4][25] ) );
  EDFQD1 \Storage_reg[4][24]  ( .D(n37), .E(n164), .CP(n264), .Q(
        \Storage[4][24] ) );
  EDFQD1 \Storage_reg[4][23]  ( .D(n33), .E(n166), .CP(n265), .Q(
        \Storage[4][23] ) );
  EDFQD1 \Storage_reg[4][22]  ( .D(n29), .E(n165), .CP(n266), .Q(
        \Storage[4][22] ) );
  EDFQD1 \Storage_reg[4][21]  ( .D(n25), .E(n164), .CP(n272), .Q(
        \Storage[4][21] ) );
  EDFQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n166), .CP(n270), .Q(
        \Storage[4][20] ) );
  EDFQD1 \Storage_reg[4][19]  ( .D(n17), .E(n164), .CP(n274), .Q(
        \Storage[4][19] ) );
  EDFQD1 \Storage_reg[4][18]  ( .D(n13), .E(n164), .CP(n259), .Q(
        \Storage[4][18] ) );
  EDFQD1 \Storage_reg[4][17]  ( .D(n9), .E(n165), .CP(n260), .Q(
        \Storage[4][17] ) );
  EDFQD1 \Storage_reg[4][16]  ( .D(n5), .E(n166), .CP(n268), .Q(
        \Storage[4][16] ) );
  EDFQD1 \Storage_reg[4][15]  ( .D(n1), .E(n166), .CP(n269), .Q(
        \Storage[4][15] ) );
  EDFQD1 \Storage_reg[4][14]  ( .D(n3), .E(n165), .CP(n265), .Q(
        \Storage[4][14] ) );
  EDFQD1 \Storage_reg[4][13]  ( .D(n7), .E(n164), .CP(n260), .Q(
        \Storage[4][13] ) );
  EDFQD1 \Storage_reg[4][12]  ( .D(n11), .E(n164), .CP(n273), .Q(
        \Storage[4][12] ) );
  EDFQD1 \Storage_reg[4][11]  ( .D(n15), .E(n165), .CP(n241), .Q(
        \Storage[4][11] ) );
  EDFQD1 \Storage_reg[4][10]  ( .D(n19), .E(n166), .CP(n224), .Q(
        \Storage[4][10] ) );
  EDFQD1 \Storage_reg[4][9]  ( .D(n23), .E(n166), .CP(n252), .Q(
        \Storage[4][9] ) );
  EDFQD1 \Storage_reg[4][8]  ( .D(n27), .E(n165), .CP(n260), .Q(
        \Storage[4][8] ) );
  EDFQD1 \Storage_reg[4][7]  ( .D(n31), .E(n164), .CP(n257), .Q(
        \Storage[4][7] ) );
  EDFQD1 \Storage_reg[4][6]  ( .D(n35), .E(n164), .CP(n245), .Q(
        \Storage[4][6] ) );
  EDFQD1 \Storage_reg[4][5]  ( .D(n39), .E(n165), .CP(n229), .Q(
        \Storage[4][5] ) );
  EDFQD1 \Storage_reg[4][4]  ( .D(n43), .E(n166), .CP(n255), .Q(
        \Storage[4][4] ) );
  EDFQD1 \Storage_reg[4][3]  ( .D(n47), .E(n166), .CP(n263), .Q(
        \Storage[4][3] ) );
  EDFQD1 \Storage_reg[4][2]  ( .D(n51), .E(n165), .CP(n254), .Q(
        \Storage[4][2] ) );
  EDFQD1 \Storage_reg[4][1]  ( .D(n55), .E(n166), .CP(n259), .Q(
        \Storage[4][1] ) );
  EDFQD1 \Storage_reg[4][0]  ( .D(n59), .E(n164), .CP(n275), .Q(
        \Storage[4][0] ) );
  EDFQD1 \Storage_reg[3][32]  ( .D(n202), .E(n173), .CP(n277), .Q(
        \Storage[3][32] ) );
  EDFQD1 \Storage_reg[3][31]  ( .D(n64), .E(n173), .CP(n258), .Q(
        \Storage[3][31] ) );
  EDFQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n174), .CP(n228), .Q(
        \Storage[3][30] ) );
  EDFQD1 \Storage_reg[3][29]  ( .D(n57), .E(n174), .CP(n271), .Q(
        \Storage[3][29] ) );
  EDFQD1 \Storage_reg[3][28]  ( .D(n54), .E(n173), .CP(n239), .Q(
        \Storage[3][28] ) );
  EDFQD1 \Storage_reg[3][27]  ( .D(n50), .E(n172), .CP(n252), .Q(
        \Storage[3][27] ) );
  EDFQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n172), .CP(ChipClock), .Q(
        \Storage[3][26] ) );
  EDFQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n173), .CP(n278), .Q(
        \Storage[3][25] ) );
  EDFQD1 \Storage_reg[3][24]  ( .D(n38), .E(n172), .CP(n276), .Q(
        \Storage[3][24] ) );
  EDFQD1 \Storage_reg[3][23]  ( .D(n34), .E(n174), .CP(n255), .Q(
        \Storage[3][23] ) );
  EDFQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n173), .CP(n256), .Q(
        \Storage[3][22] ) );
  EDFQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n172), .CP(n257), .Q(
        \Storage[3][21] ) );
  EDFQD1 \Storage_reg[3][20]  ( .D(n21), .E(n174), .CP(n261), .Q(
        \Storage[3][20] ) );
  EDFQD1 \Storage_reg[3][19]  ( .D(n18), .E(n172), .CP(n270), .Q(
        \Storage[3][19] ) );
  EDFQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n172), .CP(n255), .Q(
        \Storage[3][18] ) );
  EDFQD1 \Storage_reg[3][17]  ( .D(n9), .E(n173), .CP(n267), .Q(
        \Storage[3][17] ) );
  EDFQD1 \Storage_reg[3][16]  ( .D(n6), .E(n174), .CP(n268), .Q(
        \Storage[3][16] ) );
  EDFQD1 \Storage_reg[3][15]  ( .D(n1), .E(n174), .CP(n269), .Q(
        \Storage[3][15] ) );
  EDFQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n173), .CP(n273), .Q(
        \Storage[3][14] ) );
  EDFQD1 \Storage_reg[3][13]  ( .D(n8), .E(n172), .CP(n264), .Q(
        \Storage[3][13] ) );
  EDFQD1 \Storage_reg[3][12]  ( .D(n12), .E(n172), .CP(n265), .Q(
        \Storage[3][12] ) );
  EDFQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n173), .CP(n266), .Q(
        \Storage[3][11] ) );
  EDFQD1 \Storage_reg[3][10]  ( .D(n19), .E(n174), .CP(n263), .Q(
        \Storage[3][10] ) );
  EDFQD1 \Storage_reg[3][9]  ( .D(n24), .E(n174), .CP(n266), .Q(
        \Storage[3][9] ) );
  EDFQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n173), .CP(n256), .Q(
        \Storage[3][8] ) );
  EDFQD1 \Storage_reg[3][7]  ( .D(n31), .E(n172), .CP(n271), .Q(
        \Storage[3][7] ) );
  EDFQD1 \Storage_reg[3][6]  ( .D(n36), .E(n172), .CP(n256), .Q(
        \Storage[3][6] ) );
  EDFQD1 \Storage_reg[3][5]  ( .D(n40), .E(n173), .CP(ChipClock), .Q(
        \Storage[3][5] ) );
  EDFQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n174), .CP(n238), .Q(
        \Storage[3][4] ) );
  EDFQD1 \Storage_reg[3][3]  ( .D(n47), .E(n174), .CP(n223), .Q(
        \Storage[3][3] ) );
  EDFQD1 \Storage_reg[3][2]  ( .D(n52), .E(n173), .CP(n278), .Q(
        \Storage[3][2] ) );
  EDFQD1 \Storage_reg[3][1]  ( .D(n55), .E(n174), .CP(n276), .Q(
        \Storage[3][1] ) );
  EDFQD1 \Storage_reg[3][0]  ( .D(n60), .E(n172), .CP(n255), .Q(
        \Storage[3][0] ) );
  EDFQD1 \Storage_reg[0][32]  ( .D(n201), .E(n197), .CP(n255), .Q(
        \Storage[0][32] ) );
  EDFQD1 \Storage_reg[0][31]  ( .D(n64), .E(n197), .CP(n263), .Q(
        \Storage[0][31] ) );
  EDFQD1 \Storage_reg[0][30]  ( .D(n62), .E(n198), .CP(n270), .Q(
        \Storage[0][30] ) );
  EDFQD1 \Storage_reg[0][29]  ( .D(n57), .E(n198), .CP(n275), .Q(
        \Storage[0][29] ) );
  EDFQD1 \Storage_reg[0][28]  ( .D(n54), .E(n197), .CP(n258), .Q(
        \Storage[0][28] ) );
  EDFQD1 \Storage_reg[0][27]  ( .D(n50), .E(n196), .CP(n259), .Q(
        \Storage[0][27] ) );
  EDFQD1 \Storage_reg[0][26]  ( .D(n46), .E(n196), .CP(n260), .Q(
        \Storage[0][26] ) );
  EDFQD1 \Storage_reg[0][25]  ( .D(n42), .E(n197), .CP(n257), .Q(
        \Storage[0][25] ) );
  EDFQD1 \Storage_reg[0][24]  ( .D(n38), .E(n196), .CP(n279), .Q(
        \Storage[0][24] ) );
  EDFQD1 \Storage_reg[0][23]  ( .D(n34), .E(n198), .CP(n274), .Q(
        \Storage[0][23] ) );
  EDFQD1 \Storage_reg[0][22]  ( .D(n30), .E(n197), .CP(n261), .Q(
        \Storage[0][22] ) );
  EDFQD1 \Storage_reg[0][21]  ( .D(n26), .E(n196), .CP(n262), .Q(
        \Storage[0][21] ) );
  EDFQD1 \Storage_reg[0][20]  ( .D(n22), .E(n198), .CP(n247), .Q(
        \Storage[0][20] ) );
  EDFQD1 \Storage_reg[0][19]  ( .D(n18), .E(n196), .CP(n258), .Q(
        \Storage[0][19] ) );
  EDFQD1 \Storage_reg[0][18]  ( .D(n14), .E(n196), .CP(n273), .Q(
        \Storage[0][18] ) );
  EDFQD1 \Storage_reg[0][17]  ( .D(n9), .E(n197), .CP(n264), .Q(
        \Storage[0][17] ) );
  EDFQD1 \Storage_reg[0][16]  ( .D(n6), .E(n198), .CP(n265), .Q(
        \Storage[0][16] ) );
  EDFQD1 \Storage_reg[0][15]  ( .D(n1), .E(n198), .CP(n266), .Q(
        \Storage[0][15] ) );
  EDFQD1 \Storage_reg[0][14]  ( .D(n4), .E(n197), .CP(n272), .Q(
        \Storage[0][14] ) );
  EDFQD1 \Storage_reg[0][13]  ( .D(n8), .E(n196), .CP(n267), .Q(
        \Storage[0][13] ) );
  EDFQD1 \Storage_reg[0][12]  ( .D(n12), .E(n196), .CP(n268), .Q(
        \Storage[0][12] ) );
  EDFQD1 \Storage_reg[0][11]  ( .D(n16), .E(n197), .CP(n269), .Q(
        \Storage[0][11] ) );
  EDFQD1 \Storage_reg[0][10]  ( .D(n19), .E(n198), .CP(n276), .Q(
        \Storage[0][10] ) );
  EDFQD1 \Storage_reg[0][9]  ( .D(n24), .E(n198), .CP(ChipClock), .Q(
        \Storage[0][9] ) );
  EDFQD1 \Storage_reg[0][8]  ( .D(n28), .E(n197), .CP(n275), .Q(
        \Storage[0][8] ) );
  EDFQD1 \Storage_reg[0][7]  ( .D(n31), .E(n196), .CP(n236), .Q(
        \Storage[0][7] ) );
  EDFQD1 \Storage_reg[0][6]  ( .D(n36), .E(n196), .CP(n217), .Q(
        \Storage[0][6] ) );
  EDFQD1 \Storage_reg[0][5]  ( .D(n40), .E(n197), .CP(n262), .Q(
        \Storage[0][5] ) );
  EDFQD1 \Storage_reg[0][4]  ( .D(n44), .E(n198), .CP(n244), .Q(
        \Storage[0][4] ) );
  EDFQD1 \Storage_reg[0][3]  ( .D(n47), .E(n198), .CP(n258), .Q(
        \Storage[0][3] ) );
  EDFQD1 \Storage_reg[0][2]  ( .D(n52), .E(n197), .CP(n279), .Q(
        \Storage[0][2] ) );
  EDFQD1 \Storage_reg[0][1]  ( .D(n56), .E(n198), .CP(n277), .Q(
        \Storage[0][1] ) );
  EDFQD1 \Storage_reg[0][0]  ( .D(n60), .E(n196), .CP(n249), .Q(
        \Storage[0][0] ) );
  EDFQD1 \Storage_reg[31][32]  ( .D(n200), .E(n193), .CP(n277), .Q(
        \Storage[31][32] ) );
  EDFQD1 \Storage_reg[31][31]  ( .D(n63), .E(n193), .CP(n253), .Q(
        \Storage[31][31] ) );
  EDFQD1 \Storage_reg[31][30]  ( .D(n62), .E(n194), .CP(n253), .Q(
        \Storage[31][30] ) );
  EDFQD1 \Storage_reg[31][29]  ( .D(n58), .E(n194), .CP(n253), .Q(
        \Storage[31][29] ) );
  EDFQD1 \Storage_reg[31][28]  ( .D(n53), .E(n193), .CP(n253), .Q(
        \Storage[31][28] ) );
  EDFQD1 \Storage_reg[31][27]  ( .D(n49), .E(n192), .CP(n253), .Q(
        \Storage[31][27] ) );
  EDFQD1 \Storage_reg[31][26]  ( .D(n46), .E(n192), .CP(n253), .Q(
        \Storage[31][26] ) );
  EDFQD1 \Storage_reg[31][25]  ( .D(n42), .E(n193), .CP(n253), .Q(
        \Storage[31][25] ) );
  EDFQD1 \Storage_reg[31][24]  ( .D(n37), .E(n192), .CP(n253), .Q(
        \Storage[31][24] ) );
  EDFQD1 \Storage_reg[31][23]  ( .D(n33), .E(n194), .CP(n253), .Q(
        \Storage[31][23] ) );
  EDFQD1 \Storage_reg[31][22]  ( .D(n30), .E(n193), .CP(n253), .Q(
        \Storage[31][22] ) );
  EDFQD1 \Storage_reg[31][21]  ( .D(n26), .E(n192), .CP(n253), .Q(
        \Storage[31][21] ) );
  EDFQD1 \Storage_reg[31][20]  ( .D(n22), .E(n194), .CP(n252), .Q(
        \Storage[31][20] ) );
  EDFQD1 \Storage_reg[31][19]  ( .D(n17), .E(n192), .CP(n252), .Q(
        \Storage[31][19] ) );
  EDFQD1 \Storage_reg[31][18]  ( .D(n14), .E(n192), .CP(n252), .Q(
        \Storage[31][18] ) );
  EDFQD1 \Storage_reg[31][17]  ( .D(n10), .E(n193), .CP(n252), .Q(
        \Storage[31][17] ) );
  EDFQD1 \Storage_reg[31][16]  ( .D(n5), .E(n194), .CP(n252), .Q(
        \Storage[31][16] ) );
  EDFQD1 \Storage_reg[31][15]  ( .D(n2), .E(n194), .CP(n252), .Q(
        \Storage[31][15] ) );
  EDFQD1 \Storage_reg[31][14]  ( .D(n4), .E(n193), .CP(n252), .Q(
        \Storage[31][14] ) );
  EDFQD1 \Storage_reg[31][13]  ( .D(n7), .E(n192), .CP(n252), .Q(
        \Storage[31][13] ) );
  EDFQD1 \Storage_reg[31][12]  ( .D(n11), .E(n192), .CP(n252), .Q(
        \Storage[31][12] ) );
  EDFQD1 \Storage_reg[31][11]  ( .D(n16), .E(n193), .CP(n252), .Q(
        \Storage[31][11] ) );
  EDFQD1 \Storage_reg[31][10]  ( .D(n20), .E(n194), .CP(n252), .Q(
        \Storage[31][10] ) );
  EDFQD1 \Storage_reg[31][9]  ( .D(n23), .E(n194), .CP(n251), .Q(
        \Storage[31][9] ) );
  EDFQD1 \Storage_reg[31][8]  ( .D(n28), .E(n193), .CP(n251), .Q(
        \Storage[31][8] ) );
  EDFQD1 \Storage_reg[31][7]  ( .D(n32), .E(n192), .CP(n251), .Q(
        \Storage[31][7] ) );
  EDFQD1 \Storage_reg[31][6]  ( .D(n35), .E(n192), .CP(n251), .Q(
        \Storage[31][6] ) );
  EDFQD1 \Storage_reg[31][5]  ( .D(n39), .E(n193), .CP(n251), .Q(
        \Storage[31][5] ) );
  EDFQD1 \Storage_reg[31][4]  ( .D(n44), .E(n194), .CP(n251), .Q(
        \Storage[31][4] ) );
  EDFQD1 \Storage_reg[31][3]  ( .D(n48), .E(n194), .CP(n251), .Q(
        \Storage[31][3] ) );
  EDFQD1 \Storage_reg[31][2]  ( .D(n51), .E(n193), .CP(n251), .Q(
        \Storage[31][2] ) );
  EDFQD1 \Storage_reg[31][1]  ( .D(n56), .E(n194), .CP(n251), .Q(
        \Storage[31][1] ) );
  EDFQD1 \Storage_reg[31][0]  ( .D(n59), .E(n192), .CP(n251), .Q(
        \Storage[31][0] ) );
  EDFQD1 DreadyReg_reg ( .D(Read), .E(ChipEna), .CP(n277), .Q(DreadyReg) );
  EDFQD1 ParityReg_reg ( .D(N84), .E(N2262), .CP(n273), .Q(ParityErr) );
  EDFQD1 \DataOreg_reg[31]  ( .D(N50), .E(N2262), .CP(n254), .Q(DataOreg[31])
         );
  EDFQD1 \DataOreg_reg[30]  ( .D(N51), .E(N2262), .CP(n278), .Q(DataOreg[30])
         );
  EDFQD1 \DataOreg_reg[29]  ( .D(N52), .E(N2262), .CP(n271), .Q(DataOreg[29])
         );
  EDFQD1 \DataOreg_reg[28]  ( .D(N53), .E(N2262), .CP(n276), .Q(DataOreg[28])
         );
  EDFQD1 \DataOreg_reg[27]  ( .D(N54), .E(N2262), .CP(n254), .Q(DataOreg[27])
         );
  EDFQD1 \DataOreg_reg[5]  ( .D(N76), .E(N2262), .CP(n259), .Q(DataOreg[5]) );
  EDFQD1 \DataOreg_reg[4]  ( .D(N77), .E(N2262), .CP(n278), .Q(DataOreg[4]) );
  EDFQD1 \DataOreg_reg[3]  ( .D(N78), .E(N2262), .CP(n226), .Q(DataOreg[3]) );
  EDFQD1 \DataOreg_reg[2]  ( .D(N79), .E(N2262), .CP(n256), .Q(DataOreg[2]) );
  EDFQD1 \DataOreg_reg[1]  ( .D(N80), .E(N2262), .CP(n230), .Q(DataOreg[1]) );
  EDFQD1 \DataOreg_reg[0]  ( .D(N81), .E(N2262), .CP(n279), .Q(DataOreg[0]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOreg[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOreg[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOreg[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOreg[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOreg[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOreg[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOreg[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOreg[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOreg[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOreg[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOreg[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOreg[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOreg[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOreg[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOreg[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOreg[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOreg[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOreg[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOreg[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOreg[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOreg[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOreg[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOreg[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOreg[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOreg[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOreg[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOreg[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOreg[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOreg[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOreg[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOreg[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOreg[16]), .OE(ChipEna), .Z(DataO[16]) );
  EDFQD1 \DataOreg_reg[26]  ( .D(N55), .E(N2262), .CP(n241), .Q(DataOreg[26])
         );
  EDFQD1 \DataOreg_reg[7]  ( .D(N74), .E(N2262), .CP(n274), .Q(DataOreg[7]) );
  EDFQD1 \DataOreg_reg[6]  ( .D(N75), .E(N2262), .CP(n272), .Q(DataOreg[6]) );
  EDFQD1 \DataOreg_reg[23]  ( .D(N58), .E(N2262), .CP(n270), .Q(DataOreg[23])
         );
  EDFQD1 \DataOreg_reg[24]  ( .D(N57), .E(N2262), .CP(n257), .Q(DataOreg[24])
         );
  EDFQD1 \DataOreg_reg[25]  ( .D(N56), .E(N2262), .CP(n262), .Q(DataOreg[25])
         );
  EDFQD1 \DataOreg_reg[11]  ( .D(N70), .E(N2262), .CP(n275), .Q(DataOreg[11])
         );
  EDFQD1 \DataOreg_reg[10]  ( .D(N71), .E(N2262), .CP(n260), .Q(DataOreg[10])
         );
  EDFQD1 \DataOreg_reg[9]  ( .D(N72), .E(N2262), .CP(n258), .Q(DataOreg[9]) );
  EDFQD1 \DataOreg_reg[8]  ( .D(N73), .E(N2262), .CP(n254), .Q(DataOreg[8]) );
  EDFQD1 \DataOreg_reg[19]  ( .D(N62), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[19]) );
  EDFQD1 \DataOreg_reg[20]  ( .D(N61), .E(N2262), .CP(n254), .Q(DataOreg[20])
         );
  EDFQD1 \DataOreg_reg[21]  ( .D(N60), .E(N2262), .CP(n279), .Q(DataOreg[21])
         );
  EDFQD1 \DataOreg_reg[22]  ( .D(N59), .E(N2262), .CP(n277), .Q(DataOreg[22])
         );
  EDFQD1 \DataOreg_reg[15]  ( .D(N66), .E(N2262), .CP(n276), .Q(DataOreg[15])
         );
  EDFQD1 \DataOreg_reg[14]  ( .D(N67), .E(N2262), .CP(n278), .Q(DataOreg[14])
         );
  EDFQD1 \DataOreg_reg[13]  ( .D(N68), .E(N2262), .CP(n216), .Q(DataOreg[13])
         );
  EDFQD1 \DataOreg_reg[18]  ( .D(N63), .E(N2262), .CP(n275), .Q(DataOreg[18])
         );
  EDFQD1 \DataOreg_reg[12]  ( .D(N69), .E(N2262), .CP(n257), .Q(DataOreg[12])
         );
  EDFQD1 \DataOreg_reg[16]  ( .D(N65), .E(N2262), .CP(n256), .Q(DataOreg[16])
         );
  EDFQD1 \DataOreg_reg[17]  ( .D(N64), .E(N2262), .CP(n255), .Q(DataOreg[17])
         );
  BUFFD0 U2 ( .I(DataI[15]), .Z(n1) );
  BUFFD0 U3 ( .I(DataI[15]), .Z(n2) );
  BUFFD0 U4 ( .I(DataI[14]), .Z(n4) );
  BUFFD0 U5 ( .I(DataI[14]), .Z(n3) );
  BUFFD0 U6 ( .I(DataI[16]), .Z(n6) );
  BUFFD0 U7 ( .I(DataI[16]), .Z(n5) );
  BUFFD0 U8 ( .I(DataI[13]), .Z(n8) );
  BUFFD0 U9 ( .I(DataI[13]), .Z(n7) );
  BUFFD0 U10 ( .I(DataI[17]), .Z(n9) );
  BUFFD0 U11 ( .I(DataI[17]), .Z(n10) );
  BUFFD0 U12 ( .I(DataI[12]), .Z(n12) );
  BUFFD0 U13 ( .I(DataI[12]), .Z(n11) );
  BUFFD0 U14 ( .I(DataI[18]), .Z(n14) );
  BUFFD0 U15 ( .I(DataI[18]), .Z(n13) );
  BUFFD0 U16 ( .I(DataI[11]), .Z(n16) );
  BUFFD0 U17 ( .I(DataI[11]), .Z(n15) );
  BUFFD0 U18 ( .I(DataI[19]), .Z(n18) );
  BUFFD0 U19 ( .I(DataI[19]), .Z(n17) );
  BUFFD0 U20 ( .I(DataI[10]), .Z(n19) );
  BUFFD0 U21 ( .I(DataI[10]), .Z(n20) );
  BUFFD0 U22 ( .I(DataI[20]), .Z(n21) );
  BUFFD0 U23 ( .I(DataI[20]), .Z(n22) );
  BUFFD0 U24 ( .I(DataI[9]), .Z(n24) );
  BUFFD0 U25 ( .I(DataI[9]), .Z(n23) );
  BUFFD0 U26 ( .I(DataI[21]), .Z(n26) );
  BUFFD0 U27 ( .I(DataI[21]), .Z(n25) );
  BUFFD0 U28 ( .I(DataI[8]), .Z(n28) );
  BUFFD0 U29 ( .I(DataI[8]), .Z(n27) );
  BUFFD0 U30 ( .I(DataI[22]), .Z(n30) );
  BUFFD0 U31 ( .I(DataI[22]), .Z(n29) );
  BUFFD0 U32 ( .I(DataI[7]), .Z(n31) );
  BUFFD0 U33 ( .I(DataI[7]), .Z(n32) );
  BUFFD0 U34 ( .I(DataI[23]), .Z(n34) );
  BUFFD0 U35 ( .I(DataI[23]), .Z(n33) );
  BUFFD0 U36 ( .I(DataI[6]), .Z(n36) );
  BUFFD0 U37 ( .I(DataI[6]), .Z(n35) );
  BUFFD0 U38 ( .I(DataI[24]), .Z(n38) );
  BUFFD0 U39 ( .I(DataI[24]), .Z(n37) );
  BUFFD0 U40 ( .I(DataI[5]), .Z(n40) );
  BUFFD0 U41 ( .I(DataI[5]), .Z(n39) );
  BUFFD0 U42 ( .I(DataI[25]), .Z(n42) );
  BUFFD0 U43 ( .I(DataI[25]), .Z(n41) );
  BUFFD0 U44 ( .I(DataI[4]), .Z(n44) );
  BUFFD0 U45 ( .I(DataI[4]), .Z(n43) );
  BUFFD0 U46 ( .I(DataI[26]), .Z(n46) );
  BUFFD0 U47 ( .I(DataI[26]), .Z(n45) );
  BUFFD0 U48 ( .I(DataI[3]), .Z(n47) );
  BUFFD0 U49 ( .I(DataI[3]), .Z(n48) );
  BUFFD0 U50 ( .I(DataI[27]), .Z(n50) );
  BUFFD0 U51 ( .I(DataI[27]), .Z(n49) );
  BUFFD0 U52 ( .I(DataI[2]), .Z(n52) );
  BUFFD0 U53 ( .I(DataI[2]), .Z(n51) );
  BUFFD0 U54 ( .I(DataI[28]), .Z(n54) );
  BUFFD0 U55 ( .I(DataI[28]), .Z(n53) );
  BUFFD0 U56 ( .I(DataI[1]), .Z(n56) );
  BUFFD0 U57 ( .I(DataI[1]), .Z(n55) );
  BUFFD0 U58 ( .I(DataI[29]), .Z(n57) );
  BUFFD0 U59 ( .I(DataI[29]), .Z(n58) );
  BUFFD0 U60 ( .I(DataI[0]), .Z(n60) );
  BUFFD0 U61 ( .I(DataI[0]), .Z(n59) );
  BUFFD0 U62 ( .I(DataI[30]), .Z(n62) );
  BUFFD0 U63 ( .I(DataI[30]), .Z(n61) );
  BUFFD0 U64 ( .I(DataI[31]), .Z(n64) );
  BUFFD0 U65 ( .I(DataI[31]), .Z(n63) );
  BUFFD0 U66 ( .I(N47), .Z(n66) );
  BUFFD0 U67 ( .I(N47), .Z(n65) );
  BUFFD1 U68 ( .I(N46), .Z(n67) );
  BUFFD1 U69 ( .I(N46), .Z(n70) );
  BUFFD1 U70 ( .I(N46), .Z(n68) );
  BUFFD1 U71 ( .I(N46), .Z(n69) );
  OR2D0 U72 ( .A1(n793), .A2(n795), .Z(n71) );
  INVD0 U73 ( .I(n71), .ZN(n72) );
  INVD0 U74 ( .I(n71), .ZN(n74) );
  INVD0 U75 ( .I(n71), .ZN(n73) );
  OR2D0 U76 ( .A1(n786), .A2(n797), .Z(n75) );
  INVD0 U77 ( .I(n75), .ZN(n76) );
  INVD0 U78 ( .I(n75), .ZN(n78) );
  INVD0 U79 ( .I(n75), .ZN(n77) );
  OR2D0 U80 ( .A1(n792), .A2(n795), .Z(n79) );
  INVD0 U81 ( .I(n79), .ZN(n80) );
  INVD0 U82 ( .I(n79), .ZN(n82) );
  INVD0 U83 ( .I(n79), .ZN(n81) );
  OR2D0 U84 ( .A1(n787), .A2(n797), .Z(n83) );
  INVD0 U85 ( .I(n83), .ZN(n84) );
  INVD0 U86 ( .I(n83), .ZN(n86) );
  INVD0 U87 ( .I(n83), .ZN(n85) );
  OR2D0 U88 ( .A1(n791), .A2(n795), .Z(n87) );
  INVD0 U89 ( .I(n87), .ZN(n88) );
  INVD0 U90 ( .I(n87), .ZN(n90) );
  INVD0 U91 ( .I(n87), .ZN(n89) );
  OR2D0 U92 ( .A1(n788), .A2(n797), .Z(n91) );
  INVD0 U93 ( .I(n91), .ZN(n92) );
  INVD0 U94 ( .I(n91), .ZN(n94) );
  INVD0 U95 ( .I(n91), .ZN(n93) );
  OR2D0 U96 ( .A1(n790), .A2(n795), .Z(n95) );
  INVD0 U97 ( .I(n95), .ZN(n96) );
  INVD0 U98 ( .I(n95), .ZN(n98) );
  INVD0 U99 ( .I(n95), .ZN(n97) );
  OR2D0 U100 ( .A1(n789), .A2(n797), .Z(n99) );
  INVD0 U101 ( .I(n99), .ZN(n100) );
  INVD0 U102 ( .I(n99), .ZN(n102) );
  INVD0 U103 ( .I(n99), .ZN(n101) );
  OR2D0 U104 ( .A1(n789), .A2(n795), .Z(n103) );
  INVD0 U105 ( .I(n103), .ZN(n104) );
  INVD0 U106 ( .I(n103), .ZN(n106) );
  INVD0 U107 ( .I(n103), .ZN(n105) );
  OR2D0 U108 ( .A1(n790), .A2(n797), .Z(n107) );
  INVD0 U109 ( .I(n107), .ZN(n108) );
  INVD0 U110 ( .I(n107), .ZN(n110) );
  INVD0 U111 ( .I(n107), .ZN(n109) );
  OR2D0 U112 ( .A1(n788), .A2(n795), .Z(n111) );
  INVD0 U113 ( .I(n111), .ZN(n112) );
  INVD0 U114 ( .I(n111), .ZN(n114) );
  INVD0 U115 ( .I(n111), .ZN(n113) );
  OR2D0 U116 ( .A1(n791), .A2(n797), .Z(n115) );
  INVD0 U117 ( .I(n115), .ZN(n116) );
  INVD0 U118 ( .I(n115), .ZN(n118) );
  INVD0 U119 ( .I(n115), .ZN(n117) );
  OR2D0 U120 ( .A1(n787), .A2(n795), .Z(n119) );
  INVD0 U121 ( .I(n119), .ZN(n120) );
  INVD0 U122 ( .I(n119), .ZN(n122) );
  INVD0 U123 ( .I(n119), .ZN(n121) );
  OR2D0 U124 ( .A1(n792), .A2(n797), .Z(n123) );
  INVD0 U125 ( .I(n123), .ZN(n124) );
  INVD0 U126 ( .I(n123), .ZN(n126) );
  INVD0 U127 ( .I(n123), .ZN(n125) );
  OR2D0 U128 ( .A1(n786), .A2(n795), .Z(n127) );
  INVD0 U129 ( .I(n127), .ZN(n128) );
  INVD0 U130 ( .I(n127), .ZN(n130) );
  INVD0 U131 ( .I(n127), .ZN(n129) );
  OR2D0 U132 ( .A1(n793), .A2(n797), .Z(n131) );
  INVD0 U133 ( .I(n131), .ZN(n132) );
  INVD0 U134 ( .I(n131), .ZN(n134) );
  INVD0 U135 ( .I(n131), .ZN(n133) );
  OR2D0 U136 ( .A1(n785), .A2(n793), .Z(n135) );
  INVD0 U137 ( .I(n135), .ZN(n136) );
  INVD0 U138 ( .I(n135), .ZN(n138) );
  INVD0 U139 ( .I(n135), .ZN(n137) );
  OR2D0 U140 ( .A1(n786), .A2(n799), .Z(n139) );
  INVD0 U141 ( .I(n139), .ZN(n140) );
  INVD0 U142 ( .I(n139), .ZN(n142) );
  INVD0 U143 ( .I(n139), .ZN(n141) );
  OR2D0 U144 ( .A1(n785), .A2(n792), .Z(n143) );
  INVD0 U145 ( .I(n143), .ZN(n144) );
  INVD0 U146 ( .I(n143), .ZN(n146) );
  INVD0 U147 ( .I(n143), .ZN(n145) );
  OR2D0 U148 ( .A1(n787), .A2(n799), .Z(n147) );
  INVD0 U149 ( .I(n147), .ZN(n148) );
  INVD0 U150 ( .I(n147), .ZN(n150) );
  INVD0 U151 ( .I(n147), .ZN(n149) );
  OR2D0 U152 ( .A1(n785), .A2(n791), .Z(n151) );
  INVD0 U153 ( .I(n151), .ZN(n152) );
  INVD0 U154 ( .I(n151), .ZN(n154) );
  INVD0 U155 ( .I(n151), .ZN(n153) );
  OR2D0 U156 ( .A1(n788), .A2(n799), .Z(n155) );
  INVD0 U157 ( .I(n155), .ZN(n156) );
  INVD0 U158 ( .I(n155), .ZN(n158) );
  INVD0 U159 ( .I(n155), .ZN(n157) );
  OR2D0 U160 ( .A1(n785), .A2(n790), .Z(n159) );
  INVD0 U161 ( .I(n159), .ZN(n160) );
  INVD0 U162 ( .I(n159), .ZN(n162) );
  INVD0 U163 ( .I(n159), .ZN(n161) );
  OR2D0 U164 ( .A1(n789), .A2(n799), .Z(n163) );
  INVD0 U165 ( .I(n163), .ZN(n164) );
  INVD0 U166 ( .I(n163), .ZN(n166) );
  INVD0 U167 ( .I(n163), .ZN(n165) );
  OR2D0 U168 ( .A1(n785), .A2(n789), .Z(n167) );
  INVD0 U169 ( .I(n167), .ZN(n168) );
  INVD0 U170 ( .I(n167), .ZN(n170) );
  INVD0 U171 ( .I(n167), .ZN(n169) );
  OR2D0 U172 ( .A1(n790), .A2(n799), .Z(n171) );
  INVD0 U173 ( .I(n171), .ZN(n172) );
  INVD0 U174 ( .I(n171), .ZN(n174) );
  INVD0 U175 ( .I(n171), .ZN(n173) );
  OR2D0 U176 ( .A1(n785), .A2(n788), .Z(n175) );
  INVD0 U177 ( .I(n175), .ZN(n176) );
  INVD0 U178 ( .I(n175), .ZN(n178) );
  INVD0 U179 ( .I(n175), .ZN(n177) );
  OR2D0 U180 ( .A1(n791), .A2(n799), .Z(n179) );
  INVD0 U181 ( .I(n179), .ZN(n180) );
  INVD0 U182 ( .I(n179), .ZN(n182) );
  INVD0 U183 ( .I(n179), .ZN(n181) );
  OR2D0 U184 ( .A1(n785), .A2(n787), .Z(n183) );
  INVD0 U185 ( .I(n183), .ZN(n184) );
  INVD0 U186 ( .I(n183), .ZN(n186) );
  INVD0 U187 ( .I(n183), .ZN(n185) );
  OR2D0 U188 ( .A1(n792), .A2(n799), .Z(n187) );
  INVD0 U189 ( .I(n187), .ZN(n188) );
  INVD0 U190 ( .I(n187), .ZN(n190) );
  INVD0 U191 ( .I(n187), .ZN(n189) );
  OR2D0 U192 ( .A1(n785), .A2(n786), .Z(n191) );
  INVD0 U193 ( .I(n191), .ZN(n192) );
  INVD0 U194 ( .I(n191), .ZN(n194) );
  INVD0 U195 ( .I(n191), .ZN(n193) );
  OR2D0 U196 ( .A1(n793), .A2(n799), .Z(n195) );
  INVD0 U197 ( .I(n195), .ZN(n196) );
  INVD0 U198 ( .I(n195), .ZN(n198) );
  INVD0 U199 ( .I(n195), .ZN(n197) );
  ND3D1 U200 ( .A1(n794), .A2(n796), .A3(n66), .ZN(n795) );
  ND3D1 U201 ( .A1(n794), .A2(n798), .A3(n70), .ZN(n797) );
  ND3D1 U202 ( .A1(n796), .A2(n798), .A3(n794), .ZN(n799) );
  ND3D1 U203 ( .A1(n68), .A2(n794), .A3(N47), .ZN(n785) );
  INR2XD2 U204 ( .A1(ChipEna), .B1(n784), .ZN(N2262) );
  XNR3D0 U205 ( .A1(n52), .A2(n55), .A3(n760), .ZN(n199) );
  INVD1 U206 ( .I(n199), .ZN(n200) );
  INVD1 U207 ( .I(n199), .ZN(n202) );
  INVD1 U208 ( .I(n199), .ZN(n201) );
  BUFFD1 U209 ( .I(n271), .Z(n203) );
  BUFFD1 U210 ( .I(n271), .Z(n204) );
  BUFFD1 U211 ( .I(n271), .Z(n205) );
  BUFFD1 U212 ( .I(n270), .Z(n206) );
  BUFFD1 U213 ( .I(n269), .Z(n207) );
  BUFFD1 U214 ( .I(n269), .Z(n208) );
  BUFFD1 U215 ( .I(n269), .Z(n209) );
  BUFFD1 U216 ( .I(n268), .Z(n210) );
  BUFFD1 U217 ( .I(n268), .Z(n211) );
  BUFFD1 U218 ( .I(n268), .Z(n212) );
  BUFFD1 U219 ( .I(n267), .Z(n213) );
  BUFFD1 U220 ( .I(n267), .Z(n214) );
  BUFFD1 U221 ( .I(n267), .Z(n215) );
  BUFFD1 U222 ( .I(n266), .Z(n216) );
  BUFFD1 U223 ( .I(n266), .Z(n217) );
  BUFFD1 U224 ( .I(n266), .Z(n218) );
  BUFFD1 U225 ( .I(n265), .Z(n219) );
  BUFFD1 U226 ( .I(n265), .Z(n220) );
  BUFFD1 U227 ( .I(n265), .Z(n221) );
  BUFFD1 U228 ( .I(n264), .Z(n222) );
  BUFFD1 U229 ( .I(n264), .Z(n223) );
  BUFFD1 U230 ( .I(n264), .Z(n224) );
  BUFFD1 U231 ( .I(n263), .Z(n225) );
  BUFFD1 U232 ( .I(n263), .Z(n226) );
  BUFFD1 U233 ( .I(n263), .Z(n227) );
  BUFFD1 U234 ( .I(n262), .Z(n228) );
  BUFFD1 U235 ( .I(n262), .Z(n229) );
  BUFFD1 U236 ( .I(n262), .Z(n230) );
  BUFFD1 U237 ( .I(n261), .Z(n231) );
  BUFFD1 U238 ( .I(n261), .Z(n232) );
  BUFFD1 U239 ( .I(n261), .Z(n233) );
  BUFFD1 U240 ( .I(n260), .Z(n234) );
  BUFFD1 U241 ( .I(n260), .Z(n235) );
  BUFFD1 U242 ( .I(n260), .Z(n236) );
  BUFFD1 U243 ( .I(n259), .Z(n237) );
  BUFFD1 U244 ( .I(n259), .Z(n238) );
  BUFFD1 U245 ( .I(n259), .Z(n239) );
  BUFFD1 U246 ( .I(n258), .Z(n240) );
  BUFFD1 U247 ( .I(n258), .Z(n241) );
  BUFFD1 U248 ( .I(n258), .Z(n242) );
  BUFFD1 U249 ( .I(n257), .Z(n243) );
  BUFFD1 U250 ( .I(n257), .Z(n244) );
  BUFFD1 U251 ( .I(n257), .Z(n245) );
  BUFFD1 U252 ( .I(n256), .Z(n246) );
  BUFFD1 U253 ( .I(n256), .Z(n247) );
  BUFFD1 U254 ( .I(n256), .Z(n248) );
  BUFFD1 U255 ( .I(n255), .Z(n249) );
  BUFFD1 U256 ( .I(n255), .Z(n250) );
  BUFFD1 U257 ( .I(n255), .Z(n251) );
  INVD1 U258 ( .I(n301), .ZN(n289) );
  INVD1 U259 ( .I(n301), .ZN(n290) );
  INVD1 U260 ( .I(n300), .ZN(n291) );
  INVD1 U261 ( .I(n300), .ZN(n292) );
  INVD1 U262 ( .I(n300), .ZN(n293) );
  INVD1 U263 ( .I(n300), .ZN(n294) );
  INVD1 U264 ( .I(n301), .ZN(n295) );
  INVD1 U265 ( .I(n301), .ZN(n288) );
  INVD1 U266 ( .I(n301), .ZN(n287) );
  INVD1 U267 ( .I(n301), .ZN(n286) );
  INVD1 U268 ( .I(n300), .ZN(n285) );
  INVD1 U269 ( .I(n300), .ZN(n284) );
  INVD1 U270 ( .I(n300), .ZN(n283) );
  INVD1 U271 ( .I(n301), .ZN(n282) );
  INVD1 U272 ( .I(n300), .ZN(n281) );
  INVD1 U273 ( .I(n300), .ZN(n280) );
  INVD1 U274 ( .I(n301), .ZN(n297) );
  INVD1 U275 ( .I(n301), .ZN(n298) );
  INVD1 U276 ( .I(n300), .ZN(n296) );
  INVD1 U277 ( .I(n300), .ZN(n299) );
  INVD1 U278 ( .I(n319), .ZN(n310) );
  INVD1 U279 ( .I(n320), .ZN(n311) );
  INVD1 U280 ( .I(n319), .ZN(n312) );
  INVD1 U281 ( .I(n319), .ZN(n313) );
  INVD1 U282 ( .I(n320), .ZN(n314) );
  INVD1 U283 ( .I(n320), .ZN(n315) );
  INVD1 U284 ( .I(n319), .ZN(n305) );
  INVD1 U285 ( .I(n320), .ZN(n306) );
  INVD1 U286 ( .I(n319), .ZN(n307) );
  INVD1 U287 ( .I(n319), .ZN(n308) );
  INVD1 U288 ( .I(n319), .ZN(n309) );
  INVD1 U289 ( .I(n320), .ZN(n316) );
  INVD1 U290 ( .I(n320), .ZN(n317) );
  INVD1 U291 ( .I(n320), .ZN(n318) );
  INVD1 U292 ( .I(n320), .ZN(n304) );
  INVD1 U293 ( .I(n319), .ZN(n303) );
  INVD1 U294 ( .I(n319), .ZN(n302) );
  BUFFD1 U295 ( .I(n217), .Z(n271) );
  BUFFD1 U296 ( .I(n218), .Z(n270) );
  BUFFD1 U297 ( .I(n272), .Z(n269) );
  BUFFD1 U298 ( .I(n272), .Z(n268) );
  BUFFD1 U299 ( .I(n272), .Z(n267) );
  BUFFD1 U300 ( .I(n273), .Z(n266) );
  BUFFD1 U301 ( .I(n273), .Z(n265) );
  BUFFD1 U302 ( .I(n273), .Z(n264) );
  BUFFD1 U303 ( .I(n274), .Z(n263) );
  BUFFD1 U304 ( .I(n274), .Z(n262) );
  BUFFD1 U305 ( .I(n274), .Z(n261) );
  BUFFD1 U306 ( .I(n275), .Z(n260) );
  BUFFD1 U307 ( .I(n275), .Z(n259) );
  BUFFD1 U308 ( .I(n275), .Z(n258) );
  BUFFD1 U309 ( .I(n276), .Z(n257) );
  BUFFD1 U310 ( .I(n276), .Z(n256) );
  BUFFD1 U311 ( .I(n276), .Z(n255) );
  BUFFD1 U312 ( .I(n254), .Z(n252) );
  BUFFD1 U313 ( .I(n254), .Z(n253) );
  BUFFD1 U314 ( .I(n301), .Z(n300) );
  BUFFD1 U315 ( .I(n320), .Z(n319) );
  BUFFD1 U316 ( .I(n279), .Z(n272) );
  BUFFD1 U317 ( .I(n279), .Z(n273) );
  BUFFD1 U318 ( .I(n279), .Z(n274) );
  BUFFD1 U319 ( .I(n278), .Z(n275) );
  BUFFD1 U320 ( .I(n278), .Z(n276) );
  BUFFD1 U321 ( .I(n277), .Z(n254) );
  BUFFD1 U322 ( .I(n278), .Z(n277) );
  INVD1 U323 ( .I(n330), .ZN(n326) );
  INVD1 U324 ( .I(n330), .ZN(n325) );
  INVD1 U325 ( .I(n330), .ZN(n324) );
  INVD1 U326 ( .I(n330), .ZN(n323) );
  INVD1 U327 ( .I(n330), .ZN(n327) );
  INVD1 U328 ( .I(n330), .ZN(n329) );
  INVD1 U329 ( .I(n330), .ZN(n328) );
  INVD1 U330 ( .I(n330), .ZN(n322) );
  INVD1 U331 ( .I(n330), .ZN(n321) );
  BUFFD1 U332 ( .I(ChipClock), .Z(n279) );
  BUFFD1 U333 ( .I(ChipClock), .Z(n278) );
  MUX4ND0 U334 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n298), .S1(N44), .ZN(
        n750) );
  MUX4ND0 U335 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n296), .S1(N44), .ZN(
        n334) );
  MUX4ND0 U336 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n299), .S1(n318), .ZN(
        n347) );
  MUX4ND0 U337 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n298), .S1(n318), .ZN(
        n360) );
  MUX4ND0 U338 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n298), .S1(n318), .ZN(
        n373) );
  MUX4ND0 U339 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n298), .S1(n318), .ZN(
        n386) );
  MUX4ND0 U340 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n298), .S1(n318), .ZN(
        n399) );
  MUX4ND0 U341 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n298), .S1(n318), .ZN(
        n412) );
  MUX4ND0 U342 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n298), .S1(n316), .ZN(
        n425) );
  MUX4ND0 U343 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n298), .S1(n317), .ZN(
        n438) );
  MUX4ND0 U344 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n297), .S1(n318), .ZN(
        n451) );
  MUX4ND0 U345 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n297), .S1(n305), .ZN(
        n464) );
  MUX4ND0 U346 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n297), .S1(n306), .ZN(
        n477) );
  MUX4ND0 U347 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n297), .S1(n307), .ZN(
        n490) );
  MUX4ND0 U348 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n297), .S1(n308), .ZN(
        n503) );
  MUX4ND0 U349 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n297), .S1(n303), .ZN(
        n516) );
  MUX4ND0 U350 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n297), .S1(n310), .ZN(
        n529) );
  MUX4ND0 U351 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n297), .S1(n311), .ZN(
        n542) );
  MUX4ND0 U352 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n296), .S1(n309), .ZN(
        n555) );
  MUX4ND0 U353 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n296), .S1(N44), .ZN(
        n568) );
  MUX4ND0 U354 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n296), .S1(n313), .ZN(
        n581) );
  MUX4ND0 U355 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n298), .S1(n314), .ZN(
        n594) );
  MUX4ND0 U356 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n296), .S1(n315), .ZN(
        n607) );
  MUX4ND0 U357 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n296), .S1(n306), .ZN(
        n620) );
  MUX4ND0 U358 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n297), .S1(n312), .ZN(
        n633) );
  MUX4ND0 U359 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n297), .S1(n309), .ZN(
        n646) );
  MUX4ND0 U360 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n297), .S1(N44), .ZN(
        n659) );
  MUX4ND0 U361 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n297), .S1(N44), .ZN(
        n672) );
  MUX4ND0 U362 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n297), .S1(N44), .ZN(
        n685) );
  MUX4ND0 U363 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n298), .S1(N44), .ZN(
        n698) );
  MUX4ND0 U364 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n298), .S1(N44), .ZN(
        n711) );
  MUX4ND0 U365 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n298), .S1(n312), .ZN(
        n724) );
  MUX4ND0 U366 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n298), .S1(N44), .ZN(
        n737) );
  INVD1 U367 ( .I(N45), .ZN(n330) );
  INVD1 U368 ( .I(N43), .ZN(n301) );
  INVD1 U369 ( .I(N44), .ZN(n320) );
  MUX4D0 U370 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n280), .S1(n309), .Z(
        n751) );
  MUX4D0 U371 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n292), .S1(n305), .Z(
        n335) );
  MUX4D0 U372 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n288), .S1(n310), .Z(
        n348) );
  MUX4D0 U373 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n289), .S1(n310), .Z(
        n361) );
  MUX4D0 U374 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n289), .S1(n311), .Z(
        n374) );
  MUX4D0 U375 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n290), .S1(n311), .Z(
        n387) );
  MUX4D0 U376 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n290), .S1(n312), .Z(
        n400) );
  MUX4D0 U377 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n291), .S1(n312), .Z(
        n413) );
  MUX4D0 U378 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n291), .S1(n313), .Z(
        n426) );
  MUX4D0 U379 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n292), .S1(n313), .Z(
        n439) );
  MUX4D0 U380 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n292), .S1(n314), .Z(
        n452) );
  MUX4D0 U381 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n293), .S1(n314), .Z(
        n465) );
  MUX4D0 U382 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n293), .S1(n315), .Z(
        n478) );
  MUX4D0 U383 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n294), .S1(n315), .Z(
        n491) );
  MUX4D0 U384 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n294), .S1(n316), .Z(
        n504) );
  MUX4D0 U385 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n295), .S1(n316), .Z(
        n517) );
  MUX4D0 U386 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n295), .S1(n317), .Z(
        n530) );
  MUX4D0 U387 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n296), .S1(n317), .Z(
        n543) );
  MUX4D0 U388 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n287), .S1(n318), .Z(
        n556) );
  MUX4D0 U389 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n287), .S1(n305), .Z(
        n569) );
  MUX4D0 U390 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n286), .S1(n305), .Z(
        n582) );
  MUX4D0 U391 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n286), .S1(n305), .Z(
        n595) );
  MUX4D0 U392 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n285), .S1(n306), .Z(
        n608) );
  MUX4D0 U393 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n285), .S1(n307), .Z(
        n621) );
  MUX4D0 U394 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n284), .S1(n307), .Z(
        n634) );
  MUX4D0 U395 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n284), .S1(n308), .Z(
        n647) );
  MUX4D0 U396 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n283), .S1(n308), .Z(
        n660) );
  MUX4D0 U397 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n283), .S1(n302), .Z(
        n673) );
  MUX4D0 U398 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n282), .S1(n304), .Z(
        n686) );
  MUX4D0 U399 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n282), .S1(n307), .Z(
        n699) );
  MUX4D0 U400 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n281), .S1(n308), .Z(
        n712) );
  MUX4D0 U401 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n281), .S1(n313), .Z(
        n725) );
  MUX4D0 U402 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n280), .S1(n314), .Z(
        n738) );
  MUX4D0 U403 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n280), .S1(n309), .Z(
        n753) );
  MUX4D0 U404 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n280), .S1(n309), .Z(
        n755) );
  MUX4D0 U405 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n288), .S1(n309), .Z(
        n337) );
  MUX4D0 U406 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n288), .S1(n309), .Z(n339)
         );
  MUX4D0 U407 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n288), .S1(n310), .Z(
        n350) );
  MUX4D0 U408 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n289), .S1(n310), .Z(n352)
         );
  MUX4D0 U409 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n289), .S1(n310), .Z(
        n363) );
  MUX4D0 U410 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n289), .S1(n310), .Z(n365)
         );
  MUX4D0 U411 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n289), .S1(n311), .Z(
        n376) );
  MUX4D0 U412 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n290), .S1(n311), .Z(n378)
         );
  MUX4D0 U413 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n290), .S1(n311), .Z(
        n389) );
  MUX4D0 U414 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n290), .S1(n311), .Z(n391)
         );
  MUX4D0 U415 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n290), .S1(n312), .Z(
        n402) );
  MUX4D0 U416 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n291), .S1(n312), .Z(n404)
         );
  MUX4D0 U417 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n291), .S1(n312), .Z(
        n415) );
  MUX4D0 U418 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n291), .S1(n312), .Z(n417)
         );
  MUX4D0 U419 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n291), .S1(n313), .Z(
        n428) );
  MUX4D0 U420 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n292), .S1(n313), .Z(n430)
         );
  MUX4D0 U421 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n292), .S1(n313), .Z(
        n441) );
  MUX4D0 U422 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n292), .S1(n313), .Z(n443)
         );
  MUX4D0 U423 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n292), .S1(n314), .Z(
        n454) );
  MUX4D0 U424 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n293), .S1(n314), .Z(n456)
         );
  MUX4D0 U425 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n293), .S1(n314), .Z(
        n467) );
  MUX4D0 U426 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n293), .S1(n314), .Z(
        n469) );
  MUX4D0 U427 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n293), .S1(n315), .Z(
        n480) );
  MUX4D0 U428 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n294), .S1(n315), .Z(
        n482) );
  MUX4D0 U429 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n294), .S1(n315), .Z(
        n493) );
  MUX4D0 U430 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n294), .S1(n315), .Z(
        n495) );
  MUX4D0 U431 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n294), .S1(n316), .Z(
        n506) );
  MUX4D0 U432 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n295), .S1(n316), .Z(
        n508) );
  MUX4D0 U433 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n295), .S1(n316), .Z(
        n519) );
  MUX4D0 U434 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n295), .S1(n316), .Z(
        n521) );
  MUX4D0 U435 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n295), .S1(n317), .Z(
        n532) );
  MUX4D0 U436 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n296), .S1(n317), .Z(
        n534) );
  MUX4D0 U437 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n296), .S1(n317), .Z(
        n545) );
  MUX4D0 U438 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n288), .S1(n317), .Z(
        n547) );
  MUX4D0 U439 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n287), .S1(n318), .Z(
        n558) );
  MUX4D0 U440 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n287), .S1(n318), .Z(
        n560) );
  MUX4D0 U441 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n287), .S1(n306), .Z(
        n571) );
  MUX4D0 U442 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n287), .S1(n305), .Z(
        n573) );
  MUX4D0 U443 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n286), .S1(n305), .Z(
        n584) );
  MUX4D0 U444 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n286), .S1(n305), .Z(
        n586) );
  MUX4D0 U445 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n286), .S1(n307), .Z(
        n597) );
  MUX4D0 U446 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n286), .S1(n306), .Z(
        n599) );
  MUX4D0 U447 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n285), .S1(n306), .Z(
        n610) );
  MUX4D0 U448 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n285), .S1(n307), .Z(
        n612) );
  MUX4D0 U449 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n285), .S1(n307), .Z(
        n623) );
  MUX4D0 U450 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n285), .S1(n307), .Z(
        n625) );
  MUX4D0 U451 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n284), .S1(n307), .Z(
        n636) );
  MUX4D0 U452 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n284), .S1(n307), .Z(
        n638) );
  MUX4D0 U453 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n284), .S1(n308), .Z(
        n649) );
  MUX4D0 U454 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n284), .S1(n308), .Z(
        n651) );
  MUX4D0 U455 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n283), .S1(n308), .Z(
        n662) );
  MUX4D0 U456 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n283), .S1(n303), .Z(
        n664) );
  MUX4D0 U457 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n283), .S1(n302), .Z(
        n675) );
  MUX4D0 U458 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n283), .S1(n310), .Z(
        n677) );
  MUX4D0 U459 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n282), .S1(n311), .Z(
        n688) );
  MUX4D0 U460 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n282), .S1(n302), .Z(
        n690) );
  MUX4D0 U461 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n282), .S1(n316), .Z(
        n701) );
  MUX4D0 U462 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n282), .S1(n317), .Z(
        n703) );
  MUX4D0 U463 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n281), .S1(n318), .Z(
        n714) );
  MUX4D0 U464 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n281), .S1(n315), .Z(
        n716) );
  MUX4D0 U465 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n281), .S1(n305), .Z(
        n727) );
  MUX4D0 U466 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n281), .S1(n306), .Z(
        n729) );
  MUX4D0 U467 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n280), .S1(n307), .Z(
        n740) );
  MUX4D0 U468 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n280), .S1(n309), .Z(
        n742) );
  MUX4D0 U469 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n280), .S1(n309), .Z(
        n752) );
  MUX4D0 U470 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n288), .S1(n309), .Z(
        n336) );
  MUX4D0 U471 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n288), .S1(n310), .Z(
        n349) );
  MUX4D0 U472 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n289), .S1(n310), .Z(
        n362) );
  MUX4D0 U473 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n289), .S1(n311), .Z(
        n375) );
  MUX4D0 U474 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n290), .S1(n311), .Z(
        n388) );
  MUX4D0 U475 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n290), .S1(n312), .Z(
        n401) );
  MUX4D0 U476 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n291), .S1(n312), .Z(
        n414) );
  MUX4D0 U477 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n291), .S1(n313), .Z(
        n427) );
  MUX4D0 U478 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n292), .S1(n313), .Z(
        n440) );
  MUX4D0 U479 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n292), .S1(n314), .Z(
        n453) );
  MUX4D0 U480 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n293), .S1(n314), .Z(
        n466) );
  MUX4D0 U481 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n293), .S1(n315), .Z(
        n479) );
  MUX4D0 U482 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n294), .S1(n315), .Z(
        n492) );
  MUX4D0 U483 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n294), .S1(n316), .Z(
        n505) );
  MUX4D0 U484 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n295), .S1(n316), .Z(
        n518) );
  MUX4D0 U485 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n295), .S1(n317), .Z(
        n531) );
  MUX4D0 U486 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n296), .S1(n317), .Z(
        n544) );
  MUX4D0 U487 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n287), .S1(n318), .Z(
        n557) );
  MUX4D0 U488 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n287), .S1(n305), .Z(
        n570) );
  MUX4D0 U489 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n286), .S1(n306), .Z(
        n583) );
  MUX4D0 U490 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n286), .S1(n306), .Z(
        n596) );
  MUX4D0 U491 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n285), .S1(n306), .Z(
        n609) );
  MUX4D0 U492 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n285), .S1(n306), .Z(
        n622) );
  MUX4D0 U493 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n284), .S1(n307), .Z(
        n635) );
  MUX4D0 U494 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n284), .S1(n308), .Z(
        n648) );
  MUX4D0 U495 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n283), .S1(n308), .Z(
        n661) );
  MUX4D0 U496 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n283), .S1(n312), .Z(
        n674) );
  MUX4D0 U497 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n282), .S1(n313), .Z(
        n687) );
  MUX4D0 U498 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n282), .S1(N44), .Z(
        n700) );
  MUX4D0 U499 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n281), .S1(n304), .Z(
        n713) );
  MUX4D0 U500 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n281), .S1(n308), .Z(
        n726) );
  MUX4D0 U501 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n280), .S1(n304), .Z(
        n739) );
  MUX4D0 U502 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n280), .S1(n309), .Z(
        n754) );
  MUX4D0 U503 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n280), .S1(n309), .Z(
        n756) );
  MUX4D0 U504 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n288), .S1(n309), .Z(
        n338) );
  MUX4D0 U505 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n288), .S1(n310), .Z(n340)
         );
  MUX4D0 U506 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n288), .S1(n310), .Z(
        n351) );
  MUX4D0 U507 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n289), .S1(n310), .Z(n353)
         );
  MUX4D0 U508 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n289), .S1(n310), .Z(
        n364) );
  MUX4D0 U509 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n289), .S1(n311), .Z(n366)
         );
  MUX4D0 U510 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n289), .S1(n311), .Z(
        n377) );
  MUX4D0 U511 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n290), .S1(n311), .Z(n379)
         );
  MUX4D0 U512 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n290), .S1(n311), .Z(
        n390) );
  MUX4D0 U513 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n290), .S1(n312), .Z(n392)
         );
  MUX4D0 U514 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n290), .S1(n312), .Z(
        n403) );
  MUX4D0 U515 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n291), .S1(n312), .Z(n405)
         );
  MUX4D0 U516 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n291), .S1(n312), .Z(
        n416) );
  MUX4D0 U517 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n291), .S1(n313), .Z(n418)
         );
  MUX4D0 U518 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n291), .S1(n313), .Z(
        n429) );
  MUX4D0 U519 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n292), .S1(n313), .Z(n431)
         );
  MUX4D0 U520 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n292), .S1(n313), .Z(
        n442) );
  MUX4D0 U521 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n292), .S1(n314), .Z(n444)
         );
  MUX4D0 U522 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n293), .S1(n314), .Z(
        n455) );
  MUX4D0 U523 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n293), .S1(n314), .Z(n457)
         );
  MUX4D0 U524 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n293), .S1(n314), .Z(
        n468) );
  MUX4D0 U525 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n293), .S1(n315), .Z(
        n470) );
  MUX4D0 U526 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n294), .S1(n315), .Z(
        n481) );
  MUX4D0 U527 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n294), .S1(n315), .Z(
        n483) );
  MUX4D0 U528 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n294), .S1(n315), .Z(
        n494) );
  MUX4D0 U529 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n294), .S1(n316), .Z(
        n496) );
  MUX4D0 U530 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n295), .S1(n316), .Z(
        n507) );
  MUX4D0 U531 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n295), .S1(n316), .Z(
        n509) );
  MUX4D0 U532 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n295), .S1(n316), .Z(
        n520) );
  MUX4D0 U533 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n295), .S1(n317), .Z(
        n522) );
  MUX4D0 U534 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n296), .S1(n317), .Z(
        n533) );
  MUX4D0 U535 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n296), .S1(n317), .Z(
        n535) );
  MUX4D0 U536 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n288), .S1(n317), .Z(
        n546) );
  MUX4D0 U537 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n288), .S1(n318), .Z(
        n548) );
  MUX4D0 U538 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n287), .S1(n318), .Z(
        n559) );
  MUX4D0 U539 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n287), .S1(n308), .Z(
        n561) );
  MUX4D0 U540 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n287), .S1(n305), .Z(
        n572) );
  MUX4D0 U541 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n287), .S1(n306), .Z(
        n574) );
  MUX4D0 U542 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n286), .S1(n306), .Z(
        n585) );
  MUX4D0 U543 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n286), .S1(n305), .Z(
        n587) );
  MUX4D0 U544 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n286), .S1(n305), .Z(
        n598) );
  MUX4D0 U545 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n286), .S1(n305), .Z(
        n600) );
  MUX4D0 U546 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n285), .S1(n306), .Z(
        n611) );
  MUX4D0 U547 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n285), .S1(n306), .Z(
        n613) );
  MUX4D0 U548 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n285), .S1(n307), .Z(
        n624) );
  MUX4D0 U549 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n285), .S1(n307), .Z(
        n626) );
  MUX4D0 U550 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n284), .S1(n307), .Z(
        n637) );
  MUX4D0 U551 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n284), .S1(n308), .Z(
        n639) );
  MUX4D0 U552 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n284), .S1(n308), .Z(
        n650) );
  MUX4D0 U553 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n284), .S1(n308), .Z(
        n652) );
  MUX4D0 U554 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n283), .S1(n308), .Z(
        n663) );
  MUX4D0 U555 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n283), .S1(n314), .Z(
        n665) );
  MUX4D0 U556 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n283), .S1(n315), .Z(
        n676) );
  MUX4D0 U557 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n283), .S1(n309), .Z(
        n678) );
  MUX4D0 U558 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n282), .S1(n303), .Z(
        n689) );
  MUX4D0 U559 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n282), .S1(n303), .Z(
        n691) );
  MUX4D0 U560 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n282), .S1(n302), .Z(
        n702) );
  MUX4D0 U561 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n282), .S1(n310), .Z(
        n704) );
  MUX4D0 U562 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n281), .S1(n305), .Z(
        n715) );
  MUX4D0 U563 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n281), .S1(n316), .Z(
        n717) );
  MUX4D0 U564 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n281), .S1(n317), .Z(
        n728) );
  MUX4D0 U565 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n281), .S1(n318), .Z(
        n730) );
  MUX4D0 U566 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n280), .S1(n311), .Z(
        n741) );
  MUX4D0 U567 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n280), .S1(n309), .Z(
        n743) );
  MUX3ND0 U568 ( .I0(n332), .I1(n333), .I2(n334), .S0(n302), .S1(n322), .ZN(
        n331) );
  MUX3ND0 U569 ( .I0(n341), .I1(n342), .I2(n343), .S0(n69), .S1(n65), .ZN(N81)
         );
  MUX3ND0 U570 ( .I0(n345), .I1(n346), .I2(n347), .S0(n302), .S1(N45), .ZN(
        n344) );
  MUX3ND0 U571 ( .I0(n354), .I1(n355), .I2(n356), .S0(n70), .S1(n65), .ZN(N80)
         );
  MUX3ND0 U572 ( .I0(n358), .I1(n359), .I2(n360), .S0(n303), .S1(n328), .ZN(
        n357) );
  MUX3ND0 U573 ( .I0(n367), .I1(n368), .I2(n369), .S0(n69), .S1(n66), .ZN(N79)
         );
  MUX3ND0 U574 ( .I0(n371), .I1(n372), .I2(n373), .S0(n302), .S1(n329), .ZN(
        n370) );
  MUX3ND0 U575 ( .I0(n380), .I1(n381), .I2(n382), .S0(n70), .S1(n66), .ZN(N78)
         );
  MUX3ND0 U576 ( .I0(n384), .I1(n385), .I2(n386), .S0(n303), .S1(n329), .ZN(
        n383) );
  MUX3ND0 U577 ( .I0(n393), .I1(n394), .I2(n395), .S0(n69), .S1(n65), .ZN(N77)
         );
  MUX3ND0 U578 ( .I0(n397), .I1(n398), .I2(n399), .S0(n302), .S1(n329), .ZN(
        n396) );
  MUX3ND0 U579 ( .I0(n406), .I1(n407), .I2(n408), .S0(n70), .S1(n65), .ZN(N76)
         );
  MUX3ND0 U580 ( .I0(n410), .I1(n411), .I2(n412), .S0(n304), .S1(n329), .ZN(
        n409) );
  MUX3ND0 U581 ( .I0(n419), .I1(n420), .I2(n421), .S0(n68), .S1(n65), .ZN(N75)
         );
  MUX3ND0 U582 ( .I0(n423), .I1(n424), .I2(n425), .S0(n303), .S1(n329), .ZN(
        n422) );
  MUX3ND0 U583 ( .I0(n432), .I1(n433), .I2(n434), .S0(n67), .S1(n65), .ZN(N74)
         );
  MUX3ND0 U584 ( .I0(n436), .I1(n437), .I2(n438), .S0(n304), .S1(n329), .ZN(
        n435) );
  MUX3ND0 U585 ( .I0(n445), .I1(n446), .I2(n447), .S0(n68), .S1(n65), .ZN(N73)
         );
  MUX3ND0 U586 ( .I0(n449), .I1(n450), .I2(n451), .S0(n303), .S1(n329), .ZN(
        n448) );
  MUX3ND0 U587 ( .I0(n458), .I1(n459), .I2(n460), .S0(n67), .S1(n65), .ZN(N72)
         );
  MUX3ND0 U588 ( .I0(n462), .I1(n463), .I2(n464), .S0(n304), .S1(n329), .ZN(
        n461) );
  MUX3ND0 U589 ( .I0(n471), .I1(n472), .I2(n473), .S0(N46), .S1(n65), .ZN(N71)
         );
  MUX3ND0 U590 ( .I0(n475), .I1(n476), .I2(n477), .S0(n304), .S1(n329), .ZN(
        n474) );
  MUX3ND0 U591 ( .I0(n484), .I1(n485), .I2(n486), .S0(n70), .S1(N47), .ZN(N70)
         );
  MUX3ND0 U592 ( .I0(n488), .I1(n489), .I2(n490), .S0(n304), .S1(n329), .ZN(
        n487) );
  MUX3ND0 U593 ( .I0(n497), .I1(n498), .I2(n499), .S0(n69), .S1(n66), .ZN(N69)
         );
  MUX3ND0 U594 ( .I0(n501), .I1(n502), .I2(n503), .S0(n303), .S1(n329), .ZN(
        n500) );
  MUX3ND0 U595 ( .I0(n510), .I1(n511), .I2(n512), .S0(n68), .S1(N47), .ZN(N68)
         );
  MUX3ND0 U596 ( .I0(n514), .I1(n515), .I2(n516), .S0(n304), .S1(n329), .ZN(
        n513) );
  MUX3ND0 U597 ( .I0(n523), .I1(n524), .I2(n525), .S0(n67), .S1(n65), .ZN(N67)
         );
  MUX3ND0 U598 ( .I0(n527), .I1(n528), .I2(n529), .S0(n303), .S1(n328), .ZN(
        n526) );
  MUX3ND0 U599 ( .I0(n536), .I1(n537), .I2(n538), .S0(N46), .S1(n65), .ZN(N66)
         );
  MUX3ND0 U600 ( .I0(n540), .I1(n541), .I2(n542), .S0(n303), .S1(n328), .ZN(
        n539) );
  MUX3ND0 U601 ( .I0(n549), .I1(n550), .I2(n551), .S0(n67), .S1(n66), .ZN(N65)
         );
  MUX3ND0 U602 ( .I0(n553), .I1(n554), .I2(n555), .S0(n302), .S1(n328), .ZN(
        n552) );
  MUX3ND0 U603 ( .I0(n562), .I1(n563), .I2(n564), .S0(N46), .S1(N47), .ZN(N64)
         );
  MUX3ND0 U604 ( .I0(n566), .I1(n567), .I2(n568), .S0(n302), .S1(n328), .ZN(
        n565) );
  MUX3ND0 U605 ( .I0(n575), .I1(n576), .I2(n577), .S0(N46), .S1(n66), .ZN(N63)
         );
  MUX3ND0 U606 ( .I0(n579), .I1(n580), .I2(n581), .S0(n302), .S1(n328), .ZN(
        n578) );
  MUX3ND0 U607 ( .I0(n588), .I1(n589), .I2(n590), .S0(n68), .S1(N47), .ZN(N62)
         );
  MUX3ND0 U608 ( .I0(n592), .I1(n593), .I2(n594), .S0(n302), .S1(n328), .ZN(
        n591) );
  MUX3ND0 U609 ( .I0(n601), .I1(n602), .I2(n603), .S0(N46), .S1(n66), .ZN(N61)
         );
  MUX3ND0 U610 ( .I0(n605), .I1(n606), .I2(n607), .S0(n303), .S1(n328), .ZN(
        n604) );
  MUX3ND0 U611 ( .I0(n614), .I1(n615), .I2(n616), .S0(N46), .S1(N47), .ZN(N60)
         );
  MUX3ND0 U612 ( .I0(n618), .I1(n619), .I2(n620), .S0(n304), .S1(n328), .ZN(
        n617) );
  MUX3ND0 U613 ( .I0(n627), .I1(n628), .I2(n629), .S0(n68), .S1(n66), .ZN(N59)
         );
  MUX3ND0 U614 ( .I0(n631), .I1(n632), .I2(n633), .S0(n302), .S1(n328), .ZN(
        n630) );
  MUX3ND0 U615 ( .I0(n640), .I1(n641), .I2(n642), .S0(n70), .S1(N47), .ZN(N58)
         );
  MUX3ND0 U616 ( .I0(n644), .I1(n645), .I2(n646), .S0(n304), .S1(n328), .ZN(
        n643) );
  MUX3ND0 U617 ( .I0(n653), .I1(n654), .I2(n655), .S0(n69), .S1(n66), .ZN(N57)
         );
  MUX3ND0 U618 ( .I0(n657), .I1(n658), .I2(n659), .S0(n304), .S1(n328), .ZN(
        n656) );
  MUX3ND0 U619 ( .I0(n666), .I1(n667), .I2(n668), .S0(n67), .S1(N47), .ZN(N56)
         );
  MUX3ND0 U620 ( .I0(n670), .I1(n671), .I2(n672), .S0(n304), .S1(n328), .ZN(
        n669) );
  MUX3ND0 U621 ( .I0(n679), .I1(n680), .I2(n681), .S0(n69), .S1(n66), .ZN(N55)
         );
  MUX3ND0 U622 ( .I0(n683), .I1(n684), .I2(n685), .S0(n304), .S1(n327), .ZN(
        n682) );
  MUX3ND0 U623 ( .I0(n692), .I1(n693), .I2(n694), .S0(N46), .S1(N47), .ZN(N54)
         );
  MUX3ND0 U624 ( .I0(n696), .I1(n697), .I2(n698), .S0(n303), .S1(n327), .ZN(
        n695) );
  MUX3ND0 U625 ( .I0(n705), .I1(n706), .I2(n707), .S0(n70), .S1(n66), .ZN(N53)
         );
  MUX3ND0 U626 ( .I0(n709), .I1(n710), .I2(n711), .S0(n303), .S1(n327), .ZN(
        n708) );
  MUX3ND0 U627 ( .I0(n718), .I1(n719), .I2(n720), .S0(n69), .S1(N47), .ZN(N52)
         );
  MUX3ND0 U628 ( .I0(n722), .I1(n723), .I2(n724), .S0(n303), .S1(n327), .ZN(
        n721) );
  MUX3ND0 U629 ( .I0(n731), .I1(n732), .I2(n733), .S0(n68), .S1(n66), .ZN(N51)
         );
  MUX3ND0 U630 ( .I0(n735), .I1(n736), .I2(n737), .S0(n302), .S1(n327), .ZN(
        n734) );
  MUX3ND0 U631 ( .I0(n744), .I1(n745), .I2(n746), .S0(n67), .S1(N47), .ZN(N50)
         );
  MUX3ND0 U632 ( .I0(n748), .I1(n749), .I2(n750), .S0(n302), .S1(n327), .ZN(
        n747) );
  MUX3ND0 U633 ( .I0(n757), .I1(n758), .I2(n759), .S0(n70), .S1(n65), .ZN(N49)
         );
  MUX2ND0 U634 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n291), .ZN(
        n333) );
  MUX2ND0 U635 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n284), .ZN(
        n332) );
  MUX3ND0 U636 ( .I0(n336), .I1(n335), .I2(n331), .S0(n322), .S1(n67), .ZN(
        n343) );
  MUX2ND0 U637 ( .I0(n338), .I1(n337), .S(n327), .ZN(n342) );
  MUX2ND0 U638 ( .I0(n340), .I1(n339), .S(n327), .ZN(n341) );
  MUX2ND0 U639 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n281), .ZN(
        n346) );
  MUX2ND0 U640 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n280), .ZN(
        n345) );
  MUX3ND0 U641 ( .I0(n349), .I1(n348), .I2(n344), .S0(N45), .S1(n68), .ZN(n356) );
  MUX2ND0 U642 ( .I0(n351), .I1(n350), .S(n327), .ZN(n355) );
  MUX2ND0 U643 ( .I0(n353), .I1(n352), .S(n327), .ZN(n354) );
  MUX2ND0 U644 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n283), .ZN(
        n359) );
  MUX2ND0 U645 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n282), .ZN(
        n358) );
  MUX3ND0 U646 ( .I0(n362), .I1(n361), .I2(n357), .S0(n322), .S1(n67), .ZN(
        n369) );
  MUX2ND0 U647 ( .I0(n364), .I1(n363), .S(n327), .ZN(n368) );
  MUX2ND0 U648 ( .I0(n366), .I1(n365), .S(n327), .ZN(n367) );
  MUX2ND0 U649 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n290), .ZN(
        n372) );
  MUX2ND0 U650 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n280), .ZN(
        n371) );
  MUX3ND0 U651 ( .I0(n375), .I1(n374), .I2(n370), .S0(N45), .S1(n69), .ZN(n382) );
  MUX2ND0 U652 ( .I0(n377), .I1(n376), .S(n326), .ZN(n381) );
  MUX2ND0 U653 ( .I0(n379), .I1(n378), .S(n326), .ZN(n380) );
  MUX2ND0 U654 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n289), .ZN(
        n385) );
  MUX2ND0 U655 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n281), .ZN(
        n384) );
  MUX3ND0 U656 ( .I0(n388), .I1(n387), .I2(n383), .S0(n322), .S1(n67), .ZN(
        n395) );
  MUX2ND0 U657 ( .I0(n390), .I1(n389), .S(n326), .ZN(n394) );
  MUX2ND0 U658 ( .I0(n392), .I1(n391), .S(n326), .ZN(n393) );
  MUX2ND0 U659 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n295), .ZN(
        n398) );
  MUX2ND0 U660 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n288), .ZN(
        n397) );
  MUX3ND0 U661 ( .I0(n401), .I1(n400), .I2(n396), .S0(N45), .S1(n70), .ZN(n408) );
  MUX2ND0 U662 ( .I0(n403), .I1(n402), .S(n326), .ZN(n407) );
  MUX2ND0 U663 ( .I0(n405), .I1(n404), .S(n326), .ZN(n406) );
  MUX2ND0 U664 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n287), .ZN(
        n411) );
  MUX2ND0 U665 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n298), .ZN(
        n410) );
  MUX3ND0 U666 ( .I0(n414), .I1(n413), .I2(n409), .S0(n322), .S1(n70), .ZN(
        n421) );
  MUX2ND0 U667 ( .I0(n416), .I1(n415), .S(n326), .ZN(n420) );
  MUX2ND0 U668 ( .I0(n418), .I1(n417), .S(n326), .ZN(n419) );
  MUX2ND0 U669 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n296), .ZN(
        n424) );
  MUX2ND0 U670 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n297), .ZN(
        n423) );
  MUX3ND0 U671 ( .I0(n427), .I1(n426), .I2(n422), .S0(N45), .S1(N46), .ZN(n434) );
  MUX2ND0 U672 ( .I0(n429), .I1(n428), .S(n326), .ZN(n433) );
  MUX2ND0 U673 ( .I0(n431), .I1(n430), .S(n326), .ZN(n432) );
  MUX2ND0 U674 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n291), .ZN(
        n437) );
  MUX2ND0 U675 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n289), .ZN(
        n436) );
  MUX3ND0 U676 ( .I0(n440), .I1(n439), .I2(n435), .S0(n322), .S1(n68), .ZN(
        n447) );
  MUX2ND0 U677 ( .I0(n442), .I1(n441), .S(n326), .ZN(n446) );
  MUX2ND0 U678 ( .I0(n444), .I1(n443), .S(n326), .ZN(n445) );
  MUX2ND0 U679 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n290), .ZN(
        n450) );
  MUX2ND0 U680 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n294), .ZN(
        n449) );
  MUX3ND0 U681 ( .I0(n453), .I1(n452), .I2(n448), .S0(n321), .S1(N46), .ZN(
        n460) );
  MUX2ND0 U682 ( .I0(n455), .I1(n454), .S(n325), .ZN(n459) );
  MUX2ND0 U683 ( .I0(n457), .I1(n456), .S(n325), .ZN(n458) );
  MUX2ND0 U684 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n292), 
        .ZN(n463) );
  MUX2ND0 U685 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n293), 
        .ZN(n462) );
  MUX3ND0 U686 ( .I0(n466), .I1(n465), .I2(n461), .S0(n322), .S1(n69), .ZN(
        n473) );
  MUX2ND0 U687 ( .I0(n468), .I1(n467), .S(n325), .ZN(n472) );
  MUX2ND0 U688 ( .I0(n470), .I1(n469), .S(n325), .ZN(n471) );
  MUX2ND0 U689 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n295), 
        .ZN(n476) );
  MUX2ND0 U690 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n282), 
        .ZN(n475) );
  MUX3ND0 U691 ( .I0(n479), .I1(n478), .I2(n474), .S0(n321), .S1(n70), .ZN(
        n486) );
  MUX2ND0 U692 ( .I0(n481), .I1(n480), .S(n325), .ZN(n485) );
  MUX2ND0 U693 ( .I0(n483), .I1(n482), .S(n325), .ZN(n484) );
  MUX2ND0 U694 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n294), 
        .ZN(n489) );
  MUX2ND0 U695 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n287), 
        .ZN(n488) );
  MUX3ND0 U696 ( .I0(n492), .I1(n491), .I2(n487), .S0(n322), .S1(n68), .ZN(
        n499) );
  MUX2ND0 U697 ( .I0(n494), .I1(n493), .S(n325), .ZN(n498) );
  MUX2ND0 U698 ( .I0(n496), .I1(n495), .S(n325), .ZN(n497) );
  MUX2ND0 U699 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n296), 
        .ZN(n502) );
  MUX2ND0 U700 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n288), 
        .ZN(n501) );
  MUX3ND0 U701 ( .I0(n505), .I1(n504), .I2(n500), .S0(n321), .S1(n67), .ZN(
        n512) );
  MUX2ND0 U702 ( .I0(n507), .I1(n506), .S(n325), .ZN(n511) );
  MUX2ND0 U703 ( .I0(n509), .I1(n508), .S(n325), .ZN(n510) );
  MUX2ND0 U704 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n284), 
        .ZN(n515) );
  MUX2ND0 U705 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n286), 
        .ZN(n514) );
  MUX3ND0 U706 ( .I0(n518), .I1(n517), .I2(n513), .S0(n321), .S1(n67), .ZN(
        n525) );
  MUX2ND0 U707 ( .I0(n520), .I1(n519), .S(n325), .ZN(n524) );
  MUX2ND0 U708 ( .I0(n522), .I1(n521), .S(n324), .ZN(n523) );
  MUX2ND0 U709 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n285), 
        .ZN(n528) );
  MUX2ND0 U710 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n281), 
        .ZN(n527) );
  MUX3ND0 U711 ( .I0(n531), .I1(n530), .I2(n526), .S0(n321), .S1(n69), .ZN(
        n538) );
  MUX2ND0 U712 ( .I0(n533), .I1(n532), .S(n328), .ZN(n537) );
  MUX2ND0 U713 ( .I0(n535), .I1(n534), .S(n329), .ZN(n536) );
  MUX2ND0 U714 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n283), 
        .ZN(n541) );
  MUX2ND0 U715 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n282), 
        .ZN(n540) );
  MUX3ND0 U716 ( .I0(n544), .I1(n543), .I2(n539), .S0(n322), .S1(N46), .ZN(
        n551) );
  MUX2ND0 U717 ( .I0(n546), .I1(n545), .S(n327), .ZN(n550) );
  MUX2ND0 U718 ( .I0(n548), .I1(n547), .S(N45), .ZN(n549) );
  MUX2ND0 U719 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(N43), .ZN(
        n554) );
  MUX2ND0 U720 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n280), 
        .ZN(n553) );
  MUX3ND0 U721 ( .I0(n557), .I1(n556), .I2(n552), .S0(n322), .S1(N46), .ZN(
        n564) );
  MUX2ND0 U722 ( .I0(n559), .I1(n558), .S(n325), .ZN(n563) );
  MUX2ND0 U723 ( .I0(n561), .I1(n560), .S(n322), .ZN(n562) );
  MUX2ND0 U724 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(N43), .ZN(
        n567) );
  MUX2ND0 U725 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n285), 
        .ZN(n566) );
  MUX3ND0 U726 ( .I0(n570), .I1(n569), .I2(n565), .S0(n321), .S1(n68), .ZN(
        n577) );
  MUX2ND0 U727 ( .I0(n572), .I1(n571), .S(n324), .ZN(n576) );
  MUX2ND0 U728 ( .I0(n574), .I1(n573), .S(n324), .ZN(n575) );
  MUX2ND0 U729 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n293), 
        .ZN(n580) );
  MUX2ND0 U730 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n292), 
        .ZN(n579) );
  MUX3ND0 U731 ( .I0(n583), .I1(n582), .I2(n578), .S0(n321), .S1(n70), .ZN(
        n590) );
  MUX2ND0 U732 ( .I0(n585), .I1(n584), .S(n326), .ZN(n589) );
  MUX2ND0 U733 ( .I0(n587), .I1(n586), .S(n324), .ZN(n588) );
  MUX2ND0 U734 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(N43), .ZN(
        n593) );
  MUX2ND0 U735 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(N43), .ZN(
        n592) );
  MUX3ND0 U736 ( .I0(n596), .I1(n595), .I2(n591), .S0(n322), .S1(n70), .ZN(
        n603) );
  MUX2ND0 U737 ( .I0(n598), .I1(n597), .S(n325), .ZN(n602) );
  MUX2ND0 U738 ( .I0(n600), .I1(n599), .S(n324), .ZN(n601) );
  MUX2ND0 U739 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(N43), .ZN(
        n606) );
  MUX2ND0 U740 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(N43), .ZN(
        n605) );
  MUX3ND0 U741 ( .I0(n609), .I1(n608), .I2(n604), .S0(n322), .S1(n69), .ZN(
        n616) );
  MUX2ND0 U742 ( .I0(n611), .I1(n610), .S(n324), .ZN(n615) );
  MUX2ND0 U743 ( .I0(n613), .I1(n612), .S(n324), .ZN(n614) );
  MUX2ND0 U744 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(N43), .ZN(
        n619) );
  MUX2ND0 U745 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(N43), .ZN(
        n618) );
  MUX3ND0 U746 ( .I0(n622), .I1(n621), .I2(n617), .S0(n321), .S1(n67), .ZN(
        n629) );
  MUX2ND0 U747 ( .I0(n624), .I1(n623), .S(n323), .ZN(n628) );
  MUX2ND0 U748 ( .I0(n626), .I1(n625), .S(n325), .ZN(n627) );
  MUX2ND0 U749 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(N43), .ZN(
        n632) );
  MUX2ND0 U750 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n299), 
        .ZN(n631) );
  MUX3ND0 U751 ( .I0(n635), .I1(n634), .I2(n630), .S0(n321), .S1(n68), .ZN(
        n642) );
  MUX2ND0 U752 ( .I0(n637), .I1(n636), .S(n324), .ZN(n641) );
  MUX2ND0 U753 ( .I0(n639), .I1(n638), .S(n323), .ZN(n640) );
  MUX2ND0 U754 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n299), 
        .ZN(n645) );
  MUX2ND0 U755 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(N43), .ZN(
        n644) );
  MUX3ND0 U756 ( .I0(n648), .I1(n647), .I2(n643), .S0(n321), .S1(n70), .ZN(
        n655) );
  MUX2ND0 U757 ( .I0(n650), .I1(n649), .S(n323), .ZN(n654) );
  MUX2ND0 U758 ( .I0(n652), .I1(n651), .S(n323), .ZN(n653) );
  MUX2ND0 U759 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n299), 
        .ZN(n658) );
  MUX2ND0 U760 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n299), 
        .ZN(n657) );
  MUX3ND0 U761 ( .I0(n661), .I1(n660), .I2(n656), .S0(n321), .S1(n70), .ZN(
        n668) );
  MUX2ND0 U762 ( .I0(n663), .I1(n662), .S(n324), .ZN(n667) );
  MUX2ND0 U763 ( .I0(n665), .I1(n664), .S(n323), .ZN(n666) );
  MUX2ND0 U764 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n299), 
        .ZN(n671) );
  MUX2ND0 U765 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n299), 
        .ZN(n670) );
  MUX3ND0 U766 ( .I0(n674), .I1(n673), .I2(n669), .S0(N45), .S1(n69), .ZN(n681) );
  MUX2ND0 U767 ( .I0(n676), .I1(n675), .S(n323), .ZN(n680) );
  MUX2ND0 U768 ( .I0(n678), .I1(n677), .S(n321), .ZN(n679) );
  MUX2ND0 U769 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n299), 
        .ZN(n684) );
  MUX2ND0 U770 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n299), 
        .ZN(n683) );
  MUX3ND0 U771 ( .I0(n687), .I1(n686), .I2(n682), .S0(n321), .S1(n67), .ZN(
        n694) );
  MUX2ND0 U772 ( .I0(n689), .I1(n688), .S(n324), .ZN(n693) );
  MUX2ND0 U773 ( .I0(n691), .I1(n690), .S(n323), .ZN(n692) );
  MUX2ND0 U774 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n299), 
        .ZN(n697) );
  MUX2ND0 U775 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n299), 
        .ZN(n696) );
  MUX3ND0 U776 ( .I0(n700), .I1(n699), .I2(n695), .S0(N45), .S1(n67), .ZN(n707) );
  MUX2ND0 U777 ( .I0(n702), .I1(n701), .S(n323), .ZN(n706) );
  MUX2ND0 U778 ( .I0(n704), .I1(n703), .S(n326), .ZN(n705) );
  MUX2ND0 U779 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n299), 
        .ZN(n710) );
  MUX2ND0 U780 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n299), 
        .ZN(n709) );
  MUX3ND0 U781 ( .I0(n713), .I1(n712), .I2(n708), .S0(N45), .S1(n68), .ZN(n720) );
  MUX2ND0 U782 ( .I0(n715), .I1(n714), .S(n324), .ZN(n719) );
  MUX2ND0 U783 ( .I0(n717), .I1(n716), .S(n323), .ZN(n718) );
  MUX2ND0 U784 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n299), 
        .ZN(n723) );
  MUX2ND0 U785 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n299), 
        .ZN(n722) );
  MUX3ND0 U786 ( .I0(n726), .I1(n725), .I2(n721), .S0(N45), .S1(n68), .ZN(n733) );
  MUX2ND0 U787 ( .I0(n728), .I1(n727), .S(n323), .ZN(n732) );
  MUX2ND0 U788 ( .I0(n730), .I1(n729), .S(n324), .ZN(n731) );
  MUX2ND0 U789 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(N43), .ZN(
        n736) );
  MUX2ND0 U790 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(N43), .ZN(
        n735) );
  MUX3ND0 U791 ( .I0(n739), .I1(n738), .I2(n734), .S0(N45), .S1(n69), .ZN(n746) );
  MUX2ND0 U792 ( .I0(n741), .I1(n740), .S(n323), .ZN(n745) );
  MUX2ND0 U793 ( .I0(n743), .I1(n742), .S(n323), .ZN(n744) );
  MUX2ND0 U794 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(N43), .ZN(
        n749) );
  MUX2ND0 U795 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n286), 
        .ZN(n748) );
  MUX3ND0 U796 ( .I0(n752), .I1(n751), .I2(n747), .S0(N45), .S1(n69), .ZN(n759) );
  MUX2ND0 U797 ( .I0(n754), .I1(n753), .S(n323), .ZN(n758) );
  MUX2ND0 U798 ( .I0(n756), .I1(n755), .S(n324), .ZN(n757) );
  XOR3D0 U799 ( .A1(n60), .A2(n761), .A3(n762), .Z(n760) );
  XOR3D0 U800 ( .A1(n40), .A2(n43), .A3(n763), .Z(n762) );
  XOR3D0 U801 ( .A1(n764), .A2(DataI[3]), .A3(n765), .Z(n763) );
  XOR3D0 U802 ( .A1(n12), .A2(n15), .A3(n766), .Z(n765) );
  XOR3D0 U803 ( .A1(n767), .A2(DataI[10]), .A3(n768), .Z(n766) );
  XOR3D0 U804 ( .A1(n18), .A2(n13), .A3(n769), .Z(n768) );
  XOR3D0 U805 ( .A1(n770), .A2(DataI[17]), .A3(n771), .Z(n769) );
  XNR4D0 U806 ( .A1(n41), .A2(n38), .A3(n50), .A4(n45), .ZN(n771) );
  XOR4D0 U807 ( .A1(DataI[29]), .A2(n54), .A3(n64), .A4(n61), .Z(n770) );
  XOR4D0 U808 ( .A1(n25), .A2(n22), .A3(n34), .A4(n29), .Z(n767) );
  XOR4D0 U809 ( .A1(n3), .A2(n8), .A3(n6), .A4(DataI[15]), .Z(n764) );
  XNR4D0 U810 ( .A1(DataI[7]), .A2(n36), .A3(n24), .A4(n27), .ZN(n761) );
  XOR4D0 U811 ( .A1(n772), .A2(N78), .A3(n773), .A4(n774), .Z(N84) );
  XNR4D0 U812 ( .A1(N75), .A2(N74), .A3(N77), .A4(N76), .ZN(n774) );
  XNR3D0 U813 ( .A1(N81), .A2(N80), .A3(N79), .ZN(n773) );
  XOR3D0 U814 ( .A1(N73), .A2(N72), .A3(n775), .Z(n772) );
  XOR3D0 U815 ( .A1(N71), .A2(n776), .A3(n777), .Z(n775) );
  XOR3D0 U816 ( .A1(N66), .A2(N65), .A3(n778), .Z(n777) );
  XOR3D0 U817 ( .A1(n779), .A2(N64), .A3(n780), .Z(n778) );
  XOR3D0 U818 ( .A1(N59), .A2(N58), .A3(n781), .Z(n780) );
  XOR3D0 U819 ( .A1(n782), .A2(N57), .A3(n783), .Z(n781) );
  XNR4D0 U820 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n783) );
  XOR4D0 U821 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n782) );
  XOR4D0 U822 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .Z(n779) );
  XNR4D0 U823 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n776) );
  ND3D0 U824 ( .A1(N44), .A2(n296), .A3(n324), .ZN(n786) );
  ND3D0 U825 ( .A1(N44), .A2(n301), .A3(n329), .ZN(n787) );
  ND3D0 U826 ( .A1(n288), .A2(n319), .A3(n327), .ZN(n788) );
  ND3D0 U827 ( .A1(n300), .A2(n319), .A3(n323), .ZN(n789) );
  ND3D0 U828 ( .A1(n287), .A2(n330), .A3(N44), .ZN(n790) );
  ND3D0 U829 ( .A1(n301), .A2(n330), .A3(N44), .ZN(n791) );
  ND3D0 U830 ( .A1(n320), .A2(n330), .A3(n295), .ZN(n792) );
  AN3D0 U831 ( .A1(n784), .A2(ChipEna), .A3(Write), .Z(n794) );
  CKND0 U832 ( .CLK(Read), .CN(n784) );
  CKND0 U833 ( .CLK(n66), .CN(n798) );
  CKND0 U834 ( .CLK(n68), .CN(n796) );
  ND3D0 U835 ( .A1(n320), .A2(n330), .A3(n301), .ZN(n793) );
  AN2D0 U836 ( .A1(DreadyReg), .A2(ChipEna), .Z(Dready) );
  AN2D0 U837 ( .A1(ClockIn), .A2(ChipEna), .Z(ChipClock) );
endmodule


module FIFOStateM_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

