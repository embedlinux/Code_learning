
module FIFOTop ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, ClkW, Reseter
 );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(n1), .WriteReq(n158), .ClkR(ClkR), 
        .ClkW(ClkW), .Reset(n167) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({n200, n199, n198, 
        n197, n196, n195, n194, n193, n192, n191, n190, n189, n188, n187, n186, 
        n185, n184, n183, n182, n117, n181, n180, n179, n178, n177, n176, n175, 
        n174, n173, n172, n171, n170}), .AddrR(SM_ReadAddr), .AddrW(
        SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), .ChipEna(\*Logic1* ), .Read(
        n169), .Write(SM_MemWriteCmd), .Reset(n167) );
  CKNXD16 U2 ( .I(Din[2]), .ZN(n136) );
  BUFFD0 U3 ( .I(n148), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n167) );
  INVD16 U5 ( .I(Reseter), .ZN(n2) );
  INVD1 U6 ( .I(n2), .ZN(n3) );
  BUFFD0 U7 ( .I(n137), .Z(n172) );
  INVD0 U8 ( .I(n4), .ZN(n5) );
  CKNXD16 U9 ( .I(Din[31]), .ZN(n4) );
  BUFFD0 U10 ( .I(n5), .Z(n6) );
  BUFFD0 U11 ( .I(n6), .Z(n7) );
  BUFFD0 U12 ( .I(n7), .Z(n8) );
  BUFFD0 U13 ( .I(n8), .Z(n9) );
  BUFFD0 U14 ( .I(n9), .Z(n10) );
  BUFFD0 U15 ( .I(n10), .Z(n11) );
  BUFFD0 U16 ( .I(n11), .Z(n12) );
  BUFFD0 U17 ( .I(n12), .Z(n13) );
  BUFFD0 U18 ( .I(n13), .Z(n14) );
  BUFFD0 U19 ( .I(n14), .Z(n15) );
  BUFFD0 U20 ( .I(n15), .Z(n16) );
  BUFFD0 U21 ( .I(n16), .Z(n17) );
  BUFFD0 U22 ( .I(n17), .Z(n18) );
  BUFFD0 U23 ( .I(n18), .Z(n19) );
  BUFFD0 U24 ( .I(n19), .Z(n20) );
  BUFFD0 U25 ( .I(n20), .Z(n21) );
  BUFFD0 U26 ( .I(n21), .Z(n22) );
  BUFFD0 U27 ( .I(n22), .Z(n23) );
  BUFFD0 U28 ( .I(n23), .Z(n24) );
  BUFFD0 U29 ( .I(n24), .Z(n25) );
  BUFFD0 U30 ( .I(n25), .Z(n26) );
  BUFFD0 U31 ( .I(n26), .Z(n27) );
  BUFFD0 U32 ( .I(n27), .Z(n28) );
  BUFFD0 U33 ( .I(n28), .Z(n29) );
  BUFFD0 U34 ( .I(n29), .Z(n30) );
  BUFFD0 U35 ( .I(n30), .Z(n31) );
  BUFFD0 U36 ( .I(n31), .Z(n32) );
  BUFFD0 U37 ( .I(n32), .Z(n33) );
  BUFFD0 U38 ( .I(n33), .Z(n34) );
  BUFFD0 U39 ( .I(n34), .Z(n35) );
  BUFFD0 U40 ( .I(n35), .Z(n36) );
  BUFFD0 U41 ( .I(n36), .Z(n37) );
  BUFFD0 U42 ( .I(n37), .Z(n38) );
  BUFFD0 U43 ( .I(n38), .Z(n39) );
  BUFFD0 U44 ( .I(n39), .Z(n40) );
  BUFFD0 U45 ( .I(n40), .Z(n41) );
  BUFFD0 U46 ( .I(n41), .Z(n42) );
  BUFFD0 U47 ( .I(n42), .Z(n43) );
  BUFFD0 U48 ( .I(n43), .Z(n44) );
  BUFFD0 U49 ( .I(n44), .Z(n45) );
  BUFFD0 U50 ( .I(n45), .Z(n46) );
  BUFFD0 U51 ( .I(n46), .Z(n47) );
  BUFFD0 U52 ( .I(n47), .Z(n48) );
  BUFFD0 U53 ( .I(n48), .Z(n49) );
  BUFFD0 U54 ( .I(n49), .Z(n50) );
  BUFFD0 U55 ( .I(n50), .Z(n51) );
  BUFFD0 U56 ( .I(n51), .Z(n52) );
  BUFFD0 U57 ( .I(n52), .Z(n53) );
  BUFFD0 U58 ( .I(n53), .Z(n54) );
  BUFFD0 U59 ( .I(n54), .Z(n55) );
  BUFFD0 U60 ( .I(n55), .Z(n56) );
  BUFFD0 U61 ( .I(n56), .Z(n57) );
  BUFFD0 U62 ( .I(n57), .Z(n58) );
  BUFFD0 U63 ( .I(n58), .Z(n59) );
  BUFFD0 U64 ( .I(n59), .Z(n60) );
  BUFFD0 U65 ( .I(n60), .Z(n61) );
  BUFFD0 U66 ( .I(n61), .Z(n62) );
  BUFFD0 U67 ( .I(n62), .Z(n63) );
  BUFFD0 U68 ( .I(n63), .Z(n64) );
  BUFFD0 U69 ( .I(n64), .Z(n65) );
  BUFFD0 U70 ( .I(n65), .Z(n66) );
  BUFFD0 U71 ( .I(n66), .Z(n67) );
  BUFFD0 U72 ( .I(n67), .Z(n68) );
  BUFFD0 U73 ( .I(n68), .Z(n69) );
  BUFFD0 U74 ( .I(n69), .Z(n70) );
  BUFFD0 U75 ( .I(n70), .Z(n71) );
  BUFFD0 U76 ( .I(n71), .Z(n72) );
  BUFFD0 U77 ( .I(n72), .Z(n73) );
  BUFFD0 U78 ( .I(n73), .Z(n74) );
  BUFFD0 U79 ( .I(n74), .Z(n75) );
  BUFFD0 U80 ( .I(n75), .Z(n76) );
  BUFFD0 U81 ( .I(n76), .Z(n77) );
  BUFFD0 U82 ( .I(n77), .Z(n78) );
  BUFFD0 U83 ( .I(n78), .Z(n79) );
  BUFFD0 U84 ( .I(n79), .Z(n80) );
  BUFFD0 U85 ( .I(n80), .Z(n81) );
  BUFFD0 U86 ( .I(n81), .Z(n82) );
  BUFFD0 U87 ( .I(n82), .Z(n83) );
  BUFFD0 U88 ( .I(n83), .Z(n84) );
  BUFFD0 U89 ( .I(n84), .Z(n85) );
  BUFFD0 U90 ( .I(n87), .Z(n199) );
  INVD0 U91 ( .I(n86), .ZN(n87) );
  CKNXD16 U92 ( .I(Din[30]), .ZN(n86) );
  BUFFD0 U93 ( .I(n89), .Z(n198) );
  INVD0 U94 ( .I(n88), .ZN(n89) );
  CKNXD16 U95 ( .I(Din[29]), .ZN(n88) );
  BUFFD0 U96 ( .I(n91), .Z(n197) );
  INVD0 U97 ( .I(n90), .ZN(n91) );
  CKNXD16 U98 ( .I(Din[28]), .ZN(n90) );
  BUFFD0 U99 ( .I(n93), .Z(n193) );
  INVD0 U100 ( .I(n92), .ZN(n93) );
  CKNXD16 U101 ( .I(Din[24]), .ZN(n92) );
  BUFFD0 U102 ( .I(n95), .Z(n192) );
  INVD0 U103 ( .I(n94), .ZN(n95) );
  CKNXD16 U104 ( .I(Din[23]), .ZN(n94) );
  BUFFD0 U105 ( .I(n97), .Z(n191) );
  INVD0 U106 ( .I(n96), .ZN(n97) );
  CKNXD16 U107 ( .I(Din[22]), .ZN(n96) );
  BUFFD0 U108 ( .I(n99), .Z(n190) );
  INVD0 U109 ( .I(n98), .ZN(n99) );
  CKNXD16 U110 ( .I(Din[21]), .ZN(n98) );
  BUFFD0 U111 ( .I(n101), .Z(n189) );
  INVD0 U112 ( .I(n100), .ZN(n101) );
  CKNXD16 U113 ( .I(Din[20]), .ZN(n100) );
  INVD0 U114 ( .I(n102), .ZN(n103) );
  CKNXD16 U115 ( .I(Din[19]), .ZN(n102) );
  INVD0 U116 ( .I(n104), .ZN(n105) );
  CKNXD16 U117 ( .I(Din[18]), .ZN(n104) );
  INVD0 U118 ( .I(n106), .ZN(n107) );
  CKNXD16 U119 ( .I(Din[17]), .ZN(n106) );
  BUFFD0 U120 ( .I(n109), .Z(n185) );
  INVD0 U121 ( .I(n108), .ZN(n109) );
  CKNXD16 U122 ( .I(Din[16]), .ZN(n108) );
  BUFFD0 U123 ( .I(n111), .Z(n184) );
  INVD0 U124 ( .I(n110), .ZN(n111) );
  CKNXD16 U125 ( .I(Din[15]), .ZN(n110) );
  BUFFD0 U126 ( .I(n113), .Z(n183) );
  INVD0 U127 ( .I(n112), .ZN(n113) );
  CKNXD16 U128 ( .I(Din[14]), .ZN(n112) );
  BUFFD0 U129 ( .I(n115), .Z(n182) );
  INVD0 U130 ( .I(n114), .ZN(n115) );
  CKNXD16 U131 ( .I(Din[13]), .ZN(n114) );
  INVD0 U132 ( .I(n116), .ZN(n117) );
  CKNXD16 U133 ( .I(Din[12]), .ZN(n116) );
  INVD0 U134 ( .I(n118), .ZN(n119) );
  CKNXD16 U135 ( .I(Din[11]), .ZN(n118) );
  INVD0 U136 ( .I(n120), .ZN(n121) );
  CKNXD16 U137 ( .I(Din[10]), .ZN(n120) );
  BUFFD0 U138 ( .I(n123), .Z(n179) );
  INVD0 U139 ( .I(n122), .ZN(n123) );
  CKNXD16 U140 ( .I(Din[9]), .ZN(n122) );
  BUFFD0 U141 ( .I(n125), .Z(n178) );
  INVD0 U142 ( .I(n124), .ZN(n125) );
  CKNXD16 U143 ( .I(Din[8]), .ZN(n124) );
  BUFFD0 U144 ( .I(n127), .Z(n177) );
  INVD0 U145 ( .I(n126), .ZN(n127) );
  CKNXD16 U146 ( .I(Din[7]), .ZN(n126) );
  BUFFD0 U147 ( .I(n129), .Z(n176) );
  INVD0 U148 ( .I(n128), .ZN(n129) );
  CKNXD16 U149 ( .I(Din[6]), .ZN(n128) );
  INVD0 U150 ( .I(n130), .ZN(n131) );
  CKNXD16 U151 ( .I(Din[5]), .ZN(n130) );
  INVD0 U152 ( .I(n132), .ZN(n133) );
  CKNXD16 U153 ( .I(Din[4]), .ZN(n132) );
  INVD0 U154 ( .I(n134), .ZN(n135) );
  CKNXD16 U155 ( .I(Din[3]), .ZN(n134) );
  INVD0 U156 ( .I(n136), .ZN(n137) );
  INVD0 U157 ( .I(n138), .ZN(n139) );
  CKNXD16 U158 ( .I(Din[1]), .ZN(n138) );
  INVD0 U159 ( .I(n140), .ZN(n141) );
  CKNXD16 U160 ( .I(Din[0]), .ZN(n140) );
  BUFFD0 U161 ( .I(n143), .Z(n196) );
  INVD0 U162 ( .I(n142), .ZN(n143) );
  CKNXD16 U163 ( .I(Din[27]), .ZN(n142) );
  BUFFD0 U164 ( .I(n145), .Z(n194) );
  INVD0 U165 ( .I(n144), .ZN(n145) );
  CKNXD16 U166 ( .I(Din[25]), .ZN(n144) );
  BUFFD0 U167 ( .I(n147), .Z(n195) );
  INVD0 U168 ( .I(n146), .ZN(n147) );
  CKNXD16 U169 ( .I(Din[26]), .ZN(n146) );
  BUFFD0 U170 ( .I(n149), .Z(n148) );
  BUFFD0 U171 ( .I(n150), .Z(n149) );
  BUFFD0 U172 ( .I(n151), .Z(n150) );
  BUFFD0 U173 ( .I(n152), .Z(n151) );
  BUFFD0 U174 ( .I(n153), .Z(n152) );
  BUFFD0 U175 ( .I(n154), .Z(n153) );
  BUFFD0 U176 ( .I(n155), .Z(n154) );
  BUFFD0 U177 ( .I(n156), .Z(n155) );
  BUFFD0 U178 ( .I(n157), .Z(n156) );
  BUFFD0 U179 ( .I(n166), .Z(n157) );
  BUFFD0 U180 ( .I(n159), .Z(n158) );
  BUFFD0 U181 ( .I(n160), .Z(n159) );
  BUFFD0 U182 ( .I(n162), .Z(n160) );
  INVD0 U183 ( .I(n161), .ZN(n162) );
  CKNXD16 U184 ( .I(n163), .ZN(n161) );
  CKNXD16 U185 ( .I(n164), .ZN(n165) );
  INVD0 U186 ( .I(WriteIn), .ZN(n164) );
  BUFFD0 U187 ( .I(n165), .Z(n163) );
  CKBD0 U188 ( .CLK(SM_MemReadCmd), .C(n169) );
  BUFFD0 U189 ( .I(n168), .Z(n166) );
  BUFFD1 U190 ( .I(n85), .Z(n200) );
  BUFFD1 U191 ( .I(n141), .Z(n170) );
  BUFFD1 U192 ( .I(n139), .Z(n171) );
  BUFFD1 U193 ( .I(n135), .Z(n173) );
  BUFFD1 U194 ( .I(n133), .Z(n174) );
  BUFFD1 U195 ( .I(n131), .Z(n175) );
  BUFFD1 U196 ( .I(n121), .Z(n180) );
  BUFFD1 U197 ( .I(n119), .Z(n181) );
  BUFFD1 U198 ( .I(n107), .Z(n186) );
  BUFFD1 U199 ( .I(n105), .Z(n187) );
  BUFFD1 U200 ( .I(n103), .Z(n188) );
  BUFFD1 U201 ( .I(ReadIn), .Z(n168) );
  TIEH U202 ( .Z(\*Logic1* ) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n1397, n1398, n1399, n1400, n1401, n1402, n1403, StateClockRaw,
         StateClock, N44, N45, N46, N47, N48, N49, N51, N52, N54, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N176, N177, N178, N330, N332,
         N333, N334, n6, n8, n9, n12, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98,
         n99, n100, n103, n104, n105, n106, n107, n108, n109, n121, n123, n124,
         n127, n128, n130, n131, n132, n134, n135, n138, n139, n140, n143,
         \add_389/carry[2] , \add_389/carry[3] , \add_389/carry[4] ,
         \add_308/carry[3] , \add_308/carry[4] , n1, n2, n3, n4, n5, n7, n10,
         n11, n13, n14, n69, n70, n71, n84, n85, n92, n101, n102, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n125,
         n126, n129, n133, n136, n137, n141, n142, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1368, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1390, n1392, n1393, n1395,
         n1396;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [4:0] OldReadAr;
  wire   [4:0] OldWriteAr;
  assign WriteAddr[0] = N330;
  assign WriteAddr[1] = \add_389/carry[2] ;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  MOAI22D1 U24 ( .A1(n29), .A2(n30), .B1(n31), .B2(CurState[2]), .ZN(n27) );
  OR3D1 U41 ( .A1(n49), .A2(CurState[2]), .A3(n50), .Z(n47) );
  OA21D1 U111 ( .A1(CurState[2]), .A2(n29), .B(n83), .Z(n35) );
  FIFOStateM_AWid5_DW01_inc_0 r110 ( .A({WriteAddr[4:2], \add_389/carry[2] , 
        n747}), .SUM({N72, N71, N70, N69, N68}) );
  FIFOStateM_AWid5_DW01_inc_1 r109 ( .A({ReadAddr[4], n657, n617, n788, n821}), 
        .SUM({N48, N47, N46, N45, N44}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n2), .CPN(StateClock), .CDN(n1390), .QN(n291) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n294), .CPN(StateClock), .CDN(n143), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n3), .CPN(StateClock), .CDN(n1390), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n877), .CPN(StateClock), .CDN(n1390), .QN(
        n290) );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n4), .CPN(StateClock), .CDN(n1390), .Q(
        OldWriteAr[4]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n13), .CPN(StateClock), .CDN(n143), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n71), .CPN(StateClock), .CDN(n1390), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n327), .CPN(StateClock), .CDN(n1390), .Q(
        OldReadAr[4]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n329), .CPN(StateClock), .CDN(n1390), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n331), .CPN(StateClock), .CDN(n1390), .Q(
        OldReadAr[3]) );
  DFNCND1 \NextState_reg[1]  ( .D(n101), .CPN(StateClock), .CDN(n143), .Q(
        NextState[1]), .QN(n124) );
  DFNCND1 \NextState_reg[0]  ( .D(n115), .CPN(StateClock), .CDN(n1390), .Q(
        NextState[0]), .QN(n123) );
  DFNCND1 \NextState_reg[2]  ( .D(n340), .CPN(StateClock), .CDN(n143), .Q(
        NextState[2]), .QN(n121) );
  DFNCND1 ReadCmdr_reg ( .D(n119), .CPN(StateClock), .CDN(n143), .Q(n1402) );
  DFNCND1 WriteCmdr_reg ( .D(n125), .CPN(StateClock), .CDN(n1390), .Q(n1403)
         );
  EDFCNQD1 \WriteAr_reg[4]  ( .D(n378), .E(n1275), .CP(StateClock), .CDN(n1390), .Q(WriteAddr[4]) );
  EDFCNQD1 \WriteAr_reg[3]  ( .D(n430), .E(n1275), .CP(StateClock), .CDN(n1390), .Q(WriteAddr[3]) );
  EDFCNQD1 \ReadAr_reg[2]  ( .D(n484), .E(n1358), .CP(StateClock), .CDN(n1390), 
        .Q(n1398) );
  EDFCNQD1 \ReadAr_reg[4]  ( .D(n524), .E(n1358), .CP(StateClock), .CDN(n143), 
        .Q(n1397) );
  EDFCNQD1 \WriteAr_reg[2]  ( .D(n565), .E(n1275), .CP(StateClock), .CDN(n1390), .Q(n1399) );
  EDFCNQD1 \ReadAr_reg[3]  ( .D(n619), .E(n1358), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[3]) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(n658), .E(n1275), .CP(StateClock), .CDN(n143), 
        .Q(\add_389/carry[2] ) );
  EDFCNQD1 \WriteAr_reg[0]  ( .D(n710), .E(n1275), .CP(StateClock), .CDN(n143), 
        .Q(N330) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[2]), .QN(n96) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[1]), .QN(n29) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n143), 
        .Q(CurState[0]), .QN(n55) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n148), .E(n1358), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[1]), .QN(n1395) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n791), .E(n1358), .CP(StateClock), .CDN(n143), 
        .Q(ReadAddr[0]), .QN(n1392) );
  DFND1 FullFIFOr_reg ( .D(n161), .CPN(StateClock), .Q(n1401) );
  DFND1 EmptyFIFOr_reg ( .D(n218), .CPN(StateClock), .Q(n1400) );
  CKND12 U3 ( .CLK(n836), .CN(n837) );
  INVD0 U4 ( .I(n838), .ZN(n839) );
  CKND12 U5 ( .CLK(n843), .CN(n838) );
  INVD0 U6 ( .I(n842), .ZN(n843) );
  CKNXD16 U7 ( .I(n841), .ZN(n842) );
  CKBD0 U8 ( .CLK(n840), .C(n841) );
  CKNXD16 U9 ( .I(n279), .ZN(n840) );
  INVD1 U10 ( .I(n823), .ZN(n1) );
  INVD1 U11 ( .I(n1), .ZN(n2) );
  CKND12 U12 ( .CLK(n875), .CN(n876) );
  BUFFD0 U13 ( .I(n852), .Z(n3) );
  BUFFD0 U14 ( .I(n5), .Z(n4) );
  BUFFD0 U15 ( .I(n7), .Z(n5) );
  BUFFD0 U16 ( .I(n10), .Z(n7) );
  BUFFD0 U17 ( .I(n11), .Z(n10) );
  BUFFD0 U18 ( .I(n324), .Z(n11) );
  BUFFD0 U19 ( .I(n14), .Z(n13) );
  BUFFD0 U20 ( .I(n69), .Z(n14) );
  BUFFD0 U21 ( .I(n70), .Z(n69) );
  BUFFD0 U22 ( .I(n325), .Z(n70) );
  BUFFD0 U23 ( .I(n84), .Z(n71) );
  BUFFD0 U25 ( .I(n85), .Z(n84) );
  BUFFD0 U26 ( .I(n92), .Z(n85) );
  BUFFD0 U27 ( .I(n326), .Z(n92) );
  BUFFD0 U28 ( .I(n1194), .Z(n1195) );
  BUFFD0 U29 ( .I(n102), .Z(n101) );
  BUFFD0 U30 ( .I(n110), .Z(n102) );
  BUFFD0 U31 ( .I(n111), .Z(n110) );
  BUFFD0 U32 ( .I(n112), .Z(n111) );
  BUFFD0 U33 ( .I(n113), .Z(n112) );
  BUFFD0 U34 ( .I(n114), .Z(n113) );
  BUFFD0 U35 ( .I(n1181), .Z(n114) );
  INVD3 U36 ( .I(n277), .ZN(n140) );
  BUFFD0 U37 ( .I(n116), .Z(n115) );
  BUFFD0 U38 ( .I(n117), .Z(n116) );
  BUFFD0 U39 ( .I(n333), .Z(n117) );
  OA21D0 U40 ( .A1(n24), .A2(n123), .B(n42), .Z(n277) );
  CKXOR2D0 U42 ( .A1(ReadAddr[1]), .A2(n290), .Z(n104) );
  CKBD0 U43 ( .CLK(n291), .C(n118) );
  BUFFD0 U44 ( .I(n120), .Z(n119) );
  CKBD0 U45 ( .CLK(n1241), .C(n120) );
  OAI32D0 U46 ( .A1(n97), .A2(n98), .A3(n95), .B1(n99), .B2(n100), .ZN(n278)
         );
  ND3D0 U47 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n23) );
  BUFFD0 U48 ( .I(n346), .Z(n122) );
  BUFFD0 U49 ( .I(n145), .Z(n125) );
  BUFFD0 U50 ( .I(n136), .Z(n126) );
  BUFFD0 U51 ( .I(n137), .Z(n129) );
  CKXOR2D0 U52 ( .A1(\add_389/carry[2] ), .A2(n870), .Z(n37) );
  BUFFD0 U53 ( .I(n141), .Z(n133) );
  BUFFD0 U54 ( .I(n142), .Z(n136) );
  BUFFD0 U55 ( .I(n144), .Z(n137) );
  BUFFD0 U56 ( .I(n375), .Z(n141) );
  BUFFD0 U57 ( .I(n377), .Z(n142) );
  BUFFD0 U58 ( .I(n376), .Z(n144) );
  BUFFD0 U59 ( .I(n341), .Z(n145) );
  CKND2D0 U60 ( .A1(WriteCmd), .A2(n1288), .ZN(n34) );
  BUFFD0 U61 ( .I(n285), .Z(n146) );
  BUFFD0 U62 ( .I(n146), .Z(n147) );
  BUFFD0 U63 ( .I(n150), .Z(n148) );
  BUFFD0 U64 ( .I(n1346), .Z(n149) );
  BUFFD0 U65 ( .I(n151), .Z(n150) );
  BUFFD0 U66 ( .I(n152), .Z(n151) );
  BUFFD0 U67 ( .I(n153), .Z(n152) );
  BUFFD0 U68 ( .I(n154), .Z(n153) );
  BUFFD0 U69 ( .I(n155), .Z(n154) );
  BUFFD0 U70 ( .I(n156), .Z(n155) );
  BUFFD0 U71 ( .I(n760), .Z(n156) );
  BUFFD0 U72 ( .I(n1354), .Z(n157) );
  BUFFD0 U73 ( .I(n55), .Z(n158) );
  BUFFD0 U74 ( .I(n96), .Z(n159) );
  BUFFD0 U75 ( .I(n284), .Z(n160) );
  BUFFD0 U76 ( .I(n164), .Z(n161) );
  BUFFD0 U77 ( .I(n132), .Z(n162) );
  BUFFD0 U78 ( .I(n162), .Z(n163) );
  BUFFD0 U79 ( .I(n165), .Z(n164) );
  BUFFD0 U80 ( .I(n166), .Z(n165) );
  BUFFD0 U81 ( .I(n167), .Z(n166) );
  BUFFD0 U82 ( .I(n168), .Z(n167) );
  BUFFD0 U83 ( .I(n169), .Z(n168) );
  BUFFD0 U84 ( .I(n170), .Z(n169) );
  BUFFD0 U85 ( .I(n171), .Z(n170) );
  BUFFD0 U86 ( .I(n172), .Z(n171) );
  BUFFD0 U87 ( .I(n173), .Z(n172) );
  BUFFD0 U88 ( .I(n174), .Z(n173) );
  BUFFD0 U89 ( .I(n175), .Z(n174) );
  BUFFD0 U90 ( .I(n176), .Z(n175) );
  BUFFD0 U91 ( .I(n177), .Z(n176) );
  BUFFD0 U92 ( .I(n178), .Z(n177) );
  BUFFD0 U93 ( .I(n179), .Z(n178) );
  BUFFD0 U94 ( .I(n180), .Z(n179) );
  BUFFD0 U95 ( .I(n181), .Z(n180) );
  BUFFD0 U96 ( .I(n182), .Z(n181) );
  BUFFD0 U97 ( .I(n183), .Z(n182) );
  BUFFD0 U98 ( .I(n184), .Z(n183) );
  BUFFD0 U99 ( .I(n185), .Z(n184) );
  BUFFD0 U100 ( .I(n186), .Z(n185) );
  BUFFD0 U101 ( .I(n187), .Z(n186) );
  BUFFD0 U102 ( .I(n188), .Z(n187) );
  BUFFD0 U103 ( .I(n189), .Z(n188) );
  BUFFD0 U104 ( .I(n190), .Z(n189) );
  BUFFD0 U105 ( .I(n191), .Z(n190) );
  BUFFD0 U106 ( .I(n192), .Z(n191) );
  BUFFD0 U107 ( .I(n193), .Z(n192) );
  BUFFD0 U108 ( .I(n194), .Z(n193) );
  BUFFD0 U109 ( .I(n195), .Z(n194) );
  BUFFD0 U110 ( .I(n196), .Z(n195) );
  BUFFD0 U112 ( .I(n197), .Z(n196) );
  BUFFD0 U113 ( .I(n198), .Z(n197) );
  BUFFD0 U114 ( .I(n199), .Z(n198) );
  BUFFD0 U115 ( .I(n200), .Z(n199) );
  BUFFD0 U116 ( .I(n201), .Z(n200) );
  BUFFD0 U117 ( .I(n202), .Z(n201) );
  BUFFD0 U118 ( .I(n203), .Z(n202) );
  BUFFD0 U119 ( .I(n204), .Z(n203) );
  BUFFD0 U120 ( .I(n205), .Z(n204) );
  BUFFD0 U121 ( .I(n206), .Z(n205) );
  BUFFD0 U122 ( .I(n207), .Z(n206) );
  BUFFD0 U123 ( .I(n208), .Z(n207) );
  BUFFD0 U124 ( .I(n209), .Z(n208) );
  BUFFD0 U125 ( .I(n210), .Z(n209) );
  BUFFD0 U126 ( .I(n211), .Z(n210) );
  BUFFD0 U127 ( .I(n212), .Z(n211) );
  BUFFD0 U128 ( .I(n213), .Z(n212) );
  BUFFD0 U129 ( .I(n214), .Z(n213) );
  BUFFD0 U130 ( .I(n215), .Z(n214) );
  BUFFD0 U131 ( .I(n216), .Z(n215) );
  BUFFD0 U132 ( .I(n217), .Z(n216) );
  BUFFD0 U133 ( .I(n163), .Z(n217) );
  BUFFD0 U134 ( .I(n221), .Z(n218) );
  BUFFD0 U135 ( .I(n127), .Z(n219) );
  BUFFD0 U136 ( .I(n219), .Z(n220) );
  BUFFD0 U137 ( .I(n222), .Z(n221) );
  BUFFD0 U138 ( .I(n223), .Z(n222) );
  BUFFD0 U139 ( .I(n224), .Z(n223) );
  BUFFD0 U140 ( .I(n225), .Z(n224) );
  BUFFD0 U141 ( .I(n226), .Z(n225) );
  BUFFD0 U142 ( .I(n227), .Z(n226) );
  BUFFD0 U143 ( .I(n228), .Z(n227) );
  BUFFD0 U144 ( .I(n229), .Z(n228) );
  BUFFD0 U145 ( .I(n230), .Z(n229) );
  BUFFD0 U146 ( .I(n231), .Z(n230) );
  BUFFD0 U147 ( .I(n232), .Z(n231) );
  BUFFD0 U148 ( .I(n233), .Z(n232) );
  BUFFD0 U149 ( .I(n234), .Z(n233) );
  BUFFD0 U150 ( .I(n235), .Z(n234) );
  BUFFD0 U151 ( .I(n236), .Z(n235) );
  BUFFD0 U152 ( .I(n237), .Z(n236) );
  BUFFD0 U153 ( .I(n238), .Z(n237) );
  BUFFD0 U154 ( .I(n239), .Z(n238) );
  BUFFD0 U155 ( .I(n240), .Z(n239) );
  BUFFD0 U156 ( .I(n241), .Z(n240) );
  BUFFD0 U157 ( .I(n242), .Z(n241) );
  BUFFD0 U158 ( .I(n243), .Z(n242) );
  BUFFD0 U159 ( .I(n244), .Z(n243) );
  BUFFD0 U160 ( .I(n245), .Z(n244) );
  BUFFD0 U161 ( .I(n246), .Z(n245) );
  BUFFD0 U162 ( .I(n247), .Z(n246) );
  BUFFD0 U163 ( .I(n248), .Z(n247) );
  BUFFD0 U164 ( .I(n249), .Z(n248) );
  BUFFD0 U165 ( .I(n250), .Z(n249) );
  BUFFD0 U166 ( .I(n251), .Z(n250) );
  BUFFD0 U167 ( .I(n252), .Z(n251) );
  BUFFD0 U168 ( .I(n253), .Z(n252) );
  BUFFD0 U169 ( .I(n254), .Z(n253) );
  BUFFD0 U170 ( .I(n255), .Z(n254) );
  BUFFD0 U171 ( .I(n256), .Z(n255) );
  BUFFD0 U172 ( .I(n257), .Z(n256) );
  BUFFD0 U173 ( .I(n258), .Z(n257) );
  BUFFD0 U174 ( .I(n259), .Z(n258) );
  BUFFD0 U175 ( .I(n260), .Z(n259) );
  BUFFD0 U176 ( .I(n261), .Z(n260) );
  BUFFD0 U177 ( .I(n262), .Z(n261) );
  BUFFD0 U178 ( .I(n263), .Z(n262) );
  BUFFD0 U179 ( .I(n264), .Z(n263) );
  BUFFD0 U180 ( .I(n265), .Z(n264) );
  BUFFD0 U181 ( .I(n266), .Z(n265) );
  BUFFD0 U182 ( .I(n267), .Z(n266) );
  BUFFD0 U183 ( .I(n268), .Z(n267) );
  BUFFD0 U184 ( .I(n269), .Z(n268) );
  BUFFD0 U185 ( .I(n270), .Z(n269) );
  BUFFD0 U186 ( .I(n271), .Z(n270) );
  BUFFD0 U187 ( .I(n272), .Z(n271) );
  BUFFD0 U188 ( .I(n273), .Z(n272) );
  BUFFD0 U189 ( .I(n274), .Z(n273) );
  BUFFD0 U190 ( .I(n220), .Z(n274) );
  NR2D1 U191 ( .A1(n149), .A2(n99), .ZN(n275) );
  OA32D0 U192 ( .A1(n122), .A2(n32), .A3(n33), .B1(n34), .B2(n22), .Z(n276) );
  INVD1 U193 ( .I(n276), .ZN(n139) );
  INVD1 U194 ( .I(n1345), .ZN(n1346) );
  OA22D0 U195 ( .A1(n8), .A2(n118), .B1(n1392), .B2(n9), .Z(n279) );
  OA22D0 U196 ( .A1(n24), .A2(n124), .B1(n25), .B2(n57), .Z(n280) );
  AOI22D0 U197 ( .A1(WriteAddr[3]), .A2(n16), .B1(n17), .B2(n129), .ZN(n281)
         );
  AOI22D0 U198 ( .A1(WriteAddr[2]), .A2(n16), .B1(n17), .B2(n126), .ZN(n282)
         );
  AOI22D0 U199 ( .A1(WriteAddr[4]), .A2(n16), .B1(n17), .B2(n133), .ZN(n283)
         );
  AN2D1 U200 ( .A1(n1354), .A2(n99), .Z(n284) );
  AN3D1 U201 ( .A1(n1288), .A2(n157), .A3(n34), .Z(n285) );
  OAI31D0 U202 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(n1400), 
        .ZN(n286) );
  IND2D1 U203 ( .A1(Reset), .B1(n289), .ZN(n1372) );
  CKNXD12 U204 ( .I(OldWriteAr[1]), .ZN(n18) );
  CKND2D0 U205 ( .A1(n1372), .A2(n1401), .ZN(n287) );
  OA22D0 U206 ( .A1(n8), .A2(n290), .B1(n1395), .B2(n9), .Z(n288) );
  AO21D1 U207 ( .A1(CurState[2]), .A2(CurState[0]), .B(n15), .Z(n289) );
  BUFFD16 U208 ( .I(n848), .Z(n849) );
  BUFFD0 U209 ( .I(n295), .Z(n294) );
  BUFFD0 U210 ( .I(n296), .Z(n295) );
  BUFFD0 U211 ( .I(n297), .Z(n296) );
  BUFFD0 U212 ( .I(n298), .Z(n297) );
  BUFFD0 U213 ( .I(n299), .Z(n298) );
  BUFFD0 U214 ( .I(n300), .Z(n299) );
  BUFFD0 U215 ( .I(n302), .Z(n300) );
  BUFFD0 U216 ( .I(n305), .Z(n301) );
  BUFFD0 U217 ( .I(n303), .Z(n302) );
  BUFFD0 U218 ( .I(n304), .Z(n303) );
  BUFFD0 U219 ( .I(n308), .Z(n304) );
  BUFFD0 U220 ( .I(n306), .Z(n305) );
  BUFFD0 U221 ( .I(n307), .Z(n306) );
  ND3D0 U222 ( .A1(n22), .A2(n346), .A3(WriteReq), .ZN(n17) );
  BUFFD0 U223 ( .I(n844), .Z(n307) );
  BUFFD0 U224 ( .I(n309), .Z(n308) );
  BUFFD0 U225 ( .I(n310), .Z(n309) );
  BUFFD0 U226 ( .I(n311), .Z(n310) );
  BUFFD0 U227 ( .I(n312), .Z(n311) );
  BUFFD0 U228 ( .I(n313), .Z(n312) );
  BUFFD0 U229 ( .I(n314), .Z(n313) );
  BUFFD0 U230 ( .I(n315), .Z(n314) );
  BUFFD0 U231 ( .I(n316), .Z(n315) );
  BUFFD0 U232 ( .I(n317), .Z(n316) );
  BUFFD0 U233 ( .I(n318), .Z(n317) );
  BUFFD0 U234 ( .I(n319), .Z(n318) );
  BUFFD0 U235 ( .I(n320), .Z(n319) );
  BUFFD0 U236 ( .I(n321), .Z(n320) );
  BUFFD0 U237 ( .I(n322), .Z(n321) );
  BUFFD0 U238 ( .I(n20), .Z(n844) );
  INVD12 U239 ( .I(n135), .ZN(n847) );
  BUFFD0 U240 ( .I(n846), .Z(n322) );
  BUFFD0 U241 ( .I(OldWriteAr[0]), .Z(n323) );
  BUFFD0 U242 ( .I(n902), .Z(n324) );
  BUFFD0 U243 ( .I(n919), .Z(n325) );
  BUFFD0 U244 ( .I(n936), .Z(n326) );
  BUFFD0 U245 ( .I(n328), .Z(n327) );
  CKBD0 U246 ( .CLK(n953), .C(n328) );
  BUFFD0 U247 ( .I(n330), .Z(n329) );
  CKBD0 U248 ( .CLK(n971), .C(n330) );
  BUFFD0 U249 ( .I(n332), .Z(n331) );
  CKBD0 U250 ( .CLK(n989), .C(n332) );
  BUFFD0 U251 ( .I(n334), .Z(n333) );
  BUFFD0 U252 ( .I(n335), .Z(n334) );
  BUFFD0 U253 ( .I(n336), .Z(n335) );
  BUFFD0 U254 ( .I(n337), .Z(n336) );
  BUFFD0 U255 ( .I(n338), .Z(n337) );
  CKBD0 U256 ( .CLK(n1199), .C(n338) );
  INVD10 U257 ( .I(n339), .ZN(n340) );
  CKNXD0 U258 ( .I(n1219), .ZN(n339) );
  INVD0 U259 ( .I(n1239), .ZN(n1236) );
  INVD0 U260 ( .I(n1224), .ZN(n1225) );
  CKND8 U261 ( .CLK(n138), .CN(n1224) );
  OAI22D0 U262 ( .A1(n24), .A2(n121), .B1(n25), .B2(n26), .ZN(n138) );
  BUFFD0 U263 ( .I(n342), .Z(n341) );
  BUFFD0 U264 ( .I(n343), .Z(n342) );
  BUFFD0 U265 ( .I(n344), .Z(n343) );
  BUFFD0 U266 ( .I(n345), .Z(n344) );
  BUFFD0 U267 ( .I(n347), .Z(n345) );
  BUFFD0 U268 ( .I(n23), .Z(n346) );
  BUFFD0 U269 ( .I(n348), .Z(n347) );
  BUFFD0 U270 ( .I(n349), .Z(n348) );
  BUFFD0 U271 ( .I(n350), .Z(n349) );
  BUFFD0 U272 ( .I(n351), .Z(n350) );
  BUFFD0 U273 ( .I(n352), .Z(n351) );
  BUFFD0 U274 ( .I(n353), .Z(n352) );
  BUFFD0 U275 ( .I(n354), .Z(n353) );
  BUFFD0 U276 ( .I(n355), .Z(n354) );
  BUFFD0 U277 ( .I(n356), .Z(n355) );
  BUFFD0 U278 ( .I(n357), .Z(n356) );
  BUFFD0 U279 ( .I(n358), .Z(n357) );
  BUFFD0 U280 ( .I(n359), .Z(n358) );
  BUFFD0 U281 ( .I(n360), .Z(n359) );
  BUFFD0 U282 ( .I(n361), .Z(n360) );
  BUFFD0 U283 ( .I(n362), .Z(n361) );
  BUFFD0 U284 ( .I(n363), .Z(n362) );
  BUFFD0 U285 ( .I(n364), .Z(n363) );
  BUFFD0 U286 ( .I(n365), .Z(n364) );
  BUFFD0 U287 ( .I(n366), .Z(n365) );
  BUFFD0 U288 ( .I(n367), .Z(n366) );
  BUFFD0 U289 ( .I(n368), .Z(n367) );
  BUFFD0 U290 ( .I(n369), .Z(n368) );
  BUFFD0 U291 ( .I(n370), .Z(n369) );
  BUFFD0 U292 ( .I(n371), .Z(n370) );
  BUFFD0 U293 ( .I(n372), .Z(n371) );
  BUFFD0 U294 ( .I(n373), .Z(n372) );
  BUFFD0 U295 ( .I(n374), .Z(n373) );
  CKBD0 U296 ( .CLK(n1264), .C(n374) );
  XOR2D0 U297 ( .A1(WriteAddr[2]), .A2(n126), .Z(n40) );
  BUFFD0 U298 ( .I(OldWriteAr[4]), .Z(n375) );
  BUFFD0 U299 ( .I(OldWriteAr[3]), .Z(n376) );
  XOR2D0 U300 ( .A1(WriteAddr[4]), .A2(n133), .Z(n41) );
  BUFFD0 U301 ( .I(OldWriteAr[2]), .Z(n377) );
  XOR2D0 U302 ( .A1(WriteAddr[3]), .A2(n129), .Z(n39) );
  CKBD0 U303 ( .CLK(n379), .C(n380) );
  CKBD0 U304 ( .CLK(N77), .C(n379) );
  BUFFD0 U305 ( .I(n382), .Z(n378) );
  BUFFD0 U306 ( .I(n380), .Z(n381) );
  BUFFD0 U307 ( .I(n383), .Z(n382) );
  BUFFD0 U308 ( .I(n384), .Z(n383) );
  BUFFD0 U309 ( .I(n385), .Z(n384) );
  BUFFD0 U310 ( .I(n386), .Z(n385) );
  BUFFD0 U311 ( .I(n387), .Z(n386) );
  BUFFD0 U312 ( .I(n388), .Z(n387) );
  BUFFD0 U313 ( .I(n389), .Z(n388) );
  BUFFD0 U314 ( .I(n390), .Z(n389) );
  BUFFD0 U315 ( .I(n391), .Z(n390) );
  BUFFD0 U316 ( .I(n392), .Z(n391) );
  BUFFD0 U317 ( .I(n393), .Z(n392) );
  BUFFD0 U318 ( .I(n394), .Z(n393) );
  BUFFD0 U319 ( .I(n395), .Z(n394) );
  BUFFD0 U320 ( .I(n396), .Z(n395) );
  BUFFD0 U321 ( .I(n397), .Z(n396) );
  BUFFD0 U322 ( .I(n398), .Z(n397) );
  BUFFD0 U323 ( .I(n399), .Z(n398) );
  BUFFD0 U324 ( .I(n400), .Z(n399) );
  BUFFD0 U325 ( .I(n401), .Z(n400) );
  BUFFD0 U326 ( .I(n402), .Z(n401) );
  BUFFD0 U327 ( .I(n403), .Z(n402) );
  BUFFD0 U328 ( .I(n404), .Z(n403) );
  BUFFD0 U329 ( .I(n405), .Z(n404) );
  BUFFD0 U330 ( .I(n406), .Z(n405) );
  BUFFD0 U331 ( .I(n407), .Z(n406) );
  BUFFD0 U332 ( .I(n408), .Z(n407) );
  BUFFD0 U333 ( .I(n409), .Z(n408) );
  BUFFD0 U334 ( .I(n410), .Z(n409) );
  BUFFD0 U335 ( .I(n411), .Z(n410) );
  BUFFD0 U336 ( .I(n412), .Z(n411) );
  BUFFD0 U337 ( .I(n413), .Z(n412) );
  BUFFD0 U338 ( .I(n414), .Z(n413) );
  BUFFD0 U339 ( .I(n415), .Z(n414) );
  BUFFD0 U340 ( .I(n416), .Z(n415) );
  BUFFD0 U341 ( .I(n417), .Z(n416) );
  BUFFD0 U342 ( .I(n418), .Z(n417) );
  BUFFD0 U343 ( .I(n419), .Z(n418) );
  BUFFD0 U344 ( .I(n420), .Z(n419) );
  BUFFD0 U345 ( .I(n421), .Z(n420) );
  BUFFD0 U346 ( .I(n422), .Z(n421) );
  BUFFD0 U347 ( .I(n423), .Z(n422) );
  BUFFD0 U348 ( .I(n424), .Z(n423) );
  BUFFD0 U349 ( .I(n425), .Z(n424) );
  BUFFD0 U350 ( .I(n426), .Z(n425) );
  BUFFD0 U351 ( .I(n427), .Z(n426) );
  BUFFD0 U352 ( .I(n428), .Z(n427) );
  BUFFD0 U353 ( .I(n429), .Z(n428) );
  BUFFD0 U354 ( .I(n381), .Z(n429) );
  BUFFD0 U355 ( .I(n436), .Z(n430) );
  BUFFD0 U356 ( .I(N76), .Z(n431) );
  BUFFD0 U357 ( .I(n431), .Z(n432) );
  BUFFD0 U358 ( .I(n432), .Z(n433) );
  BUFFD0 U359 ( .I(n433), .Z(n434) );
  BUFFD0 U360 ( .I(n434), .Z(n435) );
  BUFFD0 U361 ( .I(n437), .Z(n436) );
  BUFFD0 U362 ( .I(n438), .Z(n437) );
  BUFFD0 U363 ( .I(n439), .Z(n438) );
  BUFFD0 U364 ( .I(n440), .Z(n439) );
  BUFFD0 U365 ( .I(n441), .Z(n440) );
  BUFFD0 U366 ( .I(n442), .Z(n441) );
  BUFFD0 U367 ( .I(n443), .Z(n442) );
  BUFFD0 U368 ( .I(n444), .Z(n443) );
  BUFFD0 U369 ( .I(n445), .Z(n444) );
  BUFFD0 U370 ( .I(n446), .Z(n445) );
  BUFFD0 U371 ( .I(n447), .Z(n446) );
  BUFFD0 U372 ( .I(n448), .Z(n447) );
  BUFFD0 U373 ( .I(n449), .Z(n448) );
  BUFFD0 U374 ( .I(n450), .Z(n449) );
  BUFFD0 U375 ( .I(n451), .Z(n450) );
  BUFFD0 U376 ( .I(n452), .Z(n451) );
  BUFFD0 U377 ( .I(n453), .Z(n452) );
  BUFFD0 U378 ( .I(n454), .Z(n453) );
  BUFFD0 U379 ( .I(n455), .Z(n454) );
  BUFFD0 U380 ( .I(n456), .Z(n455) );
  BUFFD0 U381 ( .I(n457), .Z(n456) );
  BUFFD0 U382 ( .I(n458), .Z(n457) );
  BUFFD0 U383 ( .I(n459), .Z(n458) );
  BUFFD0 U384 ( .I(n460), .Z(n459) );
  BUFFD0 U385 ( .I(n461), .Z(n460) );
  BUFFD0 U386 ( .I(n462), .Z(n461) );
  BUFFD0 U387 ( .I(n463), .Z(n462) );
  BUFFD0 U388 ( .I(n464), .Z(n463) );
  BUFFD0 U389 ( .I(n465), .Z(n464) );
  BUFFD0 U390 ( .I(n466), .Z(n465) );
  BUFFD0 U391 ( .I(n467), .Z(n466) );
  BUFFD0 U392 ( .I(n468), .Z(n467) );
  BUFFD0 U393 ( .I(n469), .Z(n468) );
  BUFFD0 U394 ( .I(n470), .Z(n469) );
  BUFFD0 U395 ( .I(n471), .Z(n470) );
  BUFFD0 U396 ( .I(n472), .Z(n471) );
  BUFFD0 U397 ( .I(n473), .Z(n472) );
  BUFFD0 U398 ( .I(n474), .Z(n473) );
  BUFFD0 U399 ( .I(n475), .Z(n474) );
  BUFFD0 U400 ( .I(n476), .Z(n475) );
  BUFFD0 U401 ( .I(n477), .Z(n476) );
  BUFFD0 U402 ( .I(n478), .Z(n477) );
  BUFFD0 U403 ( .I(n479), .Z(n478) );
  BUFFD0 U404 ( .I(n480), .Z(n479) );
  BUFFD0 U405 ( .I(n481), .Z(n480) );
  BUFFD0 U406 ( .I(n482), .Z(n481) );
  BUFFD0 U407 ( .I(n483), .Z(n482) );
  BUFFD0 U408 ( .I(n435), .Z(n483) );
  BUFFD0 U409 ( .I(n485), .Z(n484) );
  BUFFD0 U410 ( .I(n486), .Z(n485) );
  BUFFD0 U411 ( .I(n487), .Z(n486) );
  BUFFD0 U412 ( .I(n488), .Z(n487) );
  BUFFD0 U413 ( .I(n489), .Z(n488) );
  BUFFD0 U414 ( .I(n490), .Z(n489) );
  BUFFD0 U415 ( .I(n491), .Z(n490) );
  BUFFD0 U416 ( .I(n492), .Z(n491) );
  BUFFD0 U417 ( .I(n493), .Z(n492) );
  BUFFD0 U418 ( .I(n494), .Z(n493) );
  BUFFD0 U419 ( .I(n495), .Z(n494) );
  BUFFD0 U420 ( .I(n496), .Z(n495) );
  BUFFD0 U421 ( .I(n497), .Z(n496) );
  BUFFD0 U422 ( .I(n498), .Z(n497) );
  BUFFD0 U423 ( .I(n499), .Z(n498) );
  BUFFD0 U424 ( .I(n500), .Z(n499) );
  BUFFD0 U425 ( .I(n501), .Z(n500) );
  BUFFD0 U426 ( .I(n502), .Z(n501) );
  BUFFD0 U427 ( .I(n503), .Z(n502) );
  BUFFD0 U428 ( .I(n504), .Z(n503) );
  BUFFD0 U429 ( .I(n505), .Z(n504) );
  BUFFD0 U430 ( .I(n506), .Z(n505) );
  BUFFD0 U431 ( .I(n507), .Z(n506) );
  BUFFD0 U432 ( .I(n508), .Z(n507) );
  BUFFD0 U433 ( .I(n509), .Z(n508) );
  BUFFD0 U434 ( .I(n512), .Z(n509) );
  BUFFD0 U435 ( .I(N51), .Z(n510) );
  BUFFD0 U436 ( .I(n510), .Z(n511) );
  BUFFD0 U437 ( .I(n513), .Z(n512) );
  BUFFD0 U438 ( .I(n514), .Z(n513) );
  BUFFD0 U439 ( .I(n515), .Z(n514) );
  BUFFD0 U440 ( .I(n516), .Z(n515) );
  BUFFD0 U441 ( .I(n517), .Z(n516) );
  BUFFD0 U442 ( .I(n518), .Z(n517) );
  BUFFD0 U443 ( .I(n519), .Z(n518) );
  BUFFD0 U444 ( .I(n520), .Z(n519) );
  BUFFD0 U445 ( .I(n521), .Z(n520) );
  BUFFD0 U446 ( .I(n522), .Z(n521) );
  BUFFD0 U447 ( .I(n523), .Z(n522) );
  CKBD0 U448 ( .CLK(n1268), .C(n523) );
  BUFFD0 U449 ( .I(n525), .Z(n524) );
  BUFFD0 U450 ( .I(n526), .Z(n525) );
  BUFFD0 U451 ( .I(n527), .Z(n526) );
  BUFFD0 U452 ( .I(n528), .Z(n527) );
  BUFFD0 U453 ( .I(n529), .Z(n528) );
  BUFFD0 U454 ( .I(n530), .Z(n529) );
  BUFFD0 U455 ( .I(n531), .Z(n530) );
  BUFFD0 U456 ( .I(n532), .Z(n531) );
  BUFFD0 U457 ( .I(n533), .Z(n532) );
  BUFFD0 U458 ( .I(n534), .Z(n533) );
  BUFFD0 U459 ( .I(n535), .Z(n534) );
  BUFFD0 U460 ( .I(n536), .Z(n535) );
  BUFFD0 U461 ( .I(n537), .Z(n536) );
  BUFFD0 U462 ( .I(n540), .Z(n537) );
  BUFFD0 U463 ( .I(N54), .Z(n538) );
  BUFFD0 U464 ( .I(n538), .Z(n539) );
  BUFFD0 U465 ( .I(n541), .Z(n540) );
  BUFFD0 U466 ( .I(n542), .Z(n541) );
  BUFFD0 U467 ( .I(n543), .Z(n542) );
  BUFFD0 U468 ( .I(n544), .Z(n543) );
  BUFFD0 U469 ( .I(n545), .Z(n544) );
  BUFFD0 U470 ( .I(n546), .Z(n545) );
  BUFFD0 U471 ( .I(n547), .Z(n546) );
  BUFFD0 U472 ( .I(n548), .Z(n547) );
  BUFFD0 U473 ( .I(n549), .Z(n548) );
  BUFFD0 U474 ( .I(n550), .Z(n549) );
  BUFFD0 U475 ( .I(n551), .Z(n550) );
  BUFFD0 U476 ( .I(n552), .Z(n551) );
  BUFFD0 U477 ( .I(n553), .Z(n552) );
  BUFFD0 U478 ( .I(n554), .Z(n553) );
  BUFFD0 U479 ( .I(n555), .Z(n554) );
  BUFFD0 U480 ( .I(n556), .Z(n555) );
  BUFFD0 U481 ( .I(n557), .Z(n556) );
  BUFFD0 U482 ( .I(n558), .Z(n557) );
  BUFFD0 U483 ( .I(n559), .Z(n558) );
  BUFFD0 U484 ( .I(n560), .Z(n559) );
  BUFFD0 U485 ( .I(n561), .Z(n560) );
  BUFFD0 U486 ( .I(n564), .Z(n561) );
  BUFFD0 U487 ( .I(n1397), .Z(n562) );
  BUFFD0 U488 ( .I(n562), .Z(n563) );
  CKBD0 U489 ( .CLK(n1270), .C(n564) );
  CKBD0 U490 ( .CLK(n563), .C(ReadAddr[4]) );
  BUFFD0 U491 ( .I(n570), .Z(n565) );
  BUFFD0 U492 ( .I(N75), .Z(n566) );
  BUFFD0 U493 ( .I(n566), .Z(n567) );
  BUFFD0 U494 ( .I(n567), .Z(n568) );
  BUFFD0 U495 ( .I(n568), .Z(n569) );
  BUFFD0 U496 ( .I(n571), .Z(n570) );
  BUFFD0 U497 ( .I(n572), .Z(n571) );
  BUFFD0 U498 ( .I(n573), .Z(n572) );
  BUFFD0 U499 ( .I(n574), .Z(n573) );
  BUFFD0 U500 ( .I(n575), .Z(n574) );
  BUFFD0 U501 ( .I(n576), .Z(n575) );
  BUFFD0 U502 ( .I(n577), .Z(n576) );
  BUFFD0 U503 ( .I(n578), .Z(n577) );
  BUFFD0 U504 ( .I(n579), .Z(n578) );
  BUFFD0 U505 ( .I(n580), .Z(n579) );
  BUFFD0 U506 ( .I(n581), .Z(n580) );
  BUFFD0 U507 ( .I(n582), .Z(n581) );
  BUFFD0 U508 ( .I(n583), .Z(n582) );
  BUFFD0 U509 ( .I(n584), .Z(n583) );
  BUFFD0 U510 ( .I(n585), .Z(n584) );
  BUFFD0 U511 ( .I(n586), .Z(n585) );
  BUFFD0 U512 ( .I(n587), .Z(n586) );
  BUFFD0 U513 ( .I(n588), .Z(n587) );
  BUFFD0 U514 ( .I(n589), .Z(n588) );
  BUFFD0 U515 ( .I(n590), .Z(n589) );
  BUFFD0 U516 ( .I(n591), .Z(n590) );
  BUFFD0 U517 ( .I(n592), .Z(n591) );
  BUFFD0 U518 ( .I(n593), .Z(n592) );
  BUFFD0 U519 ( .I(n594), .Z(n593) );
  BUFFD0 U520 ( .I(n595), .Z(n594) );
  BUFFD0 U521 ( .I(n596), .Z(n595) );
  BUFFD0 U522 ( .I(n597), .Z(n596) );
  BUFFD0 U523 ( .I(n598), .Z(n597) );
  BUFFD0 U524 ( .I(n599), .Z(n598) );
  BUFFD0 U525 ( .I(n600), .Z(n599) );
  BUFFD0 U526 ( .I(n601), .Z(n600) );
  BUFFD0 U527 ( .I(n602), .Z(n601) );
  BUFFD0 U528 ( .I(n603), .Z(n602) );
  BUFFD0 U529 ( .I(n604), .Z(n603) );
  BUFFD0 U530 ( .I(n605), .Z(n604) );
  BUFFD0 U531 ( .I(n606), .Z(n605) );
  BUFFD0 U532 ( .I(n607), .Z(n606) );
  BUFFD0 U533 ( .I(n608), .Z(n607) );
  BUFFD0 U534 ( .I(n609), .Z(n608) );
  BUFFD0 U535 ( .I(n610), .Z(n609) );
  BUFFD0 U536 ( .I(n611), .Z(n610) );
  BUFFD0 U537 ( .I(n612), .Z(n611) );
  BUFFD0 U538 ( .I(n613), .Z(n612) );
  BUFFD0 U539 ( .I(n614), .Z(n613) );
  BUFFD0 U540 ( .I(n615), .Z(n614) );
  BUFFD0 U541 ( .I(n616), .Z(n615) );
  BUFFD0 U542 ( .I(n569), .Z(n616) );
  BUFFD0 U543 ( .I(ReadAddr[2]), .Z(n617) );
  BUFFD0 U544 ( .I(n620), .Z(n618) );
  BUFFD0 U545 ( .I(n621), .Z(n619) );
  BUFFD0 U546 ( .I(n622), .Z(n620) );
  BUFFD0 U547 ( .I(n623), .Z(n621) );
  BUFFD0 U548 ( .I(n624), .Z(n622) );
  BUFFD0 U549 ( .I(n625), .Z(n623) );
  BUFFD0 U550 ( .I(n626), .Z(n624) );
  BUFFD0 U551 ( .I(n627), .Z(n625) );
  BUFFD0 U552 ( .I(n628), .Z(n626) );
  BUFFD0 U553 ( .I(n629), .Z(n627) );
  BUFFD0 U554 ( .I(n630), .Z(n628) );
  BUFFD0 U555 ( .I(n631), .Z(n629) );
  BUFFD0 U556 ( .I(n632), .Z(n630) );
  BUFFD0 U557 ( .I(n633), .Z(n631) );
  BUFFD0 U558 ( .I(n634), .Z(n632) );
  BUFFD0 U559 ( .I(n635), .Z(n633) );
  BUFFD0 U560 ( .I(n73), .Z(n634) );
  BUFFD0 U561 ( .I(n636), .Z(n635) );
  BUFFD0 U562 ( .I(n637), .Z(n636) );
  BUFFD0 U563 ( .I(n638), .Z(n637) );
  BUFFD0 U564 ( .I(n639), .Z(n638) );
  BUFFD0 U565 ( .I(n640), .Z(n639) );
  BUFFD0 U566 ( .I(n641), .Z(n640) );
  BUFFD0 U567 ( .I(n642), .Z(n641) );
  BUFFD0 U568 ( .I(n643), .Z(n642) );
  BUFFD0 U569 ( .I(n644), .Z(n643) );
  BUFFD0 U570 ( .I(n645), .Z(n644) );
  BUFFD0 U571 ( .I(n646), .Z(n645) );
  BUFFD0 U572 ( .I(n647), .Z(n646) );
  BUFFD0 U573 ( .I(n648), .Z(n647) );
  BUFFD0 U574 ( .I(n649), .Z(n648) );
  BUFFD0 U575 ( .I(n650), .Z(n649) );
  BUFFD0 U576 ( .I(n651), .Z(n650) );
  BUFFD0 U577 ( .I(n652), .Z(n651) );
  BUFFD0 U578 ( .I(n653), .Z(n652) );
  BUFFD0 U579 ( .I(n654), .Z(n653) );
  BUFFD0 U580 ( .I(n655), .Z(n654) );
  BUFFD0 U581 ( .I(n656), .Z(n655) );
  CKBD0 U582 ( .CLK(n1272), .C(n656) );
  BUFFD0 U583 ( .I(ReadAddr[3]), .Z(n657) );
  CKBD0 U584 ( .CLK(n1398), .C(ReadAddr[2]) );
  BUFFD0 U585 ( .I(n662), .Z(n658) );
  BUFFD0 U586 ( .I(N74), .Z(n659) );
  BUFFD0 U587 ( .I(n659), .Z(n660) );
  BUFFD0 U588 ( .I(n660), .Z(n661) );
  BUFFD0 U589 ( .I(n663), .Z(n662) );
  BUFFD0 U590 ( .I(n664), .Z(n663) );
  BUFFD0 U591 ( .I(n665), .Z(n664) );
  BUFFD0 U592 ( .I(n666), .Z(n665) );
  BUFFD0 U593 ( .I(n667), .Z(n666) );
  BUFFD0 U594 ( .I(n668), .Z(n667) );
  BUFFD0 U595 ( .I(n669), .Z(n668) );
  BUFFD0 U596 ( .I(n670), .Z(n669) );
  BUFFD0 U597 ( .I(n671), .Z(n670) );
  BUFFD0 U598 ( .I(n672), .Z(n671) );
  BUFFD0 U599 ( .I(n673), .Z(n672) );
  BUFFD0 U600 ( .I(n674), .Z(n673) );
  BUFFD0 U601 ( .I(n675), .Z(n674) );
  BUFFD0 U602 ( .I(n676), .Z(n675) );
  BUFFD0 U603 ( .I(n677), .Z(n676) );
  BUFFD0 U604 ( .I(n678), .Z(n677) );
  BUFFD0 U605 ( .I(n679), .Z(n678) );
  BUFFD0 U606 ( .I(n680), .Z(n679) );
  BUFFD0 U607 ( .I(n681), .Z(n680) );
  BUFFD0 U608 ( .I(n682), .Z(n681) );
  BUFFD0 U609 ( .I(n683), .Z(n682) );
  BUFFD0 U610 ( .I(n684), .Z(n683) );
  BUFFD0 U611 ( .I(n685), .Z(n684) );
  BUFFD0 U612 ( .I(n686), .Z(n685) );
  BUFFD0 U613 ( .I(n687), .Z(n686) );
  BUFFD0 U614 ( .I(n688), .Z(n687) );
  BUFFD0 U615 ( .I(n689), .Z(n688) );
  BUFFD0 U616 ( .I(n690), .Z(n689) );
  BUFFD0 U617 ( .I(n691), .Z(n690) );
  BUFFD0 U618 ( .I(n692), .Z(n691) );
  BUFFD0 U619 ( .I(n693), .Z(n692) );
  BUFFD0 U620 ( .I(n694), .Z(n693) );
  BUFFD0 U621 ( .I(n695), .Z(n694) );
  BUFFD0 U622 ( .I(n696), .Z(n695) );
  BUFFD0 U623 ( .I(n697), .Z(n696) );
  BUFFD0 U624 ( .I(n698), .Z(n697) );
  BUFFD0 U625 ( .I(n699), .Z(n698) );
  BUFFD0 U626 ( .I(n700), .Z(n699) );
  BUFFD0 U627 ( .I(n701), .Z(n700) );
  BUFFD0 U628 ( .I(n702), .Z(n701) );
  BUFFD0 U629 ( .I(n703), .Z(n702) );
  BUFFD0 U630 ( .I(n704), .Z(n703) );
  BUFFD0 U631 ( .I(n705), .Z(n704) );
  BUFFD0 U632 ( .I(n706), .Z(n705) );
  BUFFD0 U633 ( .I(n707), .Z(n706) );
  BUFFD0 U634 ( .I(n708), .Z(n707) );
  BUFFD0 U635 ( .I(n709), .Z(n708) );
  BUFFD0 U636 ( .I(n661), .Z(n709) );
  BUFFD0 U637 ( .I(n713), .Z(n710) );
  BUFFD0 U638 ( .I(N73), .Z(n711) );
  BUFFD0 U639 ( .I(n711), .Z(n712) );
  BUFFD0 U640 ( .I(n714), .Z(n713) );
  BUFFD0 U641 ( .I(n715), .Z(n714) );
  BUFFD0 U642 ( .I(n716), .Z(n715) );
  BUFFD0 U643 ( .I(n717), .Z(n716) );
  BUFFD0 U644 ( .I(n718), .Z(n717) );
  BUFFD0 U645 ( .I(n719), .Z(n718) );
  BUFFD0 U646 ( .I(n720), .Z(n719) );
  BUFFD0 U647 ( .I(n721), .Z(n720) );
  BUFFD0 U648 ( .I(n722), .Z(n721) );
  BUFFD0 U649 ( .I(n723), .Z(n722) );
  BUFFD0 U650 ( .I(n724), .Z(n723) );
  BUFFD0 U651 ( .I(n725), .Z(n724) );
  BUFFD0 U652 ( .I(n726), .Z(n725) );
  BUFFD0 U653 ( .I(n727), .Z(n726) );
  BUFFD0 U654 ( .I(n728), .Z(n727) );
  BUFFD0 U655 ( .I(n729), .Z(n728) );
  BUFFD0 U656 ( .I(n730), .Z(n729) );
  BUFFD0 U657 ( .I(n731), .Z(n730) );
  BUFFD0 U658 ( .I(n732), .Z(n731) );
  BUFFD0 U659 ( .I(n733), .Z(n732) );
  BUFFD0 U660 ( .I(n734), .Z(n733) );
  BUFFD0 U661 ( .I(n735), .Z(n734) );
  BUFFD0 U662 ( .I(n736), .Z(n735) );
  BUFFD0 U663 ( .I(n737), .Z(n736) );
  BUFFD0 U664 ( .I(n738), .Z(n737) );
  BUFFD0 U665 ( .I(n739), .Z(n738) );
  BUFFD0 U666 ( .I(n740), .Z(n739) );
  BUFFD0 U667 ( .I(n741), .Z(n740) );
  BUFFD0 U668 ( .I(n742), .Z(n741) );
  BUFFD0 U669 ( .I(n743), .Z(n742) );
  BUFFD0 U670 ( .I(n744), .Z(n743) );
  BUFFD0 U671 ( .I(n745), .Z(n744) );
  BUFFD0 U672 ( .I(n746), .Z(n745) );
  BUFFD0 U673 ( .I(n748), .Z(n746) );
  BUFFD0 U674 ( .I(n753), .Z(n747) );
  BUFFD0 U675 ( .I(n749), .Z(n748) );
  BUFFD0 U676 ( .I(n750), .Z(n749) );
  BUFFD0 U677 ( .I(n751), .Z(n750) );
  BUFFD0 U678 ( .I(n752), .Z(n751) );
  BUFFD0 U679 ( .I(n754), .Z(n752) );
  BUFFD0 U680 ( .I(n759), .Z(n753) );
  BUFFD0 U681 ( .I(n755), .Z(n754) );
  BUFFD0 U682 ( .I(n756), .Z(n755) );
  BUFFD0 U683 ( .I(n757), .Z(n756) );
  BUFFD0 U684 ( .I(n758), .Z(n757) );
  BUFFD0 U685 ( .I(n712), .Z(n758) );
  CKBD0 U686 ( .CLK(N330), .C(n759) );
  BUFFD0 U687 ( .I(n761), .Z(n760) );
  BUFFD0 U688 ( .I(n762), .Z(n761) );
  BUFFD0 U689 ( .I(n763), .Z(n762) );
  BUFFD0 U690 ( .I(n764), .Z(n763) );
  BUFFD0 U691 ( .I(n765), .Z(n764) );
  BUFFD0 U692 ( .I(n766), .Z(n765) );
  BUFFD0 U693 ( .I(n767), .Z(n766) );
  BUFFD0 U694 ( .I(n768), .Z(n767) );
  BUFFD0 U695 ( .I(n769), .Z(n768) );
  BUFFD0 U696 ( .I(n770), .Z(n769) );
  BUFFD0 U697 ( .I(n771), .Z(n770) );
  BUFFD0 U698 ( .I(n772), .Z(n771) );
  BUFFD0 U699 ( .I(n773), .Z(n772) );
  BUFFD0 U700 ( .I(n774), .Z(n773) );
  BUFFD0 U701 ( .I(n775), .Z(n774) );
  BUFFD0 U702 ( .I(n776), .Z(n775) );
  BUFFD0 U703 ( .I(n777), .Z(n776) );
  BUFFD0 U704 ( .I(n778), .Z(n777) );
  BUFFD0 U705 ( .I(n779), .Z(n778) );
  BUFFD0 U706 ( .I(n780), .Z(n779) );
  BUFFD0 U707 ( .I(n781), .Z(n780) );
  BUFFD0 U708 ( .I(n782), .Z(n781) );
  BUFFD0 U709 ( .I(n783), .Z(n782) );
  BUFFD0 U710 ( .I(n784), .Z(n783) );
  BUFFD0 U711 ( .I(n785), .Z(n784) );
  BUFFD0 U712 ( .I(n786), .Z(n785) );
  CKBD0 U713 ( .CLK(n790), .C(n786) );
  BUFFD0 U714 ( .I(ReadAddr[1]), .Z(n787) );
  CKBD0 U715 ( .CLK(n787), .C(n788) );
  CKNXD16 U716 ( .I(n789), .ZN(n790) );
  INVD0 U717 ( .I(n275), .ZN(n789) );
  BUFFD0 U718 ( .I(n792), .Z(n791) );
  BUFFD0 U719 ( .I(n794), .Z(n792) );
  BUFFD0 U720 ( .I(n795), .Z(n793) );
  BUFFD0 U721 ( .I(n796), .Z(n794) );
  BUFFD0 U722 ( .I(n797), .Z(n795) );
  BUFFD0 U723 ( .I(n798), .Z(n796) );
  BUFFD0 U724 ( .I(n799), .Z(n797) );
  BUFFD0 U725 ( .I(n801), .Z(n798) );
  BUFFD0 U726 ( .I(n800), .Z(n799) );
  BUFFD0 U727 ( .I(n802), .Z(n800) );
  BUFFD0 U728 ( .I(n803), .Z(n801) );
  BUFFD0 U729 ( .I(n804), .Z(n802) );
  BUFFD0 U730 ( .I(n805), .Z(n803) );
  BUFFD0 U731 ( .I(n806), .Z(n804) );
  BUFFD0 U732 ( .I(n807), .Z(n805) );
  BUFFD0 U733 ( .I(n808), .Z(n806) );
  BUFFD0 U734 ( .I(n809), .Z(n807) );
  BUFFD0 U735 ( .I(n810), .Z(n808) );
  BUFFD0 U736 ( .I(n811), .Z(n809) );
  BUFFD0 U737 ( .I(n812), .Z(n810) );
  BUFFD0 U738 ( .I(n813), .Z(n811) );
  BUFFD0 U739 ( .I(n814), .Z(n812) );
  BUFFD0 U740 ( .I(n815), .Z(n813) );
  BUFFD0 U741 ( .I(n816), .Z(n814) );
  BUFFD0 U742 ( .I(N49), .Z(n815) );
  BUFFD0 U743 ( .I(n817), .Z(n816) );
  BUFFD0 U744 ( .I(n818), .Z(n817) );
  BUFFD0 U745 ( .I(n819), .Z(n818) );
  BUFFD0 U746 ( .I(n820), .Z(n819) );
  BUFFD0 U747 ( .I(n1348), .Z(n820) );
  NR2XD0 U748 ( .A1(n793), .A2(n99), .ZN(N49) );
  INVD0 U749 ( .I(N44), .ZN(n1393) );
  CKBD0 U750 ( .CLK(ReadAddr[0]), .C(n821) );
  CKNXD16 U751 ( .I(n822), .ZN(n823) );
  CKNXD0 U752 ( .I(n825), .ZN(n822) );
  CKNXD16 U753 ( .I(n824), .ZN(n825) );
  CKNXD0 U754 ( .I(n827), .ZN(n824) );
  CKNXD16 U755 ( .I(n826), .ZN(n827) );
  CKNXD0 U756 ( .I(n829), .ZN(n826) );
  CKNXD16 U757 ( .I(n828), .ZN(n829) );
  CKNXD0 U758 ( .I(n831), .ZN(n828) );
  INVD0 U759 ( .I(n839), .ZN(n836) );
  CKNXD16 U760 ( .I(n830), .ZN(n831) );
  CKNXD0 U761 ( .I(n833), .ZN(n830) );
  CKNXD16 U762 ( .I(n832), .ZN(n833) );
  CKNXD0 U763 ( .I(n835), .ZN(n832) );
  CKNXD16 U764 ( .I(n834), .ZN(n835) );
  CKNXD0 U765 ( .I(n837), .ZN(n834) );
  CKNXD16 U766 ( .I(n323), .ZN(n20) );
  CKNXD16 U767 ( .I(n845), .ZN(n846) );
  INVD0 U768 ( .I(n851), .ZN(n845) );
  INVD0 U769 ( .I(n847), .ZN(n848) );
  CKNXD16 U770 ( .I(n850), .ZN(n851) );
  INVD0 U771 ( .I(n849), .ZN(n850) );
  BUFFD0 U772 ( .I(n853), .Z(n852) );
  CKBD0 U773 ( .CLK(n855), .C(n853) );
  CKNXD16 U774 ( .I(n854), .ZN(n855) );
  CKNXD0 U775 ( .I(n857), .ZN(n854) );
  CKNXD16 U776 ( .I(n856), .ZN(n857) );
  CKNXD0 U777 ( .I(n859), .ZN(n856) );
  CKNXD16 U778 ( .I(n858), .ZN(n859) );
  CKNXD0 U779 ( .I(n861), .ZN(n858) );
  CKNXD16 U780 ( .I(n860), .ZN(n861) );
  INVD0 U781 ( .I(n863), .ZN(n860) );
  CKNXD16 U782 ( .I(n862), .ZN(n863) );
  CKNXD0 U783 ( .I(n865), .ZN(n862) );
  CKNXD16 U784 ( .I(n864), .ZN(n865) );
  CKNXD0 U785 ( .I(n867), .ZN(n864) );
  CKNXD16 U786 ( .I(n866), .ZN(n867) );
  CKNXD0 U787 ( .I(n869), .ZN(n866) );
  CKNXD16 U788 ( .I(n868), .ZN(n869) );
  CKNXD0 U789 ( .I(n872), .ZN(n868) );
  BUFFD0 U790 ( .I(n18), .Z(n870) );
  CKNXD16 U791 ( .I(n871), .ZN(n872) );
  CKNXD0 U792 ( .I(n874), .ZN(n871) );
  CKNXD16 U793 ( .I(n873), .ZN(n874) );
  INVD0 U794 ( .I(n876), .ZN(n873) );
  CKNXD0 U795 ( .I(n134), .ZN(n875) );
  OAI22D4 U796 ( .A1(n16), .A2(n870), .B1(n19), .B2(n17), .ZN(n134) );
  BUFFD0 U797 ( .I(n879), .Z(n877) );
  CKNXD16 U798 ( .I(n878), .ZN(n879) );
  CKNXD0 U799 ( .I(n881), .ZN(n878) );
  CKNXD16 U800 ( .I(n880), .ZN(n881) );
  INVD0 U801 ( .I(n883), .ZN(n880) );
  CKNXD16 U802 ( .I(n882), .ZN(n883) );
  CKNXD0 U803 ( .I(n885), .ZN(n882) );
  CKNXD16 U804 ( .I(n884), .ZN(n885) );
  CKNXD0 U805 ( .I(n887), .ZN(n884) );
  CKNXD16 U806 ( .I(n886), .ZN(n887) );
  CKNXD0 U807 ( .I(n889), .ZN(n886) );
  CKNXD16 U808 ( .I(n888), .ZN(n889) );
  CKNXD0 U809 ( .I(n891), .ZN(n888) );
  CKNXD16 U810 ( .I(n890), .ZN(n891) );
  CKNXD0 U811 ( .I(n893), .ZN(n890) );
  CKNXD16 U812 ( .I(n892), .ZN(n893) );
  CKNXD0 U813 ( .I(n895), .ZN(n892) );
  CKNXD16 U814 ( .I(n894), .ZN(n895) );
  CKNXD0 U815 ( .I(n897), .ZN(n894) );
  CKNXD16 U816 ( .I(n896), .ZN(n897) );
  CKNXD0 U817 ( .I(n899), .ZN(n896) );
  CKNXD16 U818 ( .I(n898), .ZN(n899) );
  INVD0 U819 ( .I(n900), .ZN(n898) );
  CKNXD16 U820 ( .I(n288), .ZN(n900) );
  CKNXD16 U821 ( .I(n901), .ZN(n902) );
  CKNXD0 U822 ( .I(n904), .ZN(n901) );
  CKNXD16 U823 ( .I(n903), .ZN(n904) );
  INVD0 U824 ( .I(n906), .ZN(n903) );
  INVD0 U825 ( .I(n908), .ZN(n905) );
  INVD0 U826 ( .I(n911), .ZN(n912) );
  CKNXD16 U827 ( .I(n914), .ZN(n911) );
  CKNXD16 U828 ( .I(n905), .ZN(n906) );
  CKNXD16 U829 ( .I(n907), .ZN(n908) );
  INVD0 U830 ( .I(n910), .ZN(n907) );
  INVD0 U831 ( .I(n912), .ZN(n909) );
  INVD0 U832 ( .I(n913), .ZN(n914) );
  CKNXD16 U833 ( .I(n916), .ZN(n913) );
  CKNXD16 U834 ( .I(n909), .ZN(n910) );
  INVD0 U835 ( .I(n915), .ZN(n916) );
  CKNXD16 U836 ( .I(n917), .ZN(n915) );
  INVD0 U837 ( .I(n283), .ZN(n917) );
  CKNXD16 U838 ( .I(n918), .ZN(n919) );
  CKNXD0 U839 ( .I(n921), .ZN(n918) );
  CKNXD16 U840 ( .I(n920), .ZN(n921) );
  INVD0 U841 ( .I(n923), .ZN(n920) );
  INVD0 U842 ( .I(n925), .ZN(n922) );
  INVD0 U843 ( .I(n928), .ZN(n929) );
  CKNXD16 U844 ( .I(n931), .ZN(n928) );
  CKNXD16 U845 ( .I(n922), .ZN(n923) );
  CKNXD16 U846 ( .I(n924), .ZN(n925) );
  INVD0 U847 ( .I(n927), .ZN(n924) );
  INVD0 U848 ( .I(n929), .ZN(n926) );
  INVD0 U849 ( .I(n930), .ZN(n931) );
  CKNXD16 U850 ( .I(n933), .ZN(n930) );
  CKNXD16 U851 ( .I(n926), .ZN(n927) );
  INVD0 U852 ( .I(n932), .ZN(n933) );
  CKNXD16 U853 ( .I(n934), .ZN(n932) );
  INVD0 U854 ( .I(n282), .ZN(n934) );
  CKNXD16 U855 ( .I(n935), .ZN(n936) );
  CKNXD0 U856 ( .I(n938), .ZN(n935) );
  CKNXD16 U857 ( .I(n937), .ZN(n938) );
  INVD0 U858 ( .I(n940), .ZN(n937) );
  INVD0 U859 ( .I(n942), .ZN(n939) );
  INVD0 U860 ( .I(n945), .ZN(n946) );
  CKNXD16 U861 ( .I(n948), .ZN(n945) );
  CKNXD16 U862 ( .I(n939), .ZN(n940) );
  CKNXD16 U863 ( .I(n941), .ZN(n942) );
  INVD0 U864 ( .I(n944), .ZN(n941) );
  INVD0 U865 ( .I(n946), .ZN(n943) );
  INVD0 U866 ( .I(n947), .ZN(n948) );
  CKNXD16 U867 ( .I(n950), .ZN(n947) );
  CKNXD16 U868 ( .I(n943), .ZN(n944) );
  INVD0 U869 ( .I(n949), .ZN(n950) );
  CKNXD16 U870 ( .I(n951), .ZN(n949) );
  INVD0 U871 ( .I(n281), .ZN(n951) );
  CKNXD16 U872 ( .I(n952), .ZN(n953) );
  CKNXD0 U873 ( .I(n955), .ZN(n952) );
  CKNXD16 U874 ( .I(n954), .ZN(n955) );
  INVD0 U875 ( .I(n957), .ZN(n954) );
  INVD0 U876 ( .I(n959), .ZN(n956) );
  INVD0 U877 ( .I(n962), .ZN(n963) );
  CKNXD16 U878 ( .I(n965), .ZN(n962) );
  CKNXD16 U879 ( .I(n956), .ZN(n957) );
  CKNXD16 U880 ( .I(n958), .ZN(n959) );
  INVD0 U881 ( .I(n961), .ZN(n958) );
  INVD0 U882 ( .I(n963), .ZN(n960) );
  INVD0 U883 ( .I(n964), .ZN(n965) );
  CKNXD16 U884 ( .I(n967), .ZN(n964) );
  CKNXD16 U885 ( .I(n960), .ZN(n961) );
  INVD0 U886 ( .I(n966), .ZN(n967) );
  CKNXD16 U887 ( .I(n969), .ZN(n966) );
  INVD0 U888 ( .I(n968), .ZN(n969) );
  CKNXD16 U889 ( .I(n131), .ZN(n968) );
  CKNXD16 U890 ( .I(n970), .ZN(n971) );
  CKNXD0 U891 ( .I(n973), .ZN(n970) );
  CKNXD16 U892 ( .I(n972), .ZN(n973) );
  INVD0 U893 ( .I(n975), .ZN(n972) );
  INVD0 U894 ( .I(n977), .ZN(n974) );
  INVD0 U895 ( .I(n980), .ZN(n981) );
  CKNXD16 U896 ( .I(n983), .ZN(n980) );
  CKNXD16 U897 ( .I(n974), .ZN(n975) );
  CKNXD16 U898 ( .I(n976), .ZN(n977) );
  INVD0 U899 ( .I(n979), .ZN(n976) );
  INVD0 U900 ( .I(n981), .ZN(n978) );
  INVD0 U901 ( .I(n982), .ZN(n983) );
  CKNXD16 U902 ( .I(n985), .ZN(n982) );
  CKNXD16 U903 ( .I(n978), .ZN(n979) );
  INVD0 U904 ( .I(n984), .ZN(n985) );
  CKNXD16 U905 ( .I(n987), .ZN(n984) );
  INVD0 U906 ( .I(n986), .ZN(n987) );
  CKNXD16 U907 ( .I(n130), .ZN(n986) );
  CKNXD16 U908 ( .I(n988), .ZN(n989) );
  CKNXD0 U909 ( .I(n991), .ZN(n988) );
  CKNXD16 U910 ( .I(n990), .ZN(n991) );
  INVD0 U911 ( .I(n993), .ZN(n990) );
  INVD0 U912 ( .I(n995), .ZN(n992) );
  INVD0 U913 ( .I(n998), .ZN(n999) );
  CKNXD16 U914 ( .I(n1001), .ZN(n998) );
  CKNXD16 U915 ( .I(n992), .ZN(n993) );
  CKNXD16 U916 ( .I(n994), .ZN(n995) );
  INVD0 U917 ( .I(n997), .ZN(n994) );
  INVD0 U918 ( .I(n999), .ZN(n996) );
  INVD0 U919 ( .I(n1000), .ZN(n1001) );
  CKNXD16 U920 ( .I(n1003), .ZN(n1000) );
  CKNXD16 U921 ( .I(n996), .ZN(n997) );
  INVD0 U922 ( .I(n1002), .ZN(n1003) );
  CKNXD16 U923 ( .I(n1005), .ZN(n1002) );
  INVD0 U924 ( .I(n1004), .ZN(n1005) );
  CKNXD16 U925 ( .I(n128), .ZN(n1004) );
  BUFFD0 U926 ( .I(n1403), .Z(n1006) );
  BUFFD0 U927 ( .I(n1006), .Z(n1007) );
  BUFFD0 U928 ( .I(n1007), .Z(n1008) );
  BUFFD0 U929 ( .I(n1008), .Z(n1009) );
  BUFFD0 U930 ( .I(n1009), .Z(n1010) );
  BUFFD0 U931 ( .I(n1010), .Z(n1011) );
  BUFFD0 U932 ( .I(n1011), .Z(n1012) );
  BUFFD0 U933 ( .I(n1012), .Z(n1013) );
  BUFFD0 U934 ( .I(n1013), .Z(n1014) );
  BUFFD0 U935 ( .I(n1014), .Z(n1015) );
  BUFFD0 U936 ( .I(n1015), .Z(n1016) );
  BUFFD0 U937 ( .I(n1016), .Z(n1017) );
  BUFFD0 U938 ( .I(n1017), .Z(n1018) );
  BUFFD0 U939 ( .I(n1018), .Z(n1019) );
  BUFFD0 U940 ( .I(n1019), .Z(n1020) );
  BUFFD0 U941 ( .I(n1020), .Z(n1021) );
  BUFFD0 U942 ( .I(n1021), .Z(n1022) );
  BUFFD0 U943 ( .I(n1022), .Z(n1023) );
  BUFFD0 U944 ( .I(n1023), .Z(n1024) );
  BUFFD0 U945 ( .I(n1024), .Z(n1025) );
  BUFFD0 U946 ( .I(n1025), .Z(n1026) );
  BUFFD0 U947 ( .I(n1026), .Z(n1027) );
  BUFFD0 U948 ( .I(n1027), .Z(n1028) );
  BUFFD0 U949 ( .I(n1028), .Z(n1029) );
  BUFFD0 U950 ( .I(n1029), .Z(n1030) );
  BUFFD0 U951 ( .I(n1030), .Z(n1031) );
  BUFFD0 U952 ( .I(n1031), .Z(n1032) );
  BUFFD0 U953 ( .I(n1032), .Z(n1033) );
  BUFFD0 U954 ( .I(n1033), .Z(n1034) );
  BUFFD0 U955 ( .I(n1034), .Z(n1035) );
  BUFFD0 U956 ( .I(n1035), .Z(n1036) );
  BUFFD0 U957 ( .I(n1036), .Z(n1037) );
  BUFFD0 U958 ( .I(n1037), .Z(n1038) );
  BUFFD0 U959 ( .I(n1038), .Z(n1039) );
  BUFFD0 U960 ( .I(n1039), .Z(n1040) );
  BUFFD0 U961 ( .I(n1040), .Z(n1041) );
  BUFFD0 U962 ( .I(n1041), .Z(n1042) );
  BUFFD0 U963 ( .I(n1042), .Z(n1043) );
  BUFFD0 U964 ( .I(n1043), .Z(n1044) );
  BUFFD0 U965 ( .I(n1044), .Z(n1045) );
  BUFFD0 U966 ( .I(n1045), .Z(n1046) );
  BUFFD0 U967 ( .I(n1046), .Z(n1047) );
  BUFFD0 U968 ( .I(n1047), .Z(n1048) );
  BUFFD0 U969 ( .I(n1048), .Z(n1049) );
  BUFFD0 U970 ( .I(n1049), .Z(n1050) );
  BUFFD0 U971 ( .I(n1050), .Z(n1051) );
  BUFFD0 U972 ( .I(n1051), .Z(n1052) );
  BUFFD0 U973 ( .I(n1052), .Z(n1053) );
  BUFFD0 U974 ( .I(n1053), .Z(n1054) );
  BUFFD0 U975 ( .I(n1054), .Z(n1055) );
  BUFFD0 U976 ( .I(n1055), .Z(n1056) );
  BUFFD0 U977 ( .I(n1056), .Z(n1057) );
  BUFFD0 U978 ( .I(n1057), .Z(n1058) );
  BUFFD0 U979 ( .I(n1058), .Z(n1059) );
  BUFFD0 U980 ( .I(n1059), .Z(n1060) );
  BUFFD0 U981 ( .I(n1060), .Z(n1061) );
  BUFFD0 U982 ( .I(n1061), .Z(n1062) );
  BUFFD0 U983 ( .I(n1062), .Z(n1063) );
  BUFFD0 U984 ( .I(n1063), .Z(n1064) );
  BUFFD0 U985 ( .I(n1064), .Z(n1065) );
  BUFFD0 U986 ( .I(n1065), .Z(n1066) );
  BUFFD0 U987 ( .I(n1066), .Z(n1067) );
  BUFFD0 U988 ( .I(n1067), .Z(n1068) );
  BUFFD0 U989 ( .I(n1068), .Z(n1069) );
  BUFFD0 U990 ( .I(n1069), .Z(n1070) );
  BUFFD0 U991 ( .I(n1070), .Z(n1071) );
  BUFFD0 U992 ( .I(n1071), .Z(n1072) );
  BUFFD0 U993 ( .I(n1072), .Z(n1073) );
  BUFFD0 U994 ( .I(n1073), .Z(n1074) );
  BUFFD0 U995 ( .I(n1074), .Z(n1075) );
  BUFFD0 U996 ( .I(n1075), .Z(n1076) );
  BUFFD0 U997 ( .I(n1076), .Z(n1077) );
  BUFFD0 U998 ( .I(n1077), .Z(n1078) );
  BUFFD0 U999 ( .I(n1078), .Z(n1079) );
  BUFFD0 U1000 ( .I(n1079), .Z(n1080) );
  BUFFD0 U1001 ( .I(n1080), .Z(n1081) );
  BUFFD0 U1002 ( .I(n1081), .Z(n1082) );
  BUFFD0 U1003 ( .I(n1082), .Z(n1083) );
  BUFFD0 U1004 ( .I(n1083), .Z(n1084) );
  BUFFD0 U1005 ( .I(n1084), .Z(n1085) );
  BUFFD0 U1006 ( .I(n1085), .Z(n1086) );
  BUFFD0 U1007 ( .I(n1086), .Z(n1087) );
  BUFFD0 U1008 ( .I(n1087), .Z(n1088) );
  BUFFD0 U1009 ( .I(n1088), .Z(n1089) );
  BUFFD0 U1010 ( .I(n1089), .Z(n1090) );
  BUFFD0 U1011 ( .I(n1090), .Z(n1091) );
  BUFFD0 U1012 ( .I(n1091), .Z(n1092) );
  BUFFD0 U1013 ( .I(n1092), .Z(n1093) );
  BUFFD0 U1014 ( .I(n1093), .Z(n1094) );
  BUFFD0 U1015 ( .I(n1094), .Z(n1095) );
  BUFFD0 U1016 ( .I(n1095), .Z(n1096) );
  BUFFD0 U1017 ( .I(n1096), .Z(n1097) );
  BUFFD0 U1018 ( .I(n1097), .Z(n1098) );
  BUFFD0 U1019 ( .I(n1098), .Z(n1099) );
  BUFFD0 U1020 ( .I(n1099), .Z(n1100) );
  BUFFD0 U1021 ( .I(n1100), .Z(n1101) );
  BUFFD0 U1022 ( .I(n1101), .Z(n1102) );
  BUFFD0 U1023 ( .I(n1102), .Z(n1103) );
  BUFFD0 U1024 ( .I(n1103), .Z(n1104) );
  BUFFD0 U1025 ( .I(n1104), .Z(n1105) );
  BUFFD0 U1026 ( .I(n1105), .Z(n1106) );
  BUFFD0 U1027 ( .I(n1106), .Z(n1107) );
  BUFFD0 U1028 ( .I(n1107), .Z(n1108) );
  BUFFD0 U1029 ( .I(n1108), .Z(n1109) );
  BUFFD0 U1030 ( .I(n1109), .Z(n1110) );
  BUFFD0 U1031 ( .I(n1110), .Z(n1111) );
  BUFFD0 U1032 ( .I(n1111), .Z(n1112) );
  BUFFD0 U1033 ( .I(n1112), .Z(n1113) );
  BUFFD0 U1034 ( .I(n1113), .Z(n1114) );
  BUFFD0 U1035 ( .I(n1114), .Z(n1115) );
  BUFFD0 U1036 ( .I(n1115), .Z(n1116) );
  BUFFD0 U1037 ( .I(n1116), .Z(n1117) );
  BUFFD0 U1038 ( .I(n1117), .Z(n1118) );
  BUFFD0 U1039 ( .I(n1118), .Z(n1119) );
  BUFFD0 U1040 ( .I(n1119), .Z(n1120) );
  BUFFD0 U1041 ( .I(n1120), .Z(n1121) );
  BUFFD0 U1042 ( .I(n1121), .Z(n1122) );
  BUFFD0 U1043 ( .I(n1122), .Z(n1123) );
  BUFFD0 U1044 ( .I(n1123), .Z(n1124) );
  BUFFD0 U1045 ( .I(n1124), .Z(n1125) );
  BUFFD0 U1046 ( .I(n1125), .Z(n1126) );
  BUFFD0 U1047 ( .I(n1126), .Z(n1127) );
  BUFFD0 U1048 ( .I(n1127), .Z(n1128) );
  BUFFD0 U1049 ( .I(n1128), .Z(n1129) );
  BUFFD0 U1050 ( .I(n1129), .Z(n1130) );
  BUFFD0 U1051 ( .I(n1130), .Z(n1131) );
  BUFFD0 U1052 ( .I(n1131), .Z(n1132) );
  BUFFD0 U1053 ( .I(n1132), .Z(n1133) );
  BUFFD0 U1054 ( .I(n1133), .Z(n1134) );
  BUFFD0 U1055 ( .I(n1134), .Z(n1135) );
  BUFFD0 U1056 ( .I(n1135), .Z(n1136) );
  BUFFD0 U1057 ( .I(n1136), .Z(n1137) );
  BUFFD0 U1058 ( .I(n1137), .Z(n1138) );
  BUFFD0 U1059 ( .I(n1138), .Z(n1139) );
  BUFFD0 U1060 ( .I(n1139), .Z(n1140) );
  BUFFD0 U1061 ( .I(n1140), .Z(n1141) );
  BUFFD0 U1062 ( .I(n1141), .Z(n1142) );
  BUFFD0 U1063 ( .I(n1142), .Z(n1143) );
  BUFFD0 U1064 ( .I(n1143), .Z(n1144) );
  BUFFD0 U1065 ( .I(n1144), .Z(n1145) );
  BUFFD0 U1066 ( .I(n1145), .Z(n1146) );
  BUFFD0 U1067 ( .I(n1146), .Z(n1147) );
  BUFFD0 U1068 ( .I(n1147), .Z(n1148) );
  BUFFD0 U1069 ( .I(n1148), .Z(n1149) );
  BUFFD0 U1070 ( .I(n1149), .Z(n1150) );
  BUFFD0 U1071 ( .I(n1150), .Z(n1151) );
  BUFFD0 U1072 ( .I(n1151), .Z(n1152) );
  BUFFD0 U1073 ( .I(n1152), .Z(n1153) );
  BUFFD0 U1074 ( .I(n1153), .Z(n1154) );
  BUFFD0 U1075 ( .I(n1154), .Z(n1155) );
  BUFFD0 U1076 ( .I(n1155), .Z(n1156) );
  BUFFD0 U1077 ( .I(n1156), .Z(n1157) );
  BUFFD0 U1078 ( .I(n1157), .Z(n1158) );
  BUFFD0 U1079 ( .I(n1158), .Z(n1159) );
  BUFFD0 U1080 ( .I(n1159), .Z(n1160) );
  BUFFD0 U1081 ( .I(n1160), .Z(n1161) );
  BUFFD0 U1082 ( .I(n1161), .Z(n1162) );
  BUFFD0 U1083 ( .I(n1162), .Z(n1163) );
  BUFFD0 U1084 ( .I(n1163), .Z(n1164) );
  BUFFD0 U1085 ( .I(n1164), .Z(n1165) );
  BUFFD0 U1086 ( .I(n1165), .Z(n1166) );
  BUFFD0 U1087 ( .I(n1166), .Z(n1167) );
  BUFFD0 U1088 ( .I(n1167), .Z(n1168) );
  BUFFD0 U1089 ( .I(n1168), .Z(n1169) );
  BUFFD0 U1090 ( .I(n1169), .Z(n1170) );
  BUFFD0 U1091 ( .I(n1170), .Z(n1171) );
  BUFFD0 U1092 ( .I(n1171), .Z(n1172) );
  BUFFD0 U1093 ( .I(n1172), .Z(n1173) );
  BUFFD0 U1094 ( .I(n1173), .Z(n1174) );
  BUFFD0 U1095 ( .I(n1174), .Z(n1175) );
  BUFFD0 U1096 ( .I(n1175), .Z(n1176) );
  BUFFD0 U1097 ( .I(n1176), .Z(n1177) );
  BUFFD0 U1098 ( .I(n1177), .Z(n1178) );
  BUFFD0 U1099 ( .I(n1178), .Z(n1179) );
  CKNXD16 U1100 ( .I(n1180), .ZN(n1181) );
  INVD0 U1101 ( .I(n1184), .ZN(n1180) );
  CKNXD16 U1102 ( .I(n1182), .ZN(n1185) );
  INVD0 U1103 ( .I(n280), .ZN(n1182) );
  CKNXD16 U1104 ( .I(n1183), .ZN(n1184) );
  INVD0 U1105 ( .I(n1188), .ZN(n1183) );
  CKNXD16 U1106 ( .I(n1186), .ZN(n1189) );
  INVD0 U1107 ( .I(n1185), .ZN(n1186) );
  CKNXD16 U1108 ( .I(n1187), .ZN(n1188) );
  INVD0 U1109 ( .I(n1192), .ZN(n1187) );
  CKNXD16 U1110 ( .I(n1190), .ZN(n1193) );
  INVD0 U1111 ( .I(n1189), .ZN(n1190) );
  CKNXD16 U1112 ( .I(n1191), .ZN(n1192) );
  INVD0 U1113 ( .I(n1197), .ZN(n1191) );
  INVD0 U1114 ( .I(n1193), .ZN(n1194) );
  CKNXD16 U1115 ( .I(n1196), .ZN(n1197) );
  INVD0 U1116 ( .I(n1195), .ZN(n1196) );
  CKNXD16 U1117 ( .I(n1198), .ZN(n1199) );
  CKNXD0 U1118 ( .I(n1201), .ZN(n1198) );
  CKNXD16 U1119 ( .I(n1200), .ZN(n1201) );
  CKNXD0 U1120 ( .I(n1203), .ZN(n1200) );
  CKNXD16 U1121 ( .I(n1202), .ZN(n1203) );
  CKNXD0 U1122 ( .I(n1205), .ZN(n1202) );
  CKNXD16 U1123 ( .I(n1204), .ZN(n1205) );
  CKNXD0 U1124 ( .I(n1207), .ZN(n1204) );
  CKNXD16 U1125 ( .I(n1206), .ZN(n1207) );
  CKNXD0 U1126 ( .I(n1209), .ZN(n1206) );
  CKNXD16 U1127 ( .I(n1208), .ZN(n1209) );
  CKNXD0 U1128 ( .I(n1211), .ZN(n1208) );
  CKNXD16 U1129 ( .I(n1210), .ZN(n1211) );
  CKNXD0 U1130 ( .I(n1213), .ZN(n1210) );
  INVD0 U1131 ( .I(n1217), .ZN(n1214) );
  CKNXD16 U1132 ( .I(n1212), .ZN(n1213) );
  CKNXD0 U1133 ( .I(n1215), .ZN(n1212) );
  CKNXD16 U1134 ( .I(n1214), .ZN(n1215) );
  CKNXD16 U1135 ( .I(n1216), .ZN(n1217) );
  INVD0 U1136 ( .I(n140), .ZN(n1216) );
  OAI211D0 U1137 ( .A1(CurState[1]), .A2(n55), .B(n35), .C(n93), .ZN(n24) );
  CKNXD16 U1138 ( .I(n1218), .ZN(n1219) );
  CKNXD0 U1139 ( .I(n1221), .ZN(n1218) );
  CKNXD16 U1140 ( .I(n1220), .ZN(n1221) );
  INVD0 U1141 ( .I(n1223), .ZN(n1220) );
  CKNXD16 U1142 ( .I(n1222), .ZN(n1223) );
  CKNXD0 U1143 ( .I(n1227), .ZN(n1222) );
  CKNXD16 U1144 ( .I(n1226), .ZN(n1227) );
  CKNXD0 U1145 ( .I(n1229), .ZN(n1226) );
  CKNXD16 U1146 ( .I(n1228), .ZN(n1229) );
  CKNXD0 U1147 ( .I(n1231), .ZN(n1228) );
  CKNXD16 U1148 ( .I(n1230), .ZN(n1231) );
  CKNXD0 U1149 ( .I(n1233), .ZN(n1230) );
  CKNXD16 U1150 ( .I(n1232), .ZN(n1233) );
  CKNXD0 U1151 ( .I(n1235), .ZN(n1232) );
  CKNXD16 U1152 ( .I(n1234), .ZN(n1235) );
  CKNXD0 U1153 ( .I(n1237), .ZN(n1234) );
  CKNXD16 U1154 ( .I(n1236), .ZN(n1237) );
  CKNXD16 U1155 ( .I(n1238), .ZN(n1239) );
  INVD0 U1156 ( .I(n1225), .ZN(n1238) );
  CKNXD16 U1157 ( .I(n1240), .ZN(n1241) );
  CKNXD0 U1158 ( .I(n1243), .ZN(n1240) );
  CKNXD16 U1159 ( .I(n1242), .ZN(n1243) );
  CKNXD0 U1160 ( .I(n1245), .ZN(n1242) );
  CKNXD16 U1161 ( .I(n1244), .ZN(n1245) );
  CKNXD0 U1162 ( .I(n1247), .ZN(n1244) );
  CKNXD16 U1163 ( .I(n1246), .ZN(n1247) );
  INVD0 U1164 ( .I(n1249), .ZN(n1246) );
  CKNXD16 U1165 ( .I(n1248), .ZN(n1249) );
  CKNXD0 U1166 ( .I(n1251), .ZN(n1248) );
  CKNXD16 U1167 ( .I(n1250), .ZN(n1251) );
  CKNXD0 U1168 ( .I(n1253), .ZN(n1250) );
  CKNXD16 U1169 ( .I(n1252), .ZN(n1253) );
  CKNXD0 U1170 ( .I(n1255), .ZN(n1252) );
  CKNXD16 U1171 ( .I(n1254), .ZN(n1255) );
  CKNXD0 U1172 ( .I(n1257), .ZN(n1254) );
  CKNXD16 U1173 ( .I(n1256), .ZN(n1257) );
  CKNXD0 U1174 ( .I(n1259), .ZN(n1256) );
  CKNXD16 U1175 ( .I(n1258), .ZN(n1259) );
  CKNXD0 U1176 ( .I(n1261), .ZN(n1258) );
  CKNXD16 U1177 ( .I(n1260), .ZN(n1261) );
  INVD0 U1178 ( .I(n278), .ZN(n1260) );
  CKND12 U1179 ( .CLK(WriteReq), .CN(n33) );
  CKBXD0 U1180 ( .I(n1179), .Z(WriteCmd) );
  CKNXD16 U1181 ( .I(n1263), .ZN(n1264) );
  INVD0 U1182 ( .I(n1266), .ZN(n1263) );
  CKNXD16 U1183 ( .I(n1265), .ZN(n1266) );
  INVD0 U1184 ( .I(n139), .ZN(n1265) );
  CKNXD16 U1185 ( .I(n1267), .ZN(n1268) );
  INVD0 U1186 ( .I(n511), .ZN(n1267) );
  INR2D0 U1187 ( .A1(N46), .B1(n99), .ZN(N51) );
  CKNXD16 U1188 ( .I(n1269), .ZN(n1270) );
  INVD0 U1189 ( .I(n539), .ZN(n1269) );
  INR2D0 U1190 ( .A1(N48), .B1(n99), .ZN(N54) );
  CKNXD16 U1191 ( .I(n1271), .ZN(n1272) );
  INVD0 U1192 ( .I(N52), .ZN(n1271) );
  NR2D0 U1193 ( .A1(n618), .A2(n99), .ZN(N52) );
  INVD0 U1194 ( .I(n1274), .ZN(n1275) );
  INVD16 U1195 ( .I(n147), .ZN(n1273) );
  CKNXD16 U1196 ( .I(n1289), .ZN(n1274) );
  INVD0 U1197 ( .I(n1276), .ZN(n1277) );
  INVD16 U1198 ( .I(n12), .ZN(n1276) );
  CKNXD0 U1199 ( .I(n1278), .ZN(n1279) );
  INVD16 U1200 ( .I(n1277), .ZN(n1278) );
  CKNXD0 U1201 ( .I(n1280), .ZN(n1281) );
  INVD16 U1202 ( .I(n1279), .ZN(n1280) );
  INVD0 U1203 ( .I(n1282), .ZN(n1283) );
  INVD16 U1204 ( .I(n1281), .ZN(n1282) );
  CKNXD0 U1205 ( .I(n1284), .ZN(n1285) );
  INVD16 U1206 ( .I(n1283), .ZN(n1284) );
  INVD0 U1207 ( .I(n1286), .ZN(n1287) );
  INVD16 U1208 ( .I(n1285), .ZN(n1286) );
  CKBXD0 U1209 ( .I(n1291), .Z(n1288) );
  BUFFD0 U1210 ( .I(n1273), .Z(n1289) );
  INVD0 U1211 ( .I(n1290), .ZN(n1291) );
  CKNXD16 U1212 ( .I(n1293), .ZN(n1290) );
  INVD0 U1213 ( .I(n1292), .ZN(n1293) );
  CKND12 U1214 ( .CLK(n1287), .CN(n1292) );
  ND3D0 U1215 ( .A1(CurState[1]), .A2(CurState[0]), .A3(CurState[2]), .ZN(n12)
         );
  BUFFD0 U1216 ( .I(n1402), .Z(n1294) );
  BUFFD0 U1217 ( .I(n1294), .Z(n1295) );
  BUFFD0 U1218 ( .I(n1295), .Z(n1296) );
  BUFFD0 U1219 ( .I(n1296), .Z(n1297) );
  BUFFD0 U1220 ( .I(n1297), .Z(n1298) );
  BUFFD0 U1221 ( .I(n1298), .Z(n1299) );
  BUFFD0 U1222 ( .I(n1299), .Z(n1300) );
  BUFFD0 U1223 ( .I(n1300), .Z(n1301) );
  BUFFD0 U1224 ( .I(n1301), .Z(n1302) );
  BUFFD0 U1225 ( .I(n1302), .Z(n1303) );
  BUFFD0 U1226 ( .I(n1303), .Z(n1304) );
  BUFFD0 U1227 ( .I(n1304), .Z(n1305) );
  BUFFD0 U1228 ( .I(n1305), .Z(n1306) );
  BUFFD0 U1229 ( .I(n1306), .Z(n1307) );
  BUFFD0 U1230 ( .I(n1307), .Z(n1308) );
  BUFFD0 U1231 ( .I(n1308), .Z(n1309) );
  BUFFD0 U1232 ( .I(n1309), .Z(n1310) );
  BUFFD0 U1233 ( .I(n1310), .Z(n1311) );
  BUFFD0 U1234 ( .I(n1311), .Z(n1312) );
  BUFFD0 U1235 ( .I(n1312), .Z(n1313) );
  BUFFD0 U1236 ( .I(n1313), .Z(n1314) );
  BUFFD0 U1237 ( .I(n1314), .Z(n1315) );
  BUFFD0 U1238 ( .I(n1315), .Z(n1316) );
  BUFFD0 U1239 ( .I(n1316), .Z(n1317) );
  BUFFD0 U1240 ( .I(n1317), .Z(n1318) );
  BUFFD0 U1241 ( .I(n1318), .Z(n1319) );
  BUFFD0 U1242 ( .I(n1319), .Z(n1320) );
  BUFFD0 U1243 ( .I(n1320), .Z(n1321) );
  BUFFD0 U1244 ( .I(n1321), .Z(n1322) );
  BUFFD0 U1245 ( .I(n1322), .Z(n1323) );
  BUFFD0 U1246 ( .I(n1323), .Z(n1324) );
  BUFFD0 U1247 ( .I(n1324), .Z(n1325) );
  BUFFD0 U1248 ( .I(n1325), .Z(n1326) );
  BUFFD0 U1249 ( .I(n1326), .Z(n1327) );
  BUFFD0 U1250 ( .I(n1327), .Z(n1328) );
  BUFFD0 U1251 ( .I(n1328), .Z(n1329) );
  BUFFD0 U1252 ( .I(n1329), .Z(n1330) );
  BUFFD0 U1253 ( .I(n1330), .Z(n1331) );
  BUFFD0 U1254 ( .I(n1331), .Z(n1332) );
  BUFFD0 U1255 ( .I(n1332), .Z(n1333) );
  BUFFD0 U1256 ( .I(n1333), .Z(n1334) );
  BUFFD0 U1257 ( .I(n1334), .Z(n1335) );
  BUFFD0 U1258 ( .I(n1335), .Z(n1336) );
  BUFFD0 U1259 ( .I(n1336), .Z(n1337) );
  BUFFD0 U1260 ( .I(n1337), .Z(n1338) );
  BUFFD0 U1261 ( .I(n1338), .Z(n1339) );
  BUFFD0 U1262 ( .I(n1339), .Z(n1340) );
  BUFFD0 U1263 ( .I(n1340), .Z(n1341) );
  BUFFD0 U1264 ( .I(n1341), .Z(n1342) );
  BUFFD0 U1265 ( .I(n1342), .Z(n1343) );
  CKBD0 U1266 ( .CLK(n1343), .C(ReadCmd) );
  INVD0 U1267 ( .I(n72), .ZN(n1345) );
  INVD0 U1268 ( .I(N45), .ZN(n72) );
  CKNXD16 U1269 ( .I(n1347), .ZN(n1348) );
  INVD0 U1270 ( .I(n1393), .ZN(n1347) );
  BUFFD0 U1271 ( .I(n1356), .Z(n1359) );
  INVD0 U1272 ( .I(n1349), .ZN(n1350) );
  INVD16 U1273 ( .I(n6), .ZN(n1349) );
  INVD0 U1274 ( .I(n1351), .ZN(n1352) );
  INVD16 U1275 ( .I(n1350), .ZN(n1351) );
  INVD0 U1276 ( .I(n1353), .ZN(n1354) );
  CKNXD16 U1277 ( .I(n1355), .ZN(n1353) );
  CKBXD0 U1278 ( .I(n1365), .Z(n1355) );
  CKNXD16 U1279 ( .I(n1364), .ZN(n1365) );
  INVD0 U1280 ( .I(n1363), .ZN(n1364) );
  CKNXD16 U1281 ( .I(n1361), .ZN(n1362) );
  CKNXD16 U1282 ( .I(n160), .ZN(n1356) );
  INVD0 U1283 ( .I(n1357), .ZN(n1358) );
  CKNXD16 U1284 ( .I(n1359), .ZN(n1357) );
  INVD0 U1285 ( .I(n1360), .ZN(n1361) );
  INVD16 U1286 ( .I(n1352), .ZN(n1360) );
  INVD0 U1287 ( .I(n1362), .ZN(n1363) );
  ND3D0 U1288 ( .A1(n29), .A2(n159), .A3(n158), .ZN(n6) );
  OAI31D4 U1289 ( .A1(n6), .A2(WriteReq), .A3(Reset), .B(n286), .ZN(n127) );
  OAI31D4 U1290 ( .A1(n12), .A2(Reset), .A3(ReadReq), .B(n287), .ZN(n132) );
  CKBXD0 U1291 ( .I(n1371), .Z(n1366) );
  CKNXD16 U1292 ( .I(n1366), .ZN(EmptyFIFO) );
  CKBXD0 U1293 ( .I(n1370), .Z(n1368) );
  CKNXD16 U1294 ( .I(n1368), .ZN(FullFIFO) );
  CKND0 U1295 ( .CLK(n1401), .CN(n1370) );
  CKND0 U1296 ( .CLK(n1400), .CN(n1371) );
  INVD1 U1297 ( .I(N47), .ZN(n73) );
  INVD1 U1298 ( .I(n6), .ZN(n15) );
  INVD1 U1299 ( .I(n17), .ZN(n16) );
  INVD1 U1300 ( .I(n9), .ZN(n8) );
  INVD1 U1301 ( .I(Reset), .ZN(n1390) );
  NR3D0 U1302 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n53) );
  ND3D1 U1303 ( .A1(n86), .A2(n87), .A3(n88), .ZN(n31) );
  XOR2D1 U1304 ( .A1(n19), .A2(n1395), .Z(n87) );
  XOR2D1 U1305 ( .A1(N333), .A2(n1396), .Z(n86) );
  NR3D0 U1306 ( .A1(n89), .A2(n90), .A3(n91), .ZN(n88) );
  ND4D1 U1307 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(n30) );
  XOR2D1 U1308 ( .A1(n657), .A2(n74), .Z(n62) );
  NR3D0 U1309 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n65) );
  XNR2D1 U1310 ( .A1(ReadAddr[4]), .A2(N72), .ZN(n64) );
  XOR2D1 U1311 ( .A1(WriteAddr[2]), .A2(N46), .Z(n54) );
  IIND4D1 U1312 ( .A1(n54), .A2(n56), .B1(n51), .B2(n52), .ZN(n63) );
  XNR2D1 U1313 ( .A1(N177), .A2(n81), .ZN(n49) );
  XOR2D1 U1314 ( .A1(ReadAddr[2]), .A2(N70), .Z(n68) );
  INVD1 U1315 ( .I(N71), .ZN(n74) );
  ND3D1 U1316 ( .A1(n100), .A2(n97), .A3(ReadReq), .ZN(n9) );
  INVD1 U1317 ( .I(n100), .ZN(n98) );
  INVD1 U1318 ( .I(n22), .ZN(n32) );
  ND2D1 U1319 ( .A1(n35), .A2(n12), .ZN(n100) );
  ND2D1 U1320 ( .A1(n35), .A2(n6), .ZN(n22) );
  INVD1 U1321 ( .I(n1288), .ZN(n28) );
  OAI22D0 U1322 ( .A1(n1396), .A2(n1288), .B1(n74), .B2(n34), .ZN(N76) );
  INVD1 U1323 ( .I(n24), .ZN(n25) );
  ND3D1 U1324 ( .A1(n103), .A2(n104), .A3(n105), .ZN(n97) );
  XOR2D1 U1325 ( .A1(ReadAddr[0]), .A2(n118), .Z(n103) );
  NR3D0 U1326 ( .A1(n106), .A2(n107), .A3(n108), .ZN(n105) );
  XOR2D1 U1327 ( .A1(ReadAddr[1]), .A2(n19), .Z(n78) );
  INVD1 U1328 ( .I(n34), .ZN(n109) );
  XOR2D1 U1329 ( .A1(N176), .A2(WriteAddr[2]), .Z(n50) );
  XOR2D1 U1330 ( .A1(n1395), .A2(n19), .Z(n45) );
  IND4D1 U1331 ( .A1(n80), .B1(n75), .B2(n76), .B3(n78), .ZN(n82) );
  XOR2D1 U1332 ( .A1(ReadAddr[0]), .A2(N68), .Z(n67) );
  XOR2D1 U1333 ( .A1(ReadAddr[1]), .A2(N69), .Z(n66) );
  NR2D1 U1334 ( .A1(n1373), .A2(n1374), .ZN(n76) );
  XNR2D1 U1335 ( .A1(n657), .A2(n81), .ZN(n1373) );
  XOR2D1 U1336 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .Z(n1374) );
  AO22D0 U1337 ( .A1(N72), .A2(n109), .B1(ReadAddr[4]), .B2(n28), .Z(N77) );
  AO22D0 U1338 ( .A1(N70), .A2(n109), .B1(n617), .B2(n28), .Z(N75) );
  AO22D0 U1339 ( .A1(n821), .A2(n28), .B1(N68), .B2(n109), .Z(N73) );
  AO22D0 U1340 ( .A1(n788), .A2(n28), .B1(N69), .B2(n109), .Z(N74) );
  INVD1 U1341 ( .I(ReadReq), .ZN(n95) );
  INVD1 U1342 ( .I(Reset), .ZN(n143) );
  AOI22D0 U1343 ( .A1(n61), .A2(n55), .B1(CurState[0]), .B2(n30), .ZN(n60) );
  ND4D1 U1344 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(n61) );
  AOI31D0 U1345 ( .A1(n46), .A2(n45), .A3(n79), .B(n80), .ZN(n77) );
  NR3D0 U1346 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n79) );
  OAI221D0 U1347 ( .A1(CurState[2]), .A2(n43), .B1(CurState[0]), .B2(n44), .C(
        n24), .ZN(n42) );
  IINR4D0 U1348 ( .A1(n45), .A2(n46), .B1(n47), .B2(n48), .ZN(n44) );
  AOI31D0 U1349 ( .A1(n51), .A2(n52), .A3(n53), .B(n29), .ZN(n43) );
  AOI21D1 U1350 ( .A1(CurState[0]), .A2(n27), .B(n28), .ZN(n26) );
  NR3D0 U1351 ( .A1(n58), .A2(n15), .A3(n59), .ZN(n57) );
  AOI21D1 U1352 ( .A1(n31), .A2(n82), .B(n83), .ZN(n58) );
  NR3D0 U1353 ( .A1(n29), .A2(CurState[2]), .A3(n60), .ZN(n59) );
  XOR2D1 U1354 ( .A1(WriteAddr[3]), .A2(n73), .Z(n51) );
  XOR2D1 U1355 ( .A1(WriteAddr[4]), .A2(N48), .Z(n56) );
  XNR2D1 U1356 ( .A1(N178), .A2(WriteAddr[4]), .ZN(n46) );
  INVD1 U1357 ( .I(n657), .ZN(n1396) );
  XOR2D1 U1358 ( .A1(ReadAddr[4]), .A2(N334), .Z(n90) );
  BUFFD1 U1359 ( .I(n1399), .Z(WriteAddr[2]) );
  NR2D1 U1360 ( .A1(n1375), .A2(n1376), .ZN(n52) );
  XNR2D1 U1361 ( .A1(\add_389/carry[2] ), .A2(n72), .ZN(n1375) );
  XNR2D1 U1362 ( .A1(N330), .A2(n1393), .ZN(n1376) );
  AOI21D1 U1363 ( .A1(WriteReq), .A2(n15), .B(n94), .ZN(n93) );
  AOI21D1 U1364 ( .A1(CurState[0]), .A2(n95), .B(n96), .ZN(n94) );
  ND2D1 U1365 ( .A1(ReadCmd), .A2(n157), .ZN(n99) );
  OAI22D0 U1366 ( .A1(n16), .A2(n301), .B1(n21), .B2(n17), .ZN(n135) );
  INVD1 U1367 ( .I(N330), .ZN(n21) );
  INVD1 U1368 ( .I(\add_389/carry[2] ), .ZN(n19) );
  XOR2D1 U1369 ( .A1(ReadAddr[0]), .A2(N330), .Z(n48) );
  XOR2D1 U1370 ( .A1(N330), .A2(n301), .Z(n36) );
  NR3D0 U1371 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n38) );
  XNR2D1 U1372 ( .A1(ReadAddr[4]), .A2(WriteAddr[4]), .ZN(n75) );
  ND3D1 U1373 ( .A1(CurState[0]), .A2(n29), .A3(CurState[2]), .ZN(n83) );
  INVD1 U1374 ( .I(WriteAddr[3]), .ZN(n81) );
  XOR2D1 U1375 ( .A1(ReadAddr[2]), .A2(N332), .Z(n89) );
  XOR2D1 U1376 ( .A1(ReadAddr[0]), .A2(N330), .Z(n80) );
  XOR2D1 U1377 ( .A1(ReadAddr[0]), .A2(N330), .Z(n91) );
  XOR2D1 U1378 ( .A1(n657), .A2(OldReadAr[3]), .Z(n106) );
  XOR2D1 U1379 ( .A1(ReadAddr[4]), .A2(OldReadAr[4]), .Z(n108) );
  XOR2D1 U1380 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .Z(n107) );
  AO22D0 U1381 ( .A1(n657), .A2(n8), .B1(n9), .B2(OldReadAr[3]), .Z(n128) );
  AO22D0 U1382 ( .A1(ReadAddr[2]), .A2(n8), .B1(n9), .B2(OldReadAr[2]), .Z(
        n130) );
  AO22D0 U1383 ( .A1(ReadAddr[4]), .A2(n8), .B1(n9), .B2(OldReadAr[4]), .Z(
        n131) );
  ND2D1 U1384 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  CKXOR2D0 U1385 ( .A1(ReadAddr[4]), .A2(\add_308/carry[4] ), .Z(N178) );
  AN2D0 U1386 ( .A1(n657), .A2(\add_308/carry[3] ), .Z(\add_308/carry[4] ) );
  CKXOR2D0 U1387 ( .A1(\add_308/carry[3] ), .A2(n657), .Z(N177) );
  AN2D0 U1388 ( .A1(ReadAddr[2]), .A2(ReadAddr[1]), .Z(\add_308/carry[3] ) );
  CKXOR2D0 U1389 ( .A1(ReadAddr[1]), .A2(ReadAddr[2]), .Z(N176) );
  CKXOR2D0 U1390 ( .A1(WriteAddr[4]), .A2(\add_389/carry[4] ), .Z(N334) );
  AN2D0 U1391 ( .A1(WriteAddr[3]), .A2(\add_389/carry[3] ), .Z(
        \add_389/carry[4] ) );
  CKXOR2D0 U1392 ( .A1(\add_389/carry[3] ), .A2(WriteAddr[3]), .Z(N333) );
  AN2D0 U1393 ( .A1(WriteAddr[2]), .A2(\add_389/carry[2] ), .Z(
        \add_389/carry[3] ) );
  CKXOR2D0 U1394 ( .A1(\add_389/carry[2] ), .A2(WriteAddr[2]), .Z(N332) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, ClockR, ClockW, Dreadyr, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N85, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n107,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  XNR4D1 U18 ( .A1(n8745), .A2(n8743), .A3(n8750), .A4(n8747), .ZN(n84) );
  XOR4D1 U19 ( .A1(n8755), .A2(n8753), .A3(n8760), .A4(n8757), .Z(n83) );
  XOR4D1 U20 ( .A1(n8735), .A2(n8733), .A3(n8740), .A4(n8737), .Z(n80) );
  XOR4D1 U21 ( .A1(n8719), .A2(n8717), .A3(n8724), .A4(n8721), .Z(n77) );
  XNR4D1 U22 ( .A1(n8703), .A2(n8701), .A3(n8708), .A4(n8705), .ZN(n74) );
  XOR4D1 U27 ( .A1(n90), .A2(n2097), .A3(n91), .A4(n2152), .Z(n89) );
  XNR4D1 U28 ( .A1(n2095), .A2(n2087), .A3(n2094), .A4(n2089), .ZN(n91) );
  XNR4D1 U33 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n97) );
  XOR4D1 U34 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n96) );
  XNR4D1 U35 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .ZN(n93) );
  XNR4D1 U36 ( .A1(n2086), .A2(n2092), .A3(n2088), .A4(n2085), .ZN(n87) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(n8527), .E(n8474), .CP(n8552), .CDN(
        n8415), .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(n2220), .E(n8474), .CP(n8552), .CDN(
        n8414), .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(n8757), .E(n8473), .CP(n8552), .CDN(
        n8414), .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(n8755), .E(n8474), .CP(n8552), .CDN(
        n8414), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(n2672), .E(n8473), .CP(n8552), .CDN(
        n8414), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(n7289), .E(n8474), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(n8747), .E(n8473), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(n8745), .E(n8474), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(n2849), .E(n8473), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(n3026), .E(n8474), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n8737), .E(n8473), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(n8735), .E(n8473), .CP(n8553), .CDN(
        n8414), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(n3561), .E(n8473), .CP(n8553), .CDN(
        n8413), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(n3880), .E(n8473), .CP(n8553), .CDN(
        n8413), .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(n8728), .E(n8473), .CP(n8553), .CDN(
        n8413), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(n8726), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(n4268), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n8721), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n8719), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(n4803), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n5122), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(n8712), .E(n8473), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(n8710), .E(n8474), .CP(n8554), .CDN(
        n8413), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n5512), .E(n8474), .CP(n8554), .CDN(n8412), .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(n8705), .E(n8474), .CP(n8554), .CDN(n8412), .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n8703), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n6047), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n6366), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n8696), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(n8694), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n6900), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(n8689), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n7255), .E(n8474), .CP(n8555), .CDN(n8412), .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(n8527), .E(n8478), .CP(n8559), .CDN(
        n8409), .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(n2220), .E(n8478), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(n8757), .E(n8477), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(n8755), .E(n8478), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(n2672), .E(n8477), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(n7289), .E(n8478), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(n8747), .E(n8477), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(n8745), .E(n8478), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(n2849), .E(n8477), .CP(n8559), .CDN(
        n8408), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(n3026), .E(n8478), .CP(n8560), .CDN(
        n8408), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n8737), .E(n8477), .CP(n8560), .CDN(
        n8408), .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(n8735), .E(n8477), .CP(n8560), .CDN(
        n8408), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(n3561), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(n3880), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(n8728), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(n8726), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(n4268), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n8721), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n8719), .E(n8477), .CP(n8560), .CDN(
        n8407), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(n4803), .E(n8477), .CP(n8561), .CDN(
        n8407), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n5122), .E(n8477), .CP(n8561), .CDN(
        n8407), .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(n8712), .E(n8477), .CP(n8561), .CDN(
        n8407), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(n8710), .E(n8478), .CP(n8561), .CDN(
        n8407), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n5512), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(n8705), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n8703), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n6047), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n6366), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n8696), .E(n8478), .CP(n8561), .CDN(n8406), .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(n8694), .E(n8478), .CP(n8562), .CDN(n8406), .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n6900), .E(n8478), .CP(n8562), .CDN(n8406), .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(n8689), .E(n8478), .CP(n8562), .CDN(n8406), .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n7255), .E(n8478), .CP(n8562), .CDN(n8406), .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(n8527), .E(n8466), .CP(n8539), .CDN(
        n8427), .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(n2220), .E(n8466), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(n2314), .E(n8465), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(n2493), .E(n8466), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(n2672), .E(n8465), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(n7289), .E(n8466), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(n2849), .E(n8465), .CP(n8540), .CDN(
        n8426), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(n3026), .E(n8466), .CP(n8540), .CDN(
        n8426), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(n3203), .E(n8465), .CP(n8540), .CDN(
        n8426), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(n3382), .E(n8465), .CP(n8540), .CDN(
        n8426), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(n3561), .E(n8465), .CP(n8540), .CDN(
        n8425), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(n3880), .E(n8465), .CP(n8540), .CDN(
        n8425), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(n3910), .E(n8465), .CP(n8540), .CDN(
        n8425), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(n4089), .E(n8465), .CP(n8540), .CDN(
        n8425), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(n4268), .E(n8465), .CP(n8540), .CDN(
        n8425), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(n4445), .E(n8465), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(n4624), .E(n8465), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(n4803), .E(n8465), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(n5122), .E(n8465), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(n5154), .E(n8465), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(n5333), .E(n8466), .CP(n8541), .CDN(
        n8425), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(n5512), .E(n8466), .CP(n8541), .CDN(n8424), .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(n5689), .E(n8466), .CP(n8541), .CDN(n8424), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(n5868), .E(n8466), .CP(n8541), .CDN(n8424), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n6047), .E(n8466), .CP(n8541), .CDN(n8424), .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(n6366), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(n6400), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(n6579), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(n6900), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(n6934), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(n7255), .E(n8466), .CP(n8542), .CDN(n8424), .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n8527), .E(n8468), .CP(n8542), .CDN(
        n8424), .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(n2220), .E(n8468), .CP(n8542), .CDN(
        n8423), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(n2314), .E(n8467), .CP(n8542), .CDN(
        n8423), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(n2493), .E(n8468), .CP(n8542), .CDN(
        n8423), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(n2672), .E(n8467), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(n7289), .E(n8468), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(n2849), .E(n8467), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(n3026), .E(n8468), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(n3203), .E(n8467), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(n3382), .E(n8467), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(n3561), .E(n8467), .CP(n8543), .CDN(
        n8422), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(n3880), .E(n8467), .CP(n8543), .CDN(
        n8422), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(n3910), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(n4089), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(n4268), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(n4445), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(n4624), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(n4803), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(n5122), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(n5154), .E(n8467), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(n5333), .E(n8468), .CP(n8544), .CDN(
        n8422), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(n5512), .E(n8468), .CP(n8544), .CDN(n8421), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(n5689), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(n5868), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(n6047), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(n6366), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(n6400), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(n6579), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(n6900), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(n6934), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(n7255), .E(n8468), .CP(n8545), .CDN(n8421), .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(n8527), .E(n8470), .CP(n8545), .CDN(
        n8421), .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(n2220), .E(n8470), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(n2314), .E(n8469), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(n2493), .E(n8470), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(n2672), .E(n8469), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(n2849), .E(n8470), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(n3026), .E(n8469), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n3203), .E(n8470), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(n3382), .E(n8469), .CP(n8547), .CDN(
        n8420), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(n3561), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(n3880), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(n3910), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(n4089), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(n4268), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(n4445), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(n4624), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(n4803), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n5122), .E(n8469), .CP(n8547), .CDN(
        n8419), .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(n5154), .E(n8469), .CP(n8548), .CDN(
        n8419), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(n5333), .E(n8470), .CP(n8548), .CDN(
        n8419), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n5512), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(n5689), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(n5868), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n6047), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n6366), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n6400), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(n6579), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n6900), .E(n8470), .CP(n8548), .CDN(n8418), .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(n6934), .E(n8470), .CP(n8549), .CDN(n8418), .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n7255), .E(n8470), .CP(n8549), .CDN(n8418), .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n8527), .E(n8472), .CP(n8549), .CDN(
        n8418), .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(n2220), .E(n8472), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(n8757), .E(n8471), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(n8755), .E(n8472), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(n2672), .E(n8471), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(n7289), .E(n8472), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(n8747), .E(n8471), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(n8745), .E(n8472), .CP(n8549), .CDN(
        n8417), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(n2849), .E(n8471), .CP(n8550), .CDN(
        n8417), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(n3026), .E(n8472), .CP(n8550), .CDN(
        n8417), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n8737), .E(n8471), .CP(n8550), .CDN(
        n8417), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(n8735), .E(n8471), .CP(n8550), .CDN(
        n8417), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(n3561), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(n3880), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(n3910), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(n4089), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(n4268), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n8721), .E(n8471), .CP(n8550), .CDN(
        n8416), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n8719), .E(n8471), .CP(n8551), .CDN(
        n8416), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(n4803), .E(n8471), .CP(n8551), .CDN(
        n8416), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n5122), .E(n8471), .CP(n8551), .CDN(
        n8416), .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(n5154), .E(n8471), .CP(n8551), .CDN(
        n8416), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(n5333), .E(n8472), .CP(n8551), .CDN(
        n8416), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n5512), .E(n8472), .CP(n8551), .CDN(n8415), .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(n8705), .E(n8472), .CP(n8551), .CDN(n8415), .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n8703), .E(n8472), .CP(n8551), .CDN(n8415), .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n6047), .E(n8472), .CP(n8551), .CDN(n8415), .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n6366), .E(n8472), .CP(n8551), .CDN(n8415), .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n6400), .E(n8472), .CP(n8552), .CDN(n8415), .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(n6579), .E(n8472), .CP(n8552), .CDN(n8415), .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n6900), .E(n8472), .CP(n8552), .CDN(n8415), .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(n6934), .E(n8472), .CP(n8552), .CDN(n8415), .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n7255), .E(n8472), .CP(n8552), .CDN(n8415), .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n8527), .E(n8476), .CP(n8555), .CDN(
        n8412), .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(n2220), .E(n8476), .CP(n8555), .CDN(
        n8411), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(n8757), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(n8755), .E(n8476), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(n2672), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(n7289), .E(n8476), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(n8747), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(n8745), .E(n8476), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(n2849), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(n3026), .E(n8476), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n8737), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(n8735), .E(n8475), .CP(n8556), .CDN(
        n8411), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(n3561), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(n3880), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(n8728), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(n8726), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(n4268), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(n8721), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(n8719), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(n4803), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n5122), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(n8712), .E(n8475), .CP(n8557), .CDN(
        n8410), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(n8710), .E(n8476), .CP(n8558), .CDN(
        n8410), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n5512), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(n8705), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(n8703), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n6047), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n6366), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n8696), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(n8694), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n6900), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(n8689), .E(n8476), .CP(n8558), .CDN(n8409), .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n7255), .E(n8476), .CP(n8559), .CDN(n8409), .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(n8527), .E(n8482), .CP(n8565), .CDN(
        n8403), .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n8759), .E(n8482), .CP(n8565), .CDN(
        n8402), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n8757), .E(n8481), .CP(n8565), .CDN(
        n8402), .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(n8755), .E(n8482), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(n8752), .E(n8481), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(n8749), .E(n8482), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n8747), .E(n8481), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(n8745), .E(n8482), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(n8742), .E(n8481), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(n8739), .E(n8482), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(n8737), .E(n8481), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(n8735), .E(n8481), .CP(n8566), .CDN(
        n8402), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(n8732), .E(n8481), .CP(n8566), .CDN(
        n8401), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(n3880), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(n8728), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n8726), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(n8723), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(n8721), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(n8719), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n8716), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(n5122), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(n8712), .E(n8481), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(n8710), .E(n8482), .CP(n8567), .CDN(
        n8401), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(n8707), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(n8705), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(n8703), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n8700), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n6366), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(n8696), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(n8694), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(n6900), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(n8689), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n7255), .E(n8482), .CP(n8568), .CDN(n8400), .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(N85), .E(n8484), .CP(n8569), .CDN(n8400), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n8759), .E(n8484), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n8757), .E(n8483), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n8755), .E(n8484), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n8752), .E(n8483), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(n8749), .E(n8484), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n8747), .E(n8483), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n8745), .E(n8484), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n8742), .E(n8483), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(n8739), .E(n8484), .CP(n8569), .CDN(
        n8399), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n8737), .E(n8483), .CP(n8570), .CDN(
        n8399), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n8735), .E(n8483), .CP(n8570), .CDN(
        n8399), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n8732), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n3880), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(n8728), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n8726), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n8723), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n8721), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n8719), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n8716), .E(n8483), .CP(n8570), .CDN(
        n8398), .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n5122), .E(n8483), .CP(n8571), .CDN(
        n8398), .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n8712), .E(n8483), .CP(n8571), .CDN(
        n8398), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n8710), .E(n8484), .CP(n8571), .CDN(
        n8398), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n8707), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n8705), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n8703), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n8700), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n6366), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n8696), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(n8694), .E(n8484), .CP(n8571), .CDN(n8397), .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n8691), .E(n8484), .CP(n8572), .CDN(n8397), .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n8689), .E(n8484), .CP(n8572), .CDN(n8397), .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n2219), .E(n8484), .CP(n8572), .CDN(n8397), .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(n8527), .E(n8490), .CP(n8578), .CDN(
        n8391), .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(n8759), .E(n8490), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(n8757), .E(n8489), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(n8755), .E(n8490), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(n8752), .E(n8489), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(n8749), .E(n8490), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(n8747), .E(n8489), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(n8745), .E(n8490), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(n8742), .E(n8489), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(n8739), .E(n8490), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n8737), .E(n8489), .CP(n8579), .CDN(
        n8390), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(n8735), .E(n8489), .CP(n8580), .CDN(
        n8390), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(n8732), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(n2215), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(n8728), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(n8726), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(n8723), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(n8721), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(n8719), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n8716), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n2216), .E(n8489), .CP(n8580), .CDN(
        n8389), .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(n8712), .E(n8489), .CP(n8581), .CDN(
        n8389), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(n8710), .E(n8490), .CP(n8581), .CDN(
        n8389), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n8707), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(n8705), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(n8703), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n8700), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n2217), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n8696), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(n8694), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n8691), .E(n8490), .CP(n8581), .CDN(n8388), .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(n8689), .E(n8490), .CP(n8677), .CDN(n8388), .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n7255), .E(n8490), .CP(n8639), .CDN(n8388), .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n8527), .E(n8492), .CP(n8630), .CDN(
        n8388), .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n8759), .E(n8492), .CP(n8631), .CDN(
        n8387), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n8757), .E(n8491), .CP(n8632), .CDN(
        n8387), .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(n8755), .E(n8492), .CP(n8633), .CDN(
        n8387), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(n8752), .E(n8491), .CP(n8634), .CDN(
        n8387), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n8749), .E(n8492), .CP(n8635), .CDN(
        n8387), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n8747), .E(n8491), .CP(n8627), .CDN(
        n8387), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(n8745), .E(n8492), .CP(n8640), .CDN(
        n8387), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(n8742), .E(n8491), .CP(n8666), .CDN(
        n8387), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n8739), .E(n8492), .CP(n8672), .CDN(
        n8387), .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n8737), .E(n8491), .CP(n8534), .CDN(
        n8387), .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(n8735), .E(n8491), .CP(n8673), .CDN(
        n8387), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(n8732), .E(n8491), .CP(ClockW), .CDN(
        n8386), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(n2215), .E(n8491), .CP(n8535), .CDN(
        n8386), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n8728), .E(n8491), .CP(n8529), .CDN(
        n8386), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n8726), .E(n8491), .CP(n8663), .CDN(
        n8386), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(n8723), .E(n8491), .CP(n8664), .CDN(
        n8386), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(n8721), .E(n8491), .CP(n8665), .CDN(
        n8386), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(n8719), .E(n8491), .CP(n8643), .CDN(
        n8386), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n8716), .E(n8491), .CP(n8650), .CDN(
        n8386), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n2216), .E(n8491), .CP(n8649), .CDN(
        n8386), .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(n8712), .E(n8491), .CP(n8648), .CDN(
        n8386), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(n8710), .E(n8492), .CP(n8647), .CDN(
        n8386), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n8707), .E(n8492), .CP(n8646), .CDN(n8385), .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(n8705), .E(n8492), .CP(n8645), .CDN(n8385), .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(n8703), .E(n8492), .CP(n8622), .CDN(n8385), .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n8700), .E(n8492), .CP(n8623), .CDN(n8385), .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n2217), .E(n8492), .CP(n8644), .CDN(n8385), .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n8696), .E(n8492), .CP(n8628), .CDN(n8385), .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n8694), .E(n8492), .CP(n8671), .CDN(n8385), .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n8691), .E(n8492), .CP(n8642), .CDN(n8385), .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(n8689), .E(n8492), .CP(n8641), .CDN(n8385), .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n7255), .E(n8492), .CP(n8638), .CDN(n8385), .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n8527), .E(n8498), .CP(n8587), .CDN(
        n8379), .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n8759), .E(n8498), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n8757), .E(n8497), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n8755), .E(n8498), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n8752), .E(n8497), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n8749), .E(n8498), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n8747), .E(n8497), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n8745), .E(n8498), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n8742), .E(n8497), .CP(n8587), .CDN(
        n8378), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n8739), .E(n8498), .CP(n8588), .CDN(
        n8378), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n8737), .E(n8497), .CP(n8588), .CDN(
        n8378), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n8735), .E(n8497), .CP(n8588), .CDN(
        n8378), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n8732), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n2215), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n8728), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n8726), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n8723), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n8721), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n8719), .E(n8497), .CP(n8588), .CDN(
        n8377), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n8716), .E(n8497), .CP(n8589), .CDN(
        n8377), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n2216), .E(n8497), .CP(n8589), .CDN(
        n8377), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n8712), .E(n8497), .CP(n8589), .CDN(
        n8377), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n8710), .E(n8498), .CP(n8589), .CDN(
        n8377), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n8707), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n8705), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n8703), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n8700), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n2217), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n8696), .E(n8498), .CP(n8589), .CDN(n8376), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n8694), .E(n8498), .CP(n8590), .CDN(n8376), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n8691), .E(n8498), .CP(n8590), .CDN(n8376), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n8689), .E(n8498), .CP(n8590), .CDN(n8376), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n2219), .E(n8498), .CP(n8590), .CDN(n8376), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n8527), .E(n8500), .CP(n8590), .CDN(
        n8376), .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n8759), .E(n8500), .CP(n8590), .CDN(
        n8375), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n8757), .E(n8499), .CP(n8590), .CDN(
        n8375), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n8755), .E(n8500), .CP(n8590), .CDN(
        n8375), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n8752), .E(n8499), .CP(n8590), .CDN(
        n8375), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n8749), .E(n8500), .CP(n8590), .CDN(
        n8375), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n8747), .E(n8499), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n8745), .E(n8500), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n8742), .E(n8499), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n8739), .E(n8500), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n8737), .E(n8499), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n8735), .E(n8499), .CP(n8591), .CDN(
        n8375), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n8732), .E(n8499), .CP(n8591), .CDN(
        n8374), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n2215), .E(n8499), .CP(n8591), .CDN(
        n8374), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n8728), .E(n8499), .CP(n8591), .CDN(
        n8374), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n8726), .E(n8499), .CP(n8591), .CDN(
        n8374), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n8723), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n8721), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n8719), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n8716), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n2216), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n8712), .E(n8499), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n8710), .E(n8500), .CP(n8592), .CDN(
        n8374), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n8707), .E(n8500), .CP(n8592), .CDN(n8373), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n8705), .E(n8500), .CP(n8592), .CDN(n8373), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n8703), .E(n8500), .CP(n8592), .CDN(n8373), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n8700), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n2217), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n8696), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n8694), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n8691), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n8689), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n2219), .E(n8500), .CP(n8593), .CDN(n8373), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N85), .E(n8506), .CP(n8530), .CDN(n8367), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n2220), .E(n8506), .CP(n8657), .CDN(
        n8366), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n2314), .E(n8505), .CP(n8658), .CDN(
        n8366), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n2493), .E(n8506), .CP(n8659), .CDN(
        n8366), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n2672), .E(n8505), .CP(n8660), .CDN(
        n8366), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n7289), .E(n8506), .CP(n8662), .CDN(
        n8366), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n7645), .E(n8505), .CP(n8661), .CDN(
        n8366), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n7466), .E(n8506), .CP(n8629), .CDN(
        n8366), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n2849), .E(n8505), .CP(n8628), .CDN(
        n8366), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n3026), .E(n8506), .CP(n8627), .CDN(
        n8366), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n3203), .E(n8505), .CP(n8626), .CDN(
        n8366), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n3382), .E(n8505), .CP(n8625), .CDN(
        n8366), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n3561), .E(n8505), .CP(n8624), .CDN(
        n8365), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n2215), .E(n8505), .CP(n8535), .CDN(
        n8365), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n3910), .E(n8505), .CP(n8623), .CDN(
        n8365), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n4089), .E(n8505), .CP(n8675), .CDN(
        n8365), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n4268), .E(n8505), .CP(n8629), .CDN(
        n8365), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n4445), .E(n8505), .CP(n8634), .CDN(
        n8365), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n4624), .E(n8505), .CP(n8633), .CDN(
        n8365), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n4803), .E(n8505), .CP(n8635), .CDN(
        n8365), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n2216), .E(n8505), .CP(n8638), .CDN(
        n8365), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n5154), .E(n8505), .CP(n8642), .CDN(
        n8365), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n5333), .E(n8506), .CP(n8643), .CDN(
        n8365), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n5512), .E(n8506), .CP(n8644), .CDN(n8364), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n5689), .E(n8506), .CP(n8637), .CDN(n8364), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n5868), .E(n8506), .CP(n8673), .CDN(n8364), .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n6047), .E(n8506), .CP(n8622), .CDN(n8364), .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n2217), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n6400), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n6579), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n8691), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n6934), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n2219), .E(n8506), .CP(n8597), .CDN(n8364), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N85), .E(n8508), .CP(n8597), .CDN(n8364), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n8759), .E(n8508), .CP(n8597), .CDN(n8363), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n2314), .E(n8507), .CP(n8597), .CDN(n8363), .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n2493), .E(n8508), .CP(n8597), .CDN(n8363), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n8752), .E(n8507), .CP(n8598), .CDN(n8363), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n8749), .E(n8508), .CP(n8598), .CDN(n8363), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n7645), .E(n8507), .CP(n8598), .CDN(n8363), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n7466), .E(n8508), .CP(n8598), .CDN(n8363), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n8742), .E(n8507), .CP(n8598), .CDN(n8363), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n8739), .E(n8508), .CP(n8598), .CDN(n8363), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n3203), .E(n8507), .CP(n8598), .CDN(n8363), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n3382), .E(n8507), .CP(n8598), .CDN(n8363), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n8732), .E(n8507), .CP(n8598), .CDN(n8362), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n2215), .E(n8507), .CP(n8598), .CDN(n8362), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n3910), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n4089), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n8723), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n4445), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n4624), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n8716), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n2216), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n5154), .E(n8507), .CP(n8599), .CDN(n8362), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n5333), .E(n8508), .CP(n8599), .CDN(n8362), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n8707), .E(n8508), .CP(n8599), .CDN(n8361), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n5689), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n5868), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n8700), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n2217), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n6400), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n6579), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n2218), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n6934), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n2219), .E(n8508), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n8527), .E(n8514), .CP(n8660), .CDN(n8355), .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n8759), .E(n8514), .CP(n8531), .CDN(n8354), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n2314), .E(n8513), .CP(n8669), .CDN(n8354), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n2493), .E(n8514), .CP(n8670), .CDN(n8354), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n8752), .E(n8513), .CP(n8675), .CDN(n8354), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n8749), .E(n8514), .CP(n8655), .CDN(n8354), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n7645), .E(n8513), .CP(n8651), .CDN(n8354), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n7466), .E(n8514), .CP(n8674), .CDN(n8354), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n8742), .E(n8513), .CP(ClockW), .CDN(
        n8354), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n8739), .E(n8514), .CP(n8661), .CDN(n8354), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n3203), .E(n8513), .CP(n8662), .CDN(n8354), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n3382), .E(n8513), .CP(n8657), .CDN(n8354), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n8732), .E(n8513), .CP(n8658), .CDN(n8353), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n2215), .E(n8513), .CP(n8659), .CDN(n8353), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n3910), .E(n8513), .CP(n8654), .CDN(n8353), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n4089), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n8723), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n4445), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n4624), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n8716), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n2216), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n5154), .E(n8513), .CP(n8604), .CDN(n8353), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n5333), .E(n8514), .CP(n8604), .CDN(n8353), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n8707), .E(n8514), .CP(n8604), .CDN(n8352), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n5689), .E(n8514), .CP(n8604), .CDN(n8352), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n5868), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n8700), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n2217), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n6400), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n6579), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n2218), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n6934), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n2219), .E(n8514), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N85), .E(n8516), .CP(n8605), .CDN(n8352), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n8759), .E(n8516), .CP(n8605), .CDN(n8351), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n2314), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n2493), .E(n8516), .CP(n8606), .CDN(n8351), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n8752), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n8749), .E(n8516), .CP(n8606), .CDN(n8351), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n7645), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n7466), .E(n8516), .CP(n8606), .CDN(n8351), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n8742), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n8739), .E(n8516), .CP(n8606), .CDN(n8351), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n3203), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n3382), .E(n8515), .CP(n8606), .CDN(n8351), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n8732), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n2215), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n3910), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n4089), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n8723), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n4445), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n4624), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n8716), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n2216), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n5154), .E(n8515), .CP(n8607), .CDN(n8350), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n5333), .E(n8516), .CP(n8608), .CDN(n8350), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n8707), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n5689), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n5868), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n8700), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n2217), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n6400), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n6579), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n2218), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n6934), .E(n8516), .CP(n8608), .CDN(n8349), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n2219), .E(n8516), .CP(n8609), .CDN(n8349), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(n8522), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n8759), .E(n8522), .CP(n8615), .CDN(n8342), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n2314), .E(n8521), .CP(n8615), .CDN(n8342), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n2493), .E(n8522), .CP(n8616), .CDN(n8342), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n8752), .E(n8521), .CP(n8616), .CDN(n8342), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n8749), .E(n8522), .CP(n8616), .CDN(n8342), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n7645), .E(n8521), .CP(n8616), .CDN(n8342), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n7466), .E(n8522), .CP(n8616), .CDN(n8342), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n8742), .E(n8521), .CP(n8616), .CDN(n8342), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n8739), .E(n8522), .CP(n8616), .CDN(n8342), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n3203), .E(n8521), .CP(n8616), .CDN(n8342), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n3382), .E(n8521), .CP(n8616), .CDN(n8342), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n8732), .E(n8521), .CP(n8616), .CDN(n8341), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n2215), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n3910), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n4089), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n8723), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n4445), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n4624), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n8716), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n2216), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n5154), .E(n8521), .CP(n8617), .CDN(n8341), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n5333), .E(n8522), .CP(n8617), .CDN(n8341), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n8707), .E(n8522), .CP(n8656), .CDN(n8340), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n5689), .E(n8522), .CP(n8638), .CDN(n8340), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n5868), .E(n8522), .CP(n8531), .CDN(n8340), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n8700), .E(n8522), .CP(n8650), .CDN(n8340), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n2217), .E(n8522), .CP(n8649), .CDN(n8340), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n6400), .E(n8522), .CP(n8648), .CDN(n8340), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n6579), .E(n8522), .CP(n8647), .CDN(n8340), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n2218), .E(n8522), .CP(n8646), .CDN(n8340), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n6934), .E(n8522), .CP(n8645), .CDN(n8340), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n2219), .E(n8522), .CP(n8530), .CDN(n8340), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N85), .E(n8524), .CP(n8653), .CDN(n8340), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n8759), .E(n8524), .CP(n8652), .CDN(n8339), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n2314), .E(n8523), .CP(n8659), .CDN(n8339), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n2493), .E(n8524), .CP(n8658), .CDN(n8339), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n8752), .E(n8523), .CP(n8657), .CDN(n8339), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n8749), .E(n8524), .CP(n8662), .CDN(n8339), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n7645), .E(n8523), .CP(n8661), .CDN(n8339), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n7466), .E(n8524), .CP(n8660), .CDN(n8339), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n8742), .E(n8523), .CP(n8655), .CDN(n8339), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n8739), .E(n8524), .CP(n8654), .CDN(n8339), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n3203), .E(n8523), .CP(n8532), .CDN(n8339), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n3382), .E(n8523), .CP(n8637), .CDN(n8339), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n8732), .E(n8523), .CP(n8651), .CDN(n8338), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n2215), .E(n8523), .CP(n8640), .CDN(n8338), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n3910), .E(n8523), .CP(n8644), .CDN(n8338), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n4089), .E(n8523), .CP(n8643), .CDN(n8338), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n8723), .E(n8523), .CP(n8642), .CDN(n8338), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n4445), .E(n8523), .CP(n8641), .CDN(n8338), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n4624), .E(n8523), .CP(n8637), .CDN(n8338), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n8716), .E(n8523), .CP(n8668), .CDN(n8338), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n2216), .E(n8523), .CP(n8640), .CDN(n8338), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n5154), .E(n8523), .CP(n8639), .CDN(n8338), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n5333), .E(n8524), .CP(n8533), .CDN(n8338), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n8707), .E(n8524), .CP(n8635), .CDN(n8337), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n5689), .E(n8524), .CP(n8634), .CDN(n8337), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n5868), .E(n8524), .CP(n8633), .CDN(n8337), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n8700), .E(n8524), .CP(n8628), .CDN(n8337), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n2217), .E(n8524), .CP(n8645), .CDN(n8337), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n6400), .E(n8524), .CP(n8673), .CDN(n8337), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n6579), .E(n8524), .CP(n8629), .CDN(n8337), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n2218), .E(n8524), .CP(n8618), .CDN(n8337), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n6934), .E(n8524), .CP(n8618), .CDN(n8337), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n2219), .E(n8524), .CP(n8618), .CDN(n8337), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n8527), .E(n8480), .CP(n8562), .CDN(
        n8406), .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(n2220), .E(n8480), .CP(n8562), .CDN(
        n8405), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(n8757), .E(n8479), .CP(n8562), .CDN(
        n8405), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(n8755), .E(n8480), .CP(n8562), .CDN(
        n8405), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(n2672), .E(n8479), .CP(n8562), .CDN(
        n8405), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(n7289), .E(n8480), .CP(n8562), .CDN(
        n8405), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(n8747), .E(n8479), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(n8745), .E(n8480), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(n2849), .E(n8479), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(n3026), .E(n8480), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n8737), .E(n8479), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(n8735), .E(n8479), .CP(n8563), .CDN(
        n8405), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(n3561), .E(n8479), .CP(n8563), .CDN(
        n8404), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(n3880), .E(n8479), .CP(n8563), .CDN(
        n8404), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(n8728), .E(n8479), .CP(n8563), .CDN(
        n8404), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(n8726), .E(n8479), .CP(n8563), .CDN(
        n8404), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(n4268), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(n8721), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(n8719), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n4803), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n5122), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(n8712), .E(n8479), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(n8710), .E(n8480), .CP(n8564), .CDN(
        n8404), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n5512), .E(n8480), .CP(n8564), .CDN(n8403), .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(n8705), .E(n8480), .CP(n8564), .CDN(n8403), .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(n8703), .E(n8480), .CP(n8564), .CDN(n8403), .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n6047), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n6366), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n8696), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(n8694), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n6900), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(n8689), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n7255), .E(n8480), .CP(n8565), .CDN(n8403), .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(n8527), .E(n8486), .CP(n8572), .CDN(
        n8397), .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(n8759), .E(n8486), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(n8757), .E(n8485), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(n8755), .E(n8486), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(n8752), .E(n8485), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(n8749), .E(n8486), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(n8747), .E(n8485), .CP(n8572), .CDN(
        n8396), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(n8745), .E(n8486), .CP(n8573), .CDN(
        n8396), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(n8742), .E(n8485), .CP(n8573), .CDN(
        n8396), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(n8739), .E(n8486), .CP(n8573), .CDN(
        n8396), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n8737), .E(n8485), .CP(n8573), .CDN(
        n8396), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(n8735), .E(n8485), .CP(n8573), .CDN(
        n8396), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(n8732), .E(n8485), .CP(n8573), .CDN(
        n8395), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(n2215), .E(n8485), .CP(n8573), .CDN(
        n8395), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(n8728), .E(n8485), .CP(n8573), .CDN(
        n8395), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(n8726), .E(n8485), .CP(n8573), .CDN(
        n8395), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(n8723), .E(n8485), .CP(n8573), .CDN(
        n8395), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(n8721), .E(n8485), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(n8719), .E(n8485), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(n8716), .E(n8485), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n2216), .E(n8485), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(n8712), .E(n8485), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(n8710), .E(n8486), .CP(n8574), .CDN(
        n8395), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n8707), .E(n8486), .CP(n8574), .CDN(n8394), .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(n8705), .E(n8486), .CP(n8574), .CDN(n8394), .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(n8703), .E(n8486), .CP(n8574), .CDN(n8394), .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n8700), .E(n8486), .CP(n8574), .CDN(n8394), .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n2217), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n8696), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(n8694), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n8691), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(n8689), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n2219), .E(n8486), .CP(n8575), .CDN(n8394), .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(N85), .E(n8488), .CP(n8575), .CDN(n8394), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(n8759), .E(n8488), .CP(n8575), .CDN(
        n8393), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(n8757), .E(n8487), .CP(n8575), .CDN(
        n8393), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(n8755), .E(n8488), .CP(n8575), .CDN(
        n8393), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(n8752), .E(n8487), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(n8749), .E(n8488), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(n8747), .E(n8487), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(n8745), .E(n8488), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(n8742), .E(n8487), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(n8739), .E(n8488), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n8737), .E(n8487), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(n8735), .E(n8487), .CP(n8576), .CDN(
        n8393), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(n8732), .E(n8487), .CP(n8576), .CDN(
        n8392), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(n2215), .E(n8487), .CP(n8576), .CDN(
        n8392), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(n8728), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(n8726), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(n8723), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(n8721), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(n8719), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(n8716), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n2216), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(n8712), .E(n8487), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(n8710), .E(n8488), .CP(n8577), .CDN(
        n8392), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n8707), .E(n8488), .CP(n8577), .CDN(n8391), .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(n8705), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(n8703), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n8700), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n2217), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n8696), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(n8694), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n8691), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(n8689), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n2219), .E(n8488), .CP(n8578), .CDN(n8391), .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(n8494), .CP(n8667), .CDN(n8385), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(n8759), .E(n8494), .CP(n8624), .CDN(
        n8384), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(n8757), .E(n8493), .CP(n8625), .CDN(
        n8384), .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(n8755), .E(n8494), .CP(n8626), .CDN(
        n8384), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(n8752), .E(n8493), .CP(n8627), .CDN(
        n8384), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(n8749), .E(n8494), .CP(n8531), .CDN(
        n8384), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(n8747), .E(n8493), .CP(n8676), .CDN(
        n8384), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(n8745), .E(n8494), .CP(n8669), .CDN(
        n8384), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(n8742), .E(n8493), .CP(n8534), .CDN(
        n8384), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(n8739), .E(n8494), .CP(n8636), .CDN(
        n8384), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n8737), .E(n8493), .CP(n8639), .CDN(
        n8384), .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(n8735), .E(n8493), .CP(n8632), .CDN(
        n8384), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(n8732), .E(n8493), .CP(n8631), .CDN(
        n8383), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(n3880), .E(n8493), .CP(n8630), .CDN(
        n8383), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(n8728), .E(n8493), .CP(n8532), .CDN(
        n8383), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(n8726), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(n8723), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(n8721), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(n8719), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(n8716), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n5122), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(n8712), .E(n8493), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(n8710), .E(n8494), .CP(n8582), .CDN(
        n8383), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n8707), .E(n8494), .CP(n8582), .CDN(n8382), .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(n8705), .E(n8494), .CP(n8582), .CDN(n8382), .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(n8703), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n8700), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n6366), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n8696), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(n8694), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n8691), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(n8689), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n7255), .E(n8494), .CP(n8583), .CDN(n8382), .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N85), .E(n8496), .CP(n8583), .CDN(n8382), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n8759), .E(n8496), .CP(n8583), .CDN(
        n8381), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n8757), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n8755), .E(n8496), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n8752), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n8749), .E(n8496), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n8747), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n8745), .E(n8496), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n8742), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n8739), .E(n8496), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n8737), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n8735), .E(n8495), .CP(n8584), .CDN(
        n8381), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n8732), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n3880), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n8728), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n8726), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n8723), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n8721), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n8719), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n8716), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n5122), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n8712), .E(n8495), .CP(n8585), .CDN(
        n8380), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n8710), .E(n8496), .CP(n8586), .CDN(
        n8380), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n8707), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n8705), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n8703), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n8700), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n6366), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n8696), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n8694), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n8691), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n8689), .E(n8496), .CP(n8586), .CDN(n8379), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n7255), .E(n8496), .CP(n8587), .CDN(n8379), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(n8502), .CP(n8593), .CDN(n8373), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n8759), .E(n8502), .CP(n8593), .CDN(
        n8372), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n2314), .E(n8501), .CP(n8593), .CDN(
        n8372), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n2493), .E(n8502), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n8752), .E(n8501), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n8749), .E(n8502), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n7645), .E(n8501), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n7466), .E(n8502), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n8742), .E(n8501), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n8739), .E(n8502), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n3203), .E(n8501), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n3382), .E(n8501), .CP(n8594), .CDN(
        n8372), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n8732), .E(n8501), .CP(n8594), .CDN(
        n8371), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n3880), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n3910), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n4089), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n8723), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n4445), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n4624), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n8716), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n5122), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n5154), .E(n8501), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n5333), .E(n8502), .CP(n8595), .CDN(
        n8371), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n8707), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n5689), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n5868), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n8700), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n6366), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n6400), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n6579), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n8691), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n6934), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n7255), .E(n8502), .CP(n8596), .CDN(n8370), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N85), .E(n8504), .CP(n8648), .CDN(n8370), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n8759), .E(n8504), .CP(n8645), .CDN(
        n8369), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n2314), .E(n8503), .CP(n8646), .CDN(
        n8369), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n2493), .E(n8504), .CP(n8647), .CDN(
        n8369), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n8752), .E(n8503), .CP(n8531), .CDN(
        n8369), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n8749), .E(n8504), .CP(n8533), .CDN(
        n8369), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n7645), .E(n8503), .CP(n8669), .CDN(
        n8369), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n7466), .E(n8504), .CP(n8670), .CDN(
        n8369), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n8742), .E(n8503), .CP(n8661), .CDN(
        n8369), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n8739), .E(n8504), .CP(n8649), .CDN(
        n8369), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n3203), .E(n8503), .CP(n8663), .CDN(
        n8369), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n3382), .E(n8503), .CP(n8666), .CDN(
        n8369), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n8732), .E(n8503), .CP(n8665), .CDN(
        n8368), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n3880), .E(n8503), .CP(n8668), .CDN(
        n8368), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n3910), .E(n8503), .CP(n8677), .CDN(
        n8368), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n4089), .E(n8503), .CP(n8672), .CDN(
        n8368), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n8723), .E(n8503), .CP(n8674), .CDN(
        n8368), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n4445), .E(n8503), .CP(n8667), .CDN(
        n8368), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n4624), .E(n8503), .CP(n8673), .CDN(
        n8368), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n8716), .E(n8503), .CP(n8676), .CDN(
        n8368), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n5122), .E(n8503), .CP(n8648), .CDN(
        n8368), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n5154), .E(n8503), .CP(n8649), .CDN(
        n8368), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n5333), .E(n8504), .CP(n8650), .CDN(
        n8368), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n8707), .E(n8504), .CP(n8651), .CDN(n8367), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n5689), .E(n8504), .CP(n8653), .CDN(n8367), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n5868), .E(n8504), .CP(n8652), .CDN(n8367), .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n8700), .E(n8504), .CP(n8654), .CDN(n8367), .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n6366), .E(n8504), .CP(n8655), .CDN(n8367), .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n6400), .E(n8504), .CP(n8641), .CDN(n8367), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n6579), .E(n8504), .CP(n8647), .CDN(n8367), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n8691), .E(n8504), .CP(n8533), .CDN(n8367), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n6934), .E(n8504), .CP(n8646), .CDN(n8367), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n2219), .E(n8504), .CP(n8656), .CDN(n8367), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(n8510), .CP(n8600), .CDN(n8361), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n8759), .E(n8510), .CP(n8601), .CDN(n8360), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n2314), .E(n8509), .CP(n8601), .CDN(n8360), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n2493), .E(n8510), .CP(n8601), .CDN(n8360), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n8752), .E(n8509), .CP(n8601), .CDN(n8360), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n8749), .E(n8510), .CP(n8601), .CDN(n8360), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n7645), .E(n8509), .CP(n8601), .CDN(n8360), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n7466), .E(n8510), .CP(n8601), .CDN(n8360), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n8742), .E(n8509), .CP(n8601), .CDN(n8360), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n8739), .E(n8510), .CP(n8601), .CDN(n8360), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n3203), .E(n8509), .CP(n8601), .CDN(n8360), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n3382), .E(n8509), .CP(n8602), .CDN(n8360), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n8732), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n2215), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n3910), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n4089), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n8723), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n4445), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n4624), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n8716), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n2216), .E(n8509), .CP(n8602), .CDN(n8359), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n5154), .E(n8509), .CP(n8603), .CDN(n8359), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n5333), .E(n8510), .CP(n8603), .CDN(n8359), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n8707), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n5689), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n5868), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n8700), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n2217), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n6400), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n6579), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n2218), .E(n8510), .CP(n8603), .CDN(n8358), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n6934), .E(n8510), .CP(n8631), .CDN(n8358), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n2219), .E(n8510), .CP(n8630), .CDN(n8358), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N85), .E(n8512), .CP(n8534), .CDN(n8358), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n8759), .E(n8512), .CP(n8624), .CDN(n8357), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n2314), .E(n8511), .CP(n8625), .CDN(n8357), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n2493), .E(n8512), .CP(n8626), .CDN(n8357), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n8752), .E(n8511), .CP(n8627), .CDN(n8357), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n8749), .E(n8512), .CP(n8628), .CDN(n8357), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n7645), .E(n8511), .CP(n8629), .CDN(n8357), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n7466), .E(n8512), .CP(n8632), .CDN(n8357), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n8742), .E(n8511), .CP(n8529), .CDN(n8357), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n8739), .E(n8512), .CP(n8671), .CDN(n8357), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n3203), .E(n8511), .CP(n8623), .CDN(n8357), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n3382), .E(n8511), .CP(n8622), .CDN(n8357), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n8732), .E(n8511), .CP(n8656), .CDN(n8356), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n2215), .E(n8511), .CP(n8653), .CDN(n8356), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n3910), .E(n8511), .CP(n8652), .CDN(n8356), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n4089), .E(n8511), .CP(n8533), .CDN(n8356), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n8723), .E(n8511), .CP(ClockW), .CDN(
        n8356), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n4445), .E(n8511), .CP(n8535), .CDN(n8356), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n4624), .E(n8511), .CP(n8670), .CDN(n8356), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n8716), .E(n8511), .CP(n8636), .CDN(n8356), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n2216), .E(n8511), .CP(n8663), .CDN(n8356), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n5154), .E(n8511), .CP(n8664), .CDN(n8356), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n5333), .E(n8512), .CP(n8665), .CDN(n8356), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n8707), .E(n8512), .CP(n8666), .CDN(n8355), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n5689), .E(n8512), .CP(n8667), .CDN(n8355), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n5868), .E(n8512), .CP(n8668), .CDN(n8355), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n8700), .E(n8512), .CP(n8672), .CDN(n8355), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n2217), .E(n8512), .CP(n8673), .CDN(n8355), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n6400), .E(n8512), .CP(n8676), .CDN(n8355), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n6579), .E(n8512), .CP(n8674), .CDN(n8355), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n2218), .E(n8512), .CP(n8677), .CDN(n8355), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n6934), .E(n8512), .CP(n8530), .CDN(n8355), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n2219), .E(n8512), .CP(n8532), .CDN(n8355), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(n8518), .CP(n8609), .CDN(n8349), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n8759), .E(n8518), .CP(n8609), .CDN(n8348), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n2314), .E(n8517), .CP(n8609), .CDN(n8348), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n2493), .E(n8518), .CP(n8609), .CDN(n8348), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n8752), .E(n8517), .CP(n8609), .CDN(n8348), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n8749), .E(n8518), .CP(n8609), .CDN(n8348), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n7645), .E(n8517), .CP(n8609), .CDN(n8348), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n7466), .E(n8518), .CP(n8609), .CDN(n8348), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n8742), .E(n8517), .CP(n8609), .CDN(n8348), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n8739), .E(n8518), .CP(n8610), .CDN(n8348), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n3203), .E(n8517), .CP(n8610), .CDN(n8348), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n3382), .E(n8517), .CP(n8610), .CDN(n8348), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n8732), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n2215), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n3910), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n4089), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n8723), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n4445), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n4624), .E(n8517), .CP(n8610), .CDN(n8347), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n8716), .E(n8517), .CP(n8611), .CDN(n8347), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n2216), .E(n8517), .CP(n8611), .CDN(n8347), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n5154), .E(n8517), .CP(n8611), .CDN(n8347), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n5333), .E(n8518), .CP(n8611), .CDN(n8347), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n8707), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n5689), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n5868), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n8700), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n2217), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n6400), .E(n8518), .CP(n8611), .CDN(n8346), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n6579), .E(n8518), .CP(n8612), .CDN(n8346), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n2218), .E(n8518), .CP(n8612), .CDN(n8346), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n6934), .E(n8518), .CP(n8612), .CDN(n8346), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n2219), .E(n8518), .CP(n8612), .CDN(n8346), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N85), .E(n8520), .CP(n8612), .CDN(n8346), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n2220), .E(n8520), .CP(n8612), .CDN(n8345), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n2314), .E(n8519), .CP(n8612), .CDN(n8345), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n2493), .E(n8520), .CP(n8612), .CDN(n8345), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n2672), .E(n8519), .CP(n8612), .CDN(n8345), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n7289), .E(n8520), .CP(n8612), .CDN(n8345), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n7645), .E(n8519), .CP(n8613), .CDN(n8345), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n7466), .E(n8520), .CP(n8613), .CDN(n8345), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n2849), .E(n8519), .CP(n8613), .CDN(n8345), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n3026), .E(n8520), .CP(n8613), .CDN(n8345), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n3203), .E(n8519), .CP(n8613), .CDN(n8345), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n3382), .E(n8519), .CP(n8613), .CDN(n8345), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n3561), .E(n8519), .CP(n8613), .CDN(n8344), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n2215), .E(n8519), .CP(n8613), .CDN(n8344), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n3910), .E(n8519), .CP(n8613), .CDN(n8344), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n4089), .E(n8519), .CP(n8613), .CDN(n8344), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n4268), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n4445), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n4624), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n4803), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n2216), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n5154), .E(n8519), .CP(n8614), .CDN(n8344), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n5333), .E(n8520), .CP(n8614), .CDN(n8344), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n5512), .E(n8520), .CP(n8614), .CDN(n8343), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n5689), .E(n8520), .CP(n8614), .CDN(n8343), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n5868), .E(n8520), .CP(n8614), .CDN(n8343), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n6047), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n2217), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n6400), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n6579), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n2218), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n6934), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n2219), .E(n8520), .CP(n8615), .CDN(n8343), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(n8526), .CP(n8618), .CDN(n8337), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n2220), .E(n8526), .CP(n8618), .CDN(n8336), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n2314), .E(n8525), .CP(n8618), .CDN(n8336), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n2493), .E(n8526), .CP(n8618), .CDN(n8336), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n2672), .E(n8525), .CP(n8618), .CDN(n8336), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n7289), .E(n8526), .CP(n8618), .CDN(n8336), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n7645), .E(n8525), .CP(n8618), .CDN(n8336), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n7466), .E(n8526), .CP(n8619), .CDN(n8336), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n2849), .E(n8525), .CP(n8619), .CDN(n8336), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n3026), .E(n8526), .CP(n8619), .CDN(n8336), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n3203), .E(n8525), .CP(n8619), .CDN(n8336), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n3382), .E(n8525), .CP(n8619), .CDN(n8336), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n3561), .E(n8525), .CP(n8619), .CDN(n8335), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n2215), .E(n8525), .CP(n8619), .CDN(n8335), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n3910), .E(n8525), .CP(n8619), .CDN(n8335), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n4089), .E(n8525), .CP(n8619), .CDN(n8335), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n4268), .E(n8525), .CP(n8619), .CDN(n8335), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n4445), .E(n8525), .CP(n8620), .CDN(n8335), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n4624), .E(n8525), .CP(n8620), .CDN(n8335), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n4803), .E(n8525), .CP(n8620), .CDN(n8335), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n2216), .E(n8525), .CP(n8620), .CDN(n8335), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n5154), .E(n8525), .CP(n8620), .CDN(n8335), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n5333), .E(n8526), .CP(n8620), .CDN(n8335), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n5512), .E(n8526), .CP(n8620), .CDN(n8334), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n5689), .E(n8526), .CP(n8620), .CDN(n8334), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n5868), .E(n8526), .CP(n8620), .CDN(n8334), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n6047), .E(n8526), .CP(n8620), .CDN(n8334), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n2217), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n6400), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n6579), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n2218), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n6934), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n2219), .E(n8526), .CP(n8621), .CDN(n8334), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n8527), .E(n8464), .CP(n8536), .CDN(
        n8349), .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(n2220), .E(n8464), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(n2314), .E(n8463), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(n2493), .E(n8464), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(n2672), .E(n8463), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(n7289), .E(n8464), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(n7466), .E(n8463), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(n2849), .E(n8464), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(n3026), .E(n8463), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(n3203), .E(n8464), .CP(n8537), .CDN(
        n8429), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(n3382), .E(n8463), .CP(n8537), .CDN(
        n8429), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(n3561), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(n3880), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(n3910), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(n4089), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(n4268), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(n4445), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(n4624), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(n4803), .E(n8463), .CP(n8537), .CDN(
        n8428), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(n5122), .E(n8463), .CP(n8538), .CDN(
        n8428), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(n5154), .E(n8463), .CP(n8538), .CDN(
        n8428), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(n5333), .E(n8464), .CP(n8538), .CDN(
        n8428), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(n5512), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(n5689), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(n5868), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n6047), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(n6366), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(n6400), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(n6579), .E(n8464), .CP(n8538), .CDN(n8427), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(n6900), .E(n8464), .CP(n8539), .CDN(n8427), .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(n6934), .E(n8464), .CP(n8539), .CDN(n8427), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(n7255), .E(n8464), .CP(n8539), .CDN(n8427), .Q(\Storage[31][0] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(n7645), .E(n8466), .CP(n8539), .CDN(
        n8426), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(n7466), .E(n8465), .CP(n8540), .CDN(
        n8426), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(n7645), .E(n8468), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(n7466), .E(n8467), .CP(n8543), .CDN(
        n8423), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(n7289), .E(n8469), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(n7645), .E(n8470), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(n7466), .E(n8469), .CP(n8546), .CDN(
        n8420), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(n7645), .E(n8463), .CP(n8536), .CDN(
        n8429), .Q(\Storage[31][26] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n4), .E(n8682), .CP(n8678), .CDN(n8423), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n112), .E(n8682), .CP(ClockR), .CDN(n8354), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n178), .E(n8682), .CP(ClockR), .CDN(n8422), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n244), .E(n8682), .CP(ClockR), .CDN(n8343), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n310), .E(n8682), .CP(ClockR), .CDN(n8347), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n376), .E(n8682), .CP(ClockR), .CDN(n8357), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n442), .E(n8682), .CP(n8678), .CDN(n8346), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n508), .E(n8682), .CP(ClockR), .CDN(n8435), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n574), .E(n8682), .CP(ClockR), .CDN(n8454), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n640), .E(n8682), .CP(n8678), .CDN(n8345), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n706), .E(n8682), .CP(n8678), .CDN(n8451), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n772), .E(n8683), .CP(ClockR), .CDN(n8452), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n838), .E(n8683), .CP(n8678), .CDN(n8429), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n904), .E(n8683), .CP(ClockR), .CDN(n8344), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n970), .E(n8683), .CP(n8678), .CDN(n8342), 
        .Q(DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n1036), .E(n8683), .CP(ClockR), .CDN(n8428), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n1100), .E(n8683), .CP(n8678), .CDN(n8412), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n1), .E(n8683), .CP(ClockR), .CDN(n8427), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n1227), .E(n8683), .CP(n8678), .CDN(n8426), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n1291), .E(n8683), .CP(ClockR), .CDN(n8413), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n1355), .E(n8683), .CP(n8678), .CDN(n8425), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n1419), .E(n8683), .CP(n8678), .CDN(n8348), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n1481), .E(n8684), .CP(n8678), .CDN(n8424), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n1540), .E(n8684), .CP(n8678), .CDN(n8333), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n1598), .E(n8684), .CP(n8678), .CDN(n8449), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n1660), .E(n8684), .CP(n8678), .CDN(n8450), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n1721), .E(n8684), .CP(n8678), .CDN(n8355), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n1781), .E(n8684), .CP(n8678), .CDN(n8354), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n2), .E(n8684), .CP(n8678), .CDN(n8334), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n1900), .E(n8684), .CP(n8678), .CDN(n8356), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n1961), .E(n8684), .CP(ClockR), .CDN(n8357), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n3), .E(n8684), .CP(ClockR), .CDN(n8355), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n2100), .E(n8684), .CP(ClockR), .CDN(n8356), .Q(
        ParityErr) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  EDFCNQD1 Dreadyr_reg ( .D(n7827), .E(n7824), .CP(ClockR), .CDN(n8453), .Q(
        Dreadyr) );
  TIEH U3 ( .Z(n7827) );
  MUX3ND1 U4 ( .I0(n8260), .I1(n8261), .I2(n177), .S0(n8293), .S1(n8291), .ZN(
        N52) );
  MUX3ND1 U5 ( .I0(n8247), .I1(n8248), .I2(n243), .S0(n8293), .S1(n8291), .ZN(
        N53) );
  MUX3ND1 U6 ( .I0(n8234), .I1(n8235), .I2(n309), .S0(n8293), .S1(n8291), .ZN(
        N54) );
  MUX3ND1 U7 ( .I0(n8221), .I1(n8222), .I2(n375), .S0(n8293), .S1(n8291), .ZN(
        N55) );
  MUX3ND1 U8 ( .I0(n8208), .I1(n8209), .I2(n441), .S0(n8293), .S1(n8291), .ZN(
        N56) );
  MUX3ND1 U9 ( .I0(n8195), .I1(n8196), .I2(n507), .S0(n8686), .S1(n8291), .ZN(
        N57) );
  MUX3ND1 U10 ( .I0(n8182), .I1(n8183), .I2(n573), .S0(n8686), .S1(n8291), 
        .ZN(N58) );
  MUX3ND1 U11 ( .I0(n8169), .I1(n8170), .I2(n639), .S0(n8293), .S1(n8291), 
        .ZN(N59) );
  MUX3ND1 U12 ( .I0(n8156), .I1(n8157), .I2(n705), .S0(N47), .S1(n8291), .ZN(
        N60) );
  MUX3ND1 U13 ( .I0(n8143), .I1(n8144), .I2(n771), .S0(n8686), .S1(n8291), 
        .ZN(N61) );
  MUX3ND1 U14 ( .I0(n8130), .I1(n8131), .I2(n837), .S0(n8686), .S1(n8291), 
        .ZN(N62) );
  MUX3ND1 U15 ( .I0(n8104), .I1(n8105), .I2(n969), .S0(n8686), .S1(n8290), 
        .ZN(N64) );
  MUX3ND1 U16 ( .I0(n8091), .I1(n8092), .I2(n1035), .S0(N47), .S1(n8290), .ZN(
        N65) );
  MUX3ND1 U17 ( .I0(n8078), .I1(n8079), .I2(n2153), .S0(n8686), .S1(n8290), 
        .ZN(N66) );
  CKBD0 U23 ( .CLK(N67), .C(n1161) );
  BUFFD0 U24 ( .I(n1164), .Z(n1) );
  MUX3ND1 U25 ( .I0(n8026), .I1(n8027), .I2(n2158), .S0(N47), .S1(n8290), .ZN(
        N70) );
  CKBD0 U26 ( .CLK(N71), .C(n1416) );
  CKBD0 U29 ( .CLK(n2177), .C(n2167) );
  CKBD0 U30 ( .CLK(n2174), .C(n2162) );
  CKBD0 U31 ( .CLK(n2176), .C(n2164) );
  CKBD0 U32 ( .CLK(n2170), .C(n2154) );
  CKBD0 U37 ( .CLK(n2175), .C(n2163) );
  BUFFD0 U38 ( .I(n1842), .Z(n2) );
  CKBD0 U39 ( .CLK(n2171), .C(n2156) );
  BUFFD0 U40 ( .I(n2022), .Z(n3) );
  XOR3D0 U41 ( .A1(n2096), .A2(n2093), .A3(n86), .Z(N83) );
  CKBD0 U42 ( .CLK(n8687), .C(n2219) );
  INVD0 U43 ( .I(n8528), .ZN(n8527) );
  INVD1 U44 ( .I(DataI[2]), .ZN(n8693) );
  CKBD0 U45 ( .CLK(n6758), .C(n2214) );
  INVD0 U46 ( .I(n6758), .ZN(n8692) );
  INVD0 U47 ( .I(n2214), .ZN(n8691) );
  BUFFD0 U48 ( .I(n5), .Z(n4) );
  BUFFD0 U49 ( .I(n6), .Z(n5) );
  BUFFD0 U50 ( .I(n7), .Z(n6) );
  BUFFD0 U51 ( .I(n8), .Z(n7) );
  BUFFD0 U52 ( .I(n9), .Z(n8) );
  BUFFD0 U53 ( .I(n10), .Z(n9) );
  BUFFD0 U54 ( .I(n11), .Z(n10) );
  BUFFD0 U55 ( .I(n12), .Z(n11) );
  BUFFD0 U56 ( .I(n13), .Z(n12) );
  BUFFD0 U57 ( .I(n14), .Z(n13) );
  BUFFD0 U58 ( .I(n15), .Z(n14) );
  BUFFD0 U59 ( .I(n16), .Z(n15) );
  BUFFD0 U60 ( .I(n17), .Z(n16) );
  BUFFD0 U61 ( .I(n18), .Z(n17) );
  BUFFD0 U62 ( .I(n19), .Z(n18) );
  BUFFD0 U63 ( .I(n20), .Z(n19) );
  BUFFD0 U64 ( .I(n21), .Z(n20) );
  BUFFD0 U65 ( .I(n22), .Z(n21) );
  BUFFD0 U66 ( .I(n23), .Z(n22) );
  BUFFD0 U67 ( .I(n24), .Z(n23) );
  BUFFD0 U68 ( .I(n25), .Z(n24) );
  BUFFD0 U69 ( .I(n26), .Z(n25) );
  BUFFD0 U70 ( .I(n27), .Z(n26) );
  BUFFD0 U71 ( .I(n28), .Z(n27) );
  BUFFD0 U72 ( .I(n29), .Z(n28) );
  BUFFD0 U73 ( .I(n30), .Z(n29) );
  BUFFD0 U74 ( .I(n31), .Z(n30) );
  BUFFD0 U75 ( .I(n32), .Z(n31) );
  BUFFD0 U76 ( .I(n33), .Z(n32) );
  BUFFD0 U77 ( .I(n34), .Z(n33) );
  BUFFD0 U78 ( .I(n35), .Z(n34) );
  BUFFD0 U79 ( .I(n36), .Z(n35) );
  BUFFD0 U80 ( .I(n37), .Z(n36) );
  BUFFD0 U81 ( .I(n38), .Z(n37) );
  BUFFD0 U82 ( .I(n39), .Z(n38) );
  BUFFD0 U83 ( .I(n40), .Z(n39) );
  BUFFD0 U84 ( .I(n41), .Z(n40) );
  BUFFD0 U85 ( .I(n42), .Z(n41) );
  BUFFD0 U86 ( .I(n43), .Z(n42) );
  BUFFD0 U87 ( .I(n44), .Z(n43) );
  BUFFD0 U88 ( .I(n45), .Z(n44) );
  BUFFD0 U89 ( .I(n46), .Z(n45) );
  BUFFD0 U90 ( .I(n47), .Z(n46) );
  BUFFD0 U91 ( .I(n48), .Z(n47) );
  BUFFD0 U92 ( .I(n49), .Z(n48) );
  BUFFD0 U93 ( .I(n50), .Z(n49) );
  BUFFD0 U94 ( .I(n51), .Z(n50) );
  BUFFD0 U95 ( .I(n52), .Z(n51) );
  BUFFD0 U96 ( .I(n53), .Z(n52) );
  BUFFD0 U97 ( .I(n54), .Z(n53) );
  BUFFD0 U98 ( .I(n55), .Z(n54) );
  BUFFD0 U99 ( .I(n56), .Z(n55) );
  BUFFD0 U100 ( .I(n57), .Z(n56) );
  BUFFD0 U101 ( .I(n58), .Z(n57) );
  BUFFD0 U102 ( .I(n59), .Z(n58) );
  BUFFD0 U103 ( .I(n60), .Z(n59) );
  BUFFD0 U104 ( .I(n61), .Z(n60) );
  BUFFD0 U105 ( .I(n62), .Z(n61) );
  BUFFD0 U106 ( .I(n63), .Z(n62) );
  BUFFD0 U107 ( .I(n64), .Z(n63) );
  BUFFD0 U108 ( .I(n65), .Z(n64) );
  BUFFD0 U109 ( .I(n107), .Z(n65) );
  BUFFD0 U110 ( .I(n109), .Z(n107) );
  BUFFD0 U111 ( .I(n110), .Z(n109) );
  BUFFD0 U112 ( .I(N51), .Z(n110) );
  BUFFD0 U113 ( .I(n8275), .Z(n111) );
  BUFFD0 U114 ( .I(n113), .Z(n112) );
  BUFFD0 U115 ( .I(n114), .Z(n113) );
  BUFFD0 U116 ( .I(n115), .Z(n114) );
  BUFFD0 U117 ( .I(n116), .Z(n115) );
  BUFFD0 U118 ( .I(n117), .Z(n116) );
  BUFFD0 U119 ( .I(n118), .Z(n117) );
  BUFFD0 U120 ( .I(n119), .Z(n118) );
  BUFFD0 U121 ( .I(n120), .Z(n119) );
  BUFFD0 U122 ( .I(n121), .Z(n120) );
  BUFFD0 U123 ( .I(n122), .Z(n121) );
  BUFFD0 U124 ( .I(n123), .Z(n122) );
  BUFFD0 U125 ( .I(n124), .Z(n123) );
  BUFFD0 U126 ( .I(n125), .Z(n124) );
  BUFFD0 U127 ( .I(n126), .Z(n125) );
  BUFFD0 U128 ( .I(n127), .Z(n126) );
  BUFFD0 U129 ( .I(n128), .Z(n127) );
  BUFFD0 U130 ( .I(n129), .Z(n128) );
  BUFFD0 U131 ( .I(n130), .Z(n129) );
  BUFFD0 U132 ( .I(n131), .Z(n130) );
  BUFFD0 U133 ( .I(n132), .Z(n131) );
  BUFFD0 U134 ( .I(n133), .Z(n132) );
  BUFFD0 U135 ( .I(n134), .Z(n133) );
  BUFFD0 U136 ( .I(n135), .Z(n134) );
  BUFFD0 U137 ( .I(n136), .Z(n135) );
  BUFFD0 U138 ( .I(n137), .Z(n136) );
  BUFFD0 U139 ( .I(n138), .Z(n137) );
  BUFFD0 U140 ( .I(n139), .Z(n138) );
  BUFFD0 U141 ( .I(n140), .Z(n139) );
  BUFFD0 U142 ( .I(n141), .Z(n140) );
  BUFFD0 U143 ( .I(n142), .Z(n141) );
  BUFFD0 U144 ( .I(n143), .Z(n142) );
  BUFFD0 U145 ( .I(n144), .Z(n143) );
  BUFFD0 U146 ( .I(n145), .Z(n144) );
  BUFFD0 U147 ( .I(n146), .Z(n145) );
  BUFFD0 U148 ( .I(n147), .Z(n146) );
  BUFFD0 U149 ( .I(n148), .Z(n147) );
  BUFFD0 U150 ( .I(n149), .Z(n148) );
  BUFFD0 U151 ( .I(n150), .Z(n149) );
  BUFFD0 U152 ( .I(n151), .Z(n150) );
  BUFFD0 U153 ( .I(n152), .Z(n151) );
  BUFFD0 U154 ( .I(n153), .Z(n152) );
  BUFFD0 U155 ( .I(n154), .Z(n153) );
  BUFFD0 U156 ( .I(n155), .Z(n154) );
  BUFFD0 U157 ( .I(n156), .Z(n155) );
  BUFFD0 U158 ( .I(n157), .Z(n156) );
  BUFFD0 U159 ( .I(n158), .Z(n157) );
  BUFFD0 U160 ( .I(n159), .Z(n158) );
  BUFFD0 U161 ( .I(n160), .Z(n159) );
  BUFFD0 U162 ( .I(n161), .Z(n160) );
  BUFFD0 U163 ( .I(n162), .Z(n161) );
  BUFFD0 U164 ( .I(n163), .Z(n162) );
  BUFFD0 U165 ( .I(n164), .Z(n163) );
  BUFFD0 U166 ( .I(n165), .Z(n164) );
  BUFFD0 U167 ( .I(n166), .Z(n165) );
  BUFFD0 U168 ( .I(n167), .Z(n166) );
  BUFFD0 U169 ( .I(n168), .Z(n167) );
  BUFFD0 U170 ( .I(n169), .Z(n168) );
  BUFFD0 U171 ( .I(n170), .Z(n169) );
  BUFFD0 U172 ( .I(n171), .Z(n170) );
  BUFFD0 U173 ( .I(n172), .Z(n171) );
  BUFFD0 U174 ( .I(n173), .Z(n172) );
  BUFFD0 U175 ( .I(n174), .Z(n173) );
  BUFFD0 U176 ( .I(n175), .Z(n174) );
  BUFFD0 U177 ( .I(n176), .Z(n175) );
  BUFFD0 U178 ( .I(N52), .Z(n176) );
  BUFFD0 U179 ( .I(n8262), .Z(n177) );
  BUFFD0 U180 ( .I(n179), .Z(n178) );
  BUFFD0 U181 ( .I(n180), .Z(n179) );
  BUFFD0 U182 ( .I(n181), .Z(n180) );
  BUFFD0 U183 ( .I(n182), .Z(n181) );
  BUFFD0 U184 ( .I(n183), .Z(n182) );
  BUFFD0 U185 ( .I(n184), .Z(n183) );
  BUFFD0 U186 ( .I(n185), .Z(n184) );
  BUFFD0 U187 ( .I(n186), .Z(n185) );
  BUFFD0 U188 ( .I(n187), .Z(n186) );
  BUFFD0 U189 ( .I(n188), .Z(n187) );
  BUFFD0 U190 ( .I(n189), .Z(n188) );
  BUFFD0 U191 ( .I(n190), .Z(n189) );
  BUFFD0 U192 ( .I(n191), .Z(n190) );
  BUFFD0 U193 ( .I(n192), .Z(n191) );
  BUFFD0 U194 ( .I(n193), .Z(n192) );
  BUFFD0 U195 ( .I(n194), .Z(n193) );
  BUFFD0 U196 ( .I(n195), .Z(n194) );
  BUFFD0 U197 ( .I(n196), .Z(n195) );
  BUFFD0 U198 ( .I(n197), .Z(n196) );
  BUFFD0 U199 ( .I(n198), .Z(n197) );
  BUFFD0 U200 ( .I(n199), .Z(n198) );
  BUFFD0 U201 ( .I(n200), .Z(n199) );
  BUFFD0 U202 ( .I(n201), .Z(n200) );
  BUFFD0 U203 ( .I(n202), .Z(n201) );
  BUFFD0 U204 ( .I(n203), .Z(n202) );
  BUFFD0 U205 ( .I(n204), .Z(n203) );
  BUFFD0 U206 ( .I(n205), .Z(n204) );
  BUFFD0 U207 ( .I(n206), .Z(n205) );
  BUFFD0 U208 ( .I(n207), .Z(n206) );
  BUFFD0 U209 ( .I(n208), .Z(n207) );
  BUFFD0 U210 ( .I(n209), .Z(n208) );
  BUFFD0 U211 ( .I(n210), .Z(n209) );
  BUFFD0 U212 ( .I(n211), .Z(n210) );
  BUFFD0 U213 ( .I(n212), .Z(n211) );
  BUFFD0 U214 ( .I(n213), .Z(n212) );
  BUFFD0 U215 ( .I(n214), .Z(n213) );
  BUFFD0 U216 ( .I(n215), .Z(n214) );
  BUFFD0 U217 ( .I(n216), .Z(n215) );
  BUFFD0 U218 ( .I(n217), .Z(n216) );
  BUFFD0 U219 ( .I(n218), .Z(n217) );
  BUFFD0 U220 ( .I(n219), .Z(n218) );
  BUFFD0 U221 ( .I(n220), .Z(n219) );
  BUFFD0 U222 ( .I(n221), .Z(n220) );
  BUFFD0 U223 ( .I(n222), .Z(n221) );
  BUFFD0 U224 ( .I(n223), .Z(n222) );
  BUFFD0 U225 ( .I(n224), .Z(n223) );
  BUFFD0 U226 ( .I(n225), .Z(n224) );
  BUFFD0 U227 ( .I(n226), .Z(n225) );
  BUFFD0 U228 ( .I(n227), .Z(n226) );
  BUFFD0 U229 ( .I(n228), .Z(n227) );
  BUFFD0 U230 ( .I(n229), .Z(n228) );
  BUFFD0 U231 ( .I(n230), .Z(n229) );
  BUFFD0 U232 ( .I(n231), .Z(n230) );
  BUFFD0 U233 ( .I(n232), .Z(n231) );
  BUFFD0 U234 ( .I(n233), .Z(n232) );
  BUFFD0 U235 ( .I(n234), .Z(n233) );
  BUFFD0 U236 ( .I(n235), .Z(n234) );
  BUFFD0 U237 ( .I(n236), .Z(n235) );
  BUFFD0 U238 ( .I(n237), .Z(n236) );
  BUFFD0 U239 ( .I(n238), .Z(n237) );
  BUFFD0 U240 ( .I(n239), .Z(n238) );
  BUFFD0 U241 ( .I(n240), .Z(n239) );
  BUFFD0 U242 ( .I(n241), .Z(n240) );
  BUFFD0 U243 ( .I(n242), .Z(n241) );
  BUFFD0 U244 ( .I(N53), .Z(n242) );
  BUFFD0 U245 ( .I(n8249), .Z(n243) );
  BUFFD0 U246 ( .I(n245), .Z(n244) );
  BUFFD0 U247 ( .I(n246), .Z(n245) );
  BUFFD0 U248 ( .I(n247), .Z(n246) );
  BUFFD0 U249 ( .I(n248), .Z(n247) );
  BUFFD0 U250 ( .I(n249), .Z(n248) );
  BUFFD0 U251 ( .I(n250), .Z(n249) );
  BUFFD0 U252 ( .I(n251), .Z(n250) );
  BUFFD0 U253 ( .I(n252), .Z(n251) );
  BUFFD0 U254 ( .I(n253), .Z(n252) );
  BUFFD0 U255 ( .I(n254), .Z(n253) );
  BUFFD0 U256 ( .I(n255), .Z(n254) );
  BUFFD0 U257 ( .I(n256), .Z(n255) );
  BUFFD0 U258 ( .I(n257), .Z(n256) );
  BUFFD0 U259 ( .I(n258), .Z(n257) );
  BUFFD0 U260 ( .I(n259), .Z(n258) );
  BUFFD0 U261 ( .I(n260), .Z(n259) );
  BUFFD0 U262 ( .I(n261), .Z(n260) );
  BUFFD0 U263 ( .I(n262), .Z(n261) );
  BUFFD0 U264 ( .I(n263), .Z(n262) );
  BUFFD0 U265 ( .I(n264), .Z(n263) );
  BUFFD0 U266 ( .I(n265), .Z(n264) );
  BUFFD0 U267 ( .I(n266), .Z(n265) );
  BUFFD0 U268 ( .I(n267), .Z(n266) );
  BUFFD0 U269 ( .I(n268), .Z(n267) );
  BUFFD0 U270 ( .I(n269), .Z(n268) );
  BUFFD0 U271 ( .I(n270), .Z(n269) );
  BUFFD0 U272 ( .I(n271), .Z(n270) );
  BUFFD0 U273 ( .I(n272), .Z(n271) );
  BUFFD0 U274 ( .I(n273), .Z(n272) );
  BUFFD0 U275 ( .I(n274), .Z(n273) );
  BUFFD0 U276 ( .I(n275), .Z(n274) );
  BUFFD0 U277 ( .I(n276), .Z(n275) );
  BUFFD0 U278 ( .I(n277), .Z(n276) );
  BUFFD0 U279 ( .I(n278), .Z(n277) );
  BUFFD0 U280 ( .I(n279), .Z(n278) );
  BUFFD0 U281 ( .I(n280), .Z(n279) );
  BUFFD0 U282 ( .I(n281), .Z(n280) );
  BUFFD0 U283 ( .I(n282), .Z(n281) );
  BUFFD0 U284 ( .I(n283), .Z(n282) );
  BUFFD0 U285 ( .I(n284), .Z(n283) );
  BUFFD0 U286 ( .I(n285), .Z(n284) );
  BUFFD0 U287 ( .I(n286), .Z(n285) );
  BUFFD0 U288 ( .I(n287), .Z(n286) );
  BUFFD0 U289 ( .I(n288), .Z(n287) );
  BUFFD0 U290 ( .I(n289), .Z(n288) );
  BUFFD0 U291 ( .I(n290), .Z(n289) );
  BUFFD0 U292 ( .I(n291), .Z(n290) );
  BUFFD0 U293 ( .I(n292), .Z(n291) );
  BUFFD0 U294 ( .I(n293), .Z(n292) );
  BUFFD0 U295 ( .I(n294), .Z(n293) );
  BUFFD0 U296 ( .I(n295), .Z(n294) );
  BUFFD0 U297 ( .I(n296), .Z(n295) );
  BUFFD0 U298 ( .I(n297), .Z(n296) );
  BUFFD0 U299 ( .I(n298), .Z(n297) );
  BUFFD0 U300 ( .I(n299), .Z(n298) );
  BUFFD0 U301 ( .I(n300), .Z(n299) );
  BUFFD0 U302 ( .I(n301), .Z(n300) );
  BUFFD0 U303 ( .I(n302), .Z(n301) );
  BUFFD0 U304 ( .I(n303), .Z(n302) );
  BUFFD0 U305 ( .I(n304), .Z(n303) );
  BUFFD0 U306 ( .I(n305), .Z(n304) );
  BUFFD0 U307 ( .I(n306), .Z(n305) );
  BUFFD0 U308 ( .I(n307), .Z(n306) );
  BUFFD0 U309 ( .I(n308), .Z(n307) );
  BUFFD0 U310 ( .I(N54), .Z(n308) );
  BUFFD0 U311 ( .I(n8236), .Z(n309) );
  BUFFD0 U312 ( .I(n311), .Z(n310) );
  BUFFD0 U313 ( .I(n312), .Z(n311) );
  BUFFD0 U314 ( .I(n313), .Z(n312) );
  BUFFD0 U315 ( .I(n314), .Z(n313) );
  BUFFD0 U316 ( .I(n315), .Z(n314) );
  BUFFD0 U317 ( .I(n316), .Z(n315) );
  BUFFD0 U318 ( .I(n317), .Z(n316) );
  BUFFD0 U319 ( .I(n318), .Z(n317) );
  BUFFD0 U320 ( .I(n319), .Z(n318) );
  BUFFD0 U321 ( .I(n320), .Z(n319) );
  BUFFD0 U322 ( .I(n321), .Z(n320) );
  BUFFD0 U323 ( .I(n322), .Z(n321) );
  BUFFD0 U324 ( .I(n323), .Z(n322) );
  BUFFD0 U325 ( .I(n324), .Z(n323) );
  BUFFD0 U326 ( .I(n325), .Z(n324) );
  BUFFD0 U327 ( .I(n326), .Z(n325) );
  BUFFD0 U328 ( .I(n327), .Z(n326) );
  BUFFD0 U329 ( .I(n328), .Z(n327) );
  BUFFD0 U330 ( .I(n329), .Z(n328) );
  BUFFD0 U331 ( .I(n330), .Z(n329) );
  BUFFD0 U332 ( .I(n331), .Z(n330) );
  BUFFD0 U333 ( .I(n332), .Z(n331) );
  BUFFD0 U334 ( .I(n333), .Z(n332) );
  BUFFD0 U335 ( .I(n334), .Z(n333) );
  BUFFD0 U336 ( .I(n335), .Z(n334) );
  BUFFD0 U337 ( .I(n336), .Z(n335) );
  BUFFD0 U338 ( .I(n337), .Z(n336) );
  BUFFD0 U339 ( .I(n338), .Z(n337) );
  BUFFD0 U340 ( .I(n339), .Z(n338) );
  BUFFD0 U341 ( .I(n340), .Z(n339) );
  BUFFD0 U342 ( .I(n341), .Z(n340) );
  BUFFD0 U343 ( .I(n342), .Z(n341) );
  BUFFD0 U344 ( .I(n343), .Z(n342) );
  BUFFD0 U345 ( .I(n344), .Z(n343) );
  BUFFD0 U346 ( .I(n345), .Z(n344) );
  BUFFD0 U347 ( .I(n346), .Z(n345) );
  BUFFD0 U348 ( .I(n347), .Z(n346) );
  BUFFD0 U349 ( .I(n348), .Z(n347) );
  BUFFD0 U350 ( .I(n349), .Z(n348) );
  BUFFD0 U351 ( .I(n350), .Z(n349) );
  BUFFD0 U352 ( .I(n351), .Z(n350) );
  BUFFD0 U353 ( .I(n352), .Z(n351) );
  BUFFD0 U354 ( .I(n353), .Z(n352) );
  BUFFD0 U355 ( .I(n354), .Z(n353) );
  BUFFD0 U356 ( .I(n355), .Z(n354) );
  BUFFD0 U357 ( .I(n356), .Z(n355) );
  BUFFD0 U358 ( .I(n357), .Z(n356) );
  BUFFD0 U359 ( .I(n358), .Z(n357) );
  BUFFD0 U360 ( .I(n359), .Z(n358) );
  BUFFD0 U361 ( .I(n360), .Z(n359) );
  BUFFD0 U362 ( .I(n361), .Z(n360) );
  BUFFD0 U363 ( .I(n362), .Z(n361) );
  BUFFD0 U364 ( .I(n363), .Z(n362) );
  BUFFD0 U365 ( .I(n364), .Z(n363) );
  BUFFD0 U366 ( .I(n365), .Z(n364) );
  BUFFD0 U367 ( .I(n366), .Z(n365) );
  BUFFD0 U368 ( .I(n367), .Z(n366) );
  BUFFD0 U369 ( .I(n368), .Z(n367) );
  BUFFD0 U370 ( .I(n369), .Z(n368) );
  BUFFD0 U371 ( .I(n370), .Z(n369) );
  BUFFD0 U372 ( .I(n371), .Z(n370) );
  BUFFD0 U373 ( .I(n372), .Z(n371) );
  BUFFD0 U374 ( .I(n373), .Z(n372) );
  BUFFD0 U375 ( .I(n374), .Z(n373) );
  BUFFD0 U376 ( .I(N55), .Z(n374) );
  BUFFD0 U377 ( .I(n8223), .Z(n375) );
  BUFFD0 U378 ( .I(n377), .Z(n376) );
  BUFFD0 U379 ( .I(n378), .Z(n377) );
  BUFFD0 U380 ( .I(n379), .Z(n378) );
  BUFFD0 U381 ( .I(n380), .Z(n379) );
  BUFFD0 U382 ( .I(n381), .Z(n380) );
  BUFFD0 U383 ( .I(n382), .Z(n381) );
  BUFFD0 U384 ( .I(n383), .Z(n382) );
  BUFFD0 U385 ( .I(n384), .Z(n383) );
  BUFFD0 U386 ( .I(n385), .Z(n384) );
  BUFFD0 U387 ( .I(n386), .Z(n385) );
  BUFFD0 U388 ( .I(n387), .Z(n386) );
  BUFFD0 U389 ( .I(n388), .Z(n387) );
  BUFFD0 U390 ( .I(n389), .Z(n388) );
  BUFFD0 U391 ( .I(n390), .Z(n389) );
  BUFFD0 U392 ( .I(n391), .Z(n390) );
  BUFFD0 U393 ( .I(n392), .Z(n391) );
  BUFFD0 U394 ( .I(n393), .Z(n392) );
  BUFFD0 U395 ( .I(n394), .Z(n393) );
  BUFFD0 U396 ( .I(n395), .Z(n394) );
  BUFFD0 U397 ( .I(n396), .Z(n395) );
  BUFFD0 U398 ( .I(n397), .Z(n396) );
  BUFFD0 U399 ( .I(n398), .Z(n397) );
  BUFFD0 U400 ( .I(n399), .Z(n398) );
  BUFFD0 U401 ( .I(n400), .Z(n399) );
  BUFFD0 U402 ( .I(n401), .Z(n400) );
  BUFFD0 U403 ( .I(n402), .Z(n401) );
  BUFFD0 U404 ( .I(n403), .Z(n402) );
  BUFFD0 U405 ( .I(n404), .Z(n403) );
  BUFFD0 U406 ( .I(n405), .Z(n404) );
  BUFFD0 U407 ( .I(n406), .Z(n405) );
  BUFFD0 U408 ( .I(n407), .Z(n406) );
  BUFFD0 U409 ( .I(n408), .Z(n407) );
  BUFFD0 U410 ( .I(n409), .Z(n408) );
  BUFFD0 U411 ( .I(n410), .Z(n409) );
  BUFFD0 U412 ( .I(n411), .Z(n410) );
  BUFFD0 U413 ( .I(n412), .Z(n411) );
  BUFFD0 U414 ( .I(n413), .Z(n412) );
  BUFFD0 U415 ( .I(n414), .Z(n413) );
  BUFFD0 U416 ( .I(n415), .Z(n414) );
  BUFFD0 U417 ( .I(n416), .Z(n415) );
  BUFFD0 U418 ( .I(n417), .Z(n416) );
  BUFFD0 U419 ( .I(n418), .Z(n417) );
  BUFFD0 U420 ( .I(n419), .Z(n418) );
  BUFFD0 U421 ( .I(n420), .Z(n419) );
  BUFFD0 U422 ( .I(n421), .Z(n420) );
  BUFFD0 U423 ( .I(n422), .Z(n421) );
  BUFFD0 U424 ( .I(n423), .Z(n422) );
  BUFFD0 U425 ( .I(n424), .Z(n423) );
  BUFFD0 U426 ( .I(n425), .Z(n424) );
  BUFFD0 U427 ( .I(n426), .Z(n425) );
  BUFFD0 U428 ( .I(n427), .Z(n426) );
  BUFFD0 U429 ( .I(n428), .Z(n427) );
  BUFFD0 U430 ( .I(n429), .Z(n428) );
  BUFFD0 U431 ( .I(n430), .Z(n429) );
  BUFFD0 U432 ( .I(n431), .Z(n430) );
  BUFFD0 U433 ( .I(n432), .Z(n431) );
  BUFFD0 U434 ( .I(n433), .Z(n432) );
  BUFFD0 U435 ( .I(n434), .Z(n433) );
  BUFFD0 U436 ( .I(n435), .Z(n434) );
  BUFFD0 U437 ( .I(n436), .Z(n435) );
  BUFFD0 U438 ( .I(n437), .Z(n436) );
  BUFFD0 U439 ( .I(n438), .Z(n437) );
  BUFFD0 U440 ( .I(n439), .Z(n438) );
  BUFFD0 U441 ( .I(n440), .Z(n439) );
  BUFFD0 U442 ( .I(N56), .Z(n440) );
  BUFFD0 U443 ( .I(n8210), .Z(n441) );
  BUFFD0 U444 ( .I(n443), .Z(n442) );
  BUFFD0 U445 ( .I(n444), .Z(n443) );
  BUFFD0 U446 ( .I(n445), .Z(n444) );
  BUFFD0 U447 ( .I(n446), .Z(n445) );
  BUFFD0 U448 ( .I(n447), .Z(n446) );
  BUFFD0 U449 ( .I(n448), .Z(n447) );
  BUFFD0 U450 ( .I(n449), .Z(n448) );
  BUFFD0 U451 ( .I(n450), .Z(n449) );
  BUFFD0 U452 ( .I(n451), .Z(n450) );
  BUFFD0 U453 ( .I(n452), .Z(n451) );
  BUFFD0 U454 ( .I(n453), .Z(n452) );
  BUFFD0 U455 ( .I(n454), .Z(n453) );
  BUFFD0 U456 ( .I(n455), .Z(n454) );
  BUFFD0 U457 ( .I(n456), .Z(n455) );
  BUFFD0 U458 ( .I(n457), .Z(n456) );
  BUFFD0 U459 ( .I(n458), .Z(n457) );
  BUFFD0 U460 ( .I(n459), .Z(n458) );
  BUFFD0 U461 ( .I(n460), .Z(n459) );
  BUFFD0 U462 ( .I(n461), .Z(n460) );
  BUFFD0 U463 ( .I(n462), .Z(n461) );
  BUFFD0 U464 ( .I(n463), .Z(n462) );
  BUFFD0 U465 ( .I(n464), .Z(n463) );
  BUFFD0 U466 ( .I(n465), .Z(n464) );
  BUFFD0 U467 ( .I(n466), .Z(n465) );
  BUFFD0 U468 ( .I(n467), .Z(n466) );
  BUFFD0 U469 ( .I(n468), .Z(n467) );
  BUFFD0 U470 ( .I(n469), .Z(n468) );
  BUFFD0 U471 ( .I(n470), .Z(n469) );
  BUFFD0 U472 ( .I(n471), .Z(n470) );
  BUFFD0 U473 ( .I(n472), .Z(n471) );
  BUFFD0 U474 ( .I(n473), .Z(n472) );
  BUFFD0 U475 ( .I(n474), .Z(n473) );
  BUFFD0 U476 ( .I(n475), .Z(n474) );
  BUFFD0 U477 ( .I(n476), .Z(n475) );
  BUFFD0 U478 ( .I(n477), .Z(n476) );
  BUFFD0 U479 ( .I(n478), .Z(n477) );
  BUFFD0 U480 ( .I(n479), .Z(n478) );
  BUFFD0 U481 ( .I(n480), .Z(n479) );
  BUFFD0 U482 ( .I(n481), .Z(n480) );
  BUFFD0 U483 ( .I(n482), .Z(n481) );
  BUFFD0 U484 ( .I(n483), .Z(n482) );
  BUFFD0 U485 ( .I(n484), .Z(n483) );
  BUFFD0 U486 ( .I(n485), .Z(n484) );
  BUFFD0 U487 ( .I(n486), .Z(n485) );
  BUFFD0 U488 ( .I(n487), .Z(n486) );
  BUFFD0 U489 ( .I(n488), .Z(n487) );
  BUFFD0 U490 ( .I(n489), .Z(n488) );
  BUFFD0 U491 ( .I(n490), .Z(n489) );
  BUFFD0 U492 ( .I(n491), .Z(n490) );
  BUFFD0 U493 ( .I(n492), .Z(n491) );
  BUFFD0 U494 ( .I(n493), .Z(n492) );
  BUFFD0 U495 ( .I(n494), .Z(n493) );
  BUFFD0 U496 ( .I(n495), .Z(n494) );
  BUFFD0 U497 ( .I(n496), .Z(n495) );
  BUFFD0 U498 ( .I(n497), .Z(n496) );
  BUFFD0 U499 ( .I(n498), .Z(n497) );
  BUFFD0 U500 ( .I(n499), .Z(n498) );
  BUFFD0 U501 ( .I(n500), .Z(n499) );
  BUFFD0 U502 ( .I(n501), .Z(n500) );
  BUFFD0 U503 ( .I(n502), .Z(n501) );
  BUFFD0 U504 ( .I(n503), .Z(n502) );
  BUFFD0 U505 ( .I(n504), .Z(n503) );
  BUFFD0 U506 ( .I(n505), .Z(n504) );
  BUFFD0 U507 ( .I(n506), .Z(n505) );
  BUFFD0 U508 ( .I(N57), .Z(n506) );
  BUFFD0 U509 ( .I(n8197), .Z(n507) );
  BUFFD0 U510 ( .I(n509), .Z(n508) );
  BUFFD0 U511 ( .I(n510), .Z(n509) );
  BUFFD0 U512 ( .I(n511), .Z(n510) );
  BUFFD0 U513 ( .I(n512), .Z(n511) );
  BUFFD0 U514 ( .I(n513), .Z(n512) );
  BUFFD0 U515 ( .I(n514), .Z(n513) );
  BUFFD0 U516 ( .I(n515), .Z(n514) );
  BUFFD0 U517 ( .I(n516), .Z(n515) );
  BUFFD0 U518 ( .I(n517), .Z(n516) );
  BUFFD0 U519 ( .I(n518), .Z(n517) );
  BUFFD0 U520 ( .I(n519), .Z(n518) );
  BUFFD0 U521 ( .I(n520), .Z(n519) );
  BUFFD0 U522 ( .I(n521), .Z(n520) );
  BUFFD0 U523 ( .I(n522), .Z(n521) );
  BUFFD0 U524 ( .I(n523), .Z(n522) );
  BUFFD0 U525 ( .I(n524), .Z(n523) );
  BUFFD0 U526 ( .I(n525), .Z(n524) );
  BUFFD0 U527 ( .I(n526), .Z(n525) );
  BUFFD0 U528 ( .I(n527), .Z(n526) );
  BUFFD0 U529 ( .I(n528), .Z(n527) );
  BUFFD0 U530 ( .I(n529), .Z(n528) );
  BUFFD0 U531 ( .I(n530), .Z(n529) );
  BUFFD0 U532 ( .I(n531), .Z(n530) );
  BUFFD0 U533 ( .I(n532), .Z(n531) );
  BUFFD0 U534 ( .I(n533), .Z(n532) );
  BUFFD0 U535 ( .I(n534), .Z(n533) );
  BUFFD0 U536 ( .I(n535), .Z(n534) );
  BUFFD0 U537 ( .I(n536), .Z(n535) );
  BUFFD0 U538 ( .I(n537), .Z(n536) );
  BUFFD0 U539 ( .I(n538), .Z(n537) );
  BUFFD0 U540 ( .I(n539), .Z(n538) );
  BUFFD0 U541 ( .I(n540), .Z(n539) );
  BUFFD0 U542 ( .I(n541), .Z(n540) );
  BUFFD0 U543 ( .I(n542), .Z(n541) );
  BUFFD0 U544 ( .I(n543), .Z(n542) );
  BUFFD0 U545 ( .I(n544), .Z(n543) );
  BUFFD0 U546 ( .I(n545), .Z(n544) );
  BUFFD0 U547 ( .I(n546), .Z(n545) );
  BUFFD0 U548 ( .I(n547), .Z(n546) );
  BUFFD0 U549 ( .I(n548), .Z(n547) );
  BUFFD0 U550 ( .I(n549), .Z(n548) );
  BUFFD0 U551 ( .I(n550), .Z(n549) );
  BUFFD0 U552 ( .I(n551), .Z(n550) );
  BUFFD0 U553 ( .I(n552), .Z(n551) );
  BUFFD0 U554 ( .I(n553), .Z(n552) );
  BUFFD0 U555 ( .I(n554), .Z(n553) );
  BUFFD0 U556 ( .I(n555), .Z(n554) );
  BUFFD0 U557 ( .I(n556), .Z(n555) );
  BUFFD0 U558 ( .I(n557), .Z(n556) );
  BUFFD0 U559 ( .I(n558), .Z(n557) );
  BUFFD0 U560 ( .I(n559), .Z(n558) );
  BUFFD0 U561 ( .I(n560), .Z(n559) );
  BUFFD0 U562 ( .I(n561), .Z(n560) );
  BUFFD0 U563 ( .I(n562), .Z(n561) );
  BUFFD0 U564 ( .I(n563), .Z(n562) );
  BUFFD0 U565 ( .I(n564), .Z(n563) );
  BUFFD0 U566 ( .I(n565), .Z(n564) );
  BUFFD0 U567 ( .I(n566), .Z(n565) );
  BUFFD0 U568 ( .I(n567), .Z(n566) );
  BUFFD0 U569 ( .I(n568), .Z(n567) );
  BUFFD0 U570 ( .I(n569), .Z(n568) );
  BUFFD0 U571 ( .I(n570), .Z(n569) );
  BUFFD0 U572 ( .I(n571), .Z(n570) );
  BUFFD0 U573 ( .I(n572), .Z(n571) );
  BUFFD0 U574 ( .I(N58), .Z(n572) );
  BUFFD0 U575 ( .I(n8184), .Z(n573) );
  BUFFD0 U576 ( .I(n575), .Z(n574) );
  BUFFD0 U577 ( .I(n576), .Z(n575) );
  BUFFD0 U578 ( .I(n577), .Z(n576) );
  BUFFD0 U579 ( .I(n578), .Z(n577) );
  BUFFD0 U580 ( .I(n579), .Z(n578) );
  BUFFD0 U581 ( .I(n580), .Z(n579) );
  BUFFD0 U582 ( .I(n581), .Z(n580) );
  BUFFD0 U583 ( .I(n582), .Z(n581) );
  BUFFD0 U584 ( .I(n583), .Z(n582) );
  BUFFD0 U585 ( .I(n584), .Z(n583) );
  BUFFD0 U586 ( .I(n585), .Z(n584) );
  BUFFD0 U587 ( .I(n586), .Z(n585) );
  BUFFD0 U588 ( .I(n587), .Z(n586) );
  BUFFD0 U589 ( .I(n588), .Z(n587) );
  BUFFD0 U590 ( .I(n589), .Z(n588) );
  BUFFD0 U591 ( .I(n590), .Z(n589) );
  BUFFD0 U592 ( .I(n591), .Z(n590) );
  BUFFD0 U593 ( .I(n592), .Z(n591) );
  BUFFD0 U594 ( .I(n593), .Z(n592) );
  BUFFD0 U595 ( .I(n594), .Z(n593) );
  BUFFD0 U596 ( .I(n595), .Z(n594) );
  BUFFD0 U597 ( .I(n596), .Z(n595) );
  BUFFD0 U598 ( .I(n597), .Z(n596) );
  BUFFD0 U599 ( .I(n598), .Z(n597) );
  BUFFD0 U600 ( .I(n599), .Z(n598) );
  BUFFD0 U601 ( .I(n600), .Z(n599) );
  BUFFD0 U602 ( .I(n601), .Z(n600) );
  BUFFD0 U603 ( .I(n602), .Z(n601) );
  BUFFD0 U604 ( .I(n603), .Z(n602) );
  BUFFD0 U605 ( .I(n604), .Z(n603) );
  BUFFD0 U606 ( .I(n605), .Z(n604) );
  BUFFD0 U607 ( .I(n606), .Z(n605) );
  BUFFD0 U608 ( .I(n607), .Z(n606) );
  BUFFD0 U609 ( .I(n608), .Z(n607) );
  BUFFD0 U610 ( .I(n609), .Z(n608) );
  BUFFD0 U611 ( .I(n610), .Z(n609) );
  BUFFD0 U612 ( .I(n611), .Z(n610) );
  BUFFD0 U613 ( .I(n612), .Z(n611) );
  BUFFD0 U614 ( .I(n613), .Z(n612) );
  BUFFD0 U615 ( .I(n614), .Z(n613) );
  BUFFD0 U616 ( .I(n615), .Z(n614) );
  BUFFD0 U617 ( .I(n616), .Z(n615) );
  BUFFD0 U618 ( .I(n617), .Z(n616) );
  BUFFD0 U619 ( .I(n618), .Z(n617) );
  BUFFD0 U620 ( .I(n619), .Z(n618) );
  BUFFD0 U621 ( .I(n620), .Z(n619) );
  BUFFD0 U622 ( .I(n621), .Z(n620) );
  BUFFD0 U623 ( .I(n622), .Z(n621) );
  BUFFD0 U624 ( .I(n623), .Z(n622) );
  BUFFD0 U625 ( .I(n624), .Z(n623) );
  BUFFD0 U626 ( .I(n625), .Z(n624) );
  BUFFD0 U627 ( .I(n626), .Z(n625) );
  BUFFD0 U628 ( .I(n627), .Z(n626) );
  BUFFD0 U629 ( .I(n628), .Z(n627) );
  BUFFD0 U630 ( .I(n629), .Z(n628) );
  BUFFD0 U631 ( .I(n630), .Z(n629) );
  BUFFD0 U632 ( .I(n631), .Z(n630) );
  BUFFD0 U633 ( .I(n632), .Z(n631) );
  BUFFD0 U634 ( .I(n633), .Z(n632) );
  BUFFD0 U635 ( .I(n634), .Z(n633) );
  BUFFD0 U636 ( .I(n635), .Z(n634) );
  BUFFD0 U637 ( .I(n636), .Z(n635) );
  BUFFD0 U638 ( .I(n637), .Z(n636) );
  BUFFD0 U639 ( .I(n638), .Z(n637) );
  BUFFD0 U640 ( .I(N59), .Z(n638) );
  BUFFD0 U641 ( .I(n8171), .Z(n639) );
  BUFFD0 U642 ( .I(n641), .Z(n640) );
  BUFFD0 U643 ( .I(n642), .Z(n641) );
  BUFFD0 U644 ( .I(n643), .Z(n642) );
  BUFFD0 U645 ( .I(n644), .Z(n643) );
  BUFFD0 U646 ( .I(n645), .Z(n644) );
  BUFFD0 U647 ( .I(n646), .Z(n645) );
  BUFFD0 U648 ( .I(n647), .Z(n646) );
  BUFFD0 U649 ( .I(n648), .Z(n647) );
  BUFFD0 U650 ( .I(n649), .Z(n648) );
  BUFFD0 U651 ( .I(n650), .Z(n649) );
  BUFFD0 U652 ( .I(n651), .Z(n650) );
  BUFFD0 U653 ( .I(n652), .Z(n651) );
  BUFFD0 U654 ( .I(n653), .Z(n652) );
  BUFFD0 U655 ( .I(n654), .Z(n653) );
  BUFFD0 U656 ( .I(n655), .Z(n654) );
  BUFFD0 U657 ( .I(n656), .Z(n655) );
  BUFFD0 U658 ( .I(n657), .Z(n656) );
  BUFFD0 U659 ( .I(n658), .Z(n657) );
  BUFFD0 U660 ( .I(n659), .Z(n658) );
  BUFFD0 U661 ( .I(n660), .Z(n659) );
  BUFFD0 U662 ( .I(n661), .Z(n660) );
  BUFFD0 U663 ( .I(n662), .Z(n661) );
  BUFFD0 U664 ( .I(n663), .Z(n662) );
  BUFFD0 U665 ( .I(n664), .Z(n663) );
  BUFFD0 U666 ( .I(n665), .Z(n664) );
  BUFFD0 U667 ( .I(n666), .Z(n665) );
  BUFFD0 U668 ( .I(n667), .Z(n666) );
  BUFFD0 U669 ( .I(n668), .Z(n667) );
  BUFFD0 U670 ( .I(n669), .Z(n668) );
  BUFFD0 U671 ( .I(n670), .Z(n669) );
  BUFFD0 U672 ( .I(n671), .Z(n670) );
  BUFFD0 U673 ( .I(n672), .Z(n671) );
  BUFFD0 U674 ( .I(n673), .Z(n672) );
  BUFFD0 U675 ( .I(n674), .Z(n673) );
  BUFFD0 U676 ( .I(n675), .Z(n674) );
  BUFFD0 U677 ( .I(n676), .Z(n675) );
  BUFFD0 U678 ( .I(n677), .Z(n676) );
  BUFFD0 U679 ( .I(n678), .Z(n677) );
  BUFFD0 U680 ( .I(n679), .Z(n678) );
  BUFFD0 U681 ( .I(n680), .Z(n679) );
  BUFFD0 U682 ( .I(n681), .Z(n680) );
  BUFFD0 U683 ( .I(n682), .Z(n681) );
  BUFFD0 U684 ( .I(n683), .Z(n682) );
  BUFFD0 U685 ( .I(n684), .Z(n683) );
  BUFFD0 U686 ( .I(n685), .Z(n684) );
  BUFFD0 U687 ( .I(n686), .Z(n685) );
  BUFFD0 U688 ( .I(n687), .Z(n686) );
  BUFFD0 U689 ( .I(n688), .Z(n687) );
  BUFFD0 U690 ( .I(n689), .Z(n688) );
  BUFFD0 U691 ( .I(n690), .Z(n689) );
  BUFFD0 U692 ( .I(n691), .Z(n690) );
  BUFFD0 U693 ( .I(n692), .Z(n691) );
  BUFFD0 U694 ( .I(n693), .Z(n692) );
  BUFFD0 U695 ( .I(n694), .Z(n693) );
  BUFFD0 U696 ( .I(n695), .Z(n694) );
  BUFFD0 U697 ( .I(n696), .Z(n695) );
  BUFFD0 U698 ( .I(n697), .Z(n696) );
  BUFFD0 U699 ( .I(n698), .Z(n697) );
  BUFFD0 U700 ( .I(n699), .Z(n698) );
  BUFFD0 U701 ( .I(n700), .Z(n699) );
  BUFFD0 U702 ( .I(n701), .Z(n700) );
  BUFFD0 U703 ( .I(n702), .Z(n701) );
  BUFFD0 U704 ( .I(n703), .Z(n702) );
  BUFFD0 U705 ( .I(n704), .Z(n703) );
  BUFFD0 U706 ( .I(N60), .Z(n704) );
  BUFFD0 U707 ( .I(n8158), .Z(n705) );
  BUFFD0 U708 ( .I(n707), .Z(n706) );
  BUFFD0 U709 ( .I(n708), .Z(n707) );
  BUFFD0 U710 ( .I(n709), .Z(n708) );
  BUFFD0 U711 ( .I(n710), .Z(n709) );
  BUFFD0 U712 ( .I(n711), .Z(n710) );
  BUFFD0 U713 ( .I(n712), .Z(n711) );
  BUFFD0 U714 ( .I(n713), .Z(n712) );
  BUFFD0 U715 ( .I(n714), .Z(n713) );
  BUFFD0 U716 ( .I(n715), .Z(n714) );
  BUFFD0 U717 ( .I(n716), .Z(n715) );
  BUFFD0 U718 ( .I(n717), .Z(n716) );
  BUFFD0 U719 ( .I(n718), .Z(n717) );
  BUFFD0 U720 ( .I(n719), .Z(n718) );
  BUFFD0 U721 ( .I(n720), .Z(n719) );
  BUFFD0 U722 ( .I(n721), .Z(n720) );
  BUFFD0 U723 ( .I(n722), .Z(n721) );
  BUFFD0 U724 ( .I(n723), .Z(n722) );
  BUFFD0 U725 ( .I(n724), .Z(n723) );
  BUFFD0 U726 ( .I(n725), .Z(n724) );
  BUFFD0 U727 ( .I(n726), .Z(n725) );
  BUFFD0 U728 ( .I(n727), .Z(n726) );
  BUFFD0 U729 ( .I(n728), .Z(n727) );
  BUFFD0 U730 ( .I(n729), .Z(n728) );
  BUFFD0 U731 ( .I(n730), .Z(n729) );
  BUFFD0 U732 ( .I(n731), .Z(n730) );
  BUFFD0 U733 ( .I(n732), .Z(n731) );
  BUFFD0 U734 ( .I(n733), .Z(n732) );
  BUFFD0 U735 ( .I(n734), .Z(n733) );
  BUFFD0 U736 ( .I(n735), .Z(n734) );
  BUFFD0 U737 ( .I(n736), .Z(n735) );
  BUFFD0 U738 ( .I(n737), .Z(n736) );
  BUFFD0 U739 ( .I(n738), .Z(n737) );
  BUFFD0 U740 ( .I(n739), .Z(n738) );
  BUFFD0 U741 ( .I(n740), .Z(n739) );
  BUFFD0 U742 ( .I(n741), .Z(n740) );
  BUFFD0 U743 ( .I(n742), .Z(n741) );
  BUFFD0 U744 ( .I(n743), .Z(n742) );
  BUFFD0 U745 ( .I(n744), .Z(n743) );
  BUFFD0 U746 ( .I(n745), .Z(n744) );
  BUFFD0 U747 ( .I(n746), .Z(n745) );
  BUFFD0 U748 ( .I(n747), .Z(n746) );
  BUFFD0 U749 ( .I(n748), .Z(n747) );
  BUFFD0 U750 ( .I(n749), .Z(n748) );
  BUFFD0 U751 ( .I(n750), .Z(n749) );
  BUFFD0 U752 ( .I(n751), .Z(n750) );
  BUFFD0 U753 ( .I(n752), .Z(n751) );
  BUFFD0 U754 ( .I(n753), .Z(n752) );
  BUFFD0 U755 ( .I(n754), .Z(n753) );
  BUFFD0 U756 ( .I(n755), .Z(n754) );
  BUFFD0 U757 ( .I(n756), .Z(n755) );
  BUFFD0 U758 ( .I(n757), .Z(n756) );
  BUFFD0 U759 ( .I(n758), .Z(n757) );
  BUFFD0 U760 ( .I(n759), .Z(n758) );
  BUFFD0 U761 ( .I(n760), .Z(n759) );
  BUFFD0 U762 ( .I(n761), .Z(n760) );
  BUFFD0 U763 ( .I(n762), .Z(n761) );
  BUFFD0 U764 ( .I(n763), .Z(n762) );
  BUFFD0 U765 ( .I(n764), .Z(n763) );
  BUFFD0 U766 ( .I(n765), .Z(n764) );
  BUFFD0 U767 ( .I(n766), .Z(n765) );
  BUFFD0 U768 ( .I(n767), .Z(n766) );
  BUFFD0 U769 ( .I(n768), .Z(n767) );
  BUFFD0 U770 ( .I(n769), .Z(n768) );
  BUFFD0 U771 ( .I(n770), .Z(n769) );
  BUFFD0 U772 ( .I(N61), .Z(n770) );
  BUFFD0 U773 ( .I(n8145), .Z(n771) );
  BUFFD0 U774 ( .I(n773), .Z(n772) );
  BUFFD0 U775 ( .I(n774), .Z(n773) );
  BUFFD0 U776 ( .I(n775), .Z(n774) );
  BUFFD0 U777 ( .I(n776), .Z(n775) );
  BUFFD0 U778 ( .I(n777), .Z(n776) );
  BUFFD0 U779 ( .I(n778), .Z(n777) );
  BUFFD0 U780 ( .I(n779), .Z(n778) );
  BUFFD0 U781 ( .I(n780), .Z(n779) );
  BUFFD0 U782 ( .I(n781), .Z(n780) );
  BUFFD0 U783 ( .I(n782), .Z(n781) );
  BUFFD0 U784 ( .I(n783), .Z(n782) );
  BUFFD0 U785 ( .I(n784), .Z(n783) );
  BUFFD0 U786 ( .I(n785), .Z(n784) );
  BUFFD0 U787 ( .I(n786), .Z(n785) );
  BUFFD0 U788 ( .I(n787), .Z(n786) );
  BUFFD0 U789 ( .I(n788), .Z(n787) );
  BUFFD0 U790 ( .I(n789), .Z(n788) );
  BUFFD0 U791 ( .I(n790), .Z(n789) );
  BUFFD0 U792 ( .I(n791), .Z(n790) );
  BUFFD0 U793 ( .I(n792), .Z(n791) );
  BUFFD0 U794 ( .I(n793), .Z(n792) );
  BUFFD0 U795 ( .I(n794), .Z(n793) );
  BUFFD0 U796 ( .I(n795), .Z(n794) );
  BUFFD0 U797 ( .I(n796), .Z(n795) );
  BUFFD0 U798 ( .I(n797), .Z(n796) );
  BUFFD0 U799 ( .I(n798), .Z(n797) );
  BUFFD0 U800 ( .I(n799), .Z(n798) );
  BUFFD0 U801 ( .I(n800), .Z(n799) );
  BUFFD0 U802 ( .I(n801), .Z(n800) );
  BUFFD0 U803 ( .I(n802), .Z(n801) );
  BUFFD0 U804 ( .I(n803), .Z(n802) );
  BUFFD0 U805 ( .I(n804), .Z(n803) );
  BUFFD0 U806 ( .I(n805), .Z(n804) );
  BUFFD0 U807 ( .I(n806), .Z(n805) );
  BUFFD0 U808 ( .I(n807), .Z(n806) );
  BUFFD0 U809 ( .I(n808), .Z(n807) );
  BUFFD0 U810 ( .I(n809), .Z(n808) );
  BUFFD0 U811 ( .I(n810), .Z(n809) );
  BUFFD0 U812 ( .I(n811), .Z(n810) );
  BUFFD0 U813 ( .I(n812), .Z(n811) );
  BUFFD0 U814 ( .I(n813), .Z(n812) );
  BUFFD0 U815 ( .I(n814), .Z(n813) );
  BUFFD0 U816 ( .I(n815), .Z(n814) );
  BUFFD0 U817 ( .I(n816), .Z(n815) );
  BUFFD0 U818 ( .I(n817), .Z(n816) );
  BUFFD0 U819 ( .I(n818), .Z(n817) );
  BUFFD0 U820 ( .I(n819), .Z(n818) );
  BUFFD0 U821 ( .I(n820), .Z(n819) );
  BUFFD0 U822 ( .I(n821), .Z(n820) );
  BUFFD0 U823 ( .I(n822), .Z(n821) );
  BUFFD0 U824 ( .I(n823), .Z(n822) );
  BUFFD0 U825 ( .I(n824), .Z(n823) );
  BUFFD0 U826 ( .I(n825), .Z(n824) );
  BUFFD0 U827 ( .I(n826), .Z(n825) );
  BUFFD0 U828 ( .I(n827), .Z(n826) );
  BUFFD0 U829 ( .I(n828), .Z(n827) );
  BUFFD0 U830 ( .I(n829), .Z(n828) );
  BUFFD0 U831 ( .I(n830), .Z(n829) );
  BUFFD0 U832 ( .I(n831), .Z(n830) );
  BUFFD0 U833 ( .I(n832), .Z(n831) );
  BUFFD0 U834 ( .I(n833), .Z(n832) );
  BUFFD0 U835 ( .I(n834), .Z(n833) );
  BUFFD0 U836 ( .I(n835), .Z(n834) );
  BUFFD0 U837 ( .I(n836), .Z(n835) );
  BUFFD0 U838 ( .I(N62), .Z(n836) );
  BUFFD0 U839 ( .I(n8132), .Z(n837) );
  BUFFD0 U840 ( .I(n839), .Z(n838) );
  BUFFD0 U841 ( .I(n840), .Z(n839) );
  BUFFD0 U842 ( .I(n841), .Z(n840) );
  BUFFD0 U843 ( .I(n842), .Z(n841) );
  BUFFD0 U844 ( .I(n843), .Z(n842) );
  BUFFD0 U845 ( .I(n844), .Z(n843) );
  BUFFD0 U846 ( .I(n845), .Z(n844) );
  BUFFD0 U847 ( .I(n846), .Z(n845) );
  BUFFD0 U848 ( .I(n847), .Z(n846) );
  BUFFD0 U849 ( .I(n848), .Z(n847) );
  BUFFD0 U850 ( .I(n849), .Z(n848) );
  BUFFD0 U851 ( .I(n850), .Z(n849) );
  BUFFD0 U852 ( .I(n851), .Z(n850) );
  BUFFD0 U853 ( .I(n852), .Z(n851) );
  BUFFD0 U854 ( .I(n853), .Z(n852) );
  BUFFD0 U855 ( .I(n854), .Z(n853) );
  BUFFD0 U856 ( .I(n855), .Z(n854) );
  BUFFD0 U857 ( .I(n856), .Z(n855) );
  BUFFD0 U858 ( .I(n857), .Z(n856) );
  BUFFD0 U859 ( .I(n858), .Z(n857) );
  BUFFD0 U860 ( .I(n859), .Z(n858) );
  BUFFD0 U861 ( .I(n860), .Z(n859) );
  BUFFD0 U862 ( .I(n861), .Z(n860) );
  BUFFD0 U863 ( .I(n862), .Z(n861) );
  BUFFD0 U864 ( .I(n863), .Z(n862) );
  BUFFD0 U865 ( .I(n864), .Z(n863) );
  BUFFD0 U866 ( .I(n865), .Z(n864) );
  BUFFD0 U867 ( .I(n866), .Z(n865) );
  BUFFD0 U868 ( .I(n867), .Z(n866) );
  BUFFD0 U869 ( .I(n868), .Z(n867) );
  BUFFD0 U870 ( .I(n869), .Z(n868) );
  BUFFD0 U871 ( .I(n870), .Z(n869) );
  BUFFD0 U872 ( .I(n871), .Z(n870) );
  BUFFD0 U873 ( .I(n872), .Z(n871) );
  BUFFD0 U874 ( .I(n873), .Z(n872) );
  BUFFD0 U875 ( .I(n874), .Z(n873) );
  BUFFD0 U876 ( .I(n875), .Z(n874) );
  BUFFD0 U877 ( .I(n876), .Z(n875) );
  BUFFD0 U878 ( .I(n877), .Z(n876) );
  BUFFD0 U879 ( .I(n878), .Z(n877) );
  BUFFD0 U880 ( .I(n879), .Z(n878) );
  BUFFD0 U881 ( .I(n880), .Z(n879) );
  BUFFD0 U882 ( .I(n881), .Z(n880) );
  BUFFD0 U883 ( .I(n882), .Z(n881) );
  BUFFD0 U884 ( .I(n883), .Z(n882) );
  BUFFD0 U885 ( .I(n884), .Z(n883) );
  BUFFD0 U886 ( .I(n885), .Z(n884) );
  BUFFD0 U887 ( .I(n886), .Z(n885) );
  BUFFD0 U888 ( .I(n887), .Z(n886) );
  BUFFD0 U889 ( .I(n888), .Z(n887) );
  BUFFD0 U890 ( .I(n889), .Z(n888) );
  BUFFD0 U891 ( .I(n890), .Z(n889) );
  BUFFD0 U892 ( .I(n891), .Z(n890) );
  BUFFD0 U893 ( .I(n892), .Z(n891) );
  BUFFD0 U894 ( .I(n893), .Z(n892) );
  BUFFD0 U895 ( .I(n894), .Z(n893) );
  BUFFD0 U896 ( .I(n895), .Z(n894) );
  BUFFD0 U897 ( .I(n896), .Z(n895) );
  BUFFD0 U898 ( .I(n897), .Z(n896) );
  BUFFD0 U899 ( .I(n898), .Z(n897) );
  BUFFD0 U900 ( .I(n899), .Z(n898) );
  BUFFD0 U901 ( .I(n900), .Z(n899) );
  BUFFD0 U902 ( .I(n901), .Z(n900) );
  BUFFD0 U903 ( .I(n902), .Z(n901) );
  BUFFD0 U904 ( .I(N63), .Z(n902) );
  BUFFD0 U905 ( .I(n8119), .Z(n903) );
  BUFFD0 U906 ( .I(n905), .Z(n904) );
  BUFFD0 U907 ( .I(n906), .Z(n905) );
  BUFFD0 U908 ( .I(n907), .Z(n906) );
  BUFFD0 U909 ( .I(n908), .Z(n907) );
  BUFFD0 U910 ( .I(n909), .Z(n908) );
  BUFFD0 U911 ( .I(n910), .Z(n909) );
  BUFFD0 U912 ( .I(n911), .Z(n910) );
  BUFFD0 U913 ( .I(n912), .Z(n911) );
  BUFFD0 U914 ( .I(n913), .Z(n912) );
  BUFFD0 U915 ( .I(n914), .Z(n913) );
  BUFFD0 U916 ( .I(n915), .Z(n914) );
  BUFFD0 U917 ( .I(n916), .Z(n915) );
  BUFFD0 U918 ( .I(n917), .Z(n916) );
  BUFFD0 U919 ( .I(n918), .Z(n917) );
  BUFFD0 U920 ( .I(n919), .Z(n918) );
  BUFFD0 U921 ( .I(n920), .Z(n919) );
  BUFFD0 U922 ( .I(n921), .Z(n920) );
  BUFFD0 U923 ( .I(n922), .Z(n921) );
  BUFFD0 U924 ( .I(n923), .Z(n922) );
  BUFFD0 U925 ( .I(n924), .Z(n923) );
  BUFFD0 U926 ( .I(n925), .Z(n924) );
  BUFFD0 U927 ( .I(n926), .Z(n925) );
  BUFFD0 U928 ( .I(n927), .Z(n926) );
  BUFFD0 U929 ( .I(n928), .Z(n927) );
  BUFFD0 U930 ( .I(n929), .Z(n928) );
  BUFFD0 U931 ( .I(n930), .Z(n929) );
  BUFFD0 U932 ( .I(n931), .Z(n930) );
  BUFFD0 U933 ( .I(n932), .Z(n931) );
  BUFFD0 U934 ( .I(n933), .Z(n932) );
  BUFFD0 U935 ( .I(n934), .Z(n933) );
  BUFFD0 U936 ( .I(n935), .Z(n934) );
  BUFFD0 U937 ( .I(n936), .Z(n935) );
  BUFFD0 U938 ( .I(n937), .Z(n936) );
  BUFFD0 U939 ( .I(n938), .Z(n937) );
  BUFFD0 U940 ( .I(n939), .Z(n938) );
  BUFFD0 U941 ( .I(n940), .Z(n939) );
  BUFFD0 U942 ( .I(n941), .Z(n940) );
  BUFFD0 U943 ( .I(n942), .Z(n941) );
  BUFFD0 U944 ( .I(n943), .Z(n942) );
  BUFFD0 U945 ( .I(n944), .Z(n943) );
  BUFFD0 U946 ( .I(n945), .Z(n944) );
  BUFFD0 U947 ( .I(n946), .Z(n945) );
  BUFFD0 U948 ( .I(n947), .Z(n946) );
  BUFFD0 U949 ( .I(n948), .Z(n947) );
  BUFFD0 U950 ( .I(n949), .Z(n948) );
  BUFFD0 U951 ( .I(n950), .Z(n949) );
  BUFFD0 U952 ( .I(n951), .Z(n950) );
  BUFFD0 U953 ( .I(n952), .Z(n951) );
  BUFFD0 U954 ( .I(n953), .Z(n952) );
  BUFFD0 U955 ( .I(n954), .Z(n953) );
  BUFFD0 U956 ( .I(n955), .Z(n954) );
  BUFFD0 U957 ( .I(n956), .Z(n955) );
  BUFFD0 U958 ( .I(n957), .Z(n956) );
  BUFFD0 U959 ( .I(n958), .Z(n957) );
  BUFFD0 U960 ( .I(n959), .Z(n958) );
  BUFFD0 U961 ( .I(n960), .Z(n959) );
  BUFFD0 U962 ( .I(n961), .Z(n960) );
  BUFFD0 U963 ( .I(n962), .Z(n961) );
  BUFFD0 U964 ( .I(n963), .Z(n962) );
  BUFFD0 U965 ( .I(n964), .Z(n963) );
  BUFFD0 U966 ( .I(n965), .Z(n964) );
  BUFFD0 U967 ( .I(n966), .Z(n965) );
  BUFFD0 U968 ( .I(n967), .Z(n966) );
  BUFFD0 U969 ( .I(n968), .Z(n967) );
  BUFFD0 U970 ( .I(N64), .Z(n968) );
  BUFFD0 U971 ( .I(n8106), .Z(n969) );
  BUFFD0 U972 ( .I(n971), .Z(n970) );
  BUFFD0 U973 ( .I(n972), .Z(n971) );
  BUFFD0 U974 ( .I(n973), .Z(n972) );
  BUFFD0 U975 ( .I(n974), .Z(n973) );
  BUFFD0 U976 ( .I(n975), .Z(n974) );
  BUFFD0 U977 ( .I(n976), .Z(n975) );
  BUFFD0 U978 ( .I(n977), .Z(n976) );
  BUFFD0 U979 ( .I(n978), .Z(n977) );
  BUFFD0 U980 ( .I(n979), .Z(n978) );
  BUFFD0 U981 ( .I(n980), .Z(n979) );
  BUFFD0 U982 ( .I(n981), .Z(n980) );
  BUFFD0 U983 ( .I(n982), .Z(n981) );
  BUFFD0 U984 ( .I(n983), .Z(n982) );
  BUFFD0 U985 ( .I(n984), .Z(n983) );
  BUFFD0 U986 ( .I(n985), .Z(n984) );
  BUFFD0 U987 ( .I(n986), .Z(n985) );
  BUFFD0 U988 ( .I(n987), .Z(n986) );
  BUFFD0 U989 ( .I(n988), .Z(n987) );
  BUFFD0 U990 ( .I(n989), .Z(n988) );
  BUFFD0 U991 ( .I(n990), .Z(n989) );
  BUFFD0 U992 ( .I(n991), .Z(n990) );
  BUFFD0 U993 ( .I(n992), .Z(n991) );
  BUFFD0 U994 ( .I(n993), .Z(n992) );
  BUFFD0 U995 ( .I(n994), .Z(n993) );
  BUFFD0 U996 ( .I(n995), .Z(n994) );
  BUFFD0 U997 ( .I(n996), .Z(n995) );
  BUFFD0 U998 ( .I(n997), .Z(n996) );
  BUFFD0 U999 ( .I(n998), .Z(n997) );
  BUFFD0 U1000 ( .I(n999), .Z(n998) );
  BUFFD0 U1001 ( .I(n1000), .Z(n999) );
  BUFFD0 U1002 ( .I(n1001), .Z(n1000) );
  BUFFD0 U1003 ( .I(n1002), .Z(n1001) );
  BUFFD0 U1004 ( .I(n1003), .Z(n1002) );
  BUFFD0 U1005 ( .I(n1004), .Z(n1003) );
  BUFFD0 U1006 ( .I(n1005), .Z(n1004) );
  BUFFD0 U1007 ( .I(n1006), .Z(n1005) );
  BUFFD0 U1008 ( .I(n1007), .Z(n1006) );
  BUFFD0 U1009 ( .I(n1008), .Z(n1007) );
  BUFFD0 U1010 ( .I(n1009), .Z(n1008) );
  BUFFD0 U1011 ( .I(n1010), .Z(n1009) );
  BUFFD0 U1012 ( .I(n1011), .Z(n1010) );
  BUFFD0 U1013 ( .I(n1012), .Z(n1011) );
  BUFFD0 U1014 ( .I(n1013), .Z(n1012) );
  BUFFD0 U1015 ( .I(n1014), .Z(n1013) );
  BUFFD0 U1016 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1017 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1018 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1019 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1020 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1021 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1022 ( .I(n1021), .Z(n1020) );
  BUFFD0 U1023 ( .I(n1022), .Z(n1021) );
  BUFFD0 U1024 ( .I(n1023), .Z(n1022) );
  BUFFD0 U1025 ( .I(n1024), .Z(n1023) );
  BUFFD0 U1026 ( .I(n1025), .Z(n1024) );
  BUFFD0 U1027 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1028 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1029 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1030 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1031 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1032 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1033 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1034 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1035 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1036 ( .I(N65), .Z(n1034) );
  BUFFD0 U1037 ( .I(n8093), .Z(n1035) );
  BUFFD0 U1038 ( .I(n1040), .Z(n1036) );
  BUFFD0 U1039 ( .I(n2083), .Z(n1037) );
  BUFFD0 U1040 ( .I(n1037), .Z(n1038) );
  BUFFD0 U1041 ( .I(n1038), .Z(n1039) );
  BUFFD0 U1042 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1043 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1044 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1045 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1046 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1047 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1048 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1049 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1050 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1051 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1052 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1053 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1054 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1055 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1056 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1057 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1058 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1059 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1060 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1061 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1062 ( .I(n1061), .Z(n1060) );
  BUFFD0 U1063 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1064 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1065 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1066 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1067 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1068 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1069 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1070 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1071 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1072 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1073 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1074 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1075 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1076 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1077 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1078 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1079 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1080 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1081 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1082 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1083 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1084 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1085 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1086 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1087 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1088 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1089 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1090 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1091 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1092 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1093 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1094 ( .I(n1093), .Z(n1092) );
  BUFFD0 U1095 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1096 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1097 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1098 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1099 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1100 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1101 ( .I(n1039), .Z(n1099) );
  BUFFD0 U1102 ( .I(n1102), .Z(n1100) );
  BUFFD0 U1103 ( .I(n2090), .Z(n1101) );
  BUFFD0 U1104 ( .I(n1104), .Z(n1102) );
  BUFFD0 U1105 ( .I(n1101), .Z(n1103) );
  BUFFD0 U1106 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1107 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1108 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1109 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1110 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1111 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1112 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1113 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1114 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1115 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1116 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1117 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1118 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1119 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1120 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1121 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1122 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1123 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1124 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1125 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1126 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1127 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1128 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1129 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1130 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1131 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1132 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1133 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1134 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1135 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1136 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1137 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1138 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1139 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1140 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1141 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1142 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1143 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1144 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1145 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1146 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1147 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1148 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1149 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1150 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1151 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1152 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1153 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1154 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1155 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1156 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1157 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1158 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1159 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1160 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1161 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1162 ( .I(n1162), .Z(n1160) );
  BUFFD0 U1163 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1164 ( .I(n1103), .Z(n1163) );
  BUFFD0 U1165 ( .I(n1166), .Z(n1164) );
  BUFFD0 U1166 ( .I(n2087), .Z(n1165) );
  BUFFD0 U1167 ( .I(n1168), .Z(n1166) );
  BUFFD0 U1168 ( .I(n1165), .Z(n1167) );
  BUFFD0 U1169 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1170 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1171 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1172 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1173 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1174 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1175 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1176 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1177 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1178 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1179 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1180 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1181 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1182 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1183 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1184 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1185 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1186 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1187 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1188 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1189 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1190 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1191 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1192 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1193 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1194 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1195 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1196 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1197 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1198 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1199 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1200 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1201 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1202 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1203 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1204 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1205 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1206 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1207 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1208 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1209 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1210 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1211 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1212 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1213 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1214 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1215 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1216 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1217 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1218 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1219 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1220 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1221 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1222 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1223 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1224 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1225 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1226 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1227 ( .I(n1167), .Z(n1226) );
  BUFFD0 U1228 ( .I(n1231), .Z(n1227) );
  BUFFD0 U1229 ( .I(n2095), .Z(n1228) );
  BUFFD0 U1230 ( .I(n1228), .Z(n1229) );
  BUFFD0 U1231 ( .I(n1229), .Z(n1230) );
  BUFFD0 U1232 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1233 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1234 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1235 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1236 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1237 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1238 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1239 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1240 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1241 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1242 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1243 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1244 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1245 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1246 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1247 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1248 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1249 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1250 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1251 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1252 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1253 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1254 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1255 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1256 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1257 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1258 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1259 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1260 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1261 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1262 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1263 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1264 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1265 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1266 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1267 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1268 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1269 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1270 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1271 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1272 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1273 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1274 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1275 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1276 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1277 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1278 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1279 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1280 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1281 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1282 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1283 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1284 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1285 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1286 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1287 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1288 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1289 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1290 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1291 ( .I(n1230), .Z(n1290) );
  BUFFD0 U1292 ( .I(n1295), .Z(n1291) );
  BUFFD0 U1293 ( .I(n2089), .Z(n1292) );
  BUFFD0 U1294 ( .I(n1292), .Z(n1293) );
  BUFFD0 U1295 ( .I(n1293), .Z(n1294) );
  BUFFD0 U1296 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1297 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1298 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1299 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1300 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1301 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1302 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1303 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1304 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1305 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1306 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1307 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1308 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1309 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1310 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1311 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1312 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1313 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1314 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1315 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1316 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1317 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1318 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1319 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1320 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1321 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1322 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1323 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1324 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1325 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1326 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1327 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1328 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1329 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1330 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1331 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1332 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1333 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1334 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1335 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1336 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1337 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1338 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1339 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1340 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1341 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1342 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1343 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1344 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1345 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1346 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1347 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1348 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1349 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1350 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1351 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1352 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1353 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1354 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1355 ( .I(n1294), .Z(n1354) );
  BUFFD0 U1356 ( .I(n1357), .Z(n1355) );
  BUFFD0 U1357 ( .I(n2094), .Z(n1356) );
  BUFFD0 U1358 ( .I(n1359), .Z(n1357) );
  BUFFD0 U1359 ( .I(n1356), .Z(n1358) );
  BUFFD0 U1360 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1361 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1362 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1363 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1364 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1365 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1366 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1367 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1368 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1369 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1370 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1371 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1372 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1373 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1374 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1375 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1376 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1377 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1378 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1379 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1380 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1381 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1382 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1383 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1384 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1385 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1386 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1387 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1388 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1389 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1390 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1391 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1392 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1393 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1394 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1395 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1396 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1397 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1398 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1399 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1400 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1401 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1402 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1403 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1404 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1405 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1406 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1407 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1408 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1409 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1410 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1411 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1412 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1413 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1414 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1415 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1416 ( .I(n1417), .Z(n1415) );
  BUFFD0 U1417 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1418 ( .I(n1358), .Z(n1418) );
  BUFFD0 U1419 ( .I(n1423), .Z(n1419) );
  BUFFD0 U1420 ( .I(n2097), .Z(n1420) );
  BUFFD0 U1421 ( .I(n1420), .Z(n1421) );
  BUFFD0 U1422 ( .I(n1421), .Z(n1422) );
  BUFFD0 U1423 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1424 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1425 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1426 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1427 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1428 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1429 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1430 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1431 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1432 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1433 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1434 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1435 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1436 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1437 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1438 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1439 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1440 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1441 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1442 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1443 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1444 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1445 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1446 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1447 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1448 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1449 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1450 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1451 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1452 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1453 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1454 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1455 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1456 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1457 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1458 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1459 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1460 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1461 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1462 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1463 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1464 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1465 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1466 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1467 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1468 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1469 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1470 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1471 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1472 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1473 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1474 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1475 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1476 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1477 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1478 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1479 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1480 ( .I(n1422), .Z(n1480) );
  BUFFD0 U1481 ( .I(n1485), .Z(n1481) );
  BUFFD0 U1482 ( .I(n2091), .Z(n1482) );
  BUFFD0 U1483 ( .I(n1482), .Z(n1483) );
  BUFFD0 U1484 ( .I(n1483), .Z(n1484) );
  BUFFD0 U1485 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1486 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1487 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1488 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1489 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1490 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1491 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1492 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1493 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1494 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1495 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1496 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1497 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1498 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1499 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1500 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1501 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1502 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1503 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1504 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1505 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1506 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1507 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1508 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1509 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1510 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1511 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1512 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1513 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1514 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1515 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1516 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1517 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1518 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1519 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1520 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1521 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1522 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1523 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1524 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1525 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1526 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1527 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1528 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1529 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1530 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1531 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1532 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1533 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1534 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1535 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1536 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1537 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1538 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1539 ( .I(n1484), .Z(n1539) );
  BUFFD0 U1540 ( .I(n1544), .Z(n1540) );
  BUFFD0 U1541 ( .I(n2093), .Z(n1541) );
  BUFFD0 U1542 ( .I(n1541), .Z(n1542) );
  BUFFD0 U1543 ( .I(n1542), .Z(n1543) );
  BUFFD0 U1544 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1545 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1546 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1547 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1548 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1549 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1550 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1551 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1552 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1553 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1554 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1555 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1556 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1557 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1558 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1559 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1560 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1561 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1562 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1563 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1564 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1565 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1566 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1567 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1568 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1569 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1570 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1571 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1572 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1573 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1574 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1575 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1576 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1577 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1578 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1579 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1580 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1581 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1582 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1583 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1584 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1585 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1586 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1587 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1588 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1589 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1590 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1591 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1592 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1593 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1594 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1595 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1596 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1597 ( .I(n1543), .Z(n1597) );
  BUFFD0 U1598 ( .I(n1602), .Z(n1598) );
  BUFFD0 U1599 ( .I(n2152), .Z(n1599) );
  BUFFD0 U1600 ( .I(n1599), .Z(n1600) );
  BUFFD0 U1601 ( .I(n1600), .Z(n1601) );
  BUFFD0 U1602 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1603 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1604 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1605 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1606 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1607 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1608 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1609 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1610 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1611 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1612 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1613 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1614 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1615 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1616 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1617 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1618 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1619 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1620 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1621 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1622 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1623 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1624 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1625 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1626 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1627 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1628 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1629 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1630 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1631 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1632 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1633 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1634 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1635 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1636 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1637 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1638 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1639 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1640 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1641 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1642 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1643 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1644 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1645 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1646 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1647 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1648 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1649 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1650 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1651 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1652 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1653 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1654 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1655 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1656 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1657 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1658 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1659 ( .I(n1601), .Z(n1659) );
  BUFFD0 U1660 ( .I(n1664), .Z(n1660) );
  BUFFD0 U1661 ( .I(n2098), .Z(n1661) );
  BUFFD0 U1662 ( .I(n1661), .Z(n1662) );
  BUFFD0 U1663 ( .I(n1662), .Z(n1663) );
  BUFFD0 U1664 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1665 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1666 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1667 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1668 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1669 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1670 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1671 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1672 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1673 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1674 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1675 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1676 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1677 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1678 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1679 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1680 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1681 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1682 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1683 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1684 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1685 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1686 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1687 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1688 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1689 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1690 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1691 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1692 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1693 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1694 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1695 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1696 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1697 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1698 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1699 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1700 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1701 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1702 ( .I(n1703), .Z(n1702) );
  BUFFD0 U1703 ( .I(n1704), .Z(n1703) );
  BUFFD0 U1704 ( .I(n1705), .Z(n1704) );
  BUFFD0 U1705 ( .I(n1706), .Z(n1705) );
  BUFFD0 U1706 ( .I(n1707), .Z(n1706) );
  BUFFD0 U1707 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1708 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1709 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1710 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1711 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1712 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1713 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1714 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1715 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1716 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1717 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1718 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1719 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1720 ( .I(n1663), .Z(n1720) );
  BUFFD0 U1721 ( .I(n1725), .Z(n1721) );
  BUFFD0 U1722 ( .I(n2084), .Z(n1722) );
  BUFFD0 U1723 ( .I(n1722), .Z(n1723) );
  BUFFD0 U1724 ( .I(n1723), .Z(n1724) );
  BUFFD0 U1725 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1726 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1727 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1728 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1729 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1730 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1731 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1732 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1733 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1734 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1735 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1736 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1737 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1738 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1739 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1740 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1741 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1742 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1743 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1744 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1745 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1746 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1747 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1748 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1749 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1750 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1751 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1752 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1753 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1754 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1755 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1756 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1757 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1758 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1759 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1760 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1761 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1762 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1763 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1764 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1765 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1766 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1767 ( .I(n1768), .Z(n1767) );
  BUFFD0 U1768 ( .I(n1769), .Z(n1768) );
  BUFFD0 U1769 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1770 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1771 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1772 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1773 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1774 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1775 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1776 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1777 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1778 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1779 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1780 ( .I(n1724), .Z(n1780) );
  BUFFD0 U1781 ( .I(n1784), .Z(n1781) );
  BUFFD0 U1782 ( .I(n2092), .Z(n1782) );
  BUFFD0 U1783 ( .I(n1782), .Z(n1783) );
  BUFFD0 U1784 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1785 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1786 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1787 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1788 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1789 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1790 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1791 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1792 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1793 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1794 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1795 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1796 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1797 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1798 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1799 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1800 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1801 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1802 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1803 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1804 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1805 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1806 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1807 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1808 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1809 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1810 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1811 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1812 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1813 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1814 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1815 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1816 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1817 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1818 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1819 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1820 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1821 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1822 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1823 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1824 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1825 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1826 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1827 ( .I(n1828), .Z(n1827) );
  BUFFD0 U1828 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1829 ( .I(n1830), .Z(n1829) );
  BUFFD0 U1830 ( .I(n1831), .Z(n1830) );
  BUFFD0 U1831 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1832 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1833 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1834 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1835 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1836 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1837 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1838 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1839 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1840 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1841 ( .I(n1783), .Z(n1841) );
  BUFFD0 U1842 ( .I(n1846), .Z(n1842) );
  BUFFD0 U1843 ( .I(n2096), .Z(n1843) );
  BUFFD0 U1844 ( .I(n1843), .Z(n1844) );
  BUFFD0 U1845 ( .I(n1844), .Z(n1845) );
  BUFFD0 U1846 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1847 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1848 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1849 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1850 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1851 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1852 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1853 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1854 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1855 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1856 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1857 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1858 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1859 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1860 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1861 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1862 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1863 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1864 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1865 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1866 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1867 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1868 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1869 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1870 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1871 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1872 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1873 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1874 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1875 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1876 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1877 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1878 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1879 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1880 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1881 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1882 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1883 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1884 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1885 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1886 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1887 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1888 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1889 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1890 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1891 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1892 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1893 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1894 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1895 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1896 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1897 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1898 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1899 ( .I(n1845), .Z(n1899) );
  BUFFD0 U1900 ( .I(n1904), .Z(n1900) );
  BUFFD0 U1901 ( .I(n2086), .Z(n1901) );
  BUFFD0 U1902 ( .I(n1901), .Z(n1902) );
  BUFFD0 U1903 ( .I(n1902), .Z(n1903) );
  BUFFD0 U1904 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1905 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1906 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1907 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1908 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1909 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1910 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1911 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1912 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1913 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1914 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1915 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1916 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1917 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1918 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1919 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1920 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1921 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1922 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1923 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1924 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1925 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1926 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1927 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1928 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1929 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1930 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1931 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1932 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1933 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1934 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1935 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1936 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1937 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1938 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1939 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1940 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1941 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1942 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1943 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1944 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1945 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1946 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1947 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1948 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1949 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1950 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1951 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1952 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1953 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1954 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1955 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1956 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1957 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1958 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1959 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1960 ( .I(n1903), .Z(n1960) );
  BUFFD0 U1961 ( .I(n1965), .Z(n1961) );
  BUFFD0 U1962 ( .I(n2085), .Z(n1962) );
  BUFFD0 U1963 ( .I(n1962), .Z(n1963) );
  BUFFD0 U1964 ( .I(n1963), .Z(n1964) );
  BUFFD0 U1965 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1966 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1967 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1968 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1969 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1970 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1971 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1972 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1973 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1974 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1975 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1976 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1977 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1978 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1979 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1980 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1981 ( .I(n1982), .Z(n1981) );
  BUFFD0 U1982 ( .I(n1983), .Z(n1982) );
  BUFFD0 U1983 ( .I(n1984), .Z(n1983) );
  BUFFD0 U1984 ( .I(n1985), .Z(n1984) );
  BUFFD0 U1985 ( .I(n1986), .Z(n1985) );
  BUFFD0 U1986 ( .I(n1987), .Z(n1986) );
  BUFFD0 U1987 ( .I(n1988), .Z(n1987) );
  BUFFD0 U1988 ( .I(n1989), .Z(n1988) );
  BUFFD0 U1989 ( .I(n1990), .Z(n1989) );
  BUFFD0 U1990 ( .I(n1991), .Z(n1990) );
  BUFFD0 U1991 ( .I(n1992), .Z(n1991) );
  BUFFD0 U1992 ( .I(n1993), .Z(n1992) );
  BUFFD0 U1993 ( .I(n1994), .Z(n1993) );
  BUFFD0 U1994 ( .I(n1995), .Z(n1994) );
  BUFFD0 U1995 ( .I(n1996), .Z(n1995) );
  BUFFD0 U1996 ( .I(n1997), .Z(n1996) );
  BUFFD0 U1997 ( .I(n1998), .Z(n1997) );
  BUFFD0 U1998 ( .I(n1999), .Z(n1998) );
  BUFFD0 U1999 ( .I(n2000), .Z(n1999) );
  BUFFD0 U2000 ( .I(n2001), .Z(n2000) );
  BUFFD0 U2001 ( .I(n2002), .Z(n2001) );
  BUFFD0 U2002 ( .I(n2003), .Z(n2002) );
  BUFFD0 U2003 ( .I(n2004), .Z(n2003) );
  BUFFD0 U2004 ( .I(n2005), .Z(n2004) );
  BUFFD0 U2005 ( .I(n2006), .Z(n2005) );
  BUFFD0 U2006 ( .I(n2007), .Z(n2006) );
  BUFFD0 U2007 ( .I(n2008), .Z(n2007) );
  BUFFD0 U2008 ( .I(n2009), .Z(n2008) );
  BUFFD0 U2009 ( .I(n2010), .Z(n2009) );
  BUFFD0 U2010 ( .I(n2011), .Z(n2010) );
  BUFFD0 U2011 ( .I(n2012), .Z(n2011) );
  BUFFD0 U2012 ( .I(n2013), .Z(n2012) );
  BUFFD0 U2013 ( .I(n2014), .Z(n2013) );
  BUFFD0 U2014 ( .I(n2015), .Z(n2014) );
  BUFFD0 U2015 ( .I(n2016), .Z(n2015) );
  BUFFD0 U2016 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2017 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2018 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2019 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2020 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2021 ( .I(n1964), .Z(n2021) );
  BUFFD0 U2022 ( .I(n2026), .Z(n2022) );
  BUFFD0 U2023 ( .I(n2088), .Z(n2023) );
  BUFFD0 U2024 ( .I(n2023), .Z(n2024) );
  BUFFD0 U2025 ( .I(n2024), .Z(n2025) );
  BUFFD0 U2026 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2027 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2028 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2029 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2030 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2031 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2032 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2033 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2034 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2035 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2036 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2037 ( .I(n2038), .Z(n2037) );
  BUFFD0 U2038 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2039 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2040 ( .I(n2041), .Z(n2040) );
  BUFFD0 U2041 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2042 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2043 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2044 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2045 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2046 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2047 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2048 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2049 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2050 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2051 ( .I(n2052), .Z(n2051) );
  BUFFD0 U2052 ( .I(n2053), .Z(n2052) );
  BUFFD0 U2053 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2054 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2055 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2056 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2057 ( .I(n2058), .Z(n2057) );
  BUFFD0 U2058 ( .I(n2059), .Z(n2058) );
  BUFFD0 U2059 ( .I(n2060), .Z(n2059) );
  BUFFD0 U2060 ( .I(n2061), .Z(n2060) );
  BUFFD0 U2061 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2062 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2063 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2064 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2065 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2066 ( .I(n2067), .Z(n2066) );
  BUFFD0 U2067 ( .I(n2068), .Z(n2067) );
  BUFFD0 U2068 ( .I(n2069), .Z(n2068) );
  BUFFD0 U2069 ( .I(n2070), .Z(n2069) );
  BUFFD0 U2070 ( .I(n2071), .Z(n2070) );
  BUFFD0 U2071 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2072 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2073 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2074 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2075 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2076 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2077 ( .I(n2079), .Z(n2077) );
  BUFFD0 U2078 ( .I(N82), .Z(n2078) );
  BUFFD0 U2079 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2080 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2081 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2082 ( .I(n2025), .Z(n2082) );
  BUFFD0 U2083 ( .I(N66), .Z(n2083) );
  BUFFD0 U2084 ( .I(n2154), .Z(n2084) );
  BUFFD0 U2085 ( .I(n2156), .Z(n2085) );
  BUFFD0 U2086 ( .I(n2157), .Z(n2086) );
  BUFFD0 U2087 ( .I(n2099), .Z(n2087) );
  BUFFD0 U2088 ( .I(n2159), .Z(n2088) );
  BUFFD0 U2089 ( .I(N70), .Z(n2089) );
  BUFFD0 U2090 ( .I(n1161), .Z(n2090) );
  BUFFD0 U2091 ( .I(n2162), .Z(n2091) );
  BUFFD0 U2092 ( .I(n2163), .Z(n2092) );
  BUFFD0 U2093 ( .I(n2164), .Z(n2093) );
  BUFFD0 U2094 ( .I(n1416), .Z(n2094) );
  BUFFD0 U2095 ( .I(N69), .Z(n2095) );
  BUFFD0 U2096 ( .I(n2165), .Z(n2096) );
  BUFFD0 U2097 ( .I(n2167), .Z(n2097) );
  BUFFD0 U2098 ( .I(n2168), .Z(n2098) );
  BUFFD0 U2099 ( .I(N68), .Z(n2099) );
  BUFFD0 U2100 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2101 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2102 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2103 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2104 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2105 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2106 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2107 ( .I(n2108), .Z(n2107) );
  BUFFD0 U2108 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2109 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2110 ( .I(n2111), .Z(n2110) );
  BUFFD0 U2111 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2112 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2113 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2114 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2115 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2116 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2117 ( .I(n2118), .Z(n2117) );
  BUFFD0 U2118 ( .I(n2119), .Z(n2118) );
  BUFFD0 U2119 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2120 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2121 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2122 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2123 ( .I(n2124), .Z(n2123) );
  BUFFD0 U2124 ( .I(n2125), .Z(n2124) );
  BUFFD0 U2125 ( .I(n2126), .Z(n2125) );
  BUFFD0 U2126 ( .I(n2127), .Z(n2126) );
  BUFFD0 U2127 ( .I(n2128), .Z(n2127) );
  BUFFD0 U2128 ( .I(n2129), .Z(n2128) );
  BUFFD0 U2129 ( .I(n2130), .Z(n2129) );
  BUFFD0 U2130 ( .I(n2131), .Z(n2130) );
  BUFFD0 U2131 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2132 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2133 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2134 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2135 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2136 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2137 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2138 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2139 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2140 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2141 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2142 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2143 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2144 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2145 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2146 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2147 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2148 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2149 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2150 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2151 ( .I(n2179), .Z(n2151) );
  BUFFD0 U2152 ( .I(n2169), .Z(n2152) );
  BUFFD0 U2153 ( .I(n8080), .Z(n2153) );
  BUFFD0 U2154 ( .I(n8067), .Z(n2155) );
  BUFFD0 U2155 ( .I(n2172), .Z(n2157) );
  BUFFD0 U2156 ( .I(n8028), .Z(n2158) );
  BUFFD0 U2157 ( .I(n2173), .Z(n2159) );
  BUFFD0 U2158 ( .I(n8015), .Z(n2160) );
  BUFFD0 U2159 ( .I(n8041), .Z(n2161) );
  BUFFD0 U2160 ( .I(n2180), .Z(n2165) );
  BUFFD0 U2161 ( .I(n8054), .Z(n2166) );
  BUFFD0 U2162 ( .I(n2185), .Z(n2168) );
  BUFFD0 U2163 ( .I(n2178), .Z(n2169) );
  BUFFD0 U2164 ( .I(n2187), .Z(n2170) );
  BUFFD0 U2165 ( .I(n2184), .Z(n2171) );
  BUFFD0 U2166 ( .I(n2182), .Z(n2172) );
  BUFFD0 U2167 ( .I(n2186), .Z(n2173) );
  BUFFD0 U2168 ( .I(n2190), .Z(n2174) );
  BUFFD0 U2169 ( .I(n2188), .Z(n2175) );
  BUFFD0 U2170 ( .I(n2192), .Z(n2176) );
  BUFFD0 U2171 ( .I(N72), .Z(n2177) );
  BUFFD0 U2172 ( .I(N75), .Z(n2178) );
  BUFFD0 U2173 ( .I(n2181), .Z(n2179) );
  BUFFD0 U2174 ( .I(n2197), .Z(n2180) );
  BUFFD0 U2175 ( .I(n2183), .Z(n2181) );
  BUFFD0 U2176 ( .I(N80), .Z(n2182) );
  BUFFD0 U2177 ( .I(n2189), .Z(n2183) );
  BUFFD0 U2178 ( .I(N81), .Z(n2184) );
  BUFFD0 U2179 ( .I(n2193), .Z(n2185) );
  BUFFD0 U2180 ( .I(n2078), .Z(n2186) );
  BUFFD0 U2181 ( .I(n2199), .Z(n2187) );
  BUFFD0 U2182 ( .I(N78), .Z(n2188) );
  BUFFD0 U2183 ( .I(N83), .Z(n2189) );
  BUFFD0 U2184 ( .I(n2201), .Z(n2190) );
  BUFFD0 U2185 ( .I(n7963), .Z(n2191) );
  BUFFD0 U2186 ( .I(n2203), .Z(n2192) );
  BUFFD0 U2187 ( .I(N76), .Z(n2193) );
  BUFFD0 U2188 ( .I(n7898), .Z(n2194) );
  BUFFD0 U2189 ( .I(n8002), .Z(n2195) );
  BUFFD0 U2190 ( .I(n7885), .Z(n2196) );
  BUFFD0 U2191 ( .I(n2205), .Z(n2197) );
  BUFFD0 U2192 ( .I(n7872), .Z(n2198) );
  BUFFD0 U2193 ( .I(N77), .Z(n2199) );
  BUFFD0 U2194 ( .I(n7924), .Z(n2200) );
  BUFFD0 U2195 ( .I(n2206), .Z(n2201) );
  BUFFD0 U2196 ( .I(n7950), .Z(n2202) );
  BUFFD0 U2197 ( .I(n2207), .Z(n2203) );
  BUFFD0 U2198 ( .I(n7937), .Z(n2204) );
  BUFFD0 U2199 ( .I(n2208), .Z(n2205) );
  BUFFD0 U2200 ( .I(N73), .Z(n2206) );
  BUFFD0 U2201 ( .I(n2210), .Z(n2207) );
  BUFFD0 U2202 ( .I(n2211), .Z(n2208) );
  BUFFD0 U2203 ( .I(n7989), .Z(n2209) );
  BUFFD0 U2204 ( .I(N74), .Z(n2210) );
  BUFFD0 U2205 ( .I(N79), .Z(n2211) );
  BUFFD0 U2206 ( .I(n7976), .Z(n2212) );
  BUFFD0 U2207 ( .I(n7911), .Z(n2213) );
  CKBD0 U2208 ( .CLK(n8693), .C(n6933) );
  XOR3D0 U2209 ( .A1(n8692), .A2(n8689), .A3(n73), .Z(N85) );
  BUFFD0 U2210 ( .I(n8730), .Z(n2215) );
  BUFFD0 U2211 ( .I(n8714), .Z(n2216) );
  BUFFD0 U2212 ( .I(n8698), .Z(n2217) );
  BUFFD0 U2213 ( .I(n8691), .Z(n2218) );
  BUFFD0 U2214 ( .I(n8760), .Z(n2220) );
  BUFFD0 U2215 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2216 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2217 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2218 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2219 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2220 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2221 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2222 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2223 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2224 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2225 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2226 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2227 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2228 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2229 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2230 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2231 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2232 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2233 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2234 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2235 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2236 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2237 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2238 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2239 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2240 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2241 ( .I(n2248), .Z(n2247) );
  BUFFD0 U2242 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2243 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2244 ( .I(n2251), .Z(n2250) );
  BUFFD0 U2245 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2246 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2247 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2248 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2249 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2250 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2251 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2252 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2253 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2254 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2255 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2256 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2257 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2258 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2259 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2260 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2261 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2262 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2263 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2264 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2265 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2266 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2267 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2268 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2269 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2270 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2271 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2272 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2273 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2274 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2275 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2276 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2277 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2278 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2279 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2280 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2281 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2282 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2283 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2284 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2285 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2286 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2287 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2288 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2289 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2290 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2291 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2292 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2293 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2294 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2295 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2296 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2297 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2298 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2299 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2300 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2301 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2302 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2303 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2304 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2305 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2306 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2307 ( .I(n8761), .Z(n2313) );
  BUFFD0 U2308 ( .I(n8757), .Z(n2314) );
  BUFFD0 U2309 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2310 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2311 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2312 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2313 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2314 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2315 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2316 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2317 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2318 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2319 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2320 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2321 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2322 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2323 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2324 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2325 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2326 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2327 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2328 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2329 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2330 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2331 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2332 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2333 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2334 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2335 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2336 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2337 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2338 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2339 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2340 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2341 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2342 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2343 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2344 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2345 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2346 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2347 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2348 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2349 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2350 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2351 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2352 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2353 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2354 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2355 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2356 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2357 ( .I(n2364), .Z(n2363) );
  BUFFD0 U2358 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2359 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2360 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2361 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2362 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2363 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2364 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2365 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2366 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2367 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2368 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2369 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2370 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2371 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2372 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2373 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2374 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2375 ( .I(n2382), .Z(n2381) );
  BUFFD0 U2376 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2377 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2378 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2379 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2380 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2381 ( .I(n2388), .Z(n2387) );
  BUFFD0 U2382 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2383 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2384 ( .I(n2391), .Z(n2390) );
  BUFFD0 U2385 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2386 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2387 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2388 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2389 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2390 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2391 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2392 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2393 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2394 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2395 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2396 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2397 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2398 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2399 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2400 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2401 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2402 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2403 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2404 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2405 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2406 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2407 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2408 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2409 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2410 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2411 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2412 ( .I(n2419), .Z(n2418) );
  BUFFD0 U2413 ( .I(n2420), .Z(n2419) );
  BUFFD0 U2414 ( .I(n2421), .Z(n2420) );
  BUFFD0 U2415 ( .I(n2422), .Z(n2421) );
  BUFFD0 U2416 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2417 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2418 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2419 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2420 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2421 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2422 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2423 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2424 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2425 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2426 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2427 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2428 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2429 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2430 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2431 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2432 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2433 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2434 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2435 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2436 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2437 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2438 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2439 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2440 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2441 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2442 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2443 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2444 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2445 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2446 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2447 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2448 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2449 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2450 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2451 ( .I(n2458), .Z(n2457) );
  BUFFD0 U2452 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2453 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2454 ( .I(n2461), .Z(n2460) );
  BUFFD0 U2455 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2456 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2457 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2458 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2459 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2460 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2461 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2462 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2463 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2464 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2465 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2466 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2467 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2468 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2469 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2470 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2471 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2472 ( .I(n2479), .Z(n2478) );
  BUFFD0 U2473 ( .I(n2480), .Z(n2479) );
  BUFFD0 U2474 ( .I(n2481), .Z(n2480) );
  BUFFD0 U2475 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2476 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2477 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2478 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2479 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2480 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2481 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2482 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2483 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2484 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2485 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2486 ( .I(n8758), .Z(n2492) );
  BUFFD0 U2487 ( .I(n8755), .Z(n2493) );
  BUFFD0 U2488 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2489 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2490 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2491 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2492 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2493 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2494 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2495 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2496 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2497 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2498 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2499 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2500 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2501 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2502 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2503 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2504 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2505 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2506 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2507 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2508 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2509 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2510 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2511 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2512 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2513 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2514 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2515 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2516 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2517 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2518 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2519 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2520 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2521 ( .I(n2528), .Z(n2527) );
  BUFFD0 U2522 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2523 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2524 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2525 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2526 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2527 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2528 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2529 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2530 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2531 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2532 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2533 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2534 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2535 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2536 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2537 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2538 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2539 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2540 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2541 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2542 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2543 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2544 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2545 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2546 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2547 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2548 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2549 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2550 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2551 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2552 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2553 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2554 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2555 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2556 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2557 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2558 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2559 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2560 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2561 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2562 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2563 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2564 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2565 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2566 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2567 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2568 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2569 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2570 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2571 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2572 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2573 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2574 ( .I(n2581), .Z(n2580) );
  BUFFD0 U2575 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2576 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2577 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2578 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2579 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2580 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2581 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2582 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2583 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2584 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2585 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2586 ( .I(n2593), .Z(n2592) );
  BUFFD0 U2587 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2588 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2589 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2590 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2591 ( .I(n2598), .Z(n2597) );
  BUFFD0 U2592 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2593 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2594 ( .I(n2601), .Z(n2600) );
  BUFFD0 U2595 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2596 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2597 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2598 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2599 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2600 ( .I(n2607), .Z(n2606) );
  BUFFD0 U2601 ( .I(n2608), .Z(n2607) );
  BUFFD0 U2602 ( .I(n2609), .Z(n2608) );
  BUFFD0 U2603 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2604 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2605 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2606 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2607 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2608 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2609 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2610 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2611 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2612 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2613 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2614 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2615 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2616 ( .I(n2623), .Z(n2622) );
  BUFFD0 U2617 ( .I(n2624), .Z(n2623) );
  BUFFD0 U2618 ( .I(n2625), .Z(n2624) );
  BUFFD0 U2619 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2620 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2621 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2622 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2623 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2624 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2625 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2626 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2627 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2628 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2629 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2630 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2631 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2632 ( .I(n2639), .Z(n2638) );
  BUFFD0 U2633 ( .I(n2640), .Z(n2639) );
  BUFFD0 U2634 ( .I(n2641), .Z(n2640) );
  BUFFD0 U2635 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2636 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2637 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2638 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2639 ( .I(n2646), .Z(n2645) );
  BUFFD0 U2640 ( .I(n2647), .Z(n2646) );
  BUFFD0 U2641 ( .I(n2648), .Z(n2647) );
  BUFFD0 U2642 ( .I(n2649), .Z(n2648) );
  BUFFD0 U2643 ( .I(n2650), .Z(n2649) );
  BUFFD0 U2644 ( .I(n2651), .Z(n2650) );
  BUFFD0 U2645 ( .I(n2652), .Z(n2651) );
  BUFFD0 U2646 ( .I(n2653), .Z(n2652) );
  BUFFD0 U2647 ( .I(n2654), .Z(n2653) );
  BUFFD0 U2648 ( .I(n2655), .Z(n2654) );
  BUFFD0 U2649 ( .I(n2656), .Z(n2655) );
  BUFFD0 U2650 ( .I(n2657), .Z(n2656) );
  BUFFD0 U2651 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2652 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2653 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2654 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2655 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2656 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2657 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2658 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2659 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2660 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2661 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2662 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2663 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2664 ( .I(n2671), .Z(n2670) );
  BUFFD0 U2665 ( .I(n8756), .Z(n2671) );
  BUFFD0 U2666 ( .I(n8753), .Z(n2672) );
  BUFFD0 U2667 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2668 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2669 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2670 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2671 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2672 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2673 ( .I(n2680), .Z(n2679) );
  BUFFD0 U2674 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2675 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2676 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2677 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2678 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2679 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2680 ( .I(n2687), .Z(n2686) );
  BUFFD0 U2681 ( .I(n2688), .Z(n2687) );
  BUFFD0 U2682 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2683 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2684 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2685 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2686 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2687 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2688 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2689 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2690 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2691 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2692 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2693 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2694 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2695 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2696 ( .I(n2703), .Z(n2702) );
  BUFFD0 U2697 ( .I(n2704), .Z(n2703) );
  BUFFD0 U2698 ( .I(n2705), .Z(n2704) );
  BUFFD0 U2699 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2700 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2701 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2702 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2703 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2704 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2705 ( .I(n2712), .Z(n2711) );
  BUFFD0 U2706 ( .I(n2713), .Z(n2712) );
  BUFFD0 U2707 ( .I(n2714), .Z(n2713) );
  BUFFD0 U2708 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2709 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2710 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2711 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2712 ( .I(n2719), .Z(n2718) );
  BUFFD0 U2713 ( .I(n2720), .Z(n2719) );
  BUFFD0 U2714 ( .I(n2721), .Z(n2720) );
  BUFFD0 U2715 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2716 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2717 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2718 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2719 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2720 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2721 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2722 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2723 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2724 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2725 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2726 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2727 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2728 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2729 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2730 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2731 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2732 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2733 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2734 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2735 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2736 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2737 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2738 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2739 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2740 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2741 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2742 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2743 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2744 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2745 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2746 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2747 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2748 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2749 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2750 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2751 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2752 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2753 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2754 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2755 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2756 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2757 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2758 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2759 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2760 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2761 ( .I(n2768), .Z(n2767) );
  BUFFD0 U2762 ( .I(n2769), .Z(n2768) );
  BUFFD0 U2763 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2764 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2765 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2766 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2767 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2768 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2769 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2770 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2771 ( .I(n2778), .Z(n2777) );
  BUFFD0 U2772 ( .I(n2779), .Z(n2778) );
  BUFFD0 U2773 ( .I(n2780), .Z(n2779) );
  BUFFD0 U2774 ( .I(n2781), .Z(n2780) );
  BUFFD0 U2775 ( .I(n2782), .Z(n2781) );
  BUFFD0 U2776 ( .I(n2783), .Z(n2782) );
  BUFFD0 U2777 ( .I(n2784), .Z(n2783) );
  BUFFD0 U2778 ( .I(n2785), .Z(n2784) );
  BUFFD0 U2779 ( .I(n2786), .Z(n2785) );
  BUFFD0 U2780 ( .I(n2787), .Z(n2786) );
  BUFFD0 U2781 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2782 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2783 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2784 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2785 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2786 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2787 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2788 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2789 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2790 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2791 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2792 ( .I(n2799), .Z(n2798) );
  BUFFD0 U2793 ( .I(n2800), .Z(n2799) );
  BUFFD0 U2794 ( .I(n2801), .Z(n2800) );
  BUFFD0 U2795 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2796 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2797 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2798 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2799 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2800 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2801 ( .I(n2808), .Z(n2807) );
  BUFFD0 U2802 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2803 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2804 ( .I(n2811), .Z(n2810) );
  BUFFD0 U2805 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2806 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2807 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2808 ( .I(n2815), .Z(n2814) );
  BUFFD0 U2809 ( .I(n2816), .Z(n2815) );
  BUFFD0 U2810 ( .I(n2817), .Z(n2816) );
  BUFFD0 U2811 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2812 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2813 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2814 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2815 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2816 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2817 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2818 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2819 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2820 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2821 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2822 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2823 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2824 ( .I(n2831), .Z(n2830) );
  BUFFD0 U2825 ( .I(n2832), .Z(n2831) );
  BUFFD0 U2826 ( .I(n2833), .Z(n2832) );
  BUFFD0 U2827 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2828 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2829 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2830 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2831 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2832 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2833 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2834 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2835 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2836 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2837 ( .I(n2844), .Z(n2843) );
  BUFFD0 U2838 ( .I(n2845), .Z(n2844) );
  BUFFD0 U2839 ( .I(n2846), .Z(n2845) );
  BUFFD0 U2840 ( .I(n2847), .Z(n2846) );
  BUFFD0 U2841 ( .I(n2848), .Z(n2847) );
  BUFFD0 U2842 ( .I(n8754), .Z(n2848) );
  BUFFD0 U2843 ( .I(n8743), .Z(n2849) );
  BUFFD0 U2844 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2845 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2846 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2847 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2848 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2849 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2850 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2851 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2852 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2853 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2854 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2855 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2856 ( .I(n2863), .Z(n2862) );
  BUFFD0 U2857 ( .I(n2864), .Z(n2863) );
  BUFFD0 U2858 ( .I(n2865), .Z(n2864) );
  BUFFD0 U2859 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2860 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2861 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2862 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2863 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2864 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2865 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2866 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2867 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2868 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2869 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2870 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2871 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2872 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2873 ( .I(n2880), .Z(n2879) );
  BUFFD0 U2874 ( .I(n2881), .Z(n2880) );
  BUFFD0 U2875 ( .I(n2882), .Z(n2881) );
  BUFFD0 U2876 ( .I(n2883), .Z(n2882) );
  BUFFD0 U2877 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2878 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2879 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2880 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2881 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2882 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2883 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2884 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2885 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2886 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2887 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2888 ( .I(n2895), .Z(n2894) );
  BUFFD0 U2889 ( .I(n2896), .Z(n2895) );
  BUFFD0 U2890 ( .I(n2897), .Z(n2896) );
  BUFFD0 U2891 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2892 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2893 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2894 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2895 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2896 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2897 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2898 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2899 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2900 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2901 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2902 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2903 ( .I(n2910), .Z(n2909) );
  BUFFD0 U2904 ( .I(n2911), .Z(n2910) );
  BUFFD0 U2905 ( .I(n2912), .Z(n2911) );
  BUFFD0 U2906 ( .I(n2913), .Z(n2912) );
  BUFFD0 U2907 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2908 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2909 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2910 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2911 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2912 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2913 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2914 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2915 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2916 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2917 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2918 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2919 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2920 ( .I(n2927), .Z(n2926) );
  BUFFD0 U2921 ( .I(n2928), .Z(n2927) );
  BUFFD0 U2922 ( .I(n2929), .Z(n2928) );
  BUFFD0 U2923 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2924 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2925 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2926 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2927 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2928 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2929 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2930 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2931 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2932 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2933 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2934 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2935 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2936 ( .I(n2943), .Z(n2942) );
  BUFFD0 U2937 ( .I(n2944), .Z(n2943) );
  BUFFD0 U2938 ( .I(n2945), .Z(n2944) );
  BUFFD0 U2939 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2940 ( .I(n2947), .Z(n2946) );
  BUFFD0 U2941 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2942 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2943 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2944 ( .I(n2951), .Z(n2950) );
  BUFFD0 U2945 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2946 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2947 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2948 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2949 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2950 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2951 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2952 ( .I(n2959), .Z(n2958) );
  BUFFD0 U2953 ( .I(n2960), .Z(n2959) );
  BUFFD0 U2954 ( .I(n2961), .Z(n2960) );
  BUFFD0 U2955 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2956 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2957 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2958 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2959 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2960 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2961 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2962 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2963 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2964 ( .I(n2971), .Z(n2970) );
  BUFFD0 U2965 ( .I(n2972), .Z(n2971) );
  BUFFD0 U2966 ( .I(n2973), .Z(n2972) );
  BUFFD0 U2967 ( .I(n2974), .Z(n2973) );
  BUFFD0 U2968 ( .I(n2975), .Z(n2974) );
  BUFFD0 U2969 ( .I(n2976), .Z(n2975) );
  BUFFD0 U2970 ( .I(n2977), .Z(n2976) );
  BUFFD0 U2971 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2972 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2973 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2974 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2975 ( .I(n2982), .Z(n2981) );
  BUFFD0 U2976 ( .I(n2983), .Z(n2982) );
  BUFFD0 U2977 ( .I(n2984), .Z(n2983) );
  BUFFD0 U2978 ( .I(n2985), .Z(n2984) );
  BUFFD0 U2979 ( .I(n2986), .Z(n2985) );
  BUFFD0 U2980 ( .I(n2987), .Z(n2986) );
  BUFFD0 U2981 ( .I(n2988), .Z(n2987) );
  BUFFD0 U2982 ( .I(n2989), .Z(n2988) );
  BUFFD0 U2983 ( .I(n2990), .Z(n2989) );
  BUFFD0 U2984 ( .I(n2991), .Z(n2990) );
  BUFFD0 U2985 ( .I(n2992), .Z(n2991) );
  BUFFD0 U2986 ( .I(n2993), .Z(n2992) );
  BUFFD0 U2987 ( .I(n2994), .Z(n2993) );
  BUFFD0 U2988 ( .I(n2995), .Z(n2994) );
  BUFFD0 U2989 ( .I(n2996), .Z(n2995) );
  BUFFD0 U2990 ( .I(n2997), .Z(n2996) );
  BUFFD0 U2991 ( .I(n2998), .Z(n2997) );
  BUFFD0 U2992 ( .I(n2999), .Z(n2998) );
  BUFFD0 U2993 ( .I(n3000), .Z(n2999) );
  BUFFD0 U2994 ( .I(n3001), .Z(n3000) );
  BUFFD0 U2995 ( .I(n3002), .Z(n3001) );
  BUFFD0 U2996 ( .I(n3003), .Z(n3002) );
  BUFFD0 U2997 ( .I(n3004), .Z(n3003) );
  BUFFD0 U2998 ( .I(n3005), .Z(n3004) );
  BUFFD0 U2999 ( .I(n3006), .Z(n3005) );
  BUFFD0 U3000 ( .I(n3007), .Z(n3006) );
  BUFFD0 U3001 ( .I(n3008), .Z(n3007) );
  BUFFD0 U3002 ( .I(n3009), .Z(n3008) );
  BUFFD0 U3003 ( .I(n3010), .Z(n3009) );
  BUFFD0 U3004 ( .I(n3011), .Z(n3010) );
  BUFFD0 U3005 ( .I(n3012), .Z(n3011) );
  BUFFD0 U3006 ( .I(n3013), .Z(n3012) );
  BUFFD0 U3007 ( .I(n3014), .Z(n3013) );
  BUFFD0 U3008 ( .I(n3015), .Z(n3014) );
  BUFFD0 U3009 ( .I(n3016), .Z(n3015) );
  BUFFD0 U3010 ( .I(n3017), .Z(n3016) );
  BUFFD0 U3011 ( .I(n3018), .Z(n3017) );
  BUFFD0 U3012 ( .I(n3019), .Z(n3018) );
  BUFFD0 U3013 ( .I(n3020), .Z(n3019) );
  BUFFD0 U3014 ( .I(n3021), .Z(n3020) );
  BUFFD0 U3015 ( .I(n3022), .Z(n3021) );
  BUFFD0 U3016 ( .I(n3023), .Z(n3022) );
  BUFFD0 U3017 ( .I(n3024), .Z(n3023) );
  BUFFD0 U3018 ( .I(n3025), .Z(n3024) );
  BUFFD0 U3019 ( .I(n8744), .Z(n3025) );
  BUFFD0 U3020 ( .I(n8740), .Z(n3026) );
  BUFFD0 U3021 ( .I(n3028), .Z(n3027) );
  BUFFD0 U3022 ( .I(n3029), .Z(n3028) );
  BUFFD0 U3023 ( .I(n3030), .Z(n3029) );
  BUFFD0 U3024 ( .I(n3031), .Z(n3030) );
  BUFFD0 U3025 ( .I(n3032), .Z(n3031) );
  BUFFD0 U3026 ( .I(n3033), .Z(n3032) );
  BUFFD0 U3027 ( .I(n3034), .Z(n3033) );
  BUFFD0 U3028 ( .I(n3035), .Z(n3034) );
  BUFFD0 U3029 ( .I(n3036), .Z(n3035) );
  BUFFD0 U3030 ( .I(n3037), .Z(n3036) );
  BUFFD0 U3031 ( .I(n3038), .Z(n3037) );
  BUFFD0 U3032 ( .I(n3039), .Z(n3038) );
  BUFFD0 U3033 ( .I(n3040), .Z(n3039) );
  BUFFD0 U3034 ( .I(n3041), .Z(n3040) );
  BUFFD0 U3035 ( .I(n3042), .Z(n3041) );
  BUFFD0 U3036 ( .I(n3043), .Z(n3042) );
  BUFFD0 U3037 ( .I(n3044), .Z(n3043) );
  BUFFD0 U3038 ( .I(n3045), .Z(n3044) );
  BUFFD0 U3039 ( .I(n3046), .Z(n3045) );
  BUFFD0 U3040 ( .I(n3047), .Z(n3046) );
  BUFFD0 U3041 ( .I(n3048), .Z(n3047) );
  BUFFD0 U3042 ( .I(n3049), .Z(n3048) );
  BUFFD0 U3043 ( .I(n3050), .Z(n3049) );
  BUFFD0 U3044 ( .I(n3051), .Z(n3050) );
  BUFFD0 U3045 ( .I(n3052), .Z(n3051) );
  BUFFD0 U3046 ( .I(n3053), .Z(n3052) );
  BUFFD0 U3047 ( .I(n3054), .Z(n3053) );
  BUFFD0 U3048 ( .I(n3055), .Z(n3054) );
  BUFFD0 U3049 ( .I(n3056), .Z(n3055) );
  BUFFD0 U3050 ( .I(n3057), .Z(n3056) );
  BUFFD0 U3051 ( .I(n3058), .Z(n3057) );
  BUFFD0 U3052 ( .I(n3059), .Z(n3058) );
  BUFFD0 U3053 ( .I(n3060), .Z(n3059) );
  BUFFD0 U3054 ( .I(n3061), .Z(n3060) );
  BUFFD0 U3055 ( .I(n3062), .Z(n3061) );
  BUFFD0 U3056 ( .I(n3063), .Z(n3062) );
  BUFFD0 U3057 ( .I(n3064), .Z(n3063) );
  BUFFD0 U3058 ( .I(n3065), .Z(n3064) );
  BUFFD0 U3059 ( .I(n3066), .Z(n3065) );
  BUFFD0 U3060 ( .I(n3067), .Z(n3066) );
  BUFFD0 U3061 ( .I(n3068), .Z(n3067) );
  BUFFD0 U3062 ( .I(n3069), .Z(n3068) );
  BUFFD0 U3063 ( .I(n3070), .Z(n3069) );
  BUFFD0 U3064 ( .I(n3071), .Z(n3070) );
  BUFFD0 U3065 ( .I(n3072), .Z(n3071) );
  BUFFD0 U3066 ( .I(n3073), .Z(n3072) );
  BUFFD0 U3067 ( .I(n3074), .Z(n3073) );
  BUFFD0 U3068 ( .I(n3075), .Z(n3074) );
  BUFFD0 U3069 ( .I(n3076), .Z(n3075) );
  BUFFD0 U3070 ( .I(n3077), .Z(n3076) );
  BUFFD0 U3071 ( .I(n3078), .Z(n3077) );
  BUFFD0 U3072 ( .I(n3079), .Z(n3078) );
  BUFFD0 U3073 ( .I(n3080), .Z(n3079) );
  BUFFD0 U3074 ( .I(n3081), .Z(n3080) );
  BUFFD0 U3075 ( .I(n3082), .Z(n3081) );
  BUFFD0 U3076 ( .I(n3083), .Z(n3082) );
  BUFFD0 U3077 ( .I(n3084), .Z(n3083) );
  BUFFD0 U3078 ( .I(n3085), .Z(n3084) );
  BUFFD0 U3079 ( .I(n3086), .Z(n3085) );
  BUFFD0 U3080 ( .I(n3087), .Z(n3086) );
  BUFFD0 U3081 ( .I(n3088), .Z(n3087) );
  BUFFD0 U3082 ( .I(n3089), .Z(n3088) );
  BUFFD0 U3083 ( .I(n3090), .Z(n3089) );
  BUFFD0 U3084 ( .I(n3091), .Z(n3090) );
  BUFFD0 U3085 ( .I(n3092), .Z(n3091) );
  BUFFD0 U3086 ( .I(n3093), .Z(n3092) );
  BUFFD0 U3087 ( .I(n3094), .Z(n3093) );
  BUFFD0 U3088 ( .I(n3095), .Z(n3094) );
  BUFFD0 U3089 ( .I(n3096), .Z(n3095) );
  BUFFD0 U3090 ( .I(n3097), .Z(n3096) );
  BUFFD0 U3091 ( .I(n3098), .Z(n3097) );
  BUFFD0 U3092 ( .I(n3099), .Z(n3098) );
  BUFFD0 U3093 ( .I(n3100), .Z(n3099) );
  BUFFD0 U3094 ( .I(n3101), .Z(n3100) );
  BUFFD0 U3095 ( .I(n3102), .Z(n3101) );
  BUFFD0 U3096 ( .I(n3103), .Z(n3102) );
  BUFFD0 U3097 ( .I(n3104), .Z(n3103) );
  BUFFD0 U3098 ( .I(n3105), .Z(n3104) );
  BUFFD0 U3099 ( .I(n3106), .Z(n3105) );
  BUFFD0 U3100 ( .I(n3107), .Z(n3106) );
  BUFFD0 U3101 ( .I(n3108), .Z(n3107) );
  BUFFD0 U3102 ( .I(n3109), .Z(n3108) );
  BUFFD0 U3103 ( .I(n3110), .Z(n3109) );
  BUFFD0 U3104 ( .I(n3111), .Z(n3110) );
  BUFFD0 U3105 ( .I(n3112), .Z(n3111) );
  BUFFD0 U3106 ( .I(n3113), .Z(n3112) );
  BUFFD0 U3107 ( .I(n3114), .Z(n3113) );
  BUFFD0 U3108 ( .I(n3115), .Z(n3114) );
  BUFFD0 U3109 ( .I(n3116), .Z(n3115) );
  BUFFD0 U3110 ( .I(n3117), .Z(n3116) );
  BUFFD0 U3111 ( .I(n3118), .Z(n3117) );
  BUFFD0 U3112 ( .I(n3119), .Z(n3118) );
  BUFFD0 U3113 ( .I(n3120), .Z(n3119) );
  BUFFD0 U3114 ( .I(n3121), .Z(n3120) );
  BUFFD0 U3115 ( .I(n3122), .Z(n3121) );
  BUFFD0 U3116 ( .I(n3123), .Z(n3122) );
  BUFFD0 U3117 ( .I(n3124), .Z(n3123) );
  BUFFD0 U3118 ( .I(n3125), .Z(n3124) );
  BUFFD0 U3119 ( .I(n3126), .Z(n3125) );
  BUFFD0 U3120 ( .I(n3127), .Z(n3126) );
  BUFFD0 U3121 ( .I(n3128), .Z(n3127) );
  BUFFD0 U3122 ( .I(n3129), .Z(n3128) );
  BUFFD0 U3123 ( .I(n3130), .Z(n3129) );
  BUFFD0 U3124 ( .I(n3131), .Z(n3130) );
  BUFFD0 U3125 ( .I(n3132), .Z(n3131) );
  BUFFD0 U3126 ( .I(n3133), .Z(n3132) );
  BUFFD0 U3127 ( .I(n3134), .Z(n3133) );
  BUFFD0 U3128 ( .I(n3135), .Z(n3134) );
  BUFFD0 U3129 ( .I(n3136), .Z(n3135) );
  BUFFD0 U3130 ( .I(n3137), .Z(n3136) );
  BUFFD0 U3131 ( .I(n3138), .Z(n3137) );
  BUFFD0 U3132 ( .I(n3139), .Z(n3138) );
  BUFFD0 U3133 ( .I(n3140), .Z(n3139) );
  BUFFD0 U3134 ( .I(n3141), .Z(n3140) );
  BUFFD0 U3135 ( .I(n3142), .Z(n3141) );
  BUFFD0 U3136 ( .I(n3143), .Z(n3142) );
  BUFFD0 U3137 ( .I(n3144), .Z(n3143) );
  BUFFD0 U3138 ( .I(n3145), .Z(n3144) );
  BUFFD0 U3139 ( .I(n3146), .Z(n3145) );
  BUFFD0 U3140 ( .I(n3147), .Z(n3146) );
  BUFFD0 U3141 ( .I(n3148), .Z(n3147) );
  BUFFD0 U3142 ( .I(n3149), .Z(n3148) );
  BUFFD0 U3143 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3144 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3145 ( .I(n3152), .Z(n3151) );
  BUFFD0 U3146 ( .I(n3153), .Z(n3152) );
  BUFFD0 U3147 ( .I(n3154), .Z(n3153) );
  BUFFD0 U3148 ( .I(n3155), .Z(n3154) );
  BUFFD0 U3149 ( .I(n3156), .Z(n3155) );
  BUFFD0 U3150 ( .I(n3157), .Z(n3156) );
  BUFFD0 U3151 ( .I(n3158), .Z(n3157) );
  BUFFD0 U3152 ( .I(n3159), .Z(n3158) );
  BUFFD0 U3153 ( .I(n3160), .Z(n3159) );
  BUFFD0 U3154 ( .I(n3161), .Z(n3160) );
  BUFFD0 U3155 ( .I(n3162), .Z(n3161) );
  BUFFD0 U3156 ( .I(n3163), .Z(n3162) );
  BUFFD0 U3157 ( .I(n3164), .Z(n3163) );
  BUFFD0 U3158 ( .I(n3165), .Z(n3164) );
  BUFFD0 U3159 ( .I(n3166), .Z(n3165) );
  BUFFD0 U3160 ( .I(n3167), .Z(n3166) );
  BUFFD0 U3161 ( .I(n3168), .Z(n3167) );
  BUFFD0 U3162 ( .I(n3169), .Z(n3168) );
  BUFFD0 U3163 ( .I(n3170), .Z(n3169) );
  BUFFD0 U3164 ( .I(n3171), .Z(n3170) );
  BUFFD0 U3165 ( .I(n3172), .Z(n3171) );
  BUFFD0 U3166 ( .I(n3173), .Z(n3172) );
  BUFFD0 U3167 ( .I(n3174), .Z(n3173) );
  BUFFD0 U3168 ( .I(n3175), .Z(n3174) );
  BUFFD0 U3169 ( .I(n3176), .Z(n3175) );
  BUFFD0 U3170 ( .I(n3177), .Z(n3176) );
  BUFFD0 U3171 ( .I(n3178), .Z(n3177) );
  BUFFD0 U3172 ( .I(n3179), .Z(n3178) );
  BUFFD0 U3173 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3174 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3175 ( .I(n3182), .Z(n3181) );
  BUFFD0 U3176 ( .I(n3183), .Z(n3182) );
  BUFFD0 U3177 ( .I(n3184), .Z(n3183) );
  BUFFD0 U3178 ( .I(n3185), .Z(n3184) );
  BUFFD0 U3179 ( .I(n3186), .Z(n3185) );
  BUFFD0 U3180 ( .I(n3187), .Z(n3186) );
  BUFFD0 U3181 ( .I(n3188), .Z(n3187) );
  BUFFD0 U3182 ( .I(n3189), .Z(n3188) );
  BUFFD0 U3183 ( .I(n3190), .Z(n3189) );
  BUFFD0 U3184 ( .I(n3191), .Z(n3190) );
  BUFFD0 U3185 ( .I(n3192), .Z(n3191) );
  BUFFD0 U3186 ( .I(n3193), .Z(n3192) );
  BUFFD0 U3187 ( .I(n3194), .Z(n3193) );
  BUFFD0 U3188 ( .I(n3195), .Z(n3194) );
  BUFFD0 U3189 ( .I(n3196), .Z(n3195) );
  BUFFD0 U3190 ( .I(n3197), .Z(n3196) );
  BUFFD0 U3191 ( .I(n3198), .Z(n3197) );
  BUFFD0 U3192 ( .I(n3199), .Z(n3198) );
  BUFFD0 U3193 ( .I(n3200), .Z(n3199) );
  BUFFD0 U3194 ( .I(n3201), .Z(n3200) );
  BUFFD0 U3195 ( .I(n3202), .Z(n3201) );
  BUFFD0 U3196 ( .I(n8741), .Z(n3202) );
  BUFFD0 U3197 ( .I(n8737), .Z(n3203) );
  BUFFD0 U3198 ( .I(n3205), .Z(n3204) );
  BUFFD0 U3199 ( .I(n3206), .Z(n3205) );
  BUFFD0 U3200 ( .I(n3207), .Z(n3206) );
  BUFFD0 U3201 ( .I(n3208), .Z(n3207) );
  BUFFD0 U3202 ( .I(n3209), .Z(n3208) );
  BUFFD0 U3203 ( .I(n3210), .Z(n3209) );
  BUFFD0 U3204 ( .I(n3211), .Z(n3210) );
  BUFFD0 U3205 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3206 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3207 ( .I(n3214), .Z(n3213) );
  BUFFD0 U3208 ( .I(n3215), .Z(n3214) );
  BUFFD0 U3209 ( .I(n3216), .Z(n3215) );
  BUFFD0 U3210 ( .I(n3217), .Z(n3216) );
  BUFFD0 U3211 ( .I(n3218), .Z(n3217) );
  BUFFD0 U3212 ( .I(n3219), .Z(n3218) );
  BUFFD0 U3213 ( .I(n3220), .Z(n3219) );
  BUFFD0 U3214 ( .I(n3221), .Z(n3220) );
  BUFFD0 U3215 ( .I(n3222), .Z(n3221) );
  BUFFD0 U3216 ( .I(n3223), .Z(n3222) );
  BUFFD0 U3217 ( .I(n3224), .Z(n3223) );
  BUFFD0 U3218 ( .I(n3225), .Z(n3224) );
  BUFFD0 U3219 ( .I(n3226), .Z(n3225) );
  BUFFD0 U3220 ( .I(n3227), .Z(n3226) );
  BUFFD0 U3221 ( .I(n3228), .Z(n3227) );
  BUFFD0 U3222 ( .I(n3229), .Z(n3228) );
  BUFFD0 U3223 ( .I(n3230), .Z(n3229) );
  BUFFD0 U3224 ( .I(n3231), .Z(n3230) );
  BUFFD0 U3225 ( .I(n3232), .Z(n3231) );
  BUFFD0 U3226 ( .I(n3233), .Z(n3232) );
  BUFFD0 U3227 ( .I(n3234), .Z(n3233) );
  BUFFD0 U3228 ( .I(n3235), .Z(n3234) );
  BUFFD0 U3229 ( .I(n3236), .Z(n3235) );
  BUFFD0 U3230 ( .I(n3237), .Z(n3236) );
  BUFFD0 U3231 ( .I(n3238), .Z(n3237) );
  BUFFD0 U3232 ( .I(n3239), .Z(n3238) );
  BUFFD0 U3233 ( .I(n3240), .Z(n3239) );
  BUFFD0 U3234 ( .I(n3241), .Z(n3240) );
  BUFFD0 U3235 ( .I(n3242), .Z(n3241) );
  BUFFD0 U3236 ( .I(n3243), .Z(n3242) );
  BUFFD0 U3237 ( .I(n3244), .Z(n3243) );
  BUFFD0 U3238 ( .I(n3245), .Z(n3244) );
  BUFFD0 U3239 ( .I(n3246), .Z(n3245) );
  BUFFD0 U3240 ( .I(n3247), .Z(n3246) );
  BUFFD0 U3241 ( .I(n3248), .Z(n3247) );
  BUFFD0 U3242 ( .I(n3249), .Z(n3248) );
  BUFFD0 U3243 ( .I(n3250), .Z(n3249) );
  BUFFD0 U3244 ( .I(n3251), .Z(n3250) );
  BUFFD0 U3245 ( .I(n3252), .Z(n3251) );
  BUFFD0 U3246 ( .I(n3253), .Z(n3252) );
  BUFFD0 U3247 ( .I(n3254), .Z(n3253) );
  BUFFD0 U3248 ( .I(n3255), .Z(n3254) );
  BUFFD0 U3249 ( .I(n3256), .Z(n3255) );
  BUFFD0 U3250 ( .I(n3257), .Z(n3256) );
  BUFFD0 U3251 ( .I(n3258), .Z(n3257) );
  BUFFD0 U3252 ( .I(n3259), .Z(n3258) );
  BUFFD0 U3253 ( .I(n3260), .Z(n3259) );
  BUFFD0 U3254 ( .I(n3261), .Z(n3260) );
  BUFFD0 U3255 ( .I(n3262), .Z(n3261) );
  BUFFD0 U3256 ( .I(n3263), .Z(n3262) );
  BUFFD0 U3257 ( .I(n3264), .Z(n3263) );
  BUFFD0 U3258 ( .I(n3265), .Z(n3264) );
  BUFFD0 U3259 ( .I(n3266), .Z(n3265) );
  BUFFD0 U3260 ( .I(n3267), .Z(n3266) );
  BUFFD0 U3261 ( .I(n3268), .Z(n3267) );
  BUFFD0 U3262 ( .I(n3269), .Z(n3268) );
  BUFFD0 U3263 ( .I(n3270), .Z(n3269) );
  BUFFD0 U3264 ( .I(n3271), .Z(n3270) );
  BUFFD0 U3265 ( .I(n3272), .Z(n3271) );
  BUFFD0 U3266 ( .I(n3273), .Z(n3272) );
  BUFFD0 U3267 ( .I(n3274), .Z(n3273) );
  BUFFD0 U3268 ( .I(n3275), .Z(n3274) );
  BUFFD0 U3269 ( .I(n3276), .Z(n3275) );
  BUFFD0 U3270 ( .I(n3277), .Z(n3276) );
  BUFFD0 U3271 ( .I(n3278), .Z(n3277) );
  BUFFD0 U3272 ( .I(n3279), .Z(n3278) );
  BUFFD0 U3273 ( .I(n3280), .Z(n3279) );
  BUFFD0 U3274 ( .I(n3281), .Z(n3280) );
  BUFFD0 U3275 ( .I(n3282), .Z(n3281) );
  BUFFD0 U3276 ( .I(n3283), .Z(n3282) );
  BUFFD0 U3277 ( .I(n3284), .Z(n3283) );
  BUFFD0 U3278 ( .I(n3285), .Z(n3284) );
  BUFFD0 U3279 ( .I(n3286), .Z(n3285) );
  BUFFD0 U3280 ( .I(n3287), .Z(n3286) );
  BUFFD0 U3281 ( .I(n3288), .Z(n3287) );
  BUFFD0 U3282 ( .I(n3289), .Z(n3288) );
  BUFFD0 U3283 ( .I(n3290), .Z(n3289) );
  BUFFD0 U3284 ( .I(n3291), .Z(n3290) );
  BUFFD0 U3285 ( .I(n3292), .Z(n3291) );
  BUFFD0 U3286 ( .I(n3293), .Z(n3292) );
  BUFFD0 U3287 ( .I(n3294), .Z(n3293) );
  BUFFD0 U3288 ( .I(n3295), .Z(n3294) );
  BUFFD0 U3289 ( .I(n3296), .Z(n3295) );
  BUFFD0 U3290 ( .I(n3297), .Z(n3296) );
  BUFFD0 U3291 ( .I(n3298), .Z(n3297) );
  BUFFD0 U3292 ( .I(n3299), .Z(n3298) );
  BUFFD0 U3293 ( .I(n3300), .Z(n3299) );
  BUFFD0 U3294 ( .I(n3301), .Z(n3300) );
  BUFFD0 U3295 ( .I(n3302), .Z(n3301) );
  BUFFD0 U3296 ( .I(n3303), .Z(n3302) );
  BUFFD0 U3297 ( .I(n3304), .Z(n3303) );
  BUFFD0 U3298 ( .I(n3305), .Z(n3304) );
  BUFFD0 U3299 ( .I(n3306), .Z(n3305) );
  BUFFD0 U3300 ( .I(n3307), .Z(n3306) );
  BUFFD0 U3301 ( .I(n3308), .Z(n3307) );
  BUFFD0 U3302 ( .I(n3309), .Z(n3308) );
  BUFFD0 U3303 ( .I(n3310), .Z(n3309) );
  BUFFD0 U3304 ( .I(n3311), .Z(n3310) );
  BUFFD0 U3305 ( .I(n3312), .Z(n3311) );
  BUFFD0 U3306 ( .I(n3313), .Z(n3312) );
  BUFFD0 U3307 ( .I(n3314), .Z(n3313) );
  BUFFD0 U3308 ( .I(n3315), .Z(n3314) );
  BUFFD0 U3309 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3310 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3311 ( .I(n3318), .Z(n3317) );
  BUFFD0 U3312 ( .I(n3319), .Z(n3318) );
  BUFFD0 U3313 ( .I(n3320), .Z(n3319) );
  BUFFD0 U3314 ( .I(n3321), .Z(n3320) );
  BUFFD0 U3315 ( .I(n3322), .Z(n3321) );
  BUFFD0 U3316 ( .I(n3323), .Z(n3322) );
  BUFFD0 U3317 ( .I(n3324), .Z(n3323) );
  BUFFD0 U3318 ( .I(n3325), .Z(n3324) );
  BUFFD0 U3319 ( .I(n3326), .Z(n3325) );
  BUFFD0 U3320 ( .I(n3327), .Z(n3326) );
  BUFFD0 U3321 ( .I(n3328), .Z(n3327) );
  BUFFD0 U3322 ( .I(n3329), .Z(n3328) );
  BUFFD0 U3323 ( .I(n3330), .Z(n3329) );
  BUFFD0 U3324 ( .I(n3331), .Z(n3330) );
  BUFFD0 U3325 ( .I(n3332), .Z(n3331) );
  BUFFD0 U3326 ( .I(n3333), .Z(n3332) );
  BUFFD0 U3327 ( .I(n3334), .Z(n3333) );
  BUFFD0 U3328 ( .I(n3335), .Z(n3334) );
  BUFFD0 U3329 ( .I(n3336), .Z(n3335) );
  BUFFD0 U3330 ( .I(n3337), .Z(n3336) );
  BUFFD0 U3331 ( .I(n3338), .Z(n3337) );
  BUFFD0 U3332 ( .I(n3339), .Z(n3338) );
  BUFFD0 U3333 ( .I(n3340), .Z(n3339) );
  BUFFD0 U3334 ( .I(n3341), .Z(n3340) );
  BUFFD0 U3335 ( .I(n3342), .Z(n3341) );
  BUFFD0 U3336 ( .I(n3343), .Z(n3342) );
  BUFFD0 U3337 ( .I(n3344), .Z(n3343) );
  BUFFD0 U3338 ( .I(n3345), .Z(n3344) );
  BUFFD0 U3339 ( .I(n3346), .Z(n3345) );
  BUFFD0 U3340 ( .I(n3347), .Z(n3346) );
  BUFFD0 U3341 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3342 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3343 ( .I(n3350), .Z(n3349) );
  BUFFD0 U3344 ( .I(n3351), .Z(n3350) );
  BUFFD0 U3345 ( .I(n3352), .Z(n3351) );
  BUFFD0 U3346 ( .I(n3353), .Z(n3352) );
  BUFFD0 U3347 ( .I(n3354), .Z(n3353) );
  BUFFD0 U3348 ( .I(n3355), .Z(n3354) );
  BUFFD0 U3349 ( .I(n3356), .Z(n3355) );
  BUFFD0 U3350 ( .I(n3357), .Z(n3356) );
  BUFFD0 U3351 ( .I(n3358), .Z(n3357) );
  BUFFD0 U3352 ( .I(n3359), .Z(n3358) );
  BUFFD0 U3353 ( .I(n3360), .Z(n3359) );
  BUFFD0 U3354 ( .I(n3361), .Z(n3360) );
  BUFFD0 U3355 ( .I(n3362), .Z(n3361) );
  BUFFD0 U3356 ( .I(n3363), .Z(n3362) );
  BUFFD0 U3357 ( .I(n3364), .Z(n3363) );
  BUFFD0 U3358 ( .I(n3365), .Z(n3364) );
  BUFFD0 U3359 ( .I(n3366), .Z(n3365) );
  BUFFD0 U3360 ( .I(n3367), .Z(n3366) );
  BUFFD0 U3361 ( .I(n3368), .Z(n3367) );
  BUFFD0 U3362 ( .I(n3369), .Z(n3368) );
  BUFFD0 U3363 ( .I(n3370), .Z(n3369) );
  BUFFD0 U3364 ( .I(n3371), .Z(n3370) );
  BUFFD0 U3365 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3366 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3367 ( .I(n3374), .Z(n3373) );
  BUFFD0 U3368 ( .I(n3375), .Z(n3374) );
  BUFFD0 U3369 ( .I(n3376), .Z(n3375) );
  BUFFD0 U3370 ( .I(n3377), .Z(n3376) );
  BUFFD0 U3371 ( .I(n3378), .Z(n3377) );
  BUFFD0 U3372 ( .I(n3379), .Z(n3378) );
  BUFFD0 U3373 ( .I(n3380), .Z(n3379) );
  BUFFD0 U3374 ( .I(n3381), .Z(n3380) );
  BUFFD0 U3375 ( .I(n8738), .Z(n3381) );
  BUFFD0 U3376 ( .I(n8735), .Z(n3382) );
  BUFFD0 U3377 ( .I(n3384), .Z(n3383) );
  BUFFD0 U3378 ( .I(n3385), .Z(n3384) );
  BUFFD0 U3379 ( .I(n3386), .Z(n3385) );
  BUFFD0 U3380 ( .I(n3387), .Z(n3386) );
  BUFFD0 U3381 ( .I(n3388), .Z(n3387) );
  BUFFD0 U3382 ( .I(n3389), .Z(n3388) );
  BUFFD0 U3383 ( .I(n3390), .Z(n3389) );
  BUFFD0 U3384 ( .I(n3391), .Z(n3390) );
  BUFFD0 U3385 ( .I(n3392), .Z(n3391) );
  BUFFD0 U3386 ( .I(n3393), .Z(n3392) );
  BUFFD0 U3387 ( .I(n3394), .Z(n3393) );
  BUFFD0 U3388 ( .I(n3395), .Z(n3394) );
  BUFFD0 U3389 ( .I(n3396), .Z(n3395) );
  BUFFD0 U3390 ( .I(n3397), .Z(n3396) );
  BUFFD0 U3391 ( .I(n3398), .Z(n3397) );
  BUFFD0 U3392 ( .I(n3399), .Z(n3398) );
  BUFFD0 U3393 ( .I(n3400), .Z(n3399) );
  BUFFD0 U3394 ( .I(n3401), .Z(n3400) );
  BUFFD0 U3395 ( .I(n3402), .Z(n3401) );
  BUFFD0 U3396 ( .I(n3403), .Z(n3402) );
  BUFFD0 U3397 ( .I(n3404), .Z(n3403) );
  BUFFD0 U3398 ( .I(n3405), .Z(n3404) );
  BUFFD0 U3399 ( .I(n3406), .Z(n3405) );
  BUFFD0 U3400 ( .I(n3407), .Z(n3406) );
  BUFFD0 U3401 ( .I(n3408), .Z(n3407) );
  BUFFD0 U3402 ( .I(n3409), .Z(n3408) );
  BUFFD0 U3403 ( .I(n3410), .Z(n3409) );
  BUFFD0 U3404 ( .I(n3411), .Z(n3410) );
  BUFFD0 U3405 ( .I(n3412), .Z(n3411) );
  BUFFD0 U3406 ( .I(n3413), .Z(n3412) );
  BUFFD0 U3407 ( .I(n3414), .Z(n3413) );
  BUFFD0 U3408 ( .I(n3415), .Z(n3414) );
  BUFFD0 U3409 ( .I(n3416), .Z(n3415) );
  BUFFD0 U3410 ( .I(n3417), .Z(n3416) );
  BUFFD0 U3411 ( .I(n3418), .Z(n3417) );
  BUFFD0 U3412 ( .I(n3419), .Z(n3418) );
  BUFFD0 U3413 ( .I(n3420), .Z(n3419) );
  BUFFD0 U3414 ( .I(n3421), .Z(n3420) );
  BUFFD0 U3415 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3416 ( .I(n3423), .Z(n3422) );
  BUFFD0 U3417 ( .I(n3424), .Z(n3423) );
  BUFFD0 U3418 ( .I(n3425), .Z(n3424) );
  BUFFD0 U3419 ( .I(n3426), .Z(n3425) );
  BUFFD0 U3420 ( .I(n3427), .Z(n3426) );
  BUFFD0 U3421 ( .I(n3428), .Z(n3427) );
  BUFFD0 U3422 ( .I(n3429), .Z(n3428) );
  BUFFD0 U3423 ( .I(n3430), .Z(n3429) );
  BUFFD0 U3424 ( .I(n3431), .Z(n3430) );
  BUFFD0 U3425 ( .I(n3432), .Z(n3431) );
  BUFFD0 U3426 ( .I(n3433), .Z(n3432) );
  BUFFD0 U3427 ( .I(n3434), .Z(n3433) );
  BUFFD0 U3428 ( .I(n3435), .Z(n3434) );
  BUFFD0 U3429 ( .I(n3436), .Z(n3435) );
  BUFFD0 U3430 ( .I(n3437), .Z(n3436) );
  BUFFD0 U3431 ( .I(n3438), .Z(n3437) );
  BUFFD0 U3432 ( .I(n3439), .Z(n3438) );
  BUFFD0 U3433 ( .I(n3440), .Z(n3439) );
  BUFFD0 U3434 ( .I(n3441), .Z(n3440) );
  BUFFD0 U3435 ( .I(n3442), .Z(n3441) );
  BUFFD0 U3436 ( .I(n3443), .Z(n3442) );
  BUFFD0 U3437 ( .I(n3444), .Z(n3443) );
  BUFFD0 U3438 ( .I(n3445), .Z(n3444) );
  BUFFD0 U3439 ( .I(n3446), .Z(n3445) );
  BUFFD0 U3440 ( .I(n3447), .Z(n3446) );
  BUFFD0 U3441 ( .I(n3448), .Z(n3447) );
  BUFFD0 U3442 ( .I(n3449), .Z(n3448) );
  BUFFD0 U3443 ( .I(n3450), .Z(n3449) );
  BUFFD0 U3444 ( .I(n3451), .Z(n3450) );
  BUFFD0 U3445 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3446 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3447 ( .I(n3454), .Z(n3453) );
  BUFFD0 U3448 ( .I(n3455), .Z(n3454) );
  BUFFD0 U3449 ( .I(n3456), .Z(n3455) );
  BUFFD0 U3450 ( .I(n3457), .Z(n3456) );
  BUFFD0 U3451 ( .I(n3458), .Z(n3457) );
  BUFFD0 U3452 ( .I(n3459), .Z(n3458) );
  BUFFD0 U3453 ( .I(n3460), .Z(n3459) );
  BUFFD0 U3454 ( .I(n3461), .Z(n3460) );
  BUFFD0 U3455 ( .I(n3462), .Z(n3461) );
  BUFFD0 U3456 ( .I(n3463), .Z(n3462) );
  BUFFD0 U3457 ( .I(n3464), .Z(n3463) );
  BUFFD0 U3458 ( .I(n3465), .Z(n3464) );
  BUFFD0 U3459 ( .I(n3466), .Z(n3465) );
  BUFFD0 U3460 ( .I(n3467), .Z(n3466) );
  BUFFD0 U3461 ( .I(n3468), .Z(n3467) );
  BUFFD0 U3462 ( .I(n3469), .Z(n3468) );
  BUFFD0 U3463 ( .I(n3470), .Z(n3469) );
  BUFFD0 U3464 ( .I(n3471), .Z(n3470) );
  BUFFD0 U3465 ( .I(n3472), .Z(n3471) );
  BUFFD0 U3466 ( .I(n3473), .Z(n3472) );
  BUFFD0 U3467 ( .I(n3474), .Z(n3473) );
  BUFFD0 U3468 ( .I(n3475), .Z(n3474) );
  BUFFD0 U3469 ( .I(n3476), .Z(n3475) );
  BUFFD0 U3470 ( .I(n3477), .Z(n3476) );
  BUFFD0 U3471 ( .I(n3478), .Z(n3477) );
  BUFFD0 U3472 ( .I(n3479), .Z(n3478) );
  BUFFD0 U3473 ( .I(n3480), .Z(n3479) );
  BUFFD0 U3474 ( .I(n3481), .Z(n3480) );
  BUFFD0 U3475 ( .I(n3482), .Z(n3481) );
  BUFFD0 U3476 ( .I(n3483), .Z(n3482) );
  BUFFD0 U3477 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3478 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3479 ( .I(n3486), .Z(n3485) );
  BUFFD0 U3480 ( .I(n3487), .Z(n3486) );
  BUFFD0 U3481 ( .I(n3488), .Z(n3487) );
  BUFFD0 U3482 ( .I(n3489), .Z(n3488) );
  BUFFD0 U3483 ( .I(n3490), .Z(n3489) );
  BUFFD0 U3484 ( .I(n3491), .Z(n3490) );
  BUFFD0 U3485 ( .I(n3492), .Z(n3491) );
  BUFFD0 U3486 ( .I(n3493), .Z(n3492) );
  BUFFD0 U3487 ( .I(n3494), .Z(n3493) );
  BUFFD0 U3488 ( .I(n3495), .Z(n3494) );
  BUFFD0 U3489 ( .I(n3496), .Z(n3495) );
  BUFFD0 U3490 ( .I(n3497), .Z(n3496) );
  BUFFD0 U3491 ( .I(n3498), .Z(n3497) );
  BUFFD0 U3492 ( .I(n3499), .Z(n3498) );
  BUFFD0 U3493 ( .I(n3500), .Z(n3499) );
  BUFFD0 U3494 ( .I(n3501), .Z(n3500) );
  BUFFD0 U3495 ( .I(n3502), .Z(n3501) );
  BUFFD0 U3496 ( .I(n3503), .Z(n3502) );
  BUFFD0 U3497 ( .I(n3504), .Z(n3503) );
  BUFFD0 U3498 ( .I(n3505), .Z(n3504) );
  BUFFD0 U3499 ( .I(n3506), .Z(n3505) );
  BUFFD0 U3500 ( .I(n3507), .Z(n3506) );
  BUFFD0 U3501 ( .I(n3508), .Z(n3507) );
  BUFFD0 U3502 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3503 ( .I(n3510), .Z(n3509) );
  BUFFD0 U3504 ( .I(n3511), .Z(n3510) );
  BUFFD0 U3505 ( .I(n3512), .Z(n3511) );
  BUFFD0 U3506 ( .I(n3513), .Z(n3512) );
  BUFFD0 U3507 ( .I(n3514), .Z(n3513) );
  BUFFD0 U3508 ( .I(n3515), .Z(n3514) );
  BUFFD0 U3509 ( .I(n3516), .Z(n3515) );
  BUFFD0 U3510 ( .I(n3517), .Z(n3516) );
  BUFFD0 U3511 ( .I(n3518), .Z(n3517) );
  BUFFD0 U3512 ( .I(n3519), .Z(n3518) );
  BUFFD0 U3513 ( .I(n3520), .Z(n3519) );
  BUFFD0 U3514 ( .I(n3521), .Z(n3520) );
  BUFFD0 U3515 ( .I(n3522), .Z(n3521) );
  BUFFD0 U3516 ( .I(n3523), .Z(n3522) );
  BUFFD0 U3517 ( .I(n3524), .Z(n3523) );
  BUFFD0 U3518 ( .I(n3525), .Z(n3524) );
  BUFFD0 U3519 ( .I(n3526), .Z(n3525) );
  BUFFD0 U3520 ( .I(n3527), .Z(n3526) );
  BUFFD0 U3521 ( .I(n3528), .Z(n3527) );
  BUFFD0 U3522 ( .I(n3529), .Z(n3528) );
  BUFFD0 U3523 ( .I(n3530), .Z(n3529) );
  BUFFD0 U3524 ( .I(n3531), .Z(n3530) );
  BUFFD0 U3525 ( .I(n3532), .Z(n3531) );
  BUFFD0 U3526 ( .I(n3533), .Z(n3532) );
  BUFFD0 U3527 ( .I(n3534), .Z(n3533) );
  BUFFD0 U3528 ( .I(n3535), .Z(n3534) );
  BUFFD0 U3529 ( .I(n3536), .Z(n3535) );
  BUFFD0 U3530 ( .I(n3537), .Z(n3536) );
  BUFFD0 U3531 ( .I(n3538), .Z(n3537) );
  BUFFD0 U3532 ( .I(n3539), .Z(n3538) );
  BUFFD0 U3533 ( .I(n3540), .Z(n3539) );
  BUFFD0 U3534 ( .I(n3541), .Z(n3540) );
  BUFFD0 U3535 ( .I(n3542), .Z(n3541) );
  BUFFD0 U3536 ( .I(n3543), .Z(n3542) );
  BUFFD0 U3537 ( .I(n3544), .Z(n3543) );
  BUFFD0 U3538 ( .I(n3545), .Z(n3544) );
  BUFFD0 U3539 ( .I(n3546), .Z(n3545) );
  BUFFD0 U3540 ( .I(n3547), .Z(n3546) );
  BUFFD0 U3541 ( .I(n3548), .Z(n3547) );
  BUFFD0 U3542 ( .I(n3549), .Z(n3548) );
  BUFFD0 U3543 ( .I(n3550), .Z(n3549) );
  BUFFD0 U3544 ( .I(n3551), .Z(n3550) );
  BUFFD0 U3545 ( .I(n3552), .Z(n3551) );
  BUFFD0 U3546 ( .I(n3553), .Z(n3552) );
  BUFFD0 U3547 ( .I(n3554), .Z(n3553) );
  BUFFD0 U3548 ( .I(n3555), .Z(n3554) );
  BUFFD0 U3549 ( .I(n3556), .Z(n3555) );
  BUFFD0 U3550 ( .I(n3557), .Z(n3556) );
  BUFFD0 U3551 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3552 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3553 ( .I(n3560), .Z(n3559) );
  BUFFD0 U3554 ( .I(n8736), .Z(n3560) );
  BUFFD0 U3555 ( .I(n8733), .Z(n3561) );
  BUFFD0 U3556 ( .I(n3563), .Z(n3562) );
  BUFFD0 U3557 ( .I(n3564), .Z(n3563) );
  BUFFD0 U3558 ( .I(n3565), .Z(n3564) );
  BUFFD0 U3559 ( .I(n3566), .Z(n3565) );
  BUFFD0 U3560 ( .I(n3567), .Z(n3566) );
  BUFFD0 U3561 ( .I(n3568), .Z(n3567) );
  BUFFD0 U3562 ( .I(n3569), .Z(n3568) );
  BUFFD0 U3563 ( .I(n3570), .Z(n3569) );
  BUFFD0 U3564 ( .I(n3571), .Z(n3570) );
  BUFFD0 U3565 ( .I(n3572), .Z(n3571) );
  BUFFD0 U3566 ( .I(n3573), .Z(n3572) );
  BUFFD0 U3567 ( .I(n3574), .Z(n3573) );
  BUFFD0 U3568 ( .I(n3575), .Z(n3574) );
  BUFFD0 U3569 ( .I(n3576), .Z(n3575) );
  BUFFD0 U3570 ( .I(n3577), .Z(n3576) );
  BUFFD0 U3571 ( .I(n3578), .Z(n3577) );
  BUFFD0 U3572 ( .I(n3579), .Z(n3578) );
  BUFFD0 U3573 ( .I(n3580), .Z(n3579) );
  BUFFD0 U3574 ( .I(n3581), .Z(n3580) );
  BUFFD0 U3575 ( .I(n3582), .Z(n3581) );
  BUFFD0 U3576 ( .I(n3583), .Z(n3582) );
  BUFFD0 U3577 ( .I(n3584), .Z(n3583) );
  BUFFD0 U3578 ( .I(n3585), .Z(n3584) );
  BUFFD0 U3579 ( .I(n3586), .Z(n3585) );
  BUFFD0 U3580 ( .I(n3587), .Z(n3586) );
  BUFFD0 U3581 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3582 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3583 ( .I(n3590), .Z(n3589) );
  BUFFD0 U3584 ( .I(n3591), .Z(n3590) );
  BUFFD0 U3585 ( .I(n3592), .Z(n3591) );
  BUFFD0 U3586 ( .I(n3593), .Z(n3592) );
  BUFFD0 U3587 ( .I(n3594), .Z(n3593) );
  BUFFD0 U3588 ( .I(n3595), .Z(n3594) );
  BUFFD0 U3589 ( .I(n3596), .Z(n3595) );
  BUFFD0 U3590 ( .I(n3597), .Z(n3596) );
  BUFFD0 U3591 ( .I(n3598), .Z(n3597) );
  BUFFD0 U3592 ( .I(n3599), .Z(n3598) );
  BUFFD0 U3593 ( .I(n3600), .Z(n3599) );
  BUFFD0 U3594 ( .I(n3601), .Z(n3600) );
  BUFFD0 U3595 ( .I(n3602), .Z(n3601) );
  BUFFD0 U3596 ( .I(n3603), .Z(n3602) );
  BUFFD0 U3597 ( .I(n3604), .Z(n3603) );
  BUFFD0 U3598 ( .I(n3605), .Z(n3604) );
  BUFFD0 U3599 ( .I(n3606), .Z(n3605) );
  BUFFD0 U3600 ( .I(n3607), .Z(n3606) );
  BUFFD0 U3601 ( .I(n3608), .Z(n3607) );
  BUFFD0 U3602 ( .I(n3609), .Z(n3608) );
  BUFFD0 U3603 ( .I(n3610), .Z(n3609) );
  BUFFD0 U3604 ( .I(n3611), .Z(n3610) );
  BUFFD0 U3605 ( .I(n3612), .Z(n3611) );
  BUFFD0 U3606 ( .I(n3613), .Z(n3612) );
  BUFFD0 U3607 ( .I(n3614), .Z(n3613) );
  BUFFD0 U3608 ( .I(n3615), .Z(n3614) );
  BUFFD0 U3609 ( .I(n3616), .Z(n3615) );
  BUFFD0 U3610 ( .I(n3617), .Z(n3616) );
  BUFFD0 U3611 ( .I(n3618), .Z(n3617) );
  BUFFD0 U3612 ( .I(n3619), .Z(n3618) );
  BUFFD0 U3613 ( .I(n3620), .Z(n3619) );
  BUFFD0 U3614 ( .I(n3621), .Z(n3620) );
  BUFFD0 U3615 ( .I(n3622), .Z(n3621) );
  BUFFD0 U3616 ( .I(n3623), .Z(n3622) );
  BUFFD0 U3617 ( .I(n3624), .Z(n3623) );
  BUFFD0 U3618 ( .I(n3625), .Z(n3624) );
  BUFFD0 U3619 ( .I(n3626), .Z(n3625) );
  BUFFD0 U3620 ( .I(n3627), .Z(n3626) );
  BUFFD0 U3621 ( .I(n3628), .Z(n3627) );
  BUFFD0 U3622 ( .I(n3629), .Z(n3628) );
  BUFFD0 U3623 ( .I(n3630), .Z(n3629) );
  BUFFD0 U3624 ( .I(n3631), .Z(n3630) );
  BUFFD0 U3625 ( .I(n3632), .Z(n3631) );
  BUFFD0 U3626 ( .I(n3633), .Z(n3632) );
  BUFFD0 U3627 ( .I(n3634), .Z(n3633) );
  BUFFD0 U3628 ( .I(n3635), .Z(n3634) );
  BUFFD0 U3629 ( .I(n3636), .Z(n3635) );
  BUFFD0 U3630 ( .I(n3637), .Z(n3636) );
  BUFFD0 U3631 ( .I(n3638), .Z(n3637) );
  BUFFD0 U3632 ( .I(n3639), .Z(n3638) );
  BUFFD0 U3633 ( .I(n3640), .Z(n3639) );
  BUFFD0 U3634 ( .I(n3641), .Z(n3640) );
  BUFFD0 U3635 ( .I(n3642), .Z(n3641) );
  BUFFD0 U3636 ( .I(n3643), .Z(n3642) );
  BUFFD0 U3637 ( .I(n3644), .Z(n3643) );
  BUFFD0 U3638 ( .I(n3645), .Z(n3644) );
  BUFFD0 U3639 ( .I(n3646), .Z(n3645) );
  BUFFD0 U3640 ( .I(n3647), .Z(n3646) );
  BUFFD0 U3641 ( .I(n3648), .Z(n3647) );
  BUFFD0 U3642 ( .I(n3649), .Z(n3648) );
  BUFFD0 U3643 ( .I(n3650), .Z(n3649) );
  BUFFD0 U3644 ( .I(n3651), .Z(n3650) );
  BUFFD0 U3645 ( .I(n3652), .Z(n3651) );
  BUFFD0 U3646 ( .I(n3653), .Z(n3652) );
  BUFFD0 U3647 ( .I(n3654), .Z(n3653) );
  BUFFD0 U3648 ( .I(n3655), .Z(n3654) );
  BUFFD0 U3649 ( .I(n3656), .Z(n3655) );
  BUFFD0 U3650 ( .I(n3657), .Z(n3656) );
  BUFFD0 U3651 ( .I(n3658), .Z(n3657) );
  BUFFD0 U3652 ( .I(n3659), .Z(n3658) );
  BUFFD0 U3653 ( .I(n3660), .Z(n3659) );
  BUFFD0 U3654 ( .I(n3661), .Z(n3660) );
  BUFFD0 U3655 ( .I(n3662), .Z(n3661) );
  BUFFD0 U3656 ( .I(n3663), .Z(n3662) );
  BUFFD0 U3657 ( .I(n3664), .Z(n3663) );
  BUFFD0 U3658 ( .I(n3665), .Z(n3664) );
  BUFFD0 U3659 ( .I(n3666), .Z(n3665) );
  BUFFD0 U3660 ( .I(n3667), .Z(n3666) );
  BUFFD0 U3661 ( .I(n3668), .Z(n3667) );
  BUFFD0 U3662 ( .I(n3669), .Z(n3668) );
  BUFFD0 U3663 ( .I(n3670), .Z(n3669) );
  BUFFD0 U3664 ( .I(n3671), .Z(n3670) );
  BUFFD0 U3665 ( .I(n3672), .Z(n3671) );
  BUFFD0 U3666 ( .I(n3673), .Z(n3672) );
  BUFFD0 U3667 ( .I(n3674), .Z(n3673) );
  BUFFD0 U3668 ( .I(n3675), .Z(n3674) );
  BUFFD0 U3669 ( .I(n3676), .Z(n3675) );
  BUFFD0 U3670 ( .I(n3677), .Z(n3676) );
  BUFFD0 U3671 ( .I(n3678), .Z(n3677) );
  BUFFD0 U3672 ( .I(n3679), .Z(n3678) );
  BUFFD0 U3673 ( .I(n3680), .Z(n3679) );
  BUFFD0 U3674 ( .I(n3681), .Z(n3680) );
  BUFFD0 U3675 ( .I(n3682), .Z(n3681) );
  BUFFD0 U3676 ( .I(n3683), .Z(n3682) );
  BUFFD0 U3677 ( .I(n3684), .Z(n3683) );
  BUFFD0 U3678 ( .I(n3685), .Z(n3684) );
  BUFFD0 U3679 ( .I(n3686), .Z(n3685) );
  BUFFD0 U3680 ( .I(n3687), .Z(n3686) );
  BUFFD0 U3681 ( .I(n3688), .Z(n3687) );
  BUFFD0 U3682 ( .I(n3689), .Z(n3688) );
  BUFFD0 U3683 ( .I(n3690), .Z(n3689) );
  BUFFD0 U3684 ( .I(n3691), .Z(n3690) );
  BUFFD0 U3685 ( .I(n3692), .Z(n3691) );
  BUFFD0 U3686 ( .I(n3693), .Z(n3692) );
  BUFFD0 U3687 ( .I(n3694), .Z(n3693) );
  BUFFD0 U3688 ( .I(n3695), .Z(n3694) );
  BUFFD0 U3689 ( .I(n3696), .Z(n3695) );
  BUFFD0 U3690 ( .I(n3697), .Z(n3696) );
  BUFFD0 U3691 ( .I(n3698), .Z(n3697) );
  BUFFD0 U3692 ( .I(n3699), .Z(n3698) );
  BUFFD0 U3693 ( .I(n3700), .Z(n3699) );
  BUFFD0 U3694 ( .I(n3701), .Z(n3700) );
  BUFFD0 U3695 ( .I(n3702), .Z(n3701) );
  BUFFD0 U3696 ( .I(n3703), .Z(n3702) );
  BUFFD0 U3697 ( .I(n3704), .Z(n3703) );
  BUFFD0 U3698 ( .I(n3705), .Z(n3704) );
  BUFFD0 U3699 ( .I(n3706), .Z(n3705) );
  BUFFD0 U3700 ( .I(n3707), .Z(n3706) );
  BUFFD0 U3701 ( .I(n3708), .Z(n3707) );
  BUFFD0 U3702 ( .I(n3709), .Z(n3708) );
  BUFFD0 U3703 ( .I(n3710), .Z(n3709) );
  BUFFD0 U3704 ( .I(n3711), .Z(n3710) );
  BUFFD0 U3705 ( .I(n3712), .Z(n3711) );
  BUFFD0 U3706 ( .I(n3713), .Z(n3712) );
  BUFFD0 U3707 ( .I(n3714), .Z(n3713) );
  BUFFD0 U3708 ( .I(n3715), .Z(n3714) );
  BUFFD0 U3709 ( .I(n3716), .Z(n3715) );
  BUFFD0 U3710 ( .I(n3717), .Z(n3716) );
  BUFFD0 U3711 ( .I(n3718), .Z(n3717) );
  BUFFD0 U3712 ( .I(n3719), .Z(n3718) );
  BUFFD0 U3713 ( .I(n3720), .Z(n3719) );
  BUFFD0 U3714 ( .I(n3721), .Z(n3720) );
  BUFFD0 U3715 ( .I(n3722), .Z(n3721) );
  BUFFD0 U3716 ( .I(n3723), .Z(n3722) );
  BUFFD0 U3717 ( .I(n3724), .Z(n3723) );
  BUFFD0 U3718 ( .I(n3725), .Z(n3724) );
  BUFFD0 U3719 ( .I(n3726), .Z(n3725) );
  BUFFD0 U3720 ( .I(n3727), .Z(n3726) );
  BUFFD0 U3721 ( .I(n3728), .Z(n3727) );
  BUFFD0 U3722 ( .I(n3729), .Z(n3728) );
  BUFFD0 U3723 ( .I(n3730), .Z(n3729) );
  BUFFD0 U3724 ( .I(n3731), .Z(n3730) );
  BUFFD0 U3725 ( .I(n3732), .Z(n3731) );
  BUFFD0 U3726 ( .I(n3733), .Z(n3732) );
  BUFFD0 U3727 ( .I(n3734), .Z(n3733) );
  BUFFD0 U3728 ( .I(n3735), .Z(n3734) );
  BUFFD0 U3729 ( .I(n3736), .Z(n3735) );
  BUFFD0 U3730 ( .I(n3737), .Z(n3736) );
  BUFFD0 U3731 ( .I(n8734), .Z(n3737) );
  BUFFD0 U3732 ( .I(n3739), .Z(n3738) );
  BUFFD0 U3733 ( .I(n3740), .Z(n3739) );
  BUFFD0 U3734 ( .I(n3741), .Z(n3740) );
  BUFFD0 U3735 ( .I(n3742), .Z(n3741) );
  BUFFD0 U3736 ( .I(n3743), .Z(n3742) );
  BUFFD0 U3737 ( .I(n3744), .Z(n3743) );
  BUFFD0 U3738 ( .I(n3745), .Z(n3744) );
  BUFFD0 U3739 ( .I(n3746), .Z(n3745) );
  BUFFD0 U3740 ( .I(n3747), .Z(n3746) );
  BUFFD0 U3741 ( .I(n3748), .Z(n3747) );
  BUFFD0 U3742 ( .I(n3749), .Z(n3748) );
  BUFFD0 U3743 ( .I(n3750), .Z(n3749) );
  BUFFD0 U3744 ( .I(n3751), .Z(n3750) );
  BUFFD0 U3745 ( .I(n3752), .Z(n3751) );
  BUFFD0 U3746 ( .I(n3753), .Z(n3752) );
  BUFFD0 U3747 ( .I(n3754), .Z(n3753) );
  BUFFD0 U3748 ( .I(n3755), .Z(n3754) );
  BUFFD0 U3749 ( .I(n3756), .Z(n3755) );
  BUFFD0 U3750 ( .I(n3757), .Z(n3756) );
  BUFFD0 U3751 ( .I(n3758), .Z(n3757) );
  BUFFD0 U3752 ( .I(n3759), .Z(n3758) );
  BUFFD0 U3753 ( .I(n3760), .Z(n3759) );
  BUFFD0 U3754 ( .I(n3761), .Z(n3760) );
  BUFFD0 U3755 ( .I(n3762), .Z(n3761) );
  BUFFD0 U3756 ( .I(n3763), .Z(n3762) );
  BUFFD0 U3757 ( .I(n3764), .Z(n3763) );
  BUFFD0 U3758 ( .I(n3765), .Z(n3764) );
  BUFFD0 U3759 ( .I(n3766), .Z(n3765) );
  BUFFD0 U3760 ( .I(n3767), .Z(n3766) );
  BUFFD0 U3761 ( .I(n3768), .Z(n3767) );
  BUFFD0 U3762 ( .I(n3769), .Z(n3768) );
  BUFFD0 U3763 ( .I(n3770), .Z(n3769) );
  BUFFD0 U3764 ( .I(n3771), .Z(n3770) );
  BUFFD0 U3765 ( .I(n3772), .Z(n3771) );
  BUFFD0 U3766 ( .I(n3773), .Z(n3772) );
  BUFFD0 U3767 ( .I(n3774), .Z(n3773) );
  BUFFD0 U3768 ( .I(n3775), .Z(n3774) );
  BUFFD0 U3769 ( .I(n3776), .Z(n3775) );
  BUFFD0 U3770 ( .I(n3777), .Z(n3776) );
  BUFFD0 U3771 ( .I(n3778), .Z(n3777) );
  BUFFD0 U3772 ( .I(n3779), .Z(n3778) );
  BUFFD0 U3773 ( .I(n3780), .Z(n3779) );
  BUFFD0 U3774 ( .I(n3781), .Z(n3780) );
  BUFFD0 U3775 ( .I(n3782), .Z(n3781) );
  BUFFD0 U3776 ( .I(n3783), .Z(n3782) );
  BUFFD0 U3777 ( .I(n3784), .Z(n3783) );
  BUFFD0 U3778 ( .I(n3785), .Z(n3784) );
  BUFFD0 U3779 ( .I(n3786), .Z(n3785) );
  BUFFD0 U3780 ( .I(n3787), .Z(n3786) );
  BUFFD0 U3781 ( .I(n3788), .Z(n3787) );
  BUFFD0 U3782 ( .I(n3789), .Z(n3788) );
  BUFFD0 U3783 ( .I(n3790), .Z(n3789) );
  BUFFD0 U3784 ( .I(n3791), .Z(n3790) );
  BUFFD0 U3785 ( .I(n3792), .Z(n3791) );
  BUFFD0 U3786 ( .I(n3793), .Z(n3792) );
  BUFFD0 U3787 ( .I(n3794), .Z(n3793) );
  BUFFD0 U3788 ( .I(n3795), .Z(n3794) );
  BUFFD0 U3789 ( .I(n3796), .Z(n3795) );
  BUFFD0 U3790 ( .I(n3797), .Z(n3796) );
  BUFFD0 U3791 ( .I(n3798), .Z(n3797) );
  BUFFD0 U3792 ( .I(n3799), .Z(n3798) );
  BUFFD0 U3793 ( .I(n3800), .Z(n3799) );
  BUFFD0 U3794 ( .I(n3801), .Z(n3800) );
  BUFFD0 U3795 ( .I(n3802), .Z(n3801) );
  BUFFD0 U3796 ( .I(n3803), .Z(n3802) );
  BUFFD0 U3797 ( .I(n3804), .Z(n3803) );
  BUFFD0 U3798 ( .I(n3805), .Z(n3804) );
  BUFFD0 U3799 ( .I(n3806), .Z(n3805) );
  BUFFD0 U3800 ( .I(n3807), .Z(n3806) );
  BUFFD0 U3801 ( .I(n3808), .Z(n3807) );
  BUFFD0 U3802 ( .I(n3809), .Z(n3808) );
  BUFFD0 U3803 ( .I(n3810), .Z(n3809) );
  BUFFD0 U3804 ( .I(n3811), .Z(n3810) );
  BUFFD0 U3805 ( .I(n3812), .Z(n3811) );
  BUFFD0 U3806 ( .I(n3813), .Z(n3812) );
  BUFFD0 U3807 ( .I(n3814), .Z(n3813) );
  BUFFD0 U3808 ( .I(n3815), .Z(n3814) );
  BUFFD0 U3809 ( .I(n3816), .Z(n3815) );
  BUFFD0 U3810 ( .I(n3817), .Z(n3816) );
  BUFFD0 U3811 ( .I(n3818), .Z(n3817) );
  BUFFD0 U3812 ( .I(n3819), .Z(n3818) );
  BUFFD0 U3813 ( .I(n3820), .Z(n3819) );
  BUFFD0 U3814 ( .I(n3821), .Z(n3820) );
  BUFFD0 U3815 ( .I(n3822), .Z(n3821) );
  BUFFD0 U3816 ( .I(n3823), .Z(n3822) );
  BUFFD0 U3817 ( .I(n3824), .Z(n3823) );
  BUFFD0 U3818 ( .I(n3825), .Z(n3824) );
  BUFFD0 U3819 ( .I(n3826), .Z(n3825) );
  BUFFD0 U3820 ( .I(n3827), .Z(n3826) );
  BUFFD0 U3821 ( .I(n3828), .Z(n3827) );
  BUFFD0 U3822 ( .I(n3829), .Z(n3828) );
  BUFFD0 U3823 ( .I(n3830), .Z(n3829) );
  BUFFD0 U3824 ( .I(n3831), .Z(n3830) );
  BUFFD0 U3825 ( .I(n3832), .Z(n3831) );
  BUFFD0 U3826 ( .I(n3833), .Z(n3832) );
  BUFFD0 U3827 ( .I(n3834), .Z(n3833) );
  BUFFD0 U3828 ( .I(n3835), .Z(n3834) );
  BUFFD0 U3829 ( .I(n3836), .Z(n3835) );
  BUFFD0 U3830 ( .I(n3837), .Z(n3836) );
  BUFFD0 U3831 ( .I(n3838), .Z(n3837) );
  BUFFD0 U3832 ( .I(n3839), .Z(n3838) );
  BUFFD0 U3833 ( .I(n3840), .Z(n3839) );
  BUFFD0 U3834 ( .I(n3841), .Z(n3840) );
  BUFFD0 U3835 ( .I(n3842), .Z(n3841) );
  BUFFD0 U3836 ( .I(n3843), .Z(n3842) );
  BUFFD0 U3837 ( .I(n3844), .Z(n3843) );
  BUFFD0 U3838 ( .I(n3845), .Z(n3844) );
  BUFFD0 U3839 ( .I(n3846), .Z(n3845) );
  BUFFD0 U3840 ( .I(n3847), .Z(n3846) );
  BUFFD0 U3841 ( .I(n3848), .Z(n3847) );
  BUFFD0 U3842 ( .I(n3849), .Z(n3848) );
  BUFFD0 U3843 ( .I(n3850), .Z(n3849) );
  BUFFD0 U3844 ( .I(n3851), .Z(n3850) );
  BUFFD0 U3845 ( .I(n3852), .Z(n3851) );
  BUFFD0 U3846 ( .I(n3853), .Z(n3852) );
  BUFFD0 U3847 ( .I(n3854), .Z(n3853) );
  BUFFD0 U3848 ( .I(n3855), .Z(n3854) );
  BUFFD0 U3849 ( .I(n3856), .Z(n3855) );
  BUFFD0 U3850 ( .I(n3857), .Z(n3856) );
  BUFFD0 U3851 ( .I(n3858), .Z(n3857) );
  BUFFD0 U3852 ( .I(n3859), .Z(n3858) );
  BUFFD0 U3853 ( .I(n3860), .Z(n3859) );
  BUFFD0 U3854 ( .I(n3861), .Z(n3860) );
  BUFFD0 U3855 ( .I(n3862), .Z(n3861) );
  BUFFD0 U3856 ( .I(n3863), .Z(n3862) );
  BUFFD0 U3857 ( .I(n3864), .Z(n3863) );
  BUFFD0 U3858 ( .I(n3865), .Z(n3864) );
  BUFFD0 U3859 ( .I(n3866), .Z(n3865) );
  BUFFD0 U3860 ( .I(n3867), .Z(n3866) );
  BUFFD0 U3861 ( .I(n3868), .Z(n3867) );
  BUFFD0 U3862 ( .I(n3869), .Z(n3868) );
  BUFFD0 U3863 ( .I(n3870), .Z(n3869) );
  BUFFD0 U3864 ( .I(n3871), .Z(n3870) );
  BUFFD0 U3865 ( .I(n3872), .Z(n3871) );
  BUFFD0 U3866 ( .I(n3873), .Z(n3872) );
  BUFFD0 U3867 ( .I(n3874), .Z(n3873) );
  BUFFD0 U3868 ( .I(n3875), .Z(n3874) );
  BUFFD0 U3869 ( .I(n3876), .Z(n3875) );
  BUFFD0 U3870 ( .I(n3877), .Z(n3876) );
  BUFFD0 U3871 ( .I(n3878), .Z(n3877) );
  BUFFD0 U3872 ( .I(n3879), .Z(n3878) );
  BUFFD0 U3873 ( .I(n3881), .Z(n3879) );
  BUFFD0 U3874 ( .I(n2215), .Z(n3880) );
  BUFFD0 U3875 ( .I(n3882), .Z(n3881) );
  BUFFD0 U3876 ( .I(n3883), .Z(n3882) );
  BUFFD0 U3877 ( .I(n3884), .Z(n3883) );
  BUFFD0 U3878 ( .I(n3885), .Z(n3884) );
  BUFFD0 U3879 ( .I(n3886), .Z(n3885) );
  BUFFD0 U3880 ( .I(n3887), .Z(n3886) );
  BUFFD0 U3881 ( .I(n3888), .Z(n3887) );
  BUFFD0 U3882 ( .I(n3889), .Z(n3888) );
  BUFFD0 U3883 ( .I(n3890), .Z(n3889) );
  BUFFD0 U3884 ( .I(n3891), .Z(n3890) );
  BUFFD0 U3885 ( .I(n3892), .Z(n3891) );
  BUFFD0 U3886 ( .I(n3893), .Z(n3892) );
  BUFFD0 U3887 ( .I(n3894), .Z(n3893) );
  BUFFD0 U3888 ( .I(n3895), .Z(n3894) );
  BUFFD0 U3889 ( .I(n3896), .Z(n3895) );
  BUFFD0 U3890 ( .I(n3897), .Z(n3896) );
  BUFFD0 U3891 ( .I(n3898), .Z(n3897) );
  BUFFD0 U3892 ( .I(n3899), .Z(n3898) );
  BUFFD0 U3893 ( .I(n3900), .Z(n3899) );
  BUFFD0 U3894 ( .I(n3901), .Z(n3900) );
  BUFFD0 U3895 ( .I(n3902), .Z(n3901) );
  BUFFD0 U3896 ( .I(n3903), .Z(n3902) );
  BUFFD0 U3897 ( .I(n3904), .Z(n3903) );
  BUFFD0 U3898 ( .I(n3905), .Z(n3904) );
  BUFFD0 U3899 ( .I(n3906), .Z(n3905) );
  BUFFD0 U3900 ( .I(n3907), .Z(n3906) );
  BUFFD0 U3901 ( .I(n3908), .Z(n3907) );
  BUFFD0 U3902 ( .I(n3909), .Z(n3908) );
  BUFFD0 U3903 ( .I(n8731), .Z(n3909) );
  BUFFD0 U3904 ( .I(n8728), .Z(n3910) );
  BUFFD0 U3905 ( .I(n3912), .Z(n3911) );
  BUFFD0 U3906 ( .I(n3913), .Z(n3912) );
  BUFFD0 U3907 ( .I(n3914), .Z(n3913) );
  BUFFD0 U3908 ( .I(n3915), .Z(n3914) );
  BUFFD0 U3909 ( .I(n3916), .Z(n3915) );
  BUFFD0 U3910 ( .I(n3917), .Z(n3916) );
  BUFFD0 U3911 ( .I(n3918), .Z(n3917) );
  BUFFD0 U3912 ( .I(n3919), .Z(n3918) );
  BUFFD0 U3913 ( .I(n3920), .Z(n3919) );
  BUFFD0 U3914 ( .I(n3921), .Z(n3920) );
  BUFFD0 U3915 ( .I(n3922), .Z(n3921) );
  BUFFD0 U3916 ( .I(n3923), .Z(n3922) );
  BUFFD0 U3917 ( .I(n3924), .Z(n3923) );
  BUFFD0 U3918 ( .I(n3925), .Z(n3924) );
  BUFFD0 U3919 ( .I(n3926), .Z(n3925) );
  BUFFD0 U3920 ( .I(n3927), .Z(n3926) );
  BUFFD0 U3921 ( .I(n3928), .Z(n3927) );
  BUFFD0 U3922 ( .I(n3929), .Z(n3928) );
  BUFFD0 U3923 ( .I(n3930), .Z(n3929) );
  BUFFD0 U3924 ( .I(n3931), .Z(n3930) );
  BUFFD0 U3925 ( .I(n3932), .Z(n3931) );
  BUFFD0 U3926 ( .I(n3933), .Z(n3932) );
  BUFFD0 U3927 ( .I(n3934), .Z(n3933) );
  BUFFD0 U3928 ( .I(n3935), .Z(n3934) );
  BUFFD0 U3929 ( .I(n3936), .Z(n3935) );
  BUFFD0 U3930 ( .I(n3937), .Z(n3936) );
  BUFFD0 U3931 ( .I(n3938), .Z(n3937) );
  BUFFD0 U3932 ( .I(n3939), .Z(n3938) );
  BUFFD0 U3933 ( .I(n3940), .Z(n3939) );
  BUFFD0 U3934 ( .I(n3941), .Z(n3940) );
  BUFFD0 U3935 ( .I(n3942), .Z(n3941) );
  BUFFD0 U3936 ( .I(n3943), .Z(n3942) );
  BUFFD0 U3937 ( .I(n3944), .Z(n3943) );
  BUFFD0 U3938 ( .I(n3945), .Z(n3944) );
  BUFFD0 U3939 ( .I(n3946), .Z(n3945) );
  BUFFD0 U3940 ( .I(n3947), .Z(n3946) );
  BUFFD0 U3941 ( .I(n3948), .Z(n3947) );
  BUFFD0 U3942 ( .I(n3949), .Z(n3948) );
  BUFFD0 U3943 ( .I(n3950), .Z(n3949) );
  BUFFD0 U3944 ( .I(n3951), .Z(n3950) );
  BUFFD0 U3945 ( .I(n3952), .Z(n3951) );
  BUFFD0 U3946 ( .I(n3953), .Z(n3952) );
  BUFFD0 U3947 ( .I(n3954), .Z(n3953) );
  BUFFD0 U3948 ( .I(n3955), .Z(n3954) );
  BUFFD0 U3949 ( .I(n3956), .Z(n3955) );
  BUFFD0 U3950 ( .I(n3957), .Z(n3956) );
  BUFFD0 U3951 ( .I(n3958), .Z(n3957) );
  BUFFD0 U3952 ( .I(n3959), .Z(n3958) );
  BUFFD0 U3953 ( .I(n3960), .Z(n3959) );
  BUFFD0 U3954 ( .I(n3961), .Z(n3960) );
  BUFFD0 U3955 ( .I(n3962), .Z(n3961) );
  BUFFD0 U3956 ( .I(n3963), .Z(n3962) );
  BUFFD0 U3957 ( .I(n3964), .Z(n3963) );
  BUFFD0 U3958 ( .I(n3965), .Z(n3964) );
  BUFFD0 U3959 ( .I(n3966), .Z(n3965) );
  BUFFD0 U3960 ( .I(n3967), .Z(n3966) );
  BUFFD0 U3961 ( .I(n3968), .Z(n3967) );
  BUFFD0 U3962 ( .I(n3969), .Z(n3968) );
  BUFFD0 U3963 ( .I(n3970), .Z(n3969) );
  BUFFD0 U3964 ( .I(n3971), .Z(n3970) );
  BUFFD0 U3965 ( .I(n3972), .Z(n3971) );
  BUFFD0 U3966 ( .I(n3973), .Z(n3972) );
  BUFFD0 U3967 ( .I(n3974), .Z(n3973) );
  BUFFD0 U3968 ( .I(n3975), .Z(n3974) );
  BUFFD0 U3969 ( .I(n3976), .Z(n3975) );
  BUFFD0 U3970 ( .I(n3977), .Z(n3976) );
  BUFFD0 U3971 ( .I(n3978), .Z(n3977) );
  BUFFD0 U3972 ( .I(n3979), .Z(n3978) );
  BUFFD0 U3973 ( .I(n3980), .Z(n3979) );
  BUFFD0 U3974 ( .I(n3981), .Z(n3980) );
  BUFFD0 U3975 ( .I(n3982), .Z(n3981) );
  BUFFD0 U3976 ( .I(n3983), .Z(n3982) );
  BUFFD0 U3977 ( .I(n3984), .Z(n3983) );
  BUFFD0 U3978 ( .I(n3985), .Z(n3984) );
  BUFFD0 U3979 ( .I(n3986), .Z(n3985) );
  BUFFD0 U3980 ( .I(n3987), .Z(n3986) );
  BUFFD0 U3981 ( .I(n3988), .Z(n3987) );
  BUFFD0 U3982 ( .I(n3989), .Z(n3988) );
  BUFFD0 U3983 ( .I(n3990), .Z(n3989) );
  BUFFD0 U3984 ( .I(n3991), .Z(n3990) );
  BUFFD0 U3985 ( .I(n3992), .Z(n3991) );
  BUFFD0 U3986 ( .I(n3993), .Z(n3992) );
  BUFFD0 U3987 ( .I(n3994), .Z(n3993) );
  BUFFD0 U3988 ( .I(n3995), .Z(n3994) );
  BUFFD0 U3989 ( .I(n3996), .Z(n3995) );
  BUFFD0 U3990 ( .I(n3997), .Z(n3996) );
  BUFFD0 U3991 ( .I(n3998), .Z(n3997) );
  BUFFD0 U3992 ( .I(n3999), .Z(n3998) );
  BUFFD0 U3993 ( .I(n4000), .Z(n3999) );
  BUFFD0 U3994 ( .I(n4001), .Z(n4000) );
  BUFFD0 U3995 ( .I(n4002), .Z(n4001) );
  BUFFD0 U3996 ( .I(n4003), .Z(n4002) );
  BUFFD0 U3997 ( .I(n4004), .Z(n4003) );
  BUFFD0 U3998 ( .I(n4005), .Z(n4004) );
  BUFFD0 U3999 ( .I(n4006), .Z(n4005) );
  BUFFD0 U4000 ( .I(n4007), .Z(n4006) );
  BUFFD0 U4001 ( .I(n4008), .Z(n4007) );
  BUFFD0 U4002 ( .I(n4009), .Z(n4008) );
  BUFFD0 U4003 ( .I(n4010), .Z(n4009) );
  BUFFD0 U4004 ( .I(n4011), .Z(n4010) );
  BUFFD0 U4005 ( .I(n4012), .Z(n4011) );
  BUFFD0 U4006 ( .I(n4013), .Z(n4012) );
  BUFFD0 U4007 ( .I(n4014), .Z(n4013) );
  BUFFD0 U4008 ( .I(n4015), .Z(n4014) );
  BUFFD0 U4009 ( .I(n4016), .Z(n4015) );
  BUFFD0 U4010 ( .I(n4017), .Z(n4016) );
  BUFFD0 U4011 ( .I(n4018), .Z(n4017) );
  BUFFD0 U4012 ( .I(n4019), .Z(n4018) );
  BUFFD0 U4013 ( .I(n4020), .Z(n4019) );
  BUFFD0 U4014 ( .I(n4021), .Z(n4020) );
  BUFFD0 U4015 ( .I(n4022), .Z(n4021) );
  BUFFD0 U4016 ( .I(n4023), .Z(n4022) );
  BUFFD0 U4017 ( .I(n4024), .Z(n4023) );
  BUFFD0 U4018 ( .I(n4025), .Z(n4024) );
  BUFFD0 U4019 ( .I(n4026), .Z(n4025) );
  BUFFD0 U4020 ( .I(n4027), .Z(n4026) );
  BUFFD0 U4021 ( .I(n4028), .Z(n4027) );
  BUFFD0 U4022 ( .I(n4029), .Z(n4028) );
  BUFFD0 U4023 ( .I(n4030), .Z(n4029) );
  BUFFD0 U4024 ( .I(n4031), .Z(n4030) );
  BUFFD0 U4025 ( .I(n4032), .Z(n4031) );
  BUFFD0 U4026 ( .I(n4033), .Z(n4032) );
  BUFFD0 U4027 ( .I(n4034), .Z(n4033) );
  BUFFD0 U4028 ( .I(n4035), .Z(n4034) );
  BUFFD0 U4029 ( .I(n4036), .Z(n4035) );
  BUFFD0 U4030 ( .I(n4037), .Z(n4036) );
  BUFFD0 U4031 ( .I(n4038), .Z(n4037) );
  BUFFD0 U4032 ( .I(n4039), .Z(n4038) );
  BUFFD0 U4033 ( .I(n4040), .Z(n4039) );
  BUFFD0 U4034 ( .I(n4041), .Z(n4040) );
  BUFFD0 U4035 ( .I(n4042), .Z(n4041) );
  BUFFD0 U4036 ( .I(n4043), .Z(n4042) );
  BUFFD0 U4037 ( .I(n4044), .Z(n4043) );
  BUFFD0 U4038 ( .I(n4045), .Z(n4044) );
  BUFFD0 U4039 ( .I(n4046), .Z(n4045) );
  BUFFD0 U4040 ( .I(n4047), .Z(n4046) );
  BUFFD0 U4041 ( .I(n4048), .Z(n4047) );
  BUFFD0 U4042 ( .I(n4049), .Z(n4048) );
  BUFFD0 U4043 ( .I(n4050), .Z(n4049) );
  BUFFD0 U4044 ( .I(n4051), .Z(n4050) );
  BUFFD0 U4045 ( .I(n4052), .Z(n4051) );
  BUFFD0 U4046 ( .I(n4053), .Z(n4052) );
  BUFFD0 U4047 ( .I(n4054), .Z(n4053) );
  BUFFD0 U4048 ( .I(n4055), .Z(n4054) );
  BUFFD0 U4049 ( .I(n4056), .Z(n4055) );
  BUFFD0 U4050 ( .I(n4057), .Z(n4056) );
  BUFFD0 U4051 ( .I(n4058), .Z(n4057) );
  BUFFD0 U4052 ( .I(n4059), .Z(n4058) );
  BUFFD0 U4053 ( .I(n4060), .Z(n4059) );
  BUFFD0 U4054 ( .I(n4061), .Z(n4060) );
  BUFFD0 U4055 ( .I(n4062), .Z(n4061) );
  BUFFD0 U4056 ( .I(n4063), .Z(n4062) );
  BUFFD0 U4057 ( .I(n4064), .Z(n4063) );
  BUFFD0 U4058 ( .I(n4065), .Z(n4064) );
  BUFFD0 U4059 ( .I(n4066), .Z(n4065) );
  BUFFD0 U4060 ( .I(n4067), .Z(n4066) );
  BUFFD0 U4061 ( .I(n4068), .Z(n4067) );
  BUFFD0 U4062 ( .I(n4069), .Z(n4068) );
  BUFFD0 U4063 ( .I(n4070), .Z(n4069) );
  BUFFD0 U4064 ( .I(n4071), .Z(n4070) );
  BUFFD0 U4065 ( .I(n4072), .Z(n4071) );
  BUFFD0 U4066 ( .I(n4073), .Z(n4072) );
  BUFFD0 U4067 ( .I(n4074), .Z(n4073) );
  BUFFD0 U4068 ( .I(n4075), .Z(n4074) );
  BUFFD0 U4069 ( .I(n4076), .Z(n4075) );
  BUFFD0 U4070 ( .I(n4077), .Z(n4076) );
  BUFFD0 U4071 ( .I(n4078), .Z(n4077) );
  BUFFD0 U4072 ( .I(n4079), .Z(n4078) );
  BUFFD0 U4073 ( .I(n4080), .Z(n4079) );
  BUFFD0 U4074 ( .I(n4081), .Z(n4080) );
  BUFFD0 U4075 ( .I(n4082), .Z(n4081) );
  BUFFD0 U4076 ( .I(n4083), .Z(n4082) );
  BUFFD0 U4077 ( .I(n4084), .Z(n4083) );
  BUFFD0 U4078 ( .I(n4085), .Z(n4084) );
  BUFFD0 U4079 ( .I(n4086), .Z(n4085) );
  BUFFD0 U4080 ( .I(n4087), .Z(n4086) );
  BUFFD0 U4081 ( .I(n4088), .Z(n4087) );
  BUFFD0 U4082 ( .I(n8729), .Z(n4088) );
  BUFFD0 U4083 ( .I(n8726), .Z(n4089) );
  BUFFD0 U4084 ( .I(n4091), .Z(n4090) );
  BUFFD0 U4085 ( .I(n4092), .Z(n4091) );
  BUFFD0 U4086 ( .I(n4093), .Z(n4092) );
  BUFFD0 U4087 ( .I(n4094), .Z(n4093) );
  BUFFD0 U4088 ( .I(n4095), .Z(n4094) );
  BUFFD0 U4089 ( .I(n4096), .Z(n4095) );
  BUFFD0 U4090 ( .I(n4097), .Z(n4096) );
  BUFFD0 U4091 ( .I(n4098), .Z(n4097) );
  BUFFD0 U4092 ( .I(n4099), .Z(n4098) );
  BUFFD0 U4093 ( .I(n4100), .Z(n4099) );
  BUFFD0 U4094 ( .I(n4101), .Z(n4100) );
  BUFFD0 U4095 ( .I(n4102), .Z(n4101) );
  BUFFD0 U4096 ( .I(n4103), .Z(n4102) );
  BUFFD0 U4097 ( .I(n4104), .Z(n4103) );
  BUFFD0 U4098 ( .I(n4105), .Z(n4104) );
  BUFFD0 U4099 ( .I(n4106), .Z(n4105) );
  BUFFD0 U4100 ( .I(n4107), .Z(n4106) );
  BUFFD0 U4101 ( .I(n4108), .Z(n4107) );
  BUFFD0 U4102 ( .I(n4109), .Z(n4108) );
  BUFFD0 U4103 ( .I(n4110), .Z(n4109) );
  BUFFD0 U4104 ( .I(n4111), .Z(n4110) );
  BUFFD0 U4105 ( .I(n4112), .Z(n4111) );
  BUFFD0 U4106 ( .I(n4113), .Z(n4112) );
  BUFFD0 U4107 ( .I(n4114), .Z(n4113) );
  BUFFD0 U4108 ( .I(n4115), .Z(n4114) );
  BUFFD0 U4109 ( .I(n4116), .Z(n4115) );
  BUFFD0 U4110 ( .I(n4117), .Z(n4116) );
  BUFFD0 U4111 ( .I(n4118), .Z(n4117) );
  BUFFD0 U4112 ( .I(n4119), .Z(n4118) );
  BUFFD0 U4113 ( .I(n4120), .Z(n4119) );
  BUFFD0 U4114 ( .I(n4121), .Z(n4120) );
  BUFFD0 U4115 ( .I(n4122), .Z(n4121) );
  BUFFD0 U4116 ( .I(n4123), .Z(n4122) );
  BUFFD0 U4117 ( .I(n4124), .Z(n4123) );
  BUFFD0 U4118 ( .I(n4125), .Z(n4124) );
  BUFFD0 U4119 ( .I(n4126), .Z(n4125) );
  BUFFD0 U4120 ( .I(n4127), .Z(n4126) );
  BUFFD0 U4121 ( .I(n4128), .Z(n4127) );
  BUFFD0 U4122 ( .I(n4129), .Z(n4128) );
  BUFFD0 U4123 ( .I(n4130), .Z(n4129) );
  BUFFD0 U4124 ( .I(n4131), .Z(n4130) );
  BUFFD0 U4125 ( .I(n4132), .Z(n4131) );
  BUFFD0 U4126 ( .I(n4133), .Z(n4132) );
  BUFFD0 U4127 ( .I(n4134), .Z(n4133) );
  BUFFD0 U4128 ( .I(n4135), .Z(n4134) );
  BUFFD0 U4129 ( .I(n4136), .Z(n4135) );
  BUFFD0 U4130 ( .I(n4137), .Z(n4136) );
  BUFFD0 U4131 ( .I(n4138), .Z(n4137) );
  BUFFD0 U4132 ( .I(n4139), .Z(n4138) );
  BUFFD0 U4133 ( .I(n4140), .Z(n4139) );
  BUFFD0 U4134 ( .I(n4141), .Z(n4140) );
  BUFFD0 U4135 ( .I(n4142), .Z(n4141) );
  BUFFD0 U4136 ( .I(n4143), .Z(n4142) );
  BUFFD0 U4137 ( .I(n4144), .Z(n4143) );
  BUFFD0 U4138 ( .I(n4145), .Z(n4144) );
  BUFFD0 U4139 ( .I(n4146), .Z(n4145) );
  BUFFD0 U4140 ( .I(n4147), .Z(n4146) );
  BUFFD0 U4141 ( .I(n4148), .Z(n4147) );
  BUFFD0 U4142 ( .I(n4149), .Z(n4148) );
  BUFFD0 U4143 ( .I(n4150), .Z(n4149) );
  BUFFD0 U4144 ( .I(n4151), .Z(n4150) );
  BUFFD0 U4145 ( .I(n4152), .Z(n4151) );
  BUFFD0 U4146 ( .I(n4153), .Z(n4152) );
  BUFFD0 U4147 ( .I(n4154), .Z(n4153) );
  BUFFD0 U4148 ( .I(n4155), .Z(n4154) );
  BUFFD0 U4149 ( .I(n4156), .Z(n4155) );
  BUFFD0 U4150 ( .I(n4157), .Z(n4156) );
  BUFFD0 U4151 ( .I(n4158), .Z(n4157) );
  BUFFD0 U4152 ( .I(n4159), .Z(n4158) );
  BUFFD0 U4153 ( .I(n4160), .Z(n4159) );
  BUFFD0 U4154 ( .I(n4161), .Z(n4160) );
  BUFFD0 U4155 ( .I(n4162), .Z(n4161) );
  BUFFD0 U4156 ( .I(n4163), .Z(n4162) );
  BUFFD0 U4157 ( .I(n4164), .Z(n4163) );
  BUFFD0 U4158 ( .I(n4165), .Z(n4164) );
  BUFFD0 U4159 ( .I(n4166), .Z(n4165) );
  BUFFD0 U4160 ( .I(n4167), .Z(n4166) );
  BUFFD0 U4161 ( .I(n4168), .Z(n4167) );
  BUFFD0 U4162 ( .I(n4169), .Z(n4168) );
  BUFFD0 U4163 ( .I(n4170), .Z(n4169) );
  BUFFD0 U4164 ( .I(n4171), .Z(n4170) );
  BUFFD0 U4165 ( .I(n4172), .Z(n4171) );
  BUFFD0 U4166 ( .I(n4173), .Z(n4172) );
  BUFFD0 U4167 ( .I(n4174), .Z(n4173) );
  BUFFD0 U4168 ( .I(n4175), .Z(n4174) );
  BUFFD0 U4169 ( .I(n4176), .Z(n4175) );
  BUFFD0 U4170 ( .I(n4177), .Z(n4176) );
  BUFFD0 U4171 ( .I(n4178), .Z(n4177) );
  BUFFD0 U4172 ( .I(n4179), .Z(n4178) );
  BUFFD0 U4173 ( .I(n4180), .Z(n4179) );
  BUFFD0 U4174 ( .I(n4181), .Z(n4180) );
  BUFFD0 U4175 ( .I(n4182), .Z(n4181) );
  BUFFD0 U4176 ( .I(n4183), .Z(n4182) );
  BUFFD0 U4177 ( .I(n4184), .Z(n4183) );
  BUFFD0 U4178 ( .I(n4185), .Z(n4184) );
  BUFFD0 U4179 ( .I(n4186), .Z(n4185) );
  BUFFD0 U4180 ( .I(n4187), .Z(n4186) );
  BUFFD0 U4181 ( .I(n4188), .Z(n4187) );
  BUFFD0 U4182 ( .I(n4189), .Z(n4188) );
  BUFFD0 U4183 ( .I(n4190), .Z(n4189) );
  BUFFD0 U4184 ( .I(n4191), .Z(n4190) );
  BUFFD0 U4185 ( .I(n4192), .Z(n4191) );
  BUFFD0 U4186 ( .I(n4193), .Z(n4192) );
  BUFFD0 U4187 ( .I(n4194), .Z(n4193) );
  BUFFD0 U4188 ( .I(n4195), .Z(n4194) );
  BUFFD0 U4189 ( .I(n4196), .Z(n4195) );
  BUFFD0 U4190 ( .I(n4197), .Z(n4196) );
  BUFFD0 U4191 ( .I(n4198), .Z(n4197) );
  BUFFD0 U4192 ( .I(n4199), .Z(n4198) );
  BUFFD0 U4193 ( .I(n4200), .Z(n4199) );
  BUFFD0 U4194 ( .I(n4201), .Z(n4200) );
  BUFFD0 U4195 ( .I(n4202), .Z(n4201) );
  BUFFD0 U4196 ( .I(n4203), .Z(n4202) );
  BUFFD0 U4197 ( .I(n4204), .Z(n4203) );
  BUFFD0 U4198 ( .I(n4205), .Z(n4204) );
  BUFFD0 U4199 ( .I(n4206), .Z(n4205) );
  BUFFD0 U4200 ( .I(n4207), .Z(n4206) );
  BUFFD0 U4201 ( .I(n4208), .Z(n4207) );
  BUFFD0 U4202 ( .I(n4209), .Z(n4208) );
  BUFFD0 U4203 ( .I(n4210), .Z(n4209) );
  BUFFD0 U4204 ( .I(n4211), .Z(n4210) );
  BUFFD0 U4205 ( .I(n4212), .Z(n4211) );
  BUFFD0 U4206 ( .I(n4213), .Z(n4212) );
  BUFFD0 U4207 ( .I(n4214), .Z(n4213) );
  BUFFD0 U4208 ( .I(n4215), .Z(n4214) );
  BUFFD0 U4209 ( .I(n4216), .Z(n4215) );
  BUFFD0 U4210 ( .I(n4217), .Z(n4216) );
  BUFFD0 U4211 ( .I(n4218), .Z(n4217) );
  BUFFD0 U4212 ( .I(n4219), .Z(n4218) );
  BUFFD0 U4213 ( .I(n4220), .Z(n4219) );
  BUFFD0 U4214 ( .I(n4221), .Z(n4220) );
  BUFFD0 U4215 ( .I(n4222), .Z(n4221) );
  BUFFD0 U4216 ( .I(n4223), .Z(n4222) );
  BUFFD0 U4217 ( .I(n4224), .Z(n4223) );
  BUFFD0 U4218 ( .I(n4225), .Z(n4224) );
  BUFFD0 U4219 ( .I(n4226), .Z(n4225) );
  BUFFD0 U4220 ( .I(n4227), .Z(n4226) );
  BUFFD0 U4221 ( .I(n4228), .Z(n4227) );
  BUFFD0 U4222 ( .I(n4229), .Z(n4228) );
  BUFFD0 U4223 ( .I(n4230), .Z(n4229) );
  BUFFD0 U4224 ( .I(n4231), .Z(n4230) );
  BUFFD0 U4225 ( .I(n4232), .Z(n4231) );
  BUFFD0 U4226 ( .I(n4233), .Z(n4232) );
  BUFFD0 U4227 ( .I(n4234), .Z(n4233) );
  BUFFD0 U4228 ( .I(n4235), .Z(n4234) );
  BUFFD0 U4229 ( .I(n4236), .Z(n4235) );
  BUFFD0 U4230 ( .I(n4237), .Z(n4236) );
  BUFFD0 U4231 ( .I(n4238), .Z(n4237) );
  BUFFD0 U4232 ( .I(n4239), .Z(n4238) );
  BUFFD0 U4233 ( .I(n4240), .Z(n4239) );
  BUFFD0 U4234 ( .I(n4241), .Z(n4240) );
  BUFFD0 U4235 ( .I(n4242), .Z(n4241) );
  BUFFD0 U4236 ( .I(n4243), .Z(n4242) );
  BUFFD0 U4237 ( .I(n4244), .Z(n4243) );
  BUFFD0 U4238 ( .I(n4245), .Z(n4244) );
  BUFFD0 U4239 ( .I(n4246), .Z(n4245) );
  BUFFD0 U4240 ( .I(n4247), .Z(n4246) );
  BUFFD0 U4241 ( .I(n4248), .Z(n4247) );
  BUFFD0 U4242 ( .I(n4249), .Z(n4248) );
  BUFFD0 U4243 ( .I(n4250), .Z(n4249) );
  BUFFD0 U4244 ( .I(n4251), .Z(n4250) );
  BUFFD0 U4245 ( .I(n4252), .Z(n4251) );
  BUFFD0 U4246 ( .I(n4253), .Z(n4252) );
  BUFFD0 U4247 ( .I(n4254), .Z(n4253) );
  BUFFD0 U4248 ( .I(n4255), .Z(n4254) );
  BUFFD0 U4249 ( .I(n4256), .Z(n4255) );
  BUFFD0 U4250 ( .I(n4257), .Z(n4256) );
  BUFFD0 U4251 ( .I(n4258), .Z(n4257) );
  BUFFD0 U4252 ( .I(n4259), .Z(n4258) );
  BUFFD0 U4253 ( .I(n4260), .Z(n4259) );
  BUFFD0 U4254 ( .I(n4261), .Z(n4260) );
  BUFFD0 U4255 ( .I(n4262), .Z(n4261) );
  BUFFD0 U4256 ( .I(n4263), .Z(n4262) );
  BUFFD0 U4257 ( .I(n4264), .Z(n4263) );
  BUFFD0 U4258 ( .I(n4265), .Z(n4264) );
  BUFFD0 U4259 ( .I(n4266), .Z(n4265) );
  BUFFD0 U4260 ( .I(n4267), .Z(n4266) );
  BUFFD0 U4261 ( .I(n8727), .Z(n4267) );
  BUFFD0 U4262 ( .I(n8724), .Z(n4268) );
  BUFFD0 U4263 ( .I(n4270), .Z(n4269) );
  BUFFD0 U4264 ( .I(n4271), .Z(n4270) );
  BUFFD0 U4265 ( .I(n4272), .Z(n4271) );
  BUFFD0 U4266 ( .I(n4273), .Z(n4272) );
  BUFFD0 U4267 ( .I(n4274), .Z(n4273) );
  BUFFD0 U4268 ( .I(n4275), .Z(n4274) );
  BUFFD0 U4269 ( .I(n4276), .Z(n4275) );
  BUFFD0 U4270 ( .I(n4277), .Z(n4276) );
  BUFFD0 U4271 ( .I(n4278), .Z(n4277) );
  BUFFD0 U4272 ( .I(n4279), .Z(n4278) );
  BUFFD0 U4273 ( .I(n4280), .Z(n4279) );
  BUFFD0 U4274 ( .I(n4281), .Z(n4280) );
  BUFFD0 U4275 ( .I(n4282), .Z(n4281) );
  BUFFD0 U4276 ( .I(n4283), .Z(n4282) );
  BUFFD0 U4277 ( .I(n4284), .Z(n4283) );
  BUFFD0 U4278 ( .I(n4285), .Z(n4284) );
  BUFFD0 U4279 ( .I(n4286), .Z(n4285) );
  BUFFD0 U4280 ( .I(n4287), .Z(n4286) );
  BUFFD0 U4281 ( .I(n4288), .Z(n4287) );
  BUFFD0 U4282 ( .I(n4289), .Z(n4288) );
  BUFFD0 U4283 ( .I(n4290), .Z(n4289) );
  BUFFD0 U4284 ( .I(n4291), .Z(n4290) );
  BUFFD0 U4285 ( .I(n4292), .Z(n4291) );
  BUFFD0 U4286 ( .I(n4293), .Z(n4292) );
  BUFFD0 U4287 ( .I(n4294), .Z(n4293) );
  BUFFD0 U4288 ( .I(n4295), .Z(n4294) );
  BUFFD0 U4289 ( .I(n4296), .Z(n4295) );
  BUFFD0 U4290 ( .I(n4297), .Z(n4296) );
  BUFFD0 U4291 ( .I(n4298), .Z(n4297) );
  BUFFD0 U4292 ( .I(n4299), .Z(n4298) );
  BUFFD0 U4293 ( .I(n4300), .Z(n4299) );
  BUFFD0 U4294 ( .I(n4301), .Z(n4300) );
  BUFFD0 U4295 ( .I(n4302), .Z(n4301) );
  BUFFD0 U4296 ( .I(n4303), .Z(n4302) );
  BUFFD0 U4297 ( .I(n4304), .Z(n4303) );
  BUFFD0 U4298 ( .I(n4305), .Z(n4304) );
  BUFFD0 U4299 ( .I(n4306), .Z(n4305) );
  BUFFD0 U4300 ( .I(n4307), .Z(n4306) );
  BUFFD0 U4301 ( .I(n4308), .Z(n4307) );
  BUFFD0 U4302 ( .I(n4309), .Z(n4308) );
  BUFFD0 U4303 ( .I(n4310), .Z(n4309) );
  BUFFD0 U4304 ( .I(n4311), .Z(n4310) );
  BUFFD0 U4305 ( .I(n4312), .Z(n4311) );
  BUFFD0 U4306 ( .I(n4313), .Z(n4312) );
  BUFFD0 U4307 ( .I(n4314), .Z(n4313) );
  BUFFD0 U4308 ( .I(n4315), .Z(n4314) );
  BUFFD0 U4309 ( .I(n4316), .Z(n4315) );
  BUFFD0 U4310 ( .I(n4317), .Z(n4316) );
  BUFFD0 U4311 ( .I(n4318), .Z(n4317) );
  BUFFD0 U4312 ( .I(n4319), .Z(n4318) );
  BUFFD0 U4313 ( .I(n4320), .Z(n4319) );
  BUFFD0 U4314 ( .I(n4321), .Z(n4320) );
  BUFFD0 U4315 ( .I(n4322), .Z(n4321) );
  BUFFD0 U4316 ( .I(n4323), .Z(n4322) );
  BUFFD0 U4317 ( .I(n4324), .Z(n4323) );
  BUFFD0 U4318 ( .I(n4325), .Z(n4324) );
  BUFFD0 U4319 ( .I(n4326), .Z(n4325) );
  BUFFD0 U4320 ( .I(n4327), .Z(n4326) );
  BUFFD0 U4321 ( .I(n4328), .Z(n4327) );
  BUFFD0 U4322 ( .I(n4329), .Z(n4328) );
  BUFFD0 U4323 ( .I(n4330), .Z(n4329) );
  BUFFD0 U4324 ( .I(n4331), .Z(n4330) );
  BUFFD0 U4325 ( .I(n4332), .Z(n4331) );
  BUFFD0 U4326 ( .I(n4333), .Z(n4332) );
  BUFFD0 U4327 ( .I(n4334), .Z(n4333) );
  BUFFD0 U4328 ( .I(n4335), .Z(n4334) );
  BUFFD0 U4329 ( .I(n4336), .Z(n4335) );
  BUFFD0 U4330 ( .I(n4337), .Z(n4336) );
  BUFFD0 U4331 ( .I(n4338), .Z(n4337) );
  BUFFD0 U4332 ( .I(n4339), .Z(n4338) );
  BUFFD0 U4333 ( .I(n4340), .Z(n4339) );
  BUFFD0 U4334 ( .I(n4341), .Z(n4340) );
  BUFFD0 U4335 ( .I(n4342), .Z(n4341) );
  BUFFD0 U4336 ( .I(n4343), .Z(n4342) );
  BUFFD0 U4337 ( .I(n4344), .Z(n4343) );
  BUFFD0 U4338 ( .I(n4345), .Z(n4344) );
  BUFFD0 U4339 ( .I(n4346), .Z(n4345) );
  BUFFD0 U4340 ( .I(n4347), .Z(n4346) );
  BUFFD0 U4341 ( .I(n4348), .Z(n4347) );
  BUFFD0 U4342 ( .I(n4349), .Z(n4348) );
  BUFFD0 U4343 ( .I(n4350), .Z(n4349) );
  BUFFD0 U4344 ( .I(n4351), .Z(n4350) );
  BUFFD0 U4345 ( .I(n4352), .Z(n4351) );
  BUFFD0 U4346 ( .I(n4353), .Z(n4352) );
  BUFFD0 U4347 ( .I(n4354), .Z(n4353) );
  BUFFD0 U4348 ( .I(n4355), .Z(n4354) );
  BUFFD0 U4349 ( .I(n4356), .Z(n4355) );
  BUFFD0 U4350 ( .I(n4357), .Z(n4356) );
  BUFFD0 U4351 ( .I(n4358), .Z(n4357) );
  BUFFD0 U4352 ( .I(n4359), .Z(n4358) );
  BUFFD0 U4353 ( .I(n4360), .Z(n4359) );
  BUFFD0 U4354 ( .I(n4361), .Z(n4360) );
  BUFFD0 U4355 ( .I(n4362), .Z(n4361) );
  BUFFD0 U4356 ( .I(n4363), .Z(n4362) );
  BUFFD0 U4357 ( .I(n4364), .Z(n4363) );
  BUFFD0 U4358 ( .I(n4365), .Z(n4364) );
  BUFFD0 U4359 ( .I(n4366), .Z(n4365) );
  BUFFD0 U4360 ( .I(n4367), .Z(n4366) );
  BUFFD0 U4361 ( .I(n4368), .Z(n4367) );
  BUFFD0 U4362 ( .I(n4369), .Z(n4368) );
  BUFFD0 U4363 ( .I(n4370), .Z(n4369) );
  BUFFD0 U4364 ( .I(n4371), .Z(n4370) );
  BUFFD0 U4365 ( .I(n4372), .Z(n4371) );
  BUFFD0 U4366 ( .I(n4373), .Z(n4372) );
  BUFFD0 U4367 ( .I(n4374), .Z(n4373) );
  BUFFD0 U4368 ( .I(n4375), .Z(n4374) );
  BUFFD0 U4369 ( .I(n4376), .Z(n4375) );
  BUFFD0 U4370 ( .I(n4377), .Z(n4376) );
  BUFFD0 U4371 ( .I(n4378), .Z(n4377) );
  BUFFD0 U4372 ( .I(n4379), .Z(n4378) );
  BUFFD0 U4373 ( .I(n4380), .Z(n4379) );
  BUFFD0 U4374 ( .I(n4381), .Z(n4380) );
  BUFFD0 U4375 ( .I(n4382), .Z(n4381) );
  BUFFD0 U4376 ( .I(n4383), .Z(n4382) );
  BUFFD0 U4377 ( .I(n4384), .Z(n4383) );
  BUFFD0 U4378 ( .I(n4385), .Z(n4384) );
  BUFFD0 U4379 ( .I(n4386), .Z(n4385) );
  BUFFD0 U4380 ( .I(n4387), .Z(n4386) );
  BUFFD0 U4381 ( .I(n4388), .Z(n4387) );
  BUFFD0 U4382 ( .I(n4389), .Z(n4388) );
  BUFFD0 U4383 ( .I(n4390), .Z(n4389) );
  BUFFD0 U4384 ( .I(n4391), .Z(n4390) );
  BUFFD0 U4385 ( .I(n4392), .Z(n4391) );
  BUFFD0 U4386 ( .I(n4393), .Z(n4392) );
  BUFFD0 U4387 ( .I(n4394), .Z(n4393) );
  BUFFD0 U4388 ( .I(n4395), .Z(n4394) );
  BUFFD0 U4389 ( .I(n4396), .Z(n4395) );
  BUFFD0 U4390 ( .I(n4397), .Z(n4396) );
  BUFFD0 U4391 ( .I(n4398), .Z(n4397) );
  BUFFD0 U4392 ( .I(n4399), .Z(n4398) );
  BUFFD0 U4393 ( .I(n4400), .Z(n4399) );
  BUFFD0 U4394 ( .I(n4401), .Z(n4400) );
  BUFFD0 U4395 ( .I(n4402), .Z(n4401) );
  BUFFD0 U4396 ( .I(n4403), .Z(n4402) );
  BUFFD0 U4397 ( .I(n4404), .Z(n4403) );
  BUFFD0 U4398 ( .I(n4405), .Z(n4404) );
  BUFFD0 U4399 ( .I(n4406), .Z(n4405) );
  BUFFD0 U4400 ( .I(n4407), .Z(n4406) );
  BUFFD0 U4401 ( .I(n4408), .Z(n4407) );
  BUFFD0 U4402 ( .I(n4409), .Z(n4408) );
  BUFFD0 U4403 ( .I(n4410), .Z(n4409) );
  BUFFD0 U4404 ( .I(n4411), .Z(n4410) );
  BUFFD0 U4405 ( .I(n4412), .Z(n4411) );
  BUFFD0 U4406 ( .I(n4413), .Z(n4412) );
  BUFFD0 U4407 ( .I(n4414), .Z(n4413) );
  BUFFD0 U4408 ( .I(n4415), .Z(n4414) );
  BUFFD0 U4409 ( .I(n4416), .Z(n4415) );
  BUFFD0 U4410 ( .I(n4417), .Z(n4416) );
  BUFFD0 U4411 ( .I(n4418), .Z(n4417) );
  BUFFD0 U4412 ( .I(n4419), .Z(n4418) );
  BUFFD0 U4413 ( .I(n4420), .Z(n4419) );
  BUFFD0 U4414 ( .I(n4421), .Z(n4420) );
  BUFFD0 U4415 ( .I(n4422), .Z(n4421) );
  BUFFD0 U4416 ( .I(n4423), .Z(n4422) );
  BUFFD0 U4417 ( .I(n4424), .Z(n4423) );
  BUFFD0 U4418 ( .I(n4425), .Z(n4424) );
  BUFFD0 U4419 ( .I(n4426), .Z(n4425) );
  BUFFD0 U4420 ( .I(n4427), .Z(n4426) );
  BUFFD0 U4421 ( .I(n4428), .Z(n4427) );
  BUFFD0 U4422 ( .I(n4429), .Z(n4428) );
  BUFFD0 U4423 ( .I(n4430), .Z(n4429) );
  BUFFD0 U4424 ( .I(n4431), .Z(n4430) );
  BUFFD0 U4425 ( .I(n4432), .Z(n4431) );
  BUFFD0 U4426 ( .I(n4433), .Z(n4432) );
  BUFFD0 U4427 ( .I(n4434), .Z(n4433) );
  BUFFD0 U4428 ( .I(n4435), .Z(n4434) );
  BUFFD0 U4429 ( .I(n4436), .Z(n4435) );
  BUFFD0 U4430 ( .I(n4437), .Z(n4436) );
  BUFFD0 U4431 ( .I(n4438), .Z(n4437) );
  BUFFD0 U4432 ( .I(n4439), .Z(n4438) );
  BUFFD0 U4433 ( .I(n4440), .Z(n4439) );
  BUFFD0 U4434 ( .I(n4441), .Z(n4440) );
  BUFFD0 U4435 ( .I(n4442), .Z(n4441) );
  BUFFD0 U4436 ( .I(n4443), .Z(n4442) );
  BUFFD0 U4437 ( .I(n4444), .Z(n4443) );
  BUFFD0 U4438 ( .I(n8725), .Z(n4444) );
  BUFFD0 U4439 ( .I(n8721), .Z(n4445) );
  BUFFD0 U4440 ( .I(n4447), .Z(n4446) );
  BUFFD0 U4441 ( .I(n4448), .Z(n4447) );
  BUFFD0 U4442 ( .I(n4449), .Z(n4448) );
  BUFFD0 U4443 ( .I(n4450), .Z(n4449) );
  BUFFD0 U4444 ( .I(n4451), .Z(n4450) );
  BUFFD0 U4445 ( .I(n4452), .Z(n4451) );
  BUFFD0 U4446 ( .I(n4453), .Z(n4452) );
  BUFFD0 U4447 ( .I(n4454), .Z(n4453) );
  BUFFD0 U4448 ( .I(n4455), .Z(n4454) );
  BUFFD0 U4449 ( .I(n4456), .Z(n4455) );
  BUFFD0 U4450 ( .I(n4457), .Z(n4456) );
  BUFFD0 U4451 ( .I(n4458), .Z(n4457) );
  BUFFD0 U4452 ( .I(n4459), .Z(n4458) );
  BUFFD0 U4453 ( .I(n4460), .Z(n4459) );
  BUFFD0 U4454 ( .I(n4461), .Z(n4460) );
  BUFFD0 U4455 ( .I(n4462), .Z(n4461) );
  BUFFD0 U4456 ( .I(n4463), .Z(n4462) );
  BUFFD0 U4457 ( .I(n4464), .Z(n4463) );
  BUFFD0 U4458 ( .I(n4465), .Z(n4464) );
  BUFFD0 U4459 ( .I(n4466), .Z(n4465) );
  BUFFD0 U4460 ( .I(n4467), .Z(n4466) );
  BUFFD0 U4461 ( .I(n4468), .Z(n4467) );
  BUFFD0 U4462 ( .I(n4469), .Z(n4468) );
  BUFFD0 U4463 ( .I(n4470), .Z(n4469) );
  BUFFD0 U4464 ( .I(n4471), .Z(n4470) );
  BUFFD0 U4465 ( .I(n4472), .Z(n4471) );
  BUFFD0 U4466 ( .I(n4473), .Z(n4472) );
  BUFFD0 U4467 ( .I(n4474), .Z(n4473) );
  BUFFD0 U4468 ( .I(n4475), .Z(n4474) );
  BUFFD0 U4469 ( .I(n4476), .Z(n4475) );
  BUFFD0 U4470 ( .I(n4477), .Z(n4476) );
  BUFFD0 U4471 ( .I(n4478), .Z(n4477) );
  BUFFD0 U4472 ( .I(n4479), .Z(n4478) );
  BUFFD0 U4473 ( .I(n4480), .Z(n4479) );
  BUFFD0 U4474 ( .I(n4481), .Z(n4480) );
  BUFFD0 U4475 ( .I(n4482), .Z(n4481) );
  BUFFD0 U4476 ( .I(n4483), .Z(n4482) );
  BUFFD0 U4477 ( .I(n4484), .Z(n4483) );
  BUFFD0 U4478 ( .I(n4485), .Z(n4484) );
  BUFFD0 U4479 ( .I(n4486), .Z(n4485) );
  BUFFD0 U4480 ( .I(n4487), .Z(n4486) );
  BUFFD0 U4481 ( .I(n4488), .Z(n4487) );
  BUFFD0 U4482 ( .I(n4489), .Z(n4488) );
  BUFFD0 U4483 ( .I(n4490), .Z(n4489) );
  BUFFD0 U4484 ( .I(n4491), .Z(n4490) );
  BUFFD0 U4485 ( .I(n4492), .Z(n4491) );
  BUFFD0 U4486 ( .I(n4493), .Z(n4492) );
  BUFFD0 U4487 ( .I(n4494), .Z(n4493) );
  BUFFD0 U4488 ( .I(n4495), .Z(n4494) );
  BUFFD0 U4489 ( .I(n4496), .Z(n4495) );
  BUFFD0 U4490 ( .I(n4497), .Z(n4496) );
  BUFFD0 U4491 ( .I(n4498), .Z(n4497) );
  BUFFD0 U4492 ( .I(n4499), .Z(n4498) );
  BUFFD0 U4493 ( .I(n4500), .Z(n4499) );
  BUFFD0 U4494 ( .I(n4501), .Z(n4500) );
  BUFFD0 U4495 ( .I(n4502), .Z(n4501) );
  BUFFD0 U4496 ( .I(n4503), .Z(n4502) );
  BUFFD0 U4497 ( .I(n4504), .Z(n4503) );
  BUFFD0 U4498 ( .I(n4505), .Z(n4504) );
  BUFFD0 U4499 ( .I(n4506), .Z(n4505) );
  BUFFD0 U4500 ( .I(n4507), .Z(n4506) );
  BUFFD0 U4501 ( .I(n4508), .Z(n4507) );
  BUFFD0 U4502 ( .I(n4509), .Z(n4508) );
  BUFFD0 U4503 ( .I(n4510), .Z(n4509) );
  BUFFD0 U4504 ( .I(n4511), .Z(n4510) );
  BUFFD0 U4505 ( .I(n4512), .Z(n4511) );
  BUFFD0 U4506 ( .I(n4513), .Z(n4512) );
  BUFFD0 U4507 ( .I(n4514), .Z(n4513) );
  BUFFD0 U4508 ( .I(n4515), .Z(n4514) );
  BUFFD0 U4509 ( .I(n4516), .Z(n4515) );
  BUFFD0 U4510 ( .I(n4517), .Z(n4516) );
  BUFFD0 U4511 ( .I(n4518), .Z(n4517) );
  BUFFD0 U4512 ( .I(n4519), .Z(n4518) );
  BUFFD0 U4513 ( .I(n4520), .Z(n4519) );
  BUFFD0 U4514 ( .I(n4521), .Z(n4520) );
  BUFFD0 U4515 ( .I(n4522), .Z(n4521) );
  BUFFD0 U4516 ( .I(n4523), .Z(n4522) );
  BUFFD0 U4517 ( .I(n4524), .Z(n4523) );
  BUFFD0 U4518 ( .I(n4525), .Z(n4524) );
  BUFFD0 U4519 ( .I(n4526), .Z(n4525) );
  BUFFD0 U4520 ( .I(n4527), .Z(n4526) );
  BUFFD0 U4521 ( .I(n4528), .Z(n4527) );
  BUFFD0 U4522 ( .I(n4529), .Z(n4528) );
  BUFFD0 U4523 ( .I(n4530), .Z(n4529) );
  BUFFD0 U4524 ( .I(n4531), .Z(n4530) );
  BUFFD0 U4525 ( .I(n4532), .Z(n4531) );
  BUFFD0 U4526 ( .I(n4533), .Z(n4532) );
  BUFFD0 U4527 ( .I(n4534), .Z(n4533) );
  BUFFD0 U4528 ( .I(n4535), .Z(n4534) );
  BUFFD0 U4529 ( .I(n4536), .Z(n4535) );
  BUFFD0 U4530 ( .I(n4537), .Z(n4536) );
  BUFFD0 U4531 ( .I(n4538), .Z(n4537) );
  BUFFD0 U4532 ( .I(n4539), .Z(n4538) );
  BUFFD0 U4533 ( .I(n4540), .Z(n4539) );
  BUFFD0 U4534 ( .I(n4541), .Z(n4540) );
  BUFFD0 U4535 ( .I(n4542), .Z(n4541) );
  BUFFD0 U4536 ( .I(n4543), .Z(n4542) );
  BUFFD0 U4537 ( .I(n4544), .Z(n4543) );
  BUFFD0 U4538 ( .I(n4545), .Z(n4544) );
  BUFFD0 U4539 ( .I(n4546), .Z(n4545) );
  BUFFD0 U4540 ( .I(n4547), .Z(n4546) );
  BUFFD0 U4541 ( .I(n4548), .Z(n4547) );
  BUFFD0 U4542 ( .I(n4549), .Z(n4548) );
  BUFFD0 U4543 ( .I(n4550), .Z(n4549) );
  BUFFD0 U4544 ( .I(n4551), .Z(n4550) );
  BUFFD0 U4545 ( .I(n4552), .Z(n4551) );
  BUFFD0 U4546 ( .I(n4553), .Z(n4552) );
  BUFFD0 U4547 ( .I(n4554), .Z(n4553) );
  BUFFD0 U4548 ( .I(n4555), .Z(n4554) );
  BUFFD0 U4549 ( .I(n4556), .Z(n4555) );
  BUFFD0 U4550 ( .I(n4557), .Z(n4556) );
  BUFFD0 U4551 ( .I(n4558), .Z(n4557) );
  BUFFD0 U4552 ( .I(n4559), .Z(n4558) );
  BUFFD0 U4553 ( .I(n4560), .Z(n4559) );
  BUFFD0 U4554 ( .I(n4561), .Z(n4560) );
  BUFFD0 U4555 ( .I(n4562), .Z(n4561) );
  BUFFD0 U4556 ( .I(n4563), .Z(n4562) );
  BUFFD0 U4557 ( .I(n4564), .Z(n4563) );
  BUFFD0 U4558 ( .I(n4565), .Z(n4564) );
  BUFFD0 U4559 ( .I(n4566), .Z(n4565) );
  BUFFD0 U4560 ( .I(n4567), .Z(n4566) );
  BUFFD0 U4561 ( .I(n4568), .Z(n4567) );
  BUFFD0 U4562 ( .I(n4569), .Z(n4568) );
  BUFFD0 U4563 ( .I(n4570), .Z(n4569) );
  BUFFD0 U4564 ( .I(n4571), .Z(n4570) );
  BUFFD0 U4565 ( .I(n4572), .Z(n4571) );
  BUFFD0 U4566 ( .I(n4573), .Z(n4572) );
  BUFFD0 U4567 ( .I(n4574), .Z(n4573) );
  BUFFD0 U4568 ( .I(n4575), .Z(n4574) );
  BUFFD0 U4569 ( .I(n4576), .Z(n4575) );
  BUFFD0 U4570 ( .I(n4577), .Z(n4576) );
  BUFFD0 U4571 ( .I(n4578), .Z(n4577) );
  BUFFD0 U4572 ( .I(n4579), .Z(n4578) );
  BUFFD0 U4573 ( .I(n4580), .Z(n4579) );
  BUFFD0 U4574 ( .I(n4581), .Z(n4580) );
  BUFFD0 U4575 ( .I(n4582), .Z(n4581) );
  BUFFD0 U4576 ( .I(n4583), .Z(n4582) );
  BUFFD0 U4577 ( .I(n4584), .Z(n4583) );
  BUFFD0 U4578 ( .I(n4585), .Z(n4584) );
  BUFFD0 U4579 ( .I(n4586), .Z(n4585) );
  BUFFD0 U4580 ( .I(n4587), .Z(n4586) );
  BUFFD0 U4581 ( .I(n4588), .Z(n4587) );
  BUFFD0 U4582 ( .I(n4589), .Z(n4588) );
  BUFFD0 U4583 ( .I(n4590), .Z(n4589) );
  BUFFD0 U4584 ( .I(n4591), .Z(n4590) );
  BUFFD0 U4585 ( .I(n4592), .Z(n4591) );
  BUFFD0 U4586 ( .I(n4593), .Z(n4592) );
  BUFFD0 U4587 ( .I(n4594), .Z(n4593) );
  BUFFD0 U4588 ( .I(n4595), .Z(n4594) );
  BUFFD0 U4589 ( .I(n4596), .Z(n4595) );
  BUFFD0 U4590 ( .I(n4597), .Z(n4596) );
  BUFFD0 U4591 ( .I(n4598), .Z(n4597) );
  BUFFD0 U4592 ( .I(n4599), .Z(n4598) );
  BUFFD0 U4593 ( .I(n4600), .Z(n4599) );
  BUFFD0 U4594 ( .I(n4601), .Z(n4600) );
  BUFFD0 U4595 ( .I(n4602), .Z(n4601) );
  BUFFD0 U4596 ( .I(n4603), .Z(n4602) );
  BUFFD0 U4597 ( .I(n4604), .Z(n4603) );
  BUFFD0 U4598 ( .I(n4605), .Z(n4604) );
  BUFFD0 U4599 ( .I(n4606), .Z(n4605) );
  BUFFD0 U4600 ( .I(n4607), .Z(n4606) );
  BUFFD0 U4601 ( .I(n4608), .Z(n4607) );
  BUFFD0 U4602 ( .I(n4609), .Z(n4608) );
  BUFFD0 U4603 ( .I(n4610), .Z(n4609) );
  BUFFD0 U4604 ( .I(n4611), .Z(n4610) );
  BUFFD0 U4605 ( .I(n4612), .Z(n4611) );
  BUFFD0 U4606 ( .I(n4613), .Z(n4612) );
  BUFFD0 U4607 ( .I(n4614), .Z(n4613) );
  BUFFD0 U4608 ( .I(n4615), .Z(n4614) );
  BUFFD0 U4609 ( .I(n4616), .Z(n4615) );
  BUFFD0 U4610 ( .I(n4617), .Z(n4616) );
  BUFFD0 U4611 ( .I(n4618), .Z(n4617) );
  BUFFD0 U4612 ( .I(n4619), .Z(n4618) );
  BUFFD0 U4613 ( .I(n4620), .Z(n4619) );
  BUFFD0 U4614 ( .I(n4621), .Z(n4620) );
  BUFFD0 U4615 ( .I(n4622), .Z(n4621) );
  BUFFD0 U4616 ( .I(n4623), .Z(n4622) );
  BUFFD0 U4617 ( .I(n8722), .Z(n4623) );
  BUFFD0 U4618 ( .I(n8719), .Z(n4624) );
  BUFFD0 U4619 ( .I(n4626), .Z(n4625) );
  BUFFD0 U4620 ( .I(n4627), .Z(n4626) );
  BUFFD0 U4621 ( .I(n4628), .Z(n4627) );
  BUFFD0 U4622 ( .I(n4629), .Z(n4628) );
  BUFFD0 U4623 ( .I(n4630), .Z(n4629) );
  BUFFD0 U4624 ( .I(n4631), .Z(n4630) );
  BUFFD0 U4625 ( .I(n4632), .Z(n4631) );
  BUFFD0 U4626 ( .I(n4633), .Z(n4632) );
  BUFFD0 U4627 ( .I(n4634), .Z(n4633) );
  BUFFD0 U4628 ( .I(n4635), .Z(n4634) );
  BUFFD0 U4629 ( .I(n4636), .Z(n4635) );
  BUFFD0 U4630 ( .I(n4637), .Z(n4636) );
  BUFFD0 U4631 ( .I(n4638), .Z(n4637) );
  BUFFD0 U4632 ( .I(n4639), .Z(n4638) );
  BUFFD0 U4633 ( .I(n4640), .Z(n4639) );
  BUFFD0 U4634 ( .I(n4641), .Z(n4640) );
  BUFFD0 U4635 ( .I(n4642), .Z(n4641) );
  BUFFD0 U4636 ( .I(n4643), .Z(n4642) );
  BUFFD0 U4637 ( .I(n4644), .Z(n4643) );
  BUFFD0 U4638 ( .I(n4645), .Z(n4644) );
  BUFFD0 U4639 ( .I(n4646), .Z(n4645) );
  BUFFD0 U4640 ( .I(n4647), .Z(n4646) );
  BUFFD0 U4641 ( .I(n4648), .Z(n4647) );
  BUFFD0 U4642 ( .I(n4649), .Z(n4648) );
  BUFFD0 U4643 ( .I(n4650), .Z(n4649) );
  BUFFD0 U4644 ( .I(n4651), .Z(n4650) );
  BUFFD0 U4645 ( .I(n4652), .Z(n4651) );
  BUFFD0 U4646 ( .I(n4653), .Z(n4652) );
  BUFFD0 U4647 ( .I(n4654), .Z(n4653) );
  BUFFD0 U4648 ( .I(n4655), .Z(n4654) );
  BUFFD0 U4649 ( .I(n4656), .Z(n4655) );
  BUFFD0 U4650 ( .I(n4657), .Z(n4656) );
  BUFFD0 U4651 ( .I(n4658), .Z(n4657) );
  BUFFD0 U4652 ( .I(n4659), .Z(n4658) );
  BUFFD0 U4653 ( .I(n4660), .Z(n4659) );
  BUFFD0 U4654 ( .I(n4661), .Z(n4660) );
  BUFFD0 U4655 ( .I(n4662), .Z(n4661) );
  BUFFD0 U4656 ( .I(n4663), .Z(n4662) );
  BUFFD0 U4657 ( .I(n4664), .Z(n4663) );
  BUFFD0 U4658 ( .I(n4665), .Z(n4664) );
  BUFFD0 U4659 ( .I(n4666), .Z(n4665) );
  BUFFD0 U4660 ( .I(n4667), .Z(n4666) );
  BUFFD0 U4661 ( .I(n4668), .Z(n4667) );
  BUFFD0 U4662 ( .I(n4669), .Z(n4668) );
  BUFFD0 U4663 ( .I(n4670), .Z(n4669) );
  BUFFD0 U4664 ( .I(n4671), .Z(n4670) );
  BUFFD0 U4665 ( .I(n4672), .Z(n4671) );
  BUFFD0 U4666 ( .I(n4673), .Z(n4672) );
  BUFFD0 U4667 ( .I(n4674), .Z(n4673) );
  BUFFD0 U4668 ( .I(n4675), .Z(n4674) );
  BUFFD0 U4669 ( .I(n4676), .Z(n4675) );
  BUFFD0 U4670 ( .I(n4677), .Z(n4676) );
  BUFFD0 U4671 ( .I(n4678), .Z(n4677) );
  BUFFD0 U4672 ( .I(n4679), .Z(n4678) );
  BUFFD0 U4673 ( .I(n4680), .Z(n4679) );
  BUFFD0 U4674 ( .I(n4681), .Z(n4680) );
  BUFFD0 U4675 ( .I(n4682), .Z(n4681) );
  BUFFD0 U4676 ( .I(n4683), .Z(n4682) );
  BUFFD0 U4677 ( .I(n4684), .Z(n4683) );
  BUFFD0 U4678 ( .I(n4685), .Z(n4684) );
  BUFFD0 U4679 ( .I(n4686), .Z(n4685) );
  BUFFD0 U4680 ( .I(n4687), .Z(n4686) );
  BUFFD0 U4681 ( .I(n4688), .Z(n4687) );
  BUFFD0 U4682 ( .I(n4689), .Z(n4688) );
  BUFFD0 U4683 ( .I(n4690), .Z(n4689) );
  BUFFD0 U4684 ( .I(n4691), .Z(n4690) );
  BUFFD0 U4685 ( .I(n4692), .Z(n4691) );
  BUFFD0 U4686 ( .I(n4693), .Z(n4692) );
  BUFFD0 U4687 ( .I(n4694), .Z(n4693) );
  BUFFD0 U4688 ( .I(n4695), .Z(n4694) );
  BUFFD0 U4689 ( .I(n4696), .Z(n4695) );
  BUFFD0 U4690 ( .I(n4697), .Z(n4696) );
  BUFFD0 U4691 ( .I(n4698), .Z(n4697) );
  BUFFD0 U4692 ( .I(n4699), .Z(n4698) );
  BUFFD0 U4693 ( .I(n4700), .Z(n4699) );
  BUFFD0 U4694 ( .I(n4701), .Z(n4700) );
  BUFFD0 U4695 ( .I(n4702), .Z(n4701) );
  BUFFD0 U4696 ( .I(n4703), .Z(n4702) );
  BUFFD0 U4697 ( .I(n4704), .Z(n4703) );
  BUFFD0 U4698 ( .I(n4705), .Z(n4704) );
  BUFFD0 U4699 ( .I(n4706), .Z(n4705) );
  BUFFD0 U4700 ( .I(n4707), .Z(n4706) );
  BUFFD0 U4701 ( .I(n4708), .Z(n4707) );
  BUFFD0 U4702 ( .I(n4709), .Z(n4708) );
  BUFFD0 U4703 ( .I(n4710), .Z(n4709) );
  BUFFD0 U4704 ( .I(n4711), .Z(n4710) );
  BUFFD0 U4705 ( .I(n4712), .Z(n4711) );
  BUFFD0 U4706 ( .I(n4713), .Z(n4712) );
  BUFFD0 U4707 ( .I(n4714), .Z(n4713) );
  BUFFD0 U4708 ( .I(n4715), .Z(n4714) );
  BUFFD0 U4709 ( .I(n4716), .Z(n4715) );
  BUFFD0 U4710 ( .I(n4717), .Z(n4716) );
  BUFFD0 U4711 ( .I(n4718), .Z(n4717) );
  BUFFD0 U4712 ( .I(n4719), .Z(n4718) );
  BUFFD0 U4713 ( .I(n4720), .Z(n4719) );
  BUFFD0 U4714 ( .I(n4721), .Z(n4720) );
  BUFFD0 U4715 ( .I(n4722), .Z(n4721) );
  BUFFD0 U4716 ( .I(n4723), .Z(n4722) );
  BUFFD0 U4717 ( .I(n4724), .Z(n4723) );
  BUFFD0 U4718 ( .I(n4725), .Z(n4724) );
  BUFFD0 U4719 ( .I(n4726), .Z(n4725) );
  BUFFD0 U4720 ( .I(n4727), .Z(n4726) );
  BUFFD0 U4721 ( .I(n4728), .Z(n4727) );
  BUFFD0 U4722 ( .I(n4729), .Z(n4728) );
  BUFFD0 U4723 ( .I(n4730), .Z(n4729) );
  BUFFD0 U4724 ( .I(n4731), .Z(n4730) );
  BUFFD0 U4725 ( .I(n4732), .Z(n4731) );
  BUFFD0 U4726 ( .I(n4733), .Z(n4732) );
  BUFFD0 U4727 ( .I(n4734), .Z(n4733) );
  BUFFD0 U4728 ( .I(n4735), .Z(n4734) );
  BUFFD0 U4729 ( .I(n4736), .Z(n4735) );
  BUFFD0 U4730 ( .I(n4737), .Z(n4736) );
  BUFFD0 U4731 ( .I(n4738), .Z(n4737) );
  BUFFD0 U4732 ( .I(n4739), .Z(n4738) );
  BUFFD0 U4733 ( .I(n4740), .Z(n4739) );
  BUFFD0 U4734 ( .I(n4741), .Z(n4740) );
  BUFFD0 U4735 ( .I(n4742), .Z(n4741) );
  BUFFD0 U4736 ( .I(n4743), .Z(n4742) );
  BUFFD0 U4737 ( .I(n4744), .Z(n4743) );
  BUFFD0 U4738 ( .I(n4745), .Z(n4744) );
  BUFFD0 U4739 ( .I(n4746), .Z(n4745) );
  BUFFD0 U4740 ( .I(n4747), .Z(n4746) );
  BUFFD0 U4741 ( .I(n4748), .Z(n4747) );
  BUFFD0 U4742 ( .I(n4749), .Z(n4748) );
  BUFFD0 U4743 ( .I(n4750), .Z(n4749) );
  BUFFD0 U4744 ( .I(n4751), .Z(n4750) );
  BUFFD0 U4745 ( .I(n4752), .Z(n4751) );
  BUFFD0 U4746 ( .I(n4753), .Z(n4752) );
  BUFFD0 U4747 ( .I(n4754), .Z(n4753) );
  BUFFD0 U4748 ( .I(n4755), .Z(n4754) );
  BUFFD0 U4749 ( .I(n4756), .Z(n4755) );
  BUFFD0 U4750 ( .I(n4757), .Z(n4756) );
  BUFFD0 U4751 ( .I(n4758), .Z(n4757) );
  BUFFD0 U4752 ( .I(n4759), .Z(n4758) );
  BUFFD0 U4753 ( .I(n4760), .Z(n4759) );
  BUFFD0 U4754 ( .I(n4761), .Z(n4760) );
  BUFFD0 U4755 ( .I(n4762), .Z(n4761) );
  BUFFD0 U4756 ( .I(n4763), .Z(n4762) );
  BUFFD0 U4757 ( .I(n4764), .Z(n4763) );
  BUFFD0 U4758 ( .I(n4765), .Z(n4764) );
  BUFFD0 U4759 ( .I(n4766), .Z(n4765) );
  BUFFD0 U4760 ( .I(n4767), .Z(n4766) );
  BUFFD0 U4761 ( .I(n4768), .Z(n4767) );
  BUFFD0 U4762 ( .I(n4769), .Z(n4768) );
  BUFFD0 U4763 ( .I(n4770), .Z(n4769) );
  BUFFD0 U4764 ( .I(n4771), .Z(n4770) );
  BUFFD0 U4765 ( .I(n4772), .Z(n4771) );
  BUFFD0 U4766 ( .I(n4773), .Z(n4772) );
  BUFFD0 U4767 ( .I(n4774), .Z(n4773) );
  BUFFD0 U4768 ( .I(n4775), .Z(n4774) );
  BUFFD0 U4769 ( .I(n4776), .Z(n4775) );
  BUFFD0 U4770 ( .I(n4777), .Z(n4776) );
  BUFFD0 U4771 ( .I(n4778), .Z(n4777) );
  BUFFD0 U4772 ( .I(n4779), .Z(n4778) );
  BUFFD0 U4773 ( .I(n4780), .Z(n4779) );
  BUFFD0 U4774 ( .I(n4781), .Z(n4780) );
  BUFFD0 U4775 ( .I(n4782), .Z(n4781) );
  BUFFD0 U4776 ( .I(n4783), .Z(n4782) );
  BUFFD0 U4777 ( .I(n4784), .Z(n4783) );
  BUFFD0 U4778 ( .I(n4785), .Z(n4784) );
  BUFFD0 U4779 ( .I(n4786), .Z(n4785) );
  BUFFD0 U4780 ( .I(n4787), .Z(n4786) );
  BUFFD0 U4781 ( .I(n4788), .Z(n4787) );
  BUFFD0 U4782 ( .I(n4789), .Z(n4788) );
  BUFFD0 U4783 ( .I(n4790), .Z(n4789) );
  BUFFD0 U4784 ( .I(n4791), .Z(n4790) );
  BUFFD0 U4785 ( .I(n4792), .Z(n4791) );
  BUFFD0 U4786 ( .I(n4793), .Z(n4792) );
  BUFFD0 U4787 ( .I(n4794), .Z(n4793) );
  BUFFD0 U4788 ( .I(n4795), .Z(n4794) );
  BUFFD0 U4789 ( .I(n4796), .Z(n4795) );
  BUFFD0 U4790 ( .I(n4797), .Z(n4796) );
  BUFFD0 U4791 ( .I(n4798), .Z(n4797) );
  BUFFD0 U4792 ( .I(n4799), .Z(n4798) );
  BUFFD0 U4793 ( .I(n4800), .Z(n4799) );
  BUFFD0 U4794 ( .I(n4801), .Z(n4800) );
  BUFFD0 U4795 ( .I(n4802), .Z(n4801) );
  BUFFD0 U4796 ( .I(n8720), .Z(n4802) );
  BUFFD0 U4797 ( .I(n8717), .Z(n4803) );
  BUFFD0 U4798 ( .I(n4805), .Z(n4804) );
  BUFFD0 U4799 ( .I(n4806), .Z(n4805) );
  BUFFD0 U4800 ( .I(n4807), .Z(n4806) );
  BUFFD0 U4801 ( .I(n4808), .Z(n4807) );
  BUFFD0 U4802 ( .I(n4809), .Z(n4808) );
  BUFFD0 U4803 ( .I(n4810), .Z(n4809) );
  BUFFD0 U4804 ( .I(n4811), .Z(n4810) );
  BUFFD0 U4805 ( .I(n4812), .Z(n4811) );
  BUFFD0 U4806 ( .I(n4813), .Z(n4812) );
  BUFFD0 U4807 ( .I(n4814), .Z(n4813) );
  BUFFD0 U4808 ( .I(n4815), .Z(n4814) );
  BUFFD0 U4809 ( .I(n4816), .Z(n4815) );
  BUFFD0 U4810 ( .I(n4817), .Z(n4816) );
  BUFFD0 U4811 ( .I(n4818), .Z(n4817) );
  BUFFD0 U4812 ( .I(n4819), .Z(n4818) );
  BUFFD0 U4813 ( .I(n4820), .Z(n4819) );
  BUFFD0 U4814 ( .I(n4821), .Z(n4820) );
  BUFFD0 U4815 ( .I(n4822), .Z(n4821) );
  BUFFD0 U4816 ( .I(n4823), .Z(n4822) );
  BUFFD0 U4817 ( .I(n4824), .Z(n4823) );
  BUFFD0 U4818 ( .I(n4825), .Z(n4824) );
  BUFFD0 U4819 ( .I(n4826), .Z(n4825) );
  BUFFD0 U4820 ( .I(n4827), .Z(n4826) );
  BUFFD0 U4821 ( .I(n4828), .Z(n4827) );
  BUFFD0 U4822 ( .I(n4829), .Z(n4828) );
  BUFFD0 U4823 ( .I(n4830), .Z(n4829) );
  BUFFD0 U4824 ( .I(n4831), .Z(n4830) );
  BUFFD0 U4825 ( .I(n4832), .Z(n4831) );
  BUFFD0 U4826 ( .I(n4833), .Z(n4832) );
  BUFFD0 U4827 ( .I(n4834), .Z(n4833) );
  BUFFD0 U4828 ( .I(n4835), .Z(n4834) );
  BUFFD0 U4829 ( .I(n4836), .Z(n4835) );
  BUFFD0 U4830 ( .I(n4837), .Z(n4836) );
  BUFFD0 U4831 ( .I(n4838), .Z(n4837) );
  BUFFD0 U4832 ( .I(n4839), .Z(n4838) );
  BUFFD0 U4833 ( .I(n4840), .Z(n4839) );
  BUFFD0 U4834 ( .I(n4841), .Z(n4840) );
  BUFFD0 U4835 ( .I(n4842), .Z(n4841) );
  BUFFD0 U4836 ( .I(n4843), .Z(n4842) );
  BUFFD0 U4837 ( .I(n4844), .Z(n4843) );
  BUFFD0 U4838 ( .I(n4845), .Z(n4844) );
  BUFFD0 U4839 ( .I(n4846), .Z(n4845) );
  BUFFD0 U4840 ( .I(n4847), .Z(n4846) );
  BUFFD0 U4841 ( .I(n4848), .Z(n4847) );
  BUFFD0 U4842 ( .I(n4849), .Z(n4848) );
  BUFFD0 U4843 ( .I(n4850), .Z(n4849) );
  BUFFD0 U4844 ( .I(n4851), .Z(n4850) );
  BUFFD0 U4845 ( .I(n4852), .Z(n4851) );
  BUFFD0 U4846 ( .I(n4853), .Z(n4852) );
  BUFFD0 U4847 ( .I(n4854), .Z(n4853) );
  BUFFD0 U4848 ( .I(n4855), .Z(n4854) );
  BUFFD0 U4849 ( .I(n4856), .Z(n4855) );
  BUFFD0 U4850 ( .I(n4857), .Z(n4856) );
  BUFFD0 U4851 ( .I(n4858), .Z(n4857) );
  BUFFD0 U4852 ( .I(n4859), .Z(n4858) );
  BUFFD0 U4853 ( .I(n4860), .Z(n4859) );
  BUFFD0 U4854 ( .I(n4861), .Z(n4860) );
  BUFFD0 U4855 ( .I(n4862), .Z(n4861) );
  BUFFD0 U4856 ( .I(n4863), .Z(n4862) );
  BUFFD0 U4857 ( .I(n4864), .Z(n4863) );
  BUFFD0 U4858 ( .I(n4865), .Z(n4864) );
  BUFFD0 U4859 ( .I(n4866), .Z(n4865) );
  BUFFD0 U4860 ( .I(n4867), .Z(n4866) );
  BUFFD0 U4861 ( .I(n4868), .Z(n4867) );
  BUFFD0 U4862 ( .I(n4869), .Z(n4868) );
  BUFFD0 U4863 ( .I(n4870), .Z(n4869) );
  BUFFD0 U4864 ( .I(n4871), .Z(n4870) );
  BUFFD0 U4865 ( .I(n4872), .Z(n4871) );
  BUFFD0 U4866 ( .I(n4873), .Z(n4872) );
  BUFFD0 U4867 ( .I(n4874), .Z(n4873) );
  BUFFD0 U4868 ( .I(n4875), .Z(n4874) );
  BUFFD0 U4869 ( .I(n4876), .Z(n4875) );
  BUFFD0 U4870 ( .I(n4877), .Z(n4876) );
  BUFFD0 U4871 ( .I(n4878), .Z(n4877) );
  BUFFD0 U4872 ( .I(n4879), .Z(n4878) );
  BUFFD0 U4873 ( .I(n4880), .Z(n4879) );
  BUFFD0 U4874 ( .I(n4881), .Z(n4880) );
  BUFFD0 U4875 ( .I(n4882), .Z(n4881) );
  BUFFD0 U4876 ( .I(n4883), .Z(n4882) );
  BUFFD0 U4877 ( .I(n4884), .Z(n4883) );
  BUFFD0 U4878 ( .I(n4885), .Z(n4884) );
  BUFFD0 U4879 ( .I(n4886), .Z(n4885) );
  BUFFD0 U4880 ( .I(n4887), .Z(n4886) );
  BUFFD0 U4881 ( .I(n4888), .Z(n4887) );
  BUFFD0 U4882 ( .I(n4889), .Z(n4888) );
  BUFFD0 U4883 ( .I(n4890), .Z(n4889) );
  BUFFD0 U4884 ( .I(n4891), .Z(n4890) );
  BUFFD0 U4885 ( .I(n4892), .Z(n4891) );
  BUFFD0 U4886 ( .I(n4893), .Z(n4892) );
  BUFFD0 U4887 ( .I(n4894), .Z(n4893) );
  BUFFD0 U4888 ( .I(n4895), .Z(n4894) );
  BUFFD0 U4889 ( .I(n4896), .Z(n4895) );
  BUFFD0 U4890 ( .I(n4897), .Z(n4896) );
  BUFFD0 U4891 ( .I(n4898), .Z(n4897) );
  BUFFD0 U4892 ( .I(n4899), .Z(n4898) );
  BUFFD0 U4893 ( .I(n4900), .Z(n4899) );
  BUFFD0 U4894 ( .I(n4901), .Z(n4900) );
  BUFFD0 U4895 ( .I(n4902), .Z(n4901) );
  BUFFD0 U4896 ( .I(n4903), .Z(n4902) );
  BUFFD0 U4897 ( .I(n4904), .Z(n4903) );
  BUFFD0 U4898 ( .I(n4905), .Z(n4904) );
  BUFFD0 U4899 ( .I(n4906), .Z(n4905) );
  BUFFD0 U4900 ( .I(n4907), .Z(n4906) );
  BUFFD0 U4901 ( .I(n4908), .Z(n4907) );
  BUFFD0 U4902 ( .I(n4909), .Z(n4908) );
  BUFFD0 U4903 ( .I(n4910), .Z(n4909) );
  BUFFD0 U4904 ( .I(n4911), .Z(n4910) );
  BUFFD0 U4905 ( .I(n4912), .Z(n4911) );
  BUFFD0 U4906 ( .I(n4913), .Z(n4912) );
  BUFFD0 U4907 ( .I(n4914), .Z(n4913) );
  BUFFD0 U4908 ( .I(n4915), .Z(n4914) );
  BUFFD0 U4909 ( .I(n4916), .Z(n4915) );
  BUFFD0 U4910 ( .I(n4917), .Z(n4916) );
  BUFFD0 U4911 ( .I(n4918), .Z(n4917) );
  BUFFD0 U4912 ( .I(n4919), .Z(n4918) );
  BUFFD0 U4913 ( .I(n4920), .Z(n4919) );
  BUFFD0 U4914 ( .I(n4921), .Z(n4920) );
  BUFFD0 U4915 ( .I(n4922), .Z(n4921) );
  BUFFD0 U4916 ( .I(n4923), .Z(n4922) );
  BUFFD0 U4917 ( .I(n4924), .Z(n4923) );
  BUFFD0 U4918 ( .I(n4925), .Z(n4924) );
  BUFFD0 U4919 ( .I(n4926), .Z(n4925) );
  BUFFD0 U4920 ( .I(n4927), .Z(n4926) );
  BUFFD0 U4921 ( .I(n4928), .Z(n4927) );
  BUFFD0 U4922 ( .I(n4929), .Z(n4928) );
  BUFFD0 U4923 ( .I(n4930), .Z(n4929) );
  BUFFD0 U4924 ( .I(n4931), .Z(n4930) );
  BUFFD0 U4925 ( .I(n4932), .Z(n4931) );
  BUFFD0 U4926 ( .I(n4933), .Z(n4932) );
  BUFFD0 U4927 ( .I(n4934), .Z(n4933) );
  BUFFD0 U4928 ( .I(n4935), .Z(n4934) );
  BUFFD0 U4929 ( .I(n4936), .Z(n4935) );
  BUFFD0 U4930 ( .I(n4937), .Z(n4936) );
  BUFFD0 U4931 ( .I(n4938), .Z(n4937) );
  BUFFD0 U4932 ( .I(n4939), .Z(n4938) );
  BUFFD0 U4933 ( .I(n4940), .Z(n4939) );
  BUFFD0 U4934 ( .I(n4941), .Z(n4940) );
  BUFFD0 U4935 ( .I(n4942), .Z(n4941) );
  BUFFD0 U4936 ( .I(n4943), .Z(n4942) );
  BUFFD0 U4937 ( .I(n4944), .Z(n4943) );
  BUFFD0 U4938 ( .I(n4945), .Z(n4944) );
  BUFFD0 U4939 ( .I(n4946), .Z(n4945) );
  BUFFD0 U4940 ( .I(n4947), .Z(n4946) );
  BUFFD0 U4941 ( .I(n4948), .Z(n4947) );
  BUFFD0 U4942 ( .I(n4949), .Z(n4948) );
  BUFFD0 U4943 ( .I(n4950), .Z(n4949) );
  BUFFD0 U4944 ( .I(n4951), .Z(n4950) );
  BUFFD0 U4945 ( .I(n4952), .Z(n4951) );
  BUFFD0 U4946 ( .I(n4953), .Z(n4952) );
  BUFFD0 U4947 ( .I(n4954), .Z(n4953) );
  BUFFD0 U4948 ( .I(n4955), .Z(n4954) );
  BUFFD0 U4949 ( .I(n4956), .Z(n4955) );
  BUFFD0 U4950 ( .I(n4957), .Z(n4956) );
  BUFFD0 U4951 ( .I(n4958), .Z(n4957) );
  BUFFD0 U4952 ( .I(n4959), .Z(n4958) );
  BUFFD0 U4953 ( .I(n4960), .Z(n4959) );
  BUFFD0 U4954 ( .I(n4961), .Z(n4960) );
  BUFFD0 U4955 ( .I(n4962), .Z(n4961) );
  BUFFD0 U4956 ( .I(n4963), .Z(n4962) );
  BUFFD0 U4957 ( .I(n4964), .Z(n4963) );
  BUFFD0 U4958 ( .I(n4965), .Z(n4964) );
  BUFFD0 U4959 ( .I(n4966), .Z(n4965) );
  BUFFD0 U4960 ( .I(n4967), .Z(n4966) );
  BUFFD0 U4961 ( .I(n4968), .Z(n4967) );
  BUFFD0 U4962 ( .I(n4969), .Z(n4968) );
  BUFFD0 U4963 ( .I(n4970), .Z(n4969) );
  BUFFD0 U4964 ( .I(n4971), .Z(n4970) );
  BUFFD0 U4965 ( .I(n4972), .Z(n4971) );
  BUFFD0 U4966 ( .I(n4973), .Z(n4972) );
  BUFFD0 U4967 ( .I(n4974), .Z(n4973) );
  BUFFD0 U4968 ( .I(n4975), .Z(n4974) );
  BUFFD0 U4969 ( .I(n4976), .Z(n4975) );
  BUFFD0 U4970 ( .I(n4977), .Z(n4976) );
  BUFFD0 U4971 ( .I(n4978), .Z(n4977) );
  BUFFD0 U4972 ( .I(n4979), .Z(n4978) );
  BUFFD0 U4973 ( .I(n8718), .Z(n4979) );
  BUFFD0 U4974 ( .I(n4981), .Z(n4980) );
  BUFFD0 U4975 ( .I(n4982), .Z(n4981) );
  BUFFD0 U4976 ( .I(n4983), .Z(n4982) );
  BUFFD0 U4977 ( .I(n4984), .Z(n4983) );
  BUFFD0 U4978 ( .I(n4985), .Z(n4984) );
  BUFFD0 U4979 ( .I(n4986), .Z(n4985) );
  BUFFD0 U4980 ( .I(n4987), .Z(n4986) );
  BUFFD0 U4981 ( .I(n4988), .Z(n4987) );
  BUFFD0 U4982 ( .I(n4989), .Z(n4988) );
  BUFFD0 U4983 ( .I(n4990), .Z(n4989) );
  BUFFD0 U4984 ( .I(n4991), .Z(n4990) );
  BUFFD0 U4985 ( .I(n4992), .Z(n4991) );
  BUFFD0 U4986 ( .I(n4993), .Z(n4992) );
  BUFFD0 U4987 ( .I(n4994), .Z(n4993) );
  BUFFD0 U4988 ( .I(n4995), .Z(n4994) );
  BUFFD0 U4989 ( .I(n4996), .Z(n4995) );
  BUFFD0 U4990 ( .I(n4997), .Z(n4996) );
  BUFFD0 U4991 ( .I(n4998), .Z(n4997) );
  BUFFD0 U4992 ( .I(n4999), .Z(n4998) );
  BUFFD0 U4993 ( .I(n5000), .Z(n4999) );
  BUFFD0 U4994 ( .I(n5001), .Z(n5000) );
  BUFFD0 U4995 ( .I(n5002), .Z(n5001) );
  BUFFD0 U4996 ( .I(n5003), .Z(n5002) );
  BUFFD0 U4997 ( .I(n5004), .Z(n5003) );
  BUFFD0 U4998 ( .I(n5005), .Z(n5004) );
  BUFFD0 U4999 ( .I(n5006), .Z(n5005) );
  BUFFD0 U5000 ( .I(n5007), .Z(n5006) );
  BUFFD0 U5001 ( .I(n5008), .Z(n5007) );
  BUFFD0 U5002 ( .I(n5009), .Z(n5008) );
  BUFFD0 U5003 ( .I(n5010), .Z(n5009) );
  BUFFD0 U5004 ( .I(n5011), .Z(n5010) );
  BUFFD0 U5005 ( .I(n5012), .Z(n5011) );
  BUFFD0 U5006 ( .I(n5013), .Z(n5012) );
  BUFFD0 U5007 ( .I(n5014), .Z(n5013) );
  BUFFD0 U5008 ( .I(n5015), .Z(n5014) );
  BUFFD0 U5009 ( .I(n5016), .Z(n5015) );
  BUFFD0 U5010 ( .I(n5017), .Z(n5016) );
  BUFFD0 U5011 ( .I(n5018), .Z(n5017) );
  BUFFD0 U5012 ( .I(n5019), .Z(n5018) );
  BUFFD0 U5013 ( .I(n5020), .Z(n5019) );
  BUFFD0 U5014 ( .I(n5021), .Z(n5020) );
  BUFFD0 U5015 ( .I(n5022), .Z(n5021) );
  BUFFD0 U5016 ( .I(n5023), .Z(n5022) );
  BUFFD0 U5017 ( .I(n5024), .Z(n5023) );
  BUFFD0 U5018 ( .I(n5025), .Z(n5024) );
  BUFFD0 U5019 ( .I(n5026), .Z(n5025) );
  BUFFD0 U5020 ( .I(n5027), .Z(n5026) );
  BUFFD0 U5021 ( .I(n5028), .Z(n5027) );
  BUFFD0 U5022 ( .I(n5029), .Z(n5028) );
  BUFFD0 U5023 ( .I(n5030), .Z(n5029) );
  BUFFD0 U5024 ( .I(n5031), .Z(n5030) );
  BUFFD0 U5025 ( .I(n5032), .Z(n5031) );
  BUFFD0 U5026 ( .I(n5033), .Z(n5032) );
  BUFFD0 U5027 ( .I(n5034), .Z(n5033) );
  BUFFD0 U5028 ( .I(n5035), .Z(n5034) );
  BUFFD0 U5029 ( .I(n5036), .Z(n5035) );
  BUFFD0 U5030 ( .I(n5037), .Z(n5036) );
  BUFFD0 U5031 ( .I(n5038), .Z(n5037) );
  BUFFD0 U5032 ( .I(n5039), .Z(n5038) );
  BUFFD0 U5033 ( .I(n5040), .Z(n5039) );
  BUFFD0 U5034 ( .I(n5041), .Z(n5040) );
  BUFFD0 U5035 ( .I(n5042), .Z(n5041) );
  BUFFD0 U5036 ( .I(n5043), .Z(n5042) );
  BUFFD0 U5037 ( .I(n5044), .Z(n5043) );
  BUFFD0 U5038 ( .I(n5045), .Z(n5044) );
  BUFFD0 U5039 ( .I(n5046), .Z(n5045) );
  BUFFD0 U5040 ( .I(n5047), .Z(n5046) );
  BUFFD0 U5041 ( .I(n5048), .Z(n5047) );
  BUFFD0 U5042 ( .I(n5049), .Z(n5048) );
  BUFFD0 U5043 ( .I(n5050), .Z(n5049) );
  BUFFD0 U5044 ( .I(n5051), .Z(n5050) );
  BUFFD0 U5045 ( .I(n5052), .Z(n5051) );
  BUFFD0 U5046 ( .I(n5053), .Z(n5052) );
  BUFFD0 U5047 ( .I(n5054), .Z(n5053) );
  BUFFD0 U5048 ( .I(n5055), .Z(n5054) );
  BUFFD0 U5049 ( .I(n5056), .Z(n5055) );
  BUFFD0 U5050 ( .I(n5057), .Z(n5056) );
  BUFFD0 U5051 ( .I(n5058), .Z(n5057) );
  BUFFD0 U5052 ( .I(n5059), .Z(n5058) );
  BUFFD0 U5053 ( .I(n5060), .Z(n5059) );
  BUFFD0 U5054 ( .I(n5061), .Z(n5060) );
  BUFFD0 U5055 ( .I(n5062), .Z(n5061) );
  BUFFD0 U5056 ( .I(n5063), .Z(n5062) );
  BUFFD0 U5057 ( .I(n5064), .Z(n5063) );
  BUFFD0 U5058 ( .I(n5065), .Z(n5064) );
  BUFFD0 U5059 ( .I(n5066), .Z(n5065) );
  BUFFD0 U5060 ( .I(n5067), .Z(n5066) );
  BUFFD0 U5061 ( .I(n5068), .Z(n5067) );
  BUFFD0 U5062 ( .I(n5069), .Z(n5068) );
  BUFFD0 U5063 ( .I(n5070), .Z(n5069) );
  BUFFD0 U5064 ( .I(n5071), .Z(n5070) );
  BUFFD0 U5065 ( .I(n5072), .Z(n5071) );
  BUFFD0 U5066 ( .I(n5073), .Z(n5072) );
  BUFFD0 U5067 ( .I(n5074), .Z(n5073) );
  BUFFD0 U5068 ( .I(n5075), .Z(n5074) );
  BUFFD0 U5069 ( .I(n5076), .Z(n5075) );
  BUFFD0 U5070 ( .I(n5077), .Z(n5076) );
  BUFFD0 U5071 ( .I(n5078), .Z(n5077) );
  BUFFD0 U5072 ( .I(n5079), .Z(n5078) );
  BUFFD0 U5073 ( .I(n5080), .Z(n5079) );
  BUFFD0 U5074 ( .I(n5081), .Z(n5080) );
  BUFFD0 U5075 ( .I(n5082), .Z(n5081) );
  BUFFD0 U5076 ( .I(n5083), .Z(n5082) );
  BUFFD0 U5077 ( .I(n5084), .Z(n5083) );
  BUFFD0 U5078 ( .I(n5085), .Z(n5084) );
  BUFFD0 U5079 ( .I(n5086), .Z(n5085) );
  BUFFD0 U5080 ( .I(n5087), .Z(n5086) );
  BUFFD0 U5081 ( .I(n5088), .Z(n5087) );
  BUFFD0 U5082 ( .I(n5089), .Z(n5088) );
  BUFFD0 U5083 ( .I(n5090), .Z(n5089) );
  BUFFD0 U5084 ( .I(n5091), .Z(n5090) );
  BUFFD0 U5085 ( .I(n5092), .Z(n5091) );
  BUFFD0 U5086 ( .I(n5093), .Z(n5092) );
  BUFFD0 U5087 ( .I(n5094), .Z(n5093) );
  BUFFD0 U5088 ( .I(n5095), .Z(n5094) );
  BUFFD0 U5089 ( .I(n5096), .Z(n5095) );
  BUFFD0 U5090 ( .I(n5097), .Z(n5096) );
  BUFFD0 U5091 ( .I(n5098), .Z(n5097) );
  BUFFD0 U5092 ( .I(n5099), .Z(n5098) );
  BUFFD0 U5093 ( .I(n5100), .Z(n5099) );
  BUFFD0 U5094 ( .I(n5101), .Z(n5100) );
  BUFFD0 U5095 ( .I(n5102), .Z(n5101) );
  BUFFD0 U5096 ( .I(n5103), .Z(n5102) );
  BUFFD0 U5097 ( .I(n5104), .Z(n5103) );
  BUFFD0 U5098 ( .I(n5105), .Z(n5104) );
  BUFFD0 U5099 ( .I(n5106), .Z(n5105) );
  BUFFD0 U5100 ( .I(n5107), .Z(n5106) );
  BUFFD0 U5101 ( .I(n5108), .Z(n5107) );
  BUFFD0 U5102 ( .I(n5109), .Z(n5108) );
  BUFFD0 U5103 ( .I(n5110), .Z(n5109) );
  BUFFD0 U5104 ( .I(n5111), .Z(n5110) );
  BUFFD0 U5105 ( .I(n5112), .Z(n5111) );
  BUFFD0 U5106 ( .I(n5113), .Z(n5112) );
  BUFFD0 U5107 ( .I(n5114), .Z(n5113) );
  BUFFD0 U5108 ( .I(n5115), .Z(n5114) );
  BUFFD0 U5109 ( .I(n5116), .Z(n5115) );
  BUFFD0 U5110 ( .I(n5117), .Z(n5116) );
  BUFFD0 U5111 ( .I(n5118), .Z(n5117) );
  BUFFD0 U5112 ( .I(n5119), .Z(n5118) );
  BUFFD0 U5113 ( .I(n5120), .Z(n5119) );
  BUFFD0 U5114 ( .I(n5121), .Z(n5120) );
  BUFFD0 U5115 ( .I(n5123), .Z(n5121) );
  BUFFD0 U5116 ( .I(n2216), .Z(n5122) );
  BUFFD0 U5117 ( .I(n5124), .Z(n5123) );
  BUFFD0 U5118 ( .I(n5125), .Z(n5124) );
  BUFFD0 U5119 ( .I(n5126), .Z(n5125) );
  BUFFD0 U5120 ( .I(n5127), .Z(n5126) );
  BUFFD0 U5121 ( .I(n5128), .Z(n5127) );
  BUFFD0 U5122 ( .I(n5129), .Z(n5128) );
  BUFFD0 U5123 ( .I(n5130), .Z(n5129) );
  BUFFD0 U5124 ( .I(n5131), .Z(n5130) );
  BUFFD0 U5125 ( .I(n5132), .Z(n5131) );
  BUFFD0 U5126 ( .I(n5133), .Z(n5132) );
  BUFFD0 U5127 ( .I(n5134), .Z(n5133) );
  BUFFD0 U5128 ( .I(n5135), .Z(n5134) );
  BUFFD0 U5129 ( .I(n5136), .Z(n5135) );
  BUFFD0 U5130 ( .I(n5137), .Z(n5136) );
  BUFFD0 U5131 ( .I(n5138), .Z(n5137) );
  BUFFD0 U5132 ( .I(n5139), .Z(n5138) );
  BUFFD0 U5133 ( .I(n5140), .Z(n5139) );
  BUFFD0 U5134 ( .I(n5141), .Z(n5140) );
  BUFFD0 U5135 ( .I(n5142), .Z(n5141) );
  BUFFD0 U5136 ( .I(n5143), .Z(n5142) );
  BUFFD0 U5137 ( .I(n5144), .Z(n5143) );
  BUFFD0 U5138 ( .I(n5145), .Z(n5144) );
  BUFFD0 U5139 ( .I(n5146), .Z(n5145) );
  BUFFD0 U5140 ( .I(n5147), .Z(n5146) );
  BUFFD0 U5141 ( .I(n5148), .Z(n5147) );
  BUFFD0 U5142 ( .I(n5149), .Z(n5148) );
  BUFFD0 U5143 ( .I(n5150), .Z(n5149) );
  BUFFD0 U5144 ( .I(n5151), .Z(n5150) );
  BUFFD0 U5145 ( .I(n5152), .Z(n5151) );
  BUFFD0 U5146 ( .I(n5153), .Z(n5152) );
  BUFFD0 U5147 ( .I(n8715), .Z(n5153) );
  BUFFD0 U5148 ( .I(n8712), .Z(n5154) );
  BUFFD0 U5149 ( .I(n5156), .Z(n5155) );
  BUFFD0 U5150 ( .I(n5157), .Z(n5156) );
  BUFFD0 U5151 ( .I(n5158), .Z(n5157) );
  BUFFD0 U5152 ( .I(n5159), .Z(n5158) );
  BUFFD0 U5153 ( .I(n5160), .Z(n5159) );
  BUFFD0 U5154 ( .I(n5161), .Z(n5160) );
  BUFFD0 U5155 ( .I(n5162), .Z(n5161) );
  BUFFD0 U5156 ( .I(n5163), .Z(n5162) );
  BUFFD0 U5157 ( .I(n5164), .Z(n5163) );
  BUFFD0 U5158 ( .I(n5165), .Z(n5164) );
  BUFFD0 U5159 ( .I(n5166), .Z(n5165) );
  BUFFD0 U5160 ( .I(n5167), .Z(n5166) );
  BUFFD0 U5161 ( .I(n5168), .Z(n5167) );
  BUFFD0 U5162 ( .I(n5169), .Z(n5168) );
  BUFFD0 U5163 ( .I(n5170), .Z(n5169) );
  BUFFD0 U5164 ( .I(n5171), .Z(n5170) );
  BUFFD0 U5165 ( .I(n5172), .Z(n5171) );
  BUFFD0 U5166 ( .I(n5173), .Z(n5172) );
  BUFFD0 U5167 ( .I(n5174), .Z(n5173) );
  BUFFD0 U5168 ( .I(n5175), .Z(n5174) );
  BUFFD0 U5169 ( .I(n5176), .Z(n5175) );
  BUFFD0 U5170 ( .I(n5177), .Z(n5176) );
  BUFFD0 U5171 ( .I(n5178), .Z(n5177) );
  BUFFD0 U5172 ( .I(n5179), .Z(n5178) );
  BUFFD0 U5173 ( .I(n5180), .Z(n5179) );
  BUFFD0 U5174 ( .I(n5181), .Z(n5180) );
  BUFFD0 U5175 ( .I(n5182), .Z(n5181) );
  BUFFD0 U5176 ( .I(n5183), .Z(n5182) );
  BUFFD0 U5177 ( .I(n5184), .Z(n5183) );
  BUFFD0 U5178 ( .I(n5185), .Z(n5184) );
  BUFFD0 U5179 ( .I(n5186), .Z(n5185) );
  BUFFD0 U5180 ( .I(n5187), .Z(n5186) );
  BUFFD0 U5181 ( .I(n5188), .Z(n5187) );
  BUFFD0 U5182 ( .I(n5189), .Z(n5188) );
  BUFFD0 U5183 ( .I(n5190), .Z(n5189) );
  BUFFD0 U5184 ( .I(n5191), .Z(n5190) );
  BUFFD0 U5185 ( .I(n5192), .Z(n5191) );
  BUFFD0 U5186 ( .I(n5193), .Z(n5192) );
  BUFFD0 U5187 ( .I(n5194), .Z(n5193) );
  BUFFD0 U5188 ( .I(n5195), .Z(n5194) );
  BUFFD0 U5189 ( .I(n5196), .Z(n5195) );
  BUFFD0 U5190 ( .I(n5197), .Z(n5196) );
  BUFFD0 U5191 ( .I(n5198), .Z(n5197) );
  BUFFD0 U5192 ( .I(n5199), .Z(n5198) );
  BUFFD0 U5193 ( .I(n5200), .Z(n5199) );
  BUFFD0 U5194 ( .I(n5201), .Z(n5200) );
  BUFFD0 U5195 ( .I(n5202), .Z(n5201) );
  BUFFD0 U5196 ( .I(n5203), .Z(n5202) );
  BUFFD0 U5197 ( .I(n5204), .Z(n5203) );
  BUFFD0 U5198 ( .I(n5205), .Z(n5204) );
  BUFFD0 U5199 ( .I(n5206), .Z(n5205) );
  BUFFD0 U5200 ( .I(n5207), .Z(n5206) );
  BUFFD0 U5201 ( .I(n5208), .Z(n5207) );
  BUFFD0 U5202 ( .I(n5209), .Z(n5208) );
  BUFFD0 U5203 ( .I(n5210), .Z(n5209) );
  BUFFD0 U5204 ( .I(n5211), .Z(n5210) );
  BUFFD0 U5205 ( .I(n5212), .Z(n5211) );
  BUFFD0 U5206 ( .I(n5213), .Z(n5212) );
  BUFFD0 U5207 ( .I(n5214), .Z(n5213) );
  BUFFD0 U5208 ( .I(n5215), .Z(n5214) );
  BUFFD0 U5209 ( .I(n5216), .Z(n5215) );
  BUFFD0 U5210 ( .I(n5217), .Z(n5216) );
  BUFFD0 U5211 ( .I(n5218), .Z(n5217) );
  BUFFD0 U5212 ( .I(n5219), .Z(n5218) );
  BUFFD0 U5213 ( .I(n5220), .Z(n5219) );
  BUFFD0 U5214 ( .I(n5221), .Z(n5220) );
  BUFFD0 U5215 ( .I(n5222), .Z(n5221) );
  BUFFD0 U5216 ( .I(n5223), .Z(n5222) );
  BUFFD0 U5217 ( .I(n5224), .Z(n5223) );
  BUFFD0 U5218 ( .I(n5225), .Z(n5224) );
  BUFFD0 U5219 ( .I(n5226), .Z(n5225) );
  BUFFD0 U5220 ( .I(n5227), .Z(n5226) );
  BUFFD0 U5221 ( .I(n5228), .Z(n5227) );
  BUFFD0 U5222 ( .I(n5229), .Z(n5228) );
  BUFFD0 U5223 ( .I(n5230), .Z(n5229) );
  BUFFD0 U5224 ( .I(n5231), .Z(n5230) );
  BUFFD0 U5225 ( .I(n5232), .Z(n5231) );
  BUFFD0 U5226 ( .I(n5233), .Z(n5232) );
  BUFFD0 U5227 ( .I(n5234), .Z(n5233) );
  BUFFD0 U5228 ( .I(n5235), .Z(n5234) );
  BUFFD0 U5229 ( .I(n5236), .Z(n5235) );
  BUFFD0 U5230 ( .I(n5237), .Z(n5236) );
  BUFFD0 U5231 ( .I(n5238), .Z(n5237) );
  BUFFD0 U5232 ( .I(n5239), .Z(n5238) );
  BUFFD0 U5233 ( .I(n5240), .Z(n5239) );
  BUFFD0 U5234 ( .I(n5241), .Z(n5240) );
  BUFFD0 U5235 ( .I(n5242), .Z(n5241) );
  BUFFD0 U5236 ( .I(n5243), .Z(n5242) );
  BUFFD0 U5237 ( .I(n5244), .Z(n5243) );
  BUFFD0 U5238 ( .I(n5245), .Z(n5244) );
  BUFFD0 U5239 ( .I(n5246), .Z(n5245) );
  BUFFD0 U5240 ( .I(n5247), .Z(n5246) );
  BUFFD0 U5241 ( .I(n5248), .Z(n5247) );
  BUFFD0 U5242 ( .I(n5249), .Z(n5248) );
  BUFFD0 U5243 ( .I(n5250), .Z(n5249) );
  BUFFD0 U5244 ( .I(n5251), .Z(n5250) );
  BUFFD0 U5245 ( .I(n5252), .Z(n5251) );
  BUFFD0 U5246 ( .I(n5253), .Z(n5252) );
  BUFFD0 U5247 ( .I(n5254), .Z(n5253) );
  BUFFD0 U5248 ( .I(n5255), .Z(n5254) );
  BUFFD0 U5249 ( .I(n5256), .Z(n5255) );
  BUFFD0 U5250 ( .I(n5257), .Z(n5256) );
  BUFFD0 U5251 ( .I(n5258), .Z(n5257) );
  BUFFD0 U5252 ( .I(n5259), .Z(n5258) );
  BUFFD0 U5253 ( .I(n5260), .Z(n5259) );
  BUFFD0 U5254 ( .I(n5261), .Z(n5260) );
  BUFFD0 U5255 ( .I(n5262), .Z(n5261) );
  BUFFD0 U5256 ( .I(n5263), .Z(n5262) );
  BUFFD0 U5257 ( .I(n5264), .Z(n5263) );
  BUFFD0 U5258 ( .I(n5265), .Z(n5264) );
  BUFFD0 U5259 ( .I(n5266), .Z(n5265) );
  BUFFD0 U5260 ( .I(n5267), .Z(n5266) );
  BUFFD0 U5261 ( .I(n5268), .Z(n5267) );
  BUFFD0 U5262 ( .I(n5269), .Z(n5268) );
  BUFFD0 U5263 ( .I(n5270), .Z(n5269) );
  BUFFD0 U5264 ( .I(n5271), .Z(n5270) );
  BUFFD0 U5265 ( .I(n5272), .Z(n5271) );
  BUFFD0 U5266 ( .I(n5273), .Z(n5272) );
  BUFFD0 U5267 ( .I(n5274), .Z(n5273) );
  BUFFD0 U5268 ( .I(n5275), .Z(n5274) );
  BUFFD0 U5269 ( .I(n5276), .Z(n5275) );
  BUFFD0 U5270 ( .I(n5277), .Z(n5276) );
  BUFFD0 U5271 ( .I(n5278), .Z(n5277) );
  BUFFD0 U5272 ( .I(n5279), .Z(n5278) );
  BUFFD0 U5273 ( .I(n5280), .Z(n5279) );
  BUFFD0 U5274 ( .I(n5281), .Z(n5280) );
  BUFFD0 U5275 ( .I(n5282), .Z(n5281) );
  BUFFD0 U5276 ( .I(n5283), .Z(n5282) );
  BUFFD0 U5277 ( .I(n5284), .Z(n5283) );
  BUFFD0 U5278 ( .I(n5285), .Z(n5284) );
  BUFFD0 U5279 ( .I(n5286), .Z(n5285) );
  BUFFD0 U5280 ( .I(n5287), .Z(n5286) );
  BUFFD0 U5281 ( .I(n5288), .Z(n5287) );
  BUFFD0 U5282 ( .I(n5289), .Z(n5288) );
  BUFFD0 U5283 ( .I(n5290), .Z(n5289) );
  BUFFD0 U5284 ( .I(n5291), .Z(n5290) );
  BUFFD0 U5285 ( .I(n5292), .Z(n5291) );
  BUFFD0 U5286 ( .I(n5293), .Z(n5292) );
  BUFFD0 U5287 ( .I(n5294), .Z(n5293) );
  BUFFD0 U5288 ( .I(n5295), .Z(n5294) );
  BUFFD0 U5289 ( .I(n5296), .Z(n5295) );
  BUFFD0 U5290 ( .I(n5297), .Z(n5296) );
  BUFFD0 U5291 ( .I(n5298), .Z(n5297) );
  BUFFD0 U5292 ( .I(n5299), .Z(n5298) );
  BUFFD0 U5293 ( .I(n5300), .Z(n5299) );
  BUFFD0 U5294 ( .I(n5301), .Z(n5300) );
  BUFFD0 U5295 ( .I(n5302), .Z(n5301) );
  BUFFD0 U5296 ( .I(n5303), .Z(n5302) );
  BUFFD0 U5297 ( .I(n5304), .Z(n5303) );
  BUFFD0 U5298 ( .I(n5305), .Z(n5304) );
  BUFFD0 U5299 ( .I(n5306), .Z(n5305) );
  BUFFD0 U5300 ( .I(n5307), .Z(n5306) );
  BUFFD0 U5301 ( .I(n5308), .Z(n5307) );
  BUFFD0 U5302 ( .I(n5309), .Z(n5308) );
  BUFFD0 U5303 ( .I(n5310), .Z(n5309) );
  BUFFD0 U5304 ( .I(n5311), .Z(n5310) );
  BUFFD0 U5305 ( .I(n5312), .Z(n5311) );
  BUFFD0 U5306 ( .I(n5313), .Z(n5312) );
  BUFFD0 U5307 ( .I(n5314), .Z(n5313) );
  BUFFD0 U5308 ( .I(n5315), .Z(n5314) );
  BUFFD0 U5309 ( .I(n5316), .Z(n5315) );
  BUFFD0 U5310 ( .I(n5317), .Z(n5316) );
  BUFFD0 U5311 ( .I(n5318), .Z(n5317) );
  BUFFD0 U5312 ( .I(n5319), .Z(n5318) );
  BUFFD0 U5313 ( .I(n5320), .Z(n5319) );
  BUFFD0 U5314 ( .I(n5321), .Z(n5320) );
  BUFFD0 U5315 ( .I(n5322), .Z(n5321) );
  BUFFD0 U5316 ( .I(n5323), .Z(n5322) );
  BUFFD0 U5317 ( .I(n5324), .Z(n5323) );
  BUFFD0 U5318 ( .I(n5325), .Z(n5324) );
  BUFFD0 U5319 ( .I(n5326), .Z(n5325) );
  BUFFD0 U5320 ( .I(n5327), .Z(n5326) );
  BUFFD0 U5321 ( .I(n5328), .Z(n5327) );
  BUFFD0 U5322 ( .I(n5329), .Z(n5328) );
  BUFFD0 U5323 ( .I(n5330), .Z(n5329) );
  BUFFD0 U5324 ( .I(n5331), .Z(n5330) );
  BUFFD0 U5325 ( .I(n5332), .Z(n5331) );
  BUFFD0 U5326 ( .I(n8713), .Z(n5332) );
  BUFFD0 U5327 ( .I(n8710), .Z(n5333) );
  BUFFD0 U5328 ( .I(n5335), .Z(n5334) );
  BUFFD0 U5329 ( .I(n5336), .Z(n5335) );
  BUFFD0 U5330 ( .I(n5337), .Z(n5336) );
  BUFFD0 U5331 ( .I(n5338), .Z(n5337) );
  BUFFD0 U5332 ( .I(n5339), .Z(n5338) );
  BUFFD0 U5333 ( .I(n5340), .Z(n5339) );
  BUFFD0 U5334 ( .I(n5341), .Z(n5340) );
  BUFFD0 U5335 ( .I(n5342), .Z(n5341) );
  BUFFD0 U5336 ( .I(n5343), .Z(n5342) );
  BUFFD0 U5337 ( .I(n5344), .Z(n5343) );
  BUFFD0 U5338 ( .I(n5345), .Z(n5344) );
  BUFFD0 U5339 ( .I(n5346), .Z(n5345) );
  BUFFD0 U5340 ( .I(n5347), .Z(n5346) );
  BUFFD0 U5341 ( .I(n5348), .Z(n5347) );
  BUFFD0 U5342 ( .I(n5349), .Z(n5348) );
  BUFFD0 U5343 ( .I(n5350), .Z(n5349) );
  BUFFD0 U5344 ( .I(n5351), .Z(n5350) );
  BUFFD0 U5345 ( .I(n5352), .Z(n5351) );
  BUFFD0 U5346 ( .I(n5353), .Z(n5352) );
  BUFFD0 U5347 ( .I(n5354), .Z(n5353) );
  BUFFD0 U5348 ( .I(n5355), .Z(n5354) );
  BUFFD0 U5349 ( .I(n5356), .Z(n5355) );
  BUFFD0 U5350 ( .I(n5357), .Z(n5356) );
  BUFFD0 U5351 ( .I(n5358), .Z(n5357) );
  BUFFD0 U5352 ( .I(n5359), .Z(n5358) );
  BUFFD0 U5353 ( .I(n5360), .Z(n5359) );
  BUFFD0 U5354 ( .I(n5361), .Z(n5360) );
  BUFFD0 U5355 ( .I(n5362), .Z(n5361) );
  BUFFD0 U5356 ( .I(n5363), .Z(n5362) );
  BUFFD0 U5357 ( .I(n5364), .Z(n5363) );
  BUFFD0 U5358 ( .I(n5365), .Z(n5364) );
  BUFFD0 U5359 ( .I(n5366), .Z(n5365) );
  BUFFD0 U5360 ( .I(n5367), .Z(n5366) );
  BUFFD0 U5361 ( .I(n5368), .Z(n5367) );
  BUFFD0 U5362 ( .I(n5369), .Z(n5368) );
  BUFFD0 U5363 ( .I(n5370), .Z(n5369) );
  BUFFD0 U5364 ( .I(n5371), .Z(n5370) );
  BUFFD0 U5365 ( .I(n5372), .Z(n5371) );
  BUFFD0 U5366 ( .I(n5373), .Z(n5372) );
  BUFFD0 U5367 ( .I(n5374), .Z(n5373) );
  BUFFD0 U5368 ( .I(n5375), .Z(n5374) );
  BUFFD0 U5369 ( .I(n5376), .Z(n5375) );
  BUFFD0 U5370 ( .I(n5377), .Z(n5376) );
  BUFFD0 U5371 ( .I(n5378), .Z(n5377) );
  BUFFD0 U5372 ( .I(n5379), .Z(n5378) );
  BUFFD0 U5373 ( .I(n5380), .Z(n5379) );
  BUFFD0 U5374 ( .I(n5381), .Z(n5380) );
  BUFFD0 U5375 ( .I(n5382), .Z(n5381) );
  BUFFD0 U5376 ( .I(n5383), .Z(n5382) );
  BUFFD0 U5377 ( .I(n5384), .Z(n5383) );
  BUFFD0 U5378 ( .I(n5385), .Z(n5384) );
  BUFFD0 U5379 ( .I(n5386), .Z(n5385) );
  BUFFD0 U5380 ( .I(n5387), .Z(n5386) );
  BUFFD0 U5381 ( .I(n5388), .Z(n5387) );
  BUFFD0 U5382 ( .I(n5389), .Z(n5388) );
  BUFFD0 U5383 ( .I(n5390), .Z(n5389) );
  BUFFD0 U5384 ( .I(n5391), .Z(n5390) );
  BUFFD0 U5385 ( .I(n5392), .Z(n5391) );
  BUFFD0 U5386 ( .I(n5393), .Z(n5392) );
  BUFFD0 U5387 ( .I(n5394), .Z(n5393) );
  BUFFD0 U5388 ( .I(n5395), .Z(n5394) );
  BUFFD0 U5389 ( .I(n5396), .Z(n5395) );
  BUFFD0 U5390 ( .I(n5397), .Z(n5396) );
  BUFFD0 U5391 ( .I(n5398), .Z(n5397) );
  BUFFD0 U5392 ( .I(n5399), .Z(n5398) );
  BUFFD0 U5393 ( .I(n5400), .Z(n5399) );
  BUFFD0 U5394 ( .I(n5401), .Z(n5400) );
  BUFFD0 U5395 ( .I(n5402), .Z(n5401) );
  BUFFD0 U5396 ( .I(n5403), .Z(n5402) );
  BUFFD0 U5397 ( .I(n5404), .Z(n5403) );
  BUFFD0 U5398 ( .I(n5405), .Z(n5404) );
  BUFFD0 U5399 ( .I(n5406), .Z(n5405) );
  BUFFD0 U5400 ( .I(n5407), .Z(n5406) );
  BUFFD0 U5401 ( .I(n5408), .Z(n5407) );
  BUFFD0 U5402 ( .I(n5409), .Z(n5408) );
  BUFFD0 U5403 ( .I(n5410), .Z(n5409) );
  BUFFD0 U5404 ( .I(n5411), .Z(n5410) );
  BUFFD0 U5405 ( .I(n5412), .Z(n5411) );
  BUFFD0 U5406 ( .I(n5413), .Z(n5412) );
  BUFFD0 U5407 ( .I(n5414), .Z(n5413) );
  BUFFD0 U5408 ( .I(n5415), .Z(n5414) );
  BUFFD0 U5409 ( .I(n5416), .Z(n5415) );
  BUFFD0 U5410 ( .I(n5417), .Z(n5416) );
  BUFFD0 U5411 ( .I(n5418), .Z(n5417) );
  BUFFD0 U5412 ( .I(n5419), .Z(n5418) );
  BUFFD0 U5413 ( .I(n5420), .Z(n5419) );
  BUFFD0 U5414 ( .I(n5421), .Z(n5420) );
  BUFFD0 U5415 ( .I(n5422), .Z(n5421) );
  BUFFD0 U5416 ( .I(n5423), .Z(n5422) );
  BUFFD0 U5417 ( .I(n5424), .Z(n5423) );
  BUFFD0 U5418 ( .I(n5425), .Z(n5424) );
  BUFFD0 U5419 ( .I(n5426), .Z(n5425) );
  BUFFD0 U5420 ( .I(n5427), .Z(n5426) );
  BUFFD0 U5421 ( .I(n5428), .Z(n5427) );
  BUFFD0 U5422 ( .I(n5429), .Z(n5428) );
  BUFFD0 U5423 ( .I(n5430), .Z(n5429) );
  BUFFD0 U5424 ( .I(n5431), .Z(n5430) );
  BUFFD0 U5425 ( .I(n5432), .Z(n5431) );
  BUFFD0 U5426 ( .I(n5433), .Z(n5432) );
  BUFFD0 U5427 ( .I(n5434), .Z(n5433) );
  BUFFD0 U5428 ( .I(n5435), .Z(n5434) );
  BUFFD0 U5429 ( .I(n5436), .Z(n5435) );
  BUFFD0 U5430 ( .I(n5437), .Z(n5436) );
  BUFFD0 U5431 ( .I(n5438), .Z(n5437) );
  BUFFD0 U5432 ( .I(n5439), .Z(n5438) );
  BUFFD0 U5433 ( .I(n5440), .Z(n5439) );
  BUFFD0 U5434 ( .I(n5441), .Z(n5440) );
  BUFFD0 U5435 ( .I(n5442), .Z(n5441) );
  BUFFD0 U5436 ( .I(n5443), .Z(n5442) );
  BUFFD0 U5437 ( .I(n5444), .Z(n5443) );
  BUFFD0 U5438 ( .I(n5445), .Z(n5444) );
  BUFFD0 U5439 ( .I(n5446), .Z(n5445) );
  BUFFD0 U5440 ( .I(n5447), .Z(n5446) );
  BUFFD0 U5441 ( .I(n5448), .Z(n5447) );
  BUFFD0 U5442 ( .I(n5449), .Z(n5448) );
  BUFFD0 U5443 ( .I(n5450), .Z(n5449) );
  BUFFD0 U5444 ( .I(n5451), .Z(n5450) );
  BUFFD0 U5445 ( .I(n5452), .Z(n5451) );
  BUFFD0 U5446 ( .I(n5453), .Z(n5452) );
  BUFFD0 U5447 ( .I(n5454), .Z(n5453) );
  BUFFD0 U5448 ( .I(n5455), .Z(n5454) );
  BUFFD0 U5449 ( .I(n5456), .Z(n5455) );
  BUFFD0 U5450 ( .I(n5457), .Z(n5456) );
  BUFFD0 U5451 ( .I(n5458), .Z(n5457) );
  BUFFD0 U5452 ( .I(n5459), .Z(n5458) );
  BUFFD0 U5453 ( .I(n5460), .Z(n5459) );
  BUFFD0 U5454 ( .I(n5461), .Z(n5460) );
  BUFFD0 U5455 ( .I(n5462), .Z(n5461) );
  BUFFD0 U5456 ( .I(n5463), .Z(n5462) );
  BUFFD0 U5457 ( .I(n5464), .Z(n5463) );
  BUFFD0 U5458 ( .I(n5465), .Z(n5464) );
  BUFFD0 U5459 ( .I(n5466), .Z(n5465) );
  BUFFD0 U5460 ( .I(n5467), .Z(n5466) );
  BUFFD0 U5461 ( .I(n5468), .Z(n5467) );
  BUFFD0 U5462 ( .I(n5469), .Z(n5468) );
  BUFFD0 U5463 ( .I(n5470), .Z(n5469) );
  BUFFD0 U5464 ( .I(n5471), .Z(n5470) );
  BUFFD0 U5465 ( .I(n5472), .Z(n5471) );
  BUFFD0 U5466 ( .I(n5473), .Z(n5472) );
  BUFFD0 U5467 ( .I(n5474), .Z(n5473) );
  BUFFD0 U5468 ( .I(n5475), .Z(n5474) );
  BUFFD0 U5469 ( .I(n5476), .Z(n5475) );
  BUFFD0 U5470 ( .I(n5477), .Z(n5476) );
  BUFFD0 U5471 ( .I(n5478), .Z(n5477) );
  BUFFD0 U5472 ( .I(n5479), .Z(n5478) );
  BUFFD0 U5473 ( .I(n5480), .Z(n5479) );
  BUFFD0 U5474 ( .I(n5481), .Z(n5480) );
  BUFFD0 U5475 ( .I(n5482), .Z(n5481) );
  BUFFD0 U5476 ( .I(n5483), .Z(n5482) );
  BUFFD0 U5477 ( .I(n5484), .Z(n5483) );
  BUFFD0 U5478 ( .I(n5485), .Z(n5484) );
  BUFFD0 U5479 ( .I(n5486), .Z(n5485) );
  BUFFD0 U5480 ( .I(n5487), .Z(n5486) );
  BUFFD0 U5481 ( .I(n5488), .Z(n5487) );
  BUFFD0 U5482 ( .I(n5489), .Z(n5488) );
  BUFFD0 U5483 ( .I(n5490), .Z(n5489) );
  BUFFD0 U5484 ( .I(n5491), .Z(n5490) );
  BUFFD0 U5485 ( .I(n5492), .Z(n5491) );
  BUFFD0 U5486 ( .I(n5493), .Z(n5492) );
  BUFFD0 U5487 ( .I(n5494), .Z(n5493) );
  BUFFD0 U5488 ( .I(n5495), .Z(n5494) );
  BUFFD0 U5489 ( .I(n5496), .Z(n5495) );
  BUFFD0 U5490 ( .I(n5497), .Z(n5496) );
  BUFFD0 U5491 ( .I(n5498), .Z(n5497) );
  BUFFD0 U5492 ( .I(n5499), .Z(n5498) );
  BUFFD0 U5493 ( .I(n5500), .Z(n5499) );
  BUFFD0 U5494 ( .I(n5501), .Z(n5500) );
  BUFFD0 U5495 ( .I(n5502), .Z(n5501) );
  BUFFD0 U5496 ( .I(n5503), .Z(n5502) );
  BUFFD0 U5497 ( .I(n5504), .Z(n5503) );
  BUFFD0 U5498 ( .I(n5505), .Z(n5504) );
  BUFFD0 U5499 ( .I(n5506), .Z(n5505) );
  BUFFD0 U5500 ( .I(n5507), .Z(n5506) );
  BUFFD0 U5501 ( .I(n5508), .Z(n5507) );
  BUFFD0 U5502 ( .I(n5509), .Z(n5508) );
  BUFFD0 U5503 ( .I(n5510), .Z(n5509) );
  BUFFD0 U5504 ( .I(n5511), .Z(n5510) );
  BUFFD0 U5505 ( .I(n8711), .Z(n5511) );
  BUFFD0 U5506 ( .I(n8708), .Z(n5512) );
  BUFFD0 U5507 ( .I(n5514), .Z(n5513) );
  BUFFD0 U5508 ( .I(n5515), .Z(n5514) );
  BUFFD0 U5509 ( .I(n5516), .Z(n5515) );
  BUFFD0 U5510 ( .I(n5517), .Z(n5516) );
  BUFFD0 U5511 ( .I(n5518), .Z(n5517) );
  BUFFD0 U5512 ( .I(n5519), .Z(n5518) );
  BUFFD0 U5513 ( .I(n5520), .Z(n5519) );
  BUFFD0 U5514 ( .I(n5521), .Z(n5520) );
  BUFFD0 U5515 ( .I(n5522), .Z(n5521) );
  BUFFD0 U5516 ( .I(n5523), .Z(n5522) );
  BUFFD0 U5517 ( .I(n5524), .Z(n5523) );
  BUFFD0 U5518 ( .I(n5525), .Z(n5524) );
  BUFFD0 U5519 ( .I(n5526), .Z(n5525) );
  BUFFD0 U5520 ( .I(n5527), .Z(n5526) );
  BUFFD0 U5521 ( .I(n5528), .Z(n5527) );
  BUFFD0 U5522 ( .I(n5529), .Z(n5528) );
  BUFFD0 U5523 ( .I(n5530), .Z(n5529) );
  BUFFD0 U5524 ( .I(n5531), .Z(n5530) );
  BUFFD0 U5525 ( .I(n5532), .Z(n5531) );
  BUFFD0 U5526 ( .I(n5533), .Z(n5532) );
  BUFFD0 U5527 ( .I(n5534), .Z(n5533) );
  BUFFD0 U5528 ( .I(n5535), .Z(n5534) );
  BUFFD0 U5529 ( .I(n5536), .Z(n5535) );
  BUFFD0 U5530 ( .I(n5537), .Z(n5536) );
  BUFFD0 U5531 ( .I(n5538), .Z(n5537) );
  BUFFD0 U5532 ( .I(n5539), .Z(n5538) );
  BUFFD0 U5533 ( .I(n5540), .Z(n5539) );
  BUFFD0 U5534 ( .I(n5541), .Z(n5540) );
  BUFFD0 U5535 ( .I(n5542), .Z(n5541) );
  BUFFD0 U5536 ( .I(n5543), .Z(n5542) );
  BUFFD0 U5537 ( .I(n5544), .Z(n5543) );
  BUFFD0 U5538 ( .I(n5545), .Z(n5544) );
  BUFFD0 U5539 ( .I(n5546), .Z(n5545) );
  BUFFD0 U5540 ( .I(n5547), .Z(n5546) );
  BUFFD0 U5541 ( .I(n5548), .Z(n5547) );
  BUFFD0 U5542 ( .I(n5549), .Z(n5548) );
  BUFFD0 U5543 ( .I(n5550), .Z(n5549) );
  BUFFD0 U5544 ( .I(n5551), .Z(n5550) );
  BUFFD0 U5545 ( .I(n5552), .Z(n5551) );
  BUFFD0 U5546 ( .I(n5553), .Z(n5552) );
  BUFFD0 U5547 ( .I(n5554), .Z(n5553) );
  BUFFD0 U5548 ( .I(n5555), .Z(n5554) );
  BUFFD0 U5549 ( .I(n5556), .Z(n5555) );
  BUFFD0 U5550 ( .I(n5557), .Z(n5556) );
  BUFFD0 U5551 ( .I(n5558), .Z(n5557) );
  BUFFD0 U5552 ( .I(n5559), .Z(n5558) );
  BUFFD0 U5553 ( .I(n5560), .Z(n5559) );
  BUFFD0 U5554 ( .I(n5561), .Z(n5560) );
  BUFFD0 U5555 ( .I(n5562), .Z(n5561) );
  BUFFD0 U5556 ( .I(n5563), .Z(n5562) );
  BUFFD0 U5557 ( .I(n5564), .Z(n5563) );
  BUFFD0 U5558 ( .I(n5565), .Z(n5564) );
  BUFFD0 U5559 ( .I(n5566), .Z(n5565) );
  BUFFD0 U5560 ( .I(n5567), .Z(n5566) );
  BUFFD0 U5561 ( .I(n5568), .Z(n5567) );
  BUFFD0 U5562 ( .I(n5569), .Z(n5568) );
  BUFFD0 U5563 ( .I(n5570), .Z(n5569) );
  BUFFD0 U5564 ( .I(n5571), .Z(n5570) );
  BUFFD0 U5565 ( .I(n5572), .Z(n5571) );
  BUFFD0 U5566 ( .I(n5573), .Z(n5572) );
  BUFFD0 U5567 ( .I(n5574), .Z(n5573) );
  BUFFD0 U5568 ( .I(n5575), .Z(n5574) );
  BUFFD0 U5569 ( .I(n5576), .Z(n5575) );
  BUFFD0 U5570 ( .I(n5577), .Z(n5576) );
  BUFFD0 U5571 ( .I(n5578), .Z(n5577) );
  BUFFD0 U5572 ( .I(n5579), .Z(n5578) );
  BUFFD0 U5573 ( .I(n5580), .Z(n5579) );
  BUFFD0 U5574 ( .I(n5581), .Z(n5580) );
  BUFFD0 U5575 ( .I(n5582), .Z(n5581) );
  BUFFD0 U5576 ( .I(n5583), .Z(n5582) );
  BUFFD0 U5577 ( .I(n5584), .Z(n5583) );
  BUFFD0 U5578 ( .I(n5585), .Z(n5584) );
  BUFFD0 U5579 ( .I(n5586), .Z(n5585) );
  BUFFD0 U5580 ( .I(n5587), .Z(n5586) );
  BUFFD0 U5581 ( .I(n5588), .Z(n5587) );
  BUFFD0 U5582 ( .I(n5589), .Z(n5588) );
  BUFFD0 U5583 ( .I(n5590), .Z(n5589) );
  BUFFD0 U5584 ( .I(n5591), .Z(n5590) );
  BUFFD0 U5585 ( .I(n5592), .Z(n5591) );
  BUFFD0 U5586 ( .I(n5593), .Z(n5592) );
  BUFFD0 U5587 ( .I(n5594), .Z(n5593) );
  BUFFD0 U5588 ( .I(n5595), .Z(n5594) );
  BUFFD0 U5589 ( .I(n5596), .Z(n5595) );
  BUFFD0 U5590 ( .I(n5597), .Z(n5596) );
  BUFFD0 U5591 ( .I(n5598), .Z(n5597) );
  BUFFD0 U5592 ( .I(n5599), .Z(n5598) );
  BUFFD0 U5593 ( .I(n5600), .Z(n5599) );
  BUFFD0 U5594 ( .I(n5601), .Z(n5600) );
  BUFFD0 U5595 ( .I(n5602), .Z(n5601) );
  BUFFD0 U5596 ( .I(n5603), .Z(n5602) );
  BUFFD0 U5597 ( .I(n5604), .Z(n5603) );
  BUFFD0 U5598 ( .I(n5605), .Z(n5604) );
  BUFFD0 U5599 ( .I(n5606), .Z(n5605) );
  BUFFD0 U5600 ( .I(n5607), .Z(n5606) );
  BUFFD0 U5601 ( .I(n5608), .Z(n5607) );
  BUFFD0 U5602 ( .I(n5609), .Z(n5608) );
  BUFFD0 U5603 ( .I(n5610), .Z(n5609) );
  BUFFD0 U5604 ( .I(n5611), .Z(n5610) );
  BUFFD0 U5605 ( .I(n5612), .Z(n5611) );
  BUFFD0 U5606 ( .I(n5613), .Z(n5612) );
  BUFFD0 U5607 ( .I(n5614), .Z(n5613) );
  BUFFD0 U5608 ( .I(n5615), .Z(n5614) );
  BUFFD0 U5609 ( .I(n5616), .Z(n5615) );
  BUFFD0 U5610 ( .I(n5617), .Z(n5616) );
  BUFFD0 U5611 ( .I(n5618), .Z(n5617) );
  BUFFD0 U5612 ( .I(n5619), .Z(n5618) );
  BUFFD0 U5613 ( .I(n5620), .Z(n5619) );
  BUFFD0 U5614 ( .I(n5621), .Z(n5620) );
  BUFFD0 U5615 ( .I(n5622), .Z(n5621) );
  BUFFD0 U5616 ( .I(n5623), .Z(n5622) );
  BUFFD0 U5617 ( .I(n5624), .Z(n5623) );
  BUFFD0 U5618 ( .I(n5625), .Z(n5624) );
  BUFFD0 U5619 ( .I(n5626), .Z(n5625) );
  BUFFD0 U5620 ( .I(n5627), .Z(n5626) );
  BUFFD0 U5621 ( .I(n5628), .Z(n5627) );
  BUFFD0 U5622 ( .I(n5629), .Z(n5628) );
  BUFFD0 U5623 ( .I(n5630), .Z(n5629) );
  BUFFD0 U5624 ( .I(n5631), .Z(n5630) );
  BUFFD0 U5625 ( .I(n5632), .Z(n5631) );
  BUFFD0 U5626 ( .I(n5633), .Z(n5632) );
  BUFFD0 U5627 ( .I(n5634), .Z(n5633) );
  BUFFD0 U5628 ( .I(n5635), .Z(n5634) );
  BUFFD0 U5629 ( .I(n5636), .Z(n5635) );
  BUFFD0 U5630 ( .I(n5637), .Z(n5636) );
  BUFFD0 U5631 ( .I(n5638), .Z(n5637) );
  BUFFD0 U5632 ( .I(n5639), .Z(n5638) );
  BUFFD0 U5633 ( .I(n5640), .Z(n5639) );
  BUFFD0 U5634 ( .I(n5641), .Z(n5640) );
  BUFFD0 U5635 ( .I(n5642), .Z(n5641) );
  BUFFD0 U5636 ( .I(n5643), .Z(n5642) );
  BUFFD0 U5637 ( .I(n5644), .Z(n5643) );
  BUFFD0 U5638 ( .I(n5645), .Z(n5644) );
  BUFFD0 U5639 ( .I(n5646), .Z(n5645) );
  BUFFD0 U5640 ( .I(n5647), .Z(n5646) );
  BUFFD0 U5641 ( .I(n5648), .Z(n5647) );
  BUFFD0 U5642 ( .I(n5649), .Z(n5648) );
  BUFFD0 U5643 ( .I(n5650), .Z(n5649) );
  BUFFD0 U5644 ( .I(n5651), .Z(n5650) );
  BUFFD0 U5645 ( .I(n5652), .Z(n5651) );
  BUFFD0 U5646 ( .I(n5653), .Z(n5652) );
  BUFFD0 U5647 ( .I(n5654), .Z(n5653) );
  BUFFD0 U5648 ( .I(n5655), .Z(n5654) );
  BUFFD0 U5649 ( .I(n5656), .Z(n5655) );
  BUFFD0 U5650 ( .I(n5657), .Z(n5656) );
  BUFFD0 U5651 ( .I(n5658), .Z(n5657) );
  BUFFD0 U5652 ( .I(n5659), .Z(n5658) );
  BUFFD0 U5653 ( .I(n5660), .Z(n5659) );
  BUFFD0 U5654 ( .I(n5661), .Z(n5660) );
  BUFFD0 U5655 ( .I(n5662), .Z(n5661) );
  BUFFD0 U5656 ( .I(n5663), .Z(n5662) );
  BUFFD0 U5657 ( .I(n5664), .Z(n5663) );
  BUFFD0 U5658 ( .I(n5665), .Z(n5664) );
  BUFFD0 U5659 ( .I(n5666), .Z(n5665) );
  BUFFD0 U5660 ( .I(n5667), .Z(n5666) );
  BUFFD0 U5661 ( .I(n5668), .Z(n5667) );
  BUFFD0 U5662 ( .I(n5669), .Z(n5668) );
  BUFFD0 U5663 ( .I(n5670), .Z(n5669) );
  BUFFD0 U5664 ( .I(n5671), .Z(n5670) );
  BUFFD0 U5665 ( .I(n5672), .Z(n5671) );
  BUFFD0 U5666 ( .I(n5673), .Z(n5672) );
  BUFFD0 U5667 ( .I(n5674), .Z(n5673) );
  BUFFD0 U5668 ( .I(n5675), .Z(n5674) );
  BUFFD0 U5669 ( .I(n5676), .Z(n5675) );
  BUFFD0 U5670 ( .I(n5677), .Z(n5676) );
  BUFFD0 U5671 ( .I(n5678), .Z(n5677) );
  BUFFD0 U5672 ( .I(n5679), .Z(n5678) );
  BUFFD0 U5673 ( .I(n5680), .Z(n5679) );
  BUFFD0 U5674 ( .I(n5681), .Z(n5680) );
  BUFFD0 U5675 ( .I(n5682), .Z(n5681) );
  BUFFD0 U5676 ( .I(n5683), .Z(n5682) );
  BUFFD0 U5677 ( .I(n5684), .Z(n5683) );
  BUFFD0 U5678 ( .I(n5685), .Z(n5684) );
  BUFFD0 U5679 ( .I(n5686), .Z(n5685) );
  BUFFD0 U5680 ( .I(n5687), .Z(n5686) );
  BUFFD0 U5681 ( .I(n5688), .Z(n5687) );
  BUFFD0 U5682 ( .I(n8709), .Z(n5688) );
  BUFFD0 U5683 ( .I(n8705), .Z(n5689) );
  BUFFD0 U5684 ( .I(n5691), .Z(n5690) );
  BUFFD0 U5685 ( .I(n5692), .Z(n5691) );
  BUFFD0 U5686 ( .I(n5693), .Z(n5692) );
  BUFFD0 U5687 ( .I(n5694), .Z(n5693) );
  BUFFD0 U5688 ( .I(n5695), .Z(n5694) );
  BUFFD0 U5689 ( .I(n5696), .Z(n5695) );
  BUFFD0 U5690 ( .I(n5697), .Z(n5696) );
  BUFFD0 U5691 ( .I(n5698), .Z(n5697) );
  BUFFD0 U5692 ( .I(n5699), .Z(n5698) );
  BUFFD0 U5693 ( .I(n5700), .Z(n5699) );
  BUFFD0 U5694 ( .I(n5701), .Z(n5700) );
  BUFFD0 U5695 ( .I(n5702), .Z(n5701) );
  BUFFD0 U5696 ( .I(n5703), .Z(n5702) );
  BUFFD0 U5697 ( .I(n5704), .Z(n5703) );
  BUFFD0 U5698 ( .I(n5705), .Z(n5704) );
  BUFFD0 U5699 ( .I(n5706), .Z(n5705) );
  BUFFD0 U5700 ( .I(n5707), .Z(n5706) );
  BUFFD0 U5701 ( .I(n5708), .Z(n5707) );
  BUFFD0 U5702 ( .I(n5709), .Z(n5708) );
  BUFFD0 U5703 ( .I(n5710), .Z(n5709) );
  BUFFD0 U5704 ( .I(n5711), .Z(n5710) );
  BUFFD0 U5705 ( .I(n5712), .Z(n5711) );
  BUFFD0 U5706 ( .I(n5713), .Z(n5712) );
  BUFFD0 U5707 ( .I(n5714), .Z(n5713) );
  BUFFD0 U5708 ( .I(n5715), .Z(n5714) );
  BUFFD0 U5709 ( .I(n5716), .Z(n5715) );
  BUFFD0 U5710 ( .I(n5717), .Z(n5716) );
  BUFFD0 U5711 ( .I(n5718), .Z(n5717) );
  BUFFD0 U5712 ( .I(n5719), .Z(n5718) );
  BUFFD0 U5713 ( .I(n5720), .Z(n5719) );
  BUFFD0 U5714 ( .I(n5721), .Z(n5720) );
  BUFFD0 U5715 ( .I(n5722), .Z(n5721) );
  BUFFD0 U5716 ( .I(n5723), .Z(n5722) );
  BUFFD0 U5717 ( .I(n5724), .Z(n5723) );
  BUFFD0 U5718 ( .I(n5725), .Z(n5724) );
  BUFFD0 U5719 ( .I(n5726), .Z(n5725) );
  BUFFD0 U5720 ( .I(n5727), .Z(n5726) );
  BUFFD0 U5721 ( .I(n5728), .Z(n5727) );
  BUFFD0 U5722 ( .I(n5729), .Z(n5728) );
  BUFFD0 U5723 ( .I(n5730), .Z(n5729) );
  BUFFD0 U5724 ( .I(n5731), .Z(n5730) );
  BUFFD0 U5725 ( .I(n5732), .Z(n5731) );
  BUFFD0 U5726 ( .I(n5733), .Z(n5732) );
  BUFFD0 U5727 ( .I(n5734), .Z(n5733) );
  BUFFD0 U5728 ( .I(n5735), .Z(n5734) );
  BUFFD0 U5729 ( .I(n5736), .Z(n5735) );
  BUFFD0 U5730 ( .I(n5737), .Z(n5736) );
  BUFFD0 U5731 ( .I(n5738), .Z(n5737) );
  BUFFD0 U5732 ( .I(n5739), .Z(n5738) );
  BUFFD0 U5733 ( .I(n5740), .Z(n5739) );
  BUFFD0 U5734 ( .I(n5741), .Z(n5740) );
  BUFFD0 U5735 ( .I(n5742), .Z(n5741) );
  BUFFD0 U5736 ( .I(n5743), .Z(n5742) );
  BUFFD0 U5737 ( .I(n5744), .Z(n5743) );
  BUFFD0 U5738 ( .I(n5745), .Z(n5744) );
  BUFFD0 U5739 ( .I(n5746), .Z(n5745) );
  BUFFD0 U5740 ( .I(n5747), .Z(n5746) );
  BUFFD0 U5741 ( .I(n5748), .Z(n5747) );
  BUFFD0 U5742 ( .I(n5749), .Z(n5748) );
  BUFFD0 U5743 ( .I(n5750), .Z(n5749) );
  BUFFD0 U5744 ( .I(n5751), .Z(n5750) );
  BUFFD0 U5745 ( .I(n5752), .Z(n5751) );
  BUFFD0 U5746 ( .I(n5753), .Z(n5752) );
  BUFFD0 U5747 ( .I(n5754), .Z(n5753) );
  BUFFD0 U5748 ( .I(n5755), .Z(n5754) );
  BUFFD0 U5749 ( .I(n5756), .Z(n5755) );
  BUFFD0 U5750 ( .I(n5757), .Z(n5756) );
  BUFFD0 U5751 ( .I(n5758), .Z(n5757) );
  BUFFD0 U5752 ( .I(n5759), .Z(n5758) );
  BUFFD0 U5753 ( .I(n5760), .Z(n5759) );
  BUFFD0 U5754 ( .I(n5761), .Z(n5760) );
  BUFFD0 U5755 ( .I(n5762), .Z(n5761) );
  BUFFD0 U5756 ( .I(n5763), .Z(n5762) );
  BUFFD0 U5757 ( .I(n5764), .Z(n5763) );
  BUFFD0 U5758 ( .I(n5765), .Z(n5764) );
  BUFFD0 U5759 ( .I(n5766), .Z(n5765) );
  BUFFD0 U5760 ( .I(n5767), .Z(n5766) );
  BUFFD0 U5761 ( .I(n5768), .Z(n5767) );
  BUFFD0 U5762 ( .I(n5769), .Z(n5768) );
  BUFFD0 U5763 ( .I(n5770), .Z(n5769) );
  BUFFD0 U5764 ( .I(n5771), .Z(n5770) );
  BUFFD0 U5765 ( .I(n5772), .Z(n5771) );
  BUFFD0 U5766 ( .I(n5773), .Z(n5772) );
  BUFFD0 U5767 ( .I(n5774), .Z(n5773) );
  BUFFD0 U5768 ( .I(n5775), .Z(n5774) );
  BUFFD0 U5769 ( .I(n5776), .Z(n5775) );
  BUFFD0 U5770 ( .I(n5777), .Z(n5776) );
  BUFFD0 U5771 ( .I(n5778), .Z(n5777) );
  BUFFD0 U5772 ( .I(n5779), .Z(n5778) );
  BUFFD0 U5773 ( .I(n5780), .Z(n5779) );
  BUFFD0 U5774 ( .I(n5781), .Z(n5780) );
  BUFFD0 U5775 ( .I(n5782), .Z(n5781) );
  BUFFD0 U5776 ( .I(n5783), .Z(n5782) );
  BUFFD0 U5777 ( .I(n5784), .Z(n5783) );
  BUFFD0 U5778 ( .I(n5785), .Z(n5784) );
  BUFFD0 U5779 ( .I(n5786), .Z(n5785) );
  BUFFD0 U5780 ( .I(n5787), .Z(n5786) );
  BUFFD0 U5781 ( .I(n5788), .Z(n5787) );
  BUFFD0 U5782 ( .I(n5789), .Z(n5788) );
  BUFFD0 U5783 ( .I(n5790), .Z(n5789) );
  BUFFD0 U5784 ( .I(n5791), .Z(n5790) );
  BUFFD0 U5785 ( .I(n5792), .Z(n5791) );
  BUFFD0 U5786 ( .I(n5793), .Z(n5792) );
  BUFFD0 U5787 ( .I(n5794), .Z(n5793) );
  BUFFD0 U5788 ( .I(n5795), .Z(n5794) );
  BUFFD0 U5789 ( .I(n5796), .Z(n5795) );
  BUFFD0 U5790 ( .I(n5797), .Z(n5796) );
  BUFFD0 U5791 ( .I(n5798), .Z(n5797) );
  BUFFD0 U5792 ( .I(n5799), .Z(n5798) );
  BUFFD0 U5793 ( .I(n5800), .Z(n5799) );
  BUFFD0 U5794 ( .I(n5801), .Z(n5800) );
  BUFFD0 U5795 ( .I(n5802), .Z(n5801) );
  BUFFD0 U5796 ( .I(n5803), .Z(n5802) );
  BUFFD0 U5797 ( .I(n5804), .Z(n5803) );
  BUFFD0 U5798 ( .I(n5805), .Z(n5804) );
  BUFFD0 U5799 ( .I(n5806), .Z(n5805) );
  BUFFD0 U5800 ( .I(n5807), .Z(n5806) );
  BUFFD0 U5801 ( .I(n5808), .Z(n5807) );
  BUFFD0 U5802 ( .I(n5809), .Z(n5808) );
  BUFFD0 U5803 ( .I(n5810), .Z(n5809) );
  BUFFD0 U5804 ( .I(n5811), .Z(n5810) );
  BUFFD0 U5805 ( .I(n5812), .Z(n5811) );
  BUFFD0 U5806 ( .I(n5813), .Z(n5812) );
  BUFFD0 U5807 ( .I(n5814), .Z(n5813) );
  BUFFD0 U5808 ( .I(n5815), .Z(n5814) );
  BUFFD0 U5809 ( .I(n5816), .Z(n5815) );
  BUFFD0 U5810 ( .I(n5817), .Z(n5816) );
  BUFFD0 U5811 ( .I(n5818), .Z(n5817) );
  BUFFD0 U5812 ( .I(n5819), .Z(n5818) );
  BUFFD0 U5813 ( .I(n5820), .Z(n5819) );
  BUFFD0 U5814 ( .I(n5821), .Z(n5820) );
  BUFFD0 U5815 ( .I(n5822), .Z(n5821) );
  BUFFD0 U5816 ( .I(n5823), .Z(n5822) );
  BUFFD0 U5817 ( .I(n5824), .Z(n5823) );
  BUFFD0 U5818 ( .I(n5825), .Z(n5824) );
  BUFFD0 U5819 ( .I(n5826), .Z(n5825) );
  BUFFD0 U5820 ( .I(n5827), .Z(n5826) );
  BUFFD0 U5821 ( .I(n5828), .Z(n5827) );
  BUFFD0 U5822 ( .I(n5829), .Z(n5828) );
  BUFFD0 U5823 ( .I(n5830), .Z(n5829) );
  BUFFD0 U5824 ( .I(n5831), .Z(n5830) );
  BUFFD0 U5825 ( .I(n5832), .Z(n5831) );
  BUFFD0 U5826 ( .I(n5833), .Z(n5832) );
  BUFFD0 U5827 ( .I(n5834), .Z(n5833) );
  BUFFD0 U5828 ( .I(n5835), .Z(n5834) );
  BUFFD0 U5829 ( .I(n5836), .Z(n5835) );
  BUFFD0 U5830 ( .I(n5837), .Z(n5836) );
  BUFFD0 U5831 ( .I(n5838), .Z(n5837) );
  BUFFD0 U5832 ( .I(n5839), .Z(n5838) );
  BUFFD0 U5833 ( .I(n5840), .Z(n5839) );
  BUFFD0 U5834 ( .I(n5841), .Z(n5840) );
  BUFFD0 U5835 ( .I(n5842), .Z(n5841) );
  BUFFD0 U5836 ( .I(n5843), .Z(n5842) );
  BUFFD0 U5837 ( .I(n5844), .Z(n5843) );
  BUFFD0 U5838 ( .I(n5845), .Z(n5844) );
  BUFFD0 U5839 ( .I(n5846), .Z(n5845) );
  BUFFD0 U5840 ( .I(n5847), .Z(n5846) );
  BUFFD0 U5841 ( .I(n5848), .Z(n5847) );
  BUFFD0 U5842 ( .I(n5849), .Z(n5848) );
  BUFFD0 U5843 ( .I(n5850), .Z(n5849) );
  BUFFD0 U5844 ( .I(n5851), .Z(n5850) );
  BUFFD0 U5845 ( .I(n5852), .Z(n5851) );
  BUFFD0 U5846 ( .I(n5853), .Z(n5852) );
  BUFFD0 U5847 ( .I(n5854), .Z(n5853) );
  BUFFD0 U5848 ( .I(n5855), .Z(n5854) );
  BUFFD0 U5849 ( .I(n5856), .Z(n5855) );
  BUFFD0 U5850 ( .I(n5857), .Z(n5856) );
  BUFFD0 U5851 ( .I(n5858), .Z(n5857) );
  BUFFD0 U5852 ( .I(n5859), .Z(n5858) );
  BUFFD0 U5853 ( .I(n5860), .Z(n5859) );
  BUFFD0 U5854 ( .I(n5861), .Z(n5860) );
  BUFFD0 U5855 ( .I(n5862), .Z(n5861) );
  BUFFD0 U5856 ( .I(n5863), .Z(n5862) );
  BUFFD0 U5857 ( .I(n5864), .Z(n5863) );
  BUFFD0 U5858 ( .I(n5865), .Z(n5864) );
  BUFFD0 U5859 ( .I(n5866), .Z(n5865) );
  BUFFD0 U5860 ( .I(n5867), .Z(n5866) );
  BUFFD0 U5861 ( .I(n8706), .Z(n5867) );
  BUFFD0 U5862 ( .I(n8703), .Z(n5868) );
  BUFFD0 U5863 ( .I(n5870), .Z(n5869) );
  BUFFD0 U5864 ( .I(n5871), .Z(n5870) );
  BUFFD0 U5865 ( .I(n5872), .Z(n5871) );
  BUFFD0 U5866 ( .I(n5873), .Z(n5872) );
  BUFFD0 U5867 ( .I(n5874), .Z(n5873) );
  BUFFD0 U5868 ( .I(n5875), .Z(n5874) );
  BUFFD0 U5869 ( .I(n5876), .Z(n5875) );
  BUFFD0 U5870 ( .I(n5877), .Z(n5876) );
  BUFFD0 U5871 ( .I(n5878), .Z(n5877) );
  BUFFD0 U5872 ( .I(n5879), .Z(n5878) );
  BUFFD0 U5873 ( .I(n5880), .Z(n5879) );
  BUFFD0 U5874 ( .I(n5881), .Z(n5880) );
  BUFFD0 U5875 ( .I(n5882), .Z(n5881) );
  BUFFD0 U5876 ( .I(n5883), .Z(n5882) );
  BUFFD0 U5877 ( .I(n5884), .Z(n5883) );
  BUFFD0 U5878 ( .I(n5885), .Z(n5884) );
  BUFFD0 U5879 ( .I(n5886), .Z(n5885) );
  BUFFD0 U5880 ( .I(n5887), .Z(n5886) );
  BUFFD0 U5881 ( .I(n5888), .Z(n5887) );
  BUFFD0 U5882 ( .I(n5889), .Z(n5888) );
  BUFFD0 U5883 ( .I(n5890), .Z(n5889) );
  BUFFD0 U5884 ( .I(n5891), .Z(n5890) );
  BUFFD0 U5885 ( .I(n5892), .Z(n5891) );
  BUFFD0 U5886 ( .I(n5893), .Z(n5892) );
  BUFFD0 U5887 ( .I(n5894), .Z(n5893) );
  BUFFD0 U5888 ( .I(n5895), .Z(n5894) );
  BUFFD0 U5889 ( .I(n5896), .Z(n5895) );
  BUFFD0 U5890 ( .I(n5897), .Z(n5896) );
  BUFFD0 U5891 ( .I(n5898), .Z(n5897) );
  BUFFD0 U5892 ( .I(n5899), .Z(n5898) );
  BUFFD0 U5893 ( .I(n5900), .Z(n5899) );
  BUFFD0 U5894 ( .I(n5901), .Z(n5900) );
  BUFFD0 U5895 ( .I(n5902), .Z(n5901) );
  BUFFD0 U5896 ( .I(n5903), .Z(n5902) );
  BUFFD0 U5897 ( .I(n5904), .Z(n5903) );
  BUFFD0 U5898 ( .I(n5905), .Z(n5904) );
  BUFFD0 U5899 ( .I(n5906), .Z(n5905) );
  BUFFD0 U5900 ( .I(n5907), .Z(n5906) );
  BUFFD0 U5901 ( .I(n5908), .Z(n5907) );
  BUFFD0 U5902 ( .I(n5909), .Z(n5908) );
  BUFFD0 U5903 ( .I(n5910), .Z(n5909) );
  BUFFD0 U5904 ( .I(n5911), .Z(n5910) );
  BUFFD0 U5905 ( .I(n5912), .Z(n5911) );
  BUFFD0 U5906 ( .I(n5913), .Z(n5912) );
  BUFFD0 U5907 ( .I(n5914), .Z(n5913) );
  BUFFD0 U5908 ( .I(n5915), .Z(n5914) );
  BUFFD0 U5909 ( .I(n5916), .Z(n5915) );
  BUFFD0 U5910 ( .I(n5917), .Z(n5916) );
  BUFFD0 U5911 ( .I(n5918), .Z(n5917) );
  BUFFD0 U5912 ( .I(n5919), .Z(n5918) );
  BUFFD0 U5913 ( .I(n5920), .Z(n5919) );
  BUFFD0 U5914 ( .I(n5921), .Z(n5920) );
  BUFFD0 U5915 ( .I(n5922), .Z(n5921) );
  BUFFD0 U5916 ( .I(n5923), .Z(n5922) );
  BUFFD0 U5917 ( .I(n5924), .Z(n5923) );
  BUFFD0 U5918 ( .I(n5925), .Z(n5924) );
  BUFFD0 U5919 ( .I(n5926), .Z(n5925) );
  BUFFD0 U5920 ( .I(n5927), .Z(n5926) );
  BUFFD0 U5921 ( .I(n5928), .Z(n5927) );
  BUFFD0 U5922 ( .I(n5929), .Z(n5928) );
  BUFFD0 U5923 ( .I(n5930), .Z(n5929) );
  BUFFD0 U5924 ( .I(n5931), .Z(n5930) );
  BUFFD0 U5925 ( .I(n5932), .Z(n5931) );
  BUFFD0 U5926 ( .I(n5933), .Z(n5932) );
  BUFFD0 U5927 ( .I(n5934), .Z(n5933) );
  BUFFD0 U5928 ( .I(n5935), .Z(n5934) );
  BUFFD0 U5929 ( .I(n5936), .Z(n5935) );
  BUFFD0 U5930 ( .I(n5937), .Z(n5936) );
  BUFFD0 U5931 ( .I(n5938), .Z(n5937) );
  BUFFD0 U5932 ( .I(n5939), .Z(n5938) );
  BUFFD0 U5933 ( .I(n5940), .Z(n5939) );
  BUFFD0 U5934 ( .I(n5941), .Z(n5940) );
  BUFFD0 U5935 ( .I(n5942), .Z(n5941) );
  BUFFD0 U5936 ( .I(n5943), .Z(n5942) );
  BUFFD0 U5937 ( .I(n5944), .Z(n5943) );
  BUFFD0 U5938 ( .I(n5945), .Z(n5944) );
  BUFFD0 U5939 ( .I(n5946), .Z(n5945) );
  BUFFD0 U5940 ( .I(n5947), .Z(n5946) );
  BUFFD0 U5941 ( .I(n5948), .Z(n5947) );
  BUFFD0 U5942 ( .I(n5949), .Z(n5948) );
  BUFFD0 U5943 ( .I(n5950), .Z(n5949) );
  BUFFD0 U5944 ( .I(n5951), .Z(n5950) );
  BUFFD0 U5945 ( .I(n5952), .Z(n5951) );
  BUFFD0 U5946 ( .I(n5953), .Z(n5952) );
  BUFFD0 U5947 ( .I(n5954), .Z(n5953) );
  BUFFD0 U5948 ( .I(n5955), .Z(n5954) );
  BUFFD0 U5949 ( .I(n5956), .Z(n5955) );
  BUFFD0 U5950 ( .I(n5957), .Z(n5956) );
  BUFFD0 U5951 ( .I(n5958), .Z(n5957) );
  BUFFD0 U5952 ( .I(n5959), .Z(n5958) );
  BUFFD0 U5953 ( .I(n5960), .Z(n5959) );
  BUFFD0 U5954 ( .I(n5961), .Z(n5960) );
  BUFFD0 U5955 ( .I(n5962), .Z(n5961) );
  BUFFD0 U5956 ( .I(n5963), .Z(n5962) );
  BUFFD0 U5957 ( .I(n5964), .Z(n5963) );
  BUFFD0 U5958 ( .I(n5965), .Z(n5964) );
  BUFFD0 U5959 ( .I(n5966), .Z(n5965) );
  BUFFD0 U5960 ( .I(n5967), .Z(n5966) );
  BUFFD0 U5961 ( .I(n5968), .Z(n5967) );
  BUFFD0 U5962 ( .I(n5969), .Z(n5968) );
  BUFFD0 U5963 ( .I(n5970), .Z(n5969) );
  BUFFD0 U5964 ( .I(n5971), .Z(n5970) );
  BUFFD0 U5965 ( .I(n5972), .Z(n5971) );
  BUFFD0 U5966 ( .I(n5973), .Z(n5972) );
  BUFFD0 U5967 ( .I(n5974), .Z(n5973) );
  BUFFD0 U5968 ( .I(n5975), .Z(n5974) );
  BUFFD0 U5969 ( .I(n5976), .Z(n5975) );
  BUFFD0 U5970 ( .I(n5977), .Z(n5976) );
  BUFFD0 U5971 ( .I(n5978), .Z(n5977) );
  BUFFD0 U5972 ( .I(n5979), .Z(n5978) );
  BUFFD0 U5973 ( .I(n5980), .Z(n5979) );
  BUFFD0 U5974 ( .I(n5981), .Z(n5980) );
  BUFFD0 U5975 ( .I(n5982), .Z(n5981) );
  BUFFD0 U5976 ( .I(n5983), .Z(n5982) );
  BUFFD0 U5977 ( .I(n5984), .Z(n5983) );
  BUFFD0 U5978 ( .I(n5985), .Z(n5984) );
  BUFFD0 U5979 ( .I(n5986), .Z(n5985) );
  BUFFD0 U5980 ( .I(n5987), .Z(n5986) );
  BUFFD0 U5981 ( .I(n5988), .Z(n5987) );
  BUFFD0 U5982 ( .I(n5989), .Z(n5988) );
  BUFFD0 U5983 ( .I(n5990), .Z(n5989) );
  BUFFD0 U5984 ( .I(n5991), .Z(n5990) );
  BUFFD0 U5985 ( .I(n5992), .Z(n5991) );
  BUFFD0 U5986 ( .I(n5993), .Z(n5992) );
  BUFFD0 U5987 ( .I(n5994), .Z(n5993) );
  BUFFD0 U5988 ( .I(n5995), .Z(n5994) );
  BUFFD0 U5989 ( .I(n5996), .Z(n5995) );
  BUFFD0 U5990 ( .I(n5997), .Z(n5996) );
  BUFFD0 U5991 ( .I(n5998), .Z(n5997) );
  BUFFD0 U5992 ( .I(n5999), .Z(n5998) );
  BUFFD0 U5993 ( .I(n6000), .Z(n5999) );
  BUFFD0 U5994 ( .I(n6001), .Z(n6000) );
  BUFFD0 U5995 ( .I(n6002), .Z(n6001) );
  BUFFD0 U5996 ( .I(n6003), .Z(n6002) );
  BUFFD0 U5997 ( .I(n6004), .Z(n6003) );
  BUFFD0 U5998 ( .I(n6005), .Z(n6004) );
  BUFFD0 U5999 ( .I(n6006), .Z(n6005) );
  BUFFD0 U6000 ( .I(n6007), .Z(n6006) );
  BUFFD0 U6001 ( .I(n6008), .Z(n6007) );
  BUFFD0 U6002 ( .I(n6009), .Z(n6008) );
  BUFFD0 U6003 ( .I(n6010), .Z(n6009) );
  BUFFD0 U6004 ( .I(n6011), .Z(n6010) );
  BUFFD0 U6005 ( .I(n6012), .Z(n6011) );
  BUFFD0 U6006 ( .I(n6013), .Z(n6012) );
  BUFFD0 U6007 ( .I(n6014), .Z(n6013) );
  BUFFD0 U6008 ( .I(n6015), .Z(n6014) );
  BUFFD0 U6009 ( .I(n6016), .Z(n6015) );
  BUFFD0 U6010 ( .I(n6017), .Z(n6016) );
  BUFFD0 U6011 ( .I(n6018), .Z(n6017) );
  BUFFD0 U6012 ( .I(n6019), .Z(n6018) );
  BUFFD0 U6013 ( .I(n6020), .Z(n6019) );
  BUFFD0 U6014 ( .I(n6021), .Z(n6020) );
  BUFFD0 U6015 ( .I(n6022), .Z(n6021) );
  BUFFD0 U6016 ( .I(n6023), .Z(n6022) );
  BUFFD0 U6017 ( .I(n6024), .Z(n6023) );
  BUFFD0 U6018 ( .I(n6025), .Z(n6024) );
  BUFFD0 U6019 ( .I(n6026), .Z(n6025) );
  BUFFD0 U6020 ( .I(n6027), .Z(n6026) );
  BUFFD0 U6021 ( .I(n6028), .Z(n6027) );
  BUFFD0 U6022 ( .I(n6029), .Z(n6028) );
  BUFFD0 U6023 ( .I(n6030), .Z(n6029) );
  BUFFD0 U6024 ( .I(n6031), .Z(n6030) );
  BUFFD0 U6025 ( .I(n6032), .Z(n6031) );
  BUFFD0 U6026 ( .I(n6033), .Z(n6032) );
  BUFFD0 U6027 ( .I(n6034), .Z(n6033) );
  BUFFD0 U6028 ( .I(n6035), .Z(n6034) );
  BUFFD0 U6029 ( .I(n6036), .Z(n6035) );
  BUFFD0 U6030 ( .I(n6037), .Z(n6036) );
  BUFFD0 U6031 ( .I(n6038), .Z(n6037) );
  BUFFD0 U6032 ( .I(n6039), .Z(n6038) );
  BUFFD0 U6033 ( .I(n6040), .Z(n6039) );
  BUFFD0 U6034 ( .I(n6041), .Z(n6040) );
  BUFFD0 U6035 ( .I(n6042), .Z(n6041) );
  BUFFD0 U6036 ( .I(n6043), .Z(n6042) );
  BUFFD0 U6037 ( .I(n6044), .Z(n6043) );
  BUFFD0 U6038 ( .I(n6045), .Z(n6044) );
  BUFFD0 U6039 ( .I(n6046), .Z(n6045) );
  BUFFD0 U6040 ( .I(n8704), .Z(n6046) );
  BUFFD0 U6041 ( .I(n8701), .Z(n6047) );
  BUFFD0 U6042 ( .I(n6049), .Z(n6048) );
  BUFFD0 U6043 ( .I(n6050), .Z(n6049) );
  BUFFD0 U6044 ( .I(n6051), .Z(n6050) );
  BUFFD0 U6045 ( .I(n6052), .Z(n6051) );
  BUFFD0 U6046 ( .I(n6053), .Z(n6052) );
  BUFFD0 U6047 ( .I(n6054), .Z(n6053) );
  BUFFD0 U6048 ( .I(n6055), .Z(n6054) );
  BUFFD0 U6049 ( .I(n6056), .Z(n6055) );
  BUFFD0 U6050 ( .I(n6057), .Z(n6056) );
  BUFFD0 U6051 ( .I(n6058), .Z(n6057) );
  BUFFD0 U6052 ( .I(n6059), .Z(n6058) );
  BUFFD0 U6053 ( .I(n6060), .Z(n6059) );
  BUFFD0 U6054 ( .I(n6061), .Z(n6060) );
  BUFFD0 U6055 ( .I(n6062), .Z(n6061) );
  BUFFD0 U6056 ( .I(n6063), .Z(n6062) );
  BUFFD0 U6057 ( .I(n6064), .Z(n6063) );
  BUFFD0 U6058 ( .I(n6065), .Z(n6064) );
  BUFFD0 U6059 ( .I(n6066), .Z(n6065) );
  BUFFD0 U6060 ( .I(n6067), .Z(n6066) );
  BUFFD0 U6061 ( .I(n6068), .Z(n6067) );
  BUFFD0 U6062 ( .I(n6069), .Z(n6068) );
  BUFFD0 U6063 ( .I(n6070), .Z(n6069) );
  BUFFD0 U6064 ( .I(n6071), .Z(n6070) );
  BUFFD0 U6065 ( .I(n6072), .Z(n6071) );
  BUFFD0 U6066 ( .I(n6073), .Z(n6072) );
  BUFFD0 U6067 ( .I(n6074), .Z(n6073) );
  BUFFD0 U6068 ( .I(n6075), .Z(n6074) );
  BUFFD0 U6069 ( .I(n6076), .Z(n6075) );
  BUFFD0 U6070 ( .I(n6077), .Z(n6076) );
  BUFFD0 U6071 ( .I(n6078), .Z(n6077) );
  BUFFD0 U6072 ( .I(n6079), .Z(n6078) );
  BUFFD0 U6073 ( .I(n6080), .Z(n6079) );
  BUFFD0 U6074 ( .I(n6081), .Z(n6080) );
  BUFFD0 U6075 ( .I(n6082), .Z(n6081) );
  BUFFD0 U6076 ( .I(n6083), .Z(n6082) );
  BUFFD0 U6077 ( .I(n6084), .Z(n6083) );
  BUFFD0 U6078 ( .I(n6085), .Z(n6084) );
  BUFFD0 U6079 ( .I(n6086), .Z(n6085) );
  BUFFD0 U6080 ( .I(n6087), .Z(n6086) );
  BUFFD0 U6081 ( .I(n6088), .Z(n6087) );
  BUFFD0 U6082 ( .I(n6089), .Z(n6088) );
  BUFFD0 U6083 ( .I(n6090), .Z(n6089) );
  BUFFD0 U6084 ( .I(n6091), .Z(n6090) );
  BUFFD0 U6085 ( .I(n6092), .Z(n6091) );
  BUFFD0 U6086 ( .I(n6093), .Z(n6092) );
  BUFFD0 U6087 ( .I(n6094), .Z(n6093) );
  BUFFD0 U6088 ( .I(n6095), .Z(n6094) );
  BUFFD0 U6089 ( .I(n6096), .Z(n6095) );
  BUFFD0 U6090 ( .I(n6097), .Z(n6096) );
  BUFFD0 U6091 ( .I(n6098), .Z(n6097) );
  BUFFD0 U6092 ( .I(n6099), .Z(n6098) );
  BUFFD0 U6093 ( .I(n6100), .Z(n6099) );
  BUFFD0 U6094 ( .I(n6101), .Z(n6100) );
  BUFFD0 U6095 ( .I(n6102), .Z(n6101) );
  BUFFD0 U6096 ( .I(n6103), .Z(n6102) );
  BUFFD0 U6097 ( .I(n6104), .Z(n6103) );
  BUFFD0 U6098 ( .I(n6105), .Z(n6104) );
  BUFFD0 U6099 ( .I(n6106), .Z(n6105) );
  BUFFD0 U6100 ( .I(n6107), .Z(n6106) );
  BUFFD0 U6101 ( .I(n6108), .Z(n6107) );
  BUFFD0 U6102 ( .I(n6109), .Z(n6108) );
  BUFFD0 U6103 ( .I(n6110), .Z(n6109) );
  BUFFD0 U6104 ( .I(n6111), .Z(n6110) );
  BUFFD0 U6105 ( .I(n6112), .Z(n6111) );
  BUFFD0 U6106 ( .I(n6113), .Z(n6112) );
  BUFFD0 U6107 ( .I(n6114), .Z(n6113) );
  BUFFD0 U6108 ( .I(n6115), .Z(n6114) );
  BUFFD0 U6109 ( .I(n6116), .Z(n6115) );
  BUFFD0 U6110 ( .I(n6117), .Z(n6116) );
  BUFFD0 U6111 ( .I(n6118), .Z(n6117) );
  BUFFD0 U6112 ( .I(n6119), .Z(n6118) );
  BUFFD0 U6113 ( .I(n6120), .Z(n6119) );
  BUFFD0 U6114 ( .I(n6121), .Z(n6120) );
  BUFFD0 U6115 ( .I(n6122), .Z(n6121) );
  BUFFD0 U6116 ( .I(n6123), .Z(n6122) );
  BUFFD0 U6117 ( .I(n6124), .Z(n6123) );
  BUFFD0 U6118 ( .I(n6125), .Z(n6124) );
  BUFFD0 U6119 ( .I(n6126), .Z(n6125) );
  BUFFD0 U6120 ( .I(n6127), .Z(n6126) );
  BUFFD0 U6121 ( .I(n6128), .Z(n6127) );
  BUFFD0 U6122 ( .I(n6129), .Z(n6128) );
  BUFFD0 U6123 ( .I(n6130), .Z(n6129) );
  BUFFD0 U6124 ( .I(n6131), .Z(n6130) );
  BUFFD0 U6125 ( .I(n6132), .Z(n6131) );
  BUFFD0 U6126 ( .I(n6133), .Z(n6132) );
  BUFFD0 U6127 ( .I(n6134), .Z(n6133) );
  BUFFD0 U6128 ( .I(n6135), .Z(n6134) );
  BUFFD0 U6129 ( .I(n6136), .Z(n6135) );
  BUFFD0 U6130 ( .I(n6137), .Z(n6136) );
  BUFFD0 U6131 ( .I(n6138), .Z(n6137) );
  BUFFD0 U6132 ( .I(n6139), .Z(n6138) );
  BUFFD0 U6133 ( .I(n6140), .Z(n6139) );
  BUFFD0 U6134 ( .I(n6141), .Z(n6140) );
  BUFFD0 U6135 ( .I(n6142), .Z(n6141) );
  BUFFD0 U6136 ( .I(n6143), .Z(n6142) );
  BUFFD0 U6137 ( .I(n6144), .Z(n6143) );
  BUFFD0 U6138 ( .I(n6145), .Z(n6144) );
  BUFFD0 U6139 ( .I(n6146), .Z(n6145) );
  BUFFD0 U6140 ( .I(n6147), .Z(n6146) );
  BUFFD0 U6141 ( .I(n6148), .Z(n6147) );
  BUFFD0 U6142 ( .I(n6149), .Z(n6148) );
  BUFFD0 U6143 ( .I(n6150), .Z(n6149) );
  BUFFD0 U6144 ( .I(n6151), .Z(n6150) );
  BUFFD0 U6145 ( .I(n6152), .Z(n6151) );
  BUFFD0 U6146 ( .I(n6153), .Z(n6152) );
  BUFFD0 U6147 ( .I(n6154), .Z(n6153) );
  BUFFD0 U6148 ( .I(n6155), .Z(n6154) );
  BUFFD0 U6149 ( .I(n6156), .Z(n6155) );
  BUFFD0 U6150 ( .I(n6157), .Z(n6156) );
  BUFFD0 U6151 ( .I(n6158), .Z(n6157) );
  BUFFD0 U6152 ( .I(n6159), .Z(n6158) );
  BUFFD0 U6153 ( .I(n6160), .Z(n6159) );
  BUFFD0 U6154 ( .I(n6161), .Z(n6160) );
  BUFFD0 U6155 ( .I(n6162), .Z(n6161) );
  BUFFD0 U6156 ( .I(n6163), .Z(n6162) );
  BUFFD0 U6157 ( .I(n6164), .Z(n6163) );
  BUFFD0 U6158 ( .I(n6165), .Z(n6164) );
  BUFFD0 U6159 ( .I(n6166), .Z(n6165) );
  BUFFD0 U6160 ( .I(n6167), .Z(n6166) );
  BUFFD0 U6161 ( .I(n6168), .Z(n6167) );
  BUFFD0 U6162 ( .I(n6169), .Z(n6168) );
  BUFFD0 U6163 ( .I(n6170), .Z(n6169) );
  BUFFD0 U6164 ( .I(n6171), .Z(n6170) );
  BUFFD0 U6165 ( .I(n6172), .Z(n6171) );
  BUFFD0 U6166 ( .I(n6173), .Z(n6172) );
  BUFFD0 U6167 ( .I(n6174), .Z(n6173) );
  BUFFD0 U6168 ( .I(n6175), .Z(n6174) );
  BUFFD0 U6169 ( .I(n6176), .Z(n6175) );
  BUFFD0 U6170 ( .I(n6177), .Z(n6176) );
  BUFFD0 U6171 ( .I(n6178), .Z(n6177) );
  BUFFD0 U6172 ( .I(n6179), .Z(n6178) );
  BUFFD0 U6173 ( .I(n6180), .Z(n6179) );
  BUFFD0 U6174 ( .I(n6181), .Z(n6180) );
  BUFFD0 U6175 ( .I(n6182), .Z(n6181) );
  BUFFD0 U6176 ( .I(n6183), .Z(n6182) );
  BUFFD0 U6177 ( .I(n6184), .Z(n6183) );
  BUFFD0 U6178 ( .I(n6185), .Z(n6184) );
  BUFFD0 U6179 ( .I(n6186), .Z(n6185) );
  BUFFD0 U6180 ( .I(n6187), .Z(n6186) );
  BUFFD0 U6181 ( .I(n6188), .Z(n6187) );
  BUFFD0 U6182 ( .I(n6189), .Z(n6188) );
  BUFFD0 U6183 ( .I(n6190), .Z(n6189) );
  BUFFD0 U6184 ( .I(n6191), .Z(n6190) );
  BUFFD0 U6185 ( .I(n6192), .Z(n6191) );
  BUFFD0 U6186 ( .I(n6193), .Z(n6192) );
  BUFFD0 U6187 ( .I(n6194), .Z(n6193) );
  BUFFD0 U6188 ( .I(n6195), .Z(n6194) );
  BUFFD0 U6189 ( .I(n6196), .Z(n6195) );
  BUFFD0 U6190 ( .I(n6197), .Z(n6196) );
  BUFFD0 U6191 ( .I(n6198), .Z(n6197) );
  BUFFD0 U6192 ( .I(n6199), .Z(n6198) );
  BUFFD0 U6193 ( .I(n6200), .Z(n6199) );
  BUFFD0 U6194 ( .I(n6201), .Z(n6200) );
  BUFFD0 U6195 ( .I(n6202), .Z(n6201) );
  BUFFD0 U6196 ( .I(n6203), .Z(n6202) );
  BUFFD0 U6197 ( .I(n6204), .Z(n6203) );
  BUFFD0 U6198 ( .I(n6205), .Z(n6204) );
  BUFFD0 U6199 ( .I(n6206), .Z(n6205) );
  BUFFD0 U6200 ( .I(n6207), .Z(n6206) );
  BUFFD0 U6201 ( .I(n6208), .Z(n6207) );
  BUFFD0 U6202 ( .I(n6209), .Z(n6208) );
  BUFFD0 U6203 ( .I(n6210), .Z(n6209) );
  BUFFD0 U6204 ( .I(n6211), .Z(n6210) );
  BUFFD0 U6205 ( .I(n6212), .Z(n6211) );
  BUFFD0 U6206 ( .I(n6213), .Z(n6212) );
  BUFFD0 U6207 ( .I(n6214), .Z(n6213) );
  BUFFD0 U6208 ( .I(n6215), .Z(n6214) );
  BUFFD0 U6209 ( .I(n6216), .Z(n6215) );
  BUFFD0 U6210 ( .I(n6217), .Z(n6216) );
  BUFFD0 U6211 ( .I(n6218), .Z(n6217) );
  BUFFD0 U6212 ( .I(n6219), .Z(n6218) );
  BUFFD0 U6213 ( .I(n6220), .Z(n6219) );
  BUFFD0 U6214 ( .I(n6221), .Z(n6220) );
  BUFFD0 U6215 ( .I(n6222), .Z(n6221) );
  BUFFD0 U6216 ( .I(n6223), .Z(n6222) );
  BUFFD0 U6217 ( .I(n8702), .Z(n6223) );
  BUFFD0 U6218 ( .I(n6225), .Z(n6224) );
  BUFFD0 U6219 ( .I(n6226), .Z(n6225) );
  BUFFD0 U6220 ( .I(n6227), .Z(n6226) );
  BUFFD0 U6221 ( .I(n6228), .Z(n6227) );
  BUFFD0 U6222 ( .I(n6229), .Z(n6228) );
  BUFFD0 U6223 ( .I(n6230), .Z(n6229) );
  BUFFD0 U6224 ( .I(n6231), .Z(n6230) );
  BUFFD0 U6225 ( .I(n6232), .Z(n6231) );
  BUFFD0 U6226 ( .I(n6233), .Z(n6232) );
  BUFFD0 U6227 ( .I(n6234), .Z(n6233) );
  BUFFD0 U6228 ( .I(n6235), .Z(n6234) );
  BUFFD0 U6229 ( .I(n6236), .Z(n6235) );
  BUFFD0 U6230 ( .I(n6237), .Z(n6236) );
  BUFFD0 U6231 ( .I(n6238), .Z(n6237) );
  BUFFD0 U6232 ( .I(n6239), .Z(n6238) );
  BUFFD0 U6233 ( .I(n6240), .Z(n6239) );
  BUFFD0 U6234 ( .I(n6241), .Z(n6240) );
  BUFFD0 U6235 ( .I(n6242), .Z(n6241) );
  BUFFD0 U6236 ( .I(n6243), .Z(n6242) );
  BUFFD0 U6237 ( .I(n6244), .Z(n6243) );
  BUFFD0 U6238 ( .I(n6245), .Z(n6244) );
  BUFFD0 U6239 ( .I(n6246), .Z(n6245) );
  BUFFD0 U6240 ( .I(n6247), .Z(n6246) );
  BUFFD0 U6241 ( .I(n6248), .Z(n6247) );
  BUFFD0 U6242 ( .I(n6249), .Z(n6248) );
  BUFFD0 U6243 ( .I(n6250), .Z(n6249) );
  BUFFD0 U6244 ( .I(n6251), .Z(n6250) );
  BUFFD0 U6245 ( .I(n6252), .Z(n6251) );
  BUFFD0 U6246 ( .I(n6253), .Z(n6252) );
  BUFFD0 U6247 ( .I(n6254), .Z(n6253) );
  BUFFD0 U6248 ( .I(n6255), .Z(n6254) );
  BUFFD0 U6249 ( .I(n6256), .Z(n6255) );
  BUFFD0 U6250 ( .I(n6257), .Z(n6256) );
  BUFFD0 U6251 ( .I(n6258), .Z(n6257) );
  BUFFD0 U6252 ( .I(n6259), .Z(n6258) );
  BUFFD0 U6253 ( .I(n6260), .Z(n6259) );
  BUFFD0 U6254 ( .I(n6261), .Z(n6260) );
  BUFFD0 U6255 ( .I(n6262), .Z(n6261) );
  BUFFD0 U6256 ( .I(n6263), .Z(n6262) );
  BUFFD0 U6257 ( .I(n6264), .Z(n6263) );
  BUFFD0 U6258 ( .I(n6265), .Z(n6264) );
  BUFFD0 U6259 ( .I(n6266), .Z(n6265) );
  BUFFD0 U6260 ( .I(n6267), .Z(n6266) );
  BUFFD0 U6261 ( .I(n6268), .Z(n6267) );
  BUFFD0 U6262 ( .I(n6269), .Z(n6268) );
  BUFFD0 U6263 ( .I(n6270), .Z(n6269) );
  BUFFD0 U6264 ( .I(n6271), .Z(n6270) );
  BUFFD0 U6265 ( .I(n6272), .Z(n6271) );
  BUFFD0 U6266 ( .I(n6273), .Z(n6272) );
  BUFFD0 U6267 ( .I(n6274), .Z(n6273) );
  BUFFD0 U6268 ( .I(n6275), .Z(n6274) );
  BUFFD0 U6269 ( .I(n6276), .Z(n6275) );
  BUFFD0 U6270 ( .I(n6277), .Z(n6276) );
  BUFFD0 U6271 ( .I(n6278), .Z(n6277) );
  BUFFD0 U6272 ( .I(n6279), .Z(n6278) );
  BUFFD0 U6273 ( .I(n6280), .Z(n6279) );
  BUFFD0 U6274 ( .I(n6281), .Z(n6280) );
  BUFFD0 U6275 ( .I(n6282), .Z(n6281) );
  BUFFD0 U6276 ( .I(n6283), .Z(n6282) );
  BUFFD0 U6277 ( .I(n6284), .Z(n6283) );
  BUFFD0 U6278 ( .I(n6285), .Z(n6284) );
  BUFFD0 U6279 ( .I(n6286), .Z(n6285) );
  BUFFD0 U6280 ( .I(n6287), .Z(n6286) );
  BUFFD0 U6281 ( .I(n6288), .Z(n6287) );
  BUFFD0 U6282 ( .I(n6289), .Z(n6288) );
  BUFFD0 U6283 ( .I(n6290), .Z(n6289) );
  BUFFD0 U6284 ( .I(n6291), .Z(n6290) );
  BUFFD0 U6285 ( .I(n6292), .Z(n6291) );
  BUFFD0 U6286 ( .I(n6293), .Z(n6292) );
  BUFFD0 U6287 ( .I(n6294), .Z(n6293) );
  BUFFD0 U6288 ( .I(n6295), .Z(n6294) );
  BUFFD0 U6289 ( .I(n6296), .Z(n6295) );
  BUFFD0 U6290 ( .I(n6297), .Z(n6296) );
  BUFFD0 U6291 ( .I(n6298), .Z(n6297) );
  BUFFD0 U6292 ( .I(n6299), .Z(n6298) );
  BUFFD0 U6293 ( .I(n6300), .Z(n6299) );
  BUFFD0 U6294 ( .I(n6301), .Z(n6300) );
  BUFFD0 U6295 ( .I(n6302), .Z(n6301) );
  BUFFD0 U6296 ( .I(n6303), .Z(n6302) );
  BUFFD0 U6297 ( .I(n6304), .Z(n6303) );
  BUFFD0 U6298 ( .I(n6305), .Z(n6304) );
  BUFFD0 U6299 ( .I(n6306), .Z(n6305) );
  BUFFD0 U6300 ( .I(n6307), .Z(n6306) );
  BUFFD0 U6301 ( .I(n6308), .Z(n6307) );
  BUFFD0 U6302 ( .I(n6309), .Z(n6308) );
  BUFFD0 U6303 ( .I(n6310), .Z(n6309) );
  BUFFD0 U6304 ( .I(n6311), .Z(n6310) );
  BUFFD0 U6305 ( .I(n6312), .Z(n6311) );
  BUFFD0 U6306 ( .I(n6313), .Z(n6312) );
  BUFFD0 U6307 ( .I(n6314), .Z(n6313) );
  BUFFD0 U6308 ( .I(n6315), .Z(n6314) );
  BUFFD0 U6309 ( .I(n6316), .Z(n6315) );
  BUFFD0 U6310 ( .I(n6317), .Z(n6316) );
  BUFFD0 U6311 ( .I(n6318), .Z(n6317) );
  BUFFD0 U6312 ( .I(n6319), .Z(n6318) );
  BUFFD0 U6313 ( .I(n6320), .Z(n6319) );
  BUFFD0 U6314 ( .I(n6321), .Z(n6320) );
  BUFFD0 U6315 ( .I(n6322), .Z(n6321) );
  BUFFD0 U6316 ( .I(n6323), .Z(n6322) );
  BUFFD0 U6317 ( .I(n6324), .Z(n6323) );
  BUFFD0 U6318 ( .I(n6325), .Z(n6324) );
  BUFFD0 U6319 ( .I(n6326), .Z(n6325) );
  BUFFD0 U6320 ( .I(n6327), .Z(n6326) );
  BUFFD0 U6321 ( .I(n6328), .Z(n6327) );
  BUFFD0 U6322 ( .I(n6329), .Z(n6328) );
  BUFFD0 U6323 ( .I(n6330), .Z(n6329) );
  BUFFD0 U6324 ( .I(n6331), .Z(n6330) );
  BUFFD0 U6325 ( .I(n6332), .Z(n6331) );
  BUFFD0 U6326 ( .I(n6333), .Z(n6332) );
  BUFFD0 U6327 ( .I(n6334), .Z(n6333) );
  BUFFD0 U6328 ( .I(n6335), .Z(n6334) );
  BUFFD0 U6329 ( .I(n6336), .Z(n6335) );
  BUFFD0 U6330 ( .I(n6337), .Z(n6336) );
  BUFFD0 U6331 ( .I(n6338), .Z(n6337) );
  BUFFD0 U6332 ( .I(n6339), .Z(n6338) );
  BUFFD0 U6333 ( .I(n6340), .Z(n6339) );
  BUFFD0 U6334 ( .I(n6341), .Z(n6340) );
  BUFFD0 U6335 ( .I(n6342), .Z(n6341) );
  BUFFD0 U6336 ( .I(n6343), .Z(n6342) );
  BUFFD0 U6337 ( .I(n6344), .Z(n6343) );
  BUFFD0 U6338 ( .I(n6345), .Z(n6344) );
  BUFFD0 U6339 ( .I(n6346), .Z(n6345) );
  BUFFD0 U6340 ( .I(n6347), .Z(n6346) );
  BUFFD0 U6341 ( .I(n6348), .Z(n6347) );
  BUFFD0 U6342 ( .I(n6349), .Z(n6348) );
  BUFFD0 U6343 ( .I(n6350), .Z(n6349) );
  BUFFD0 U6344 ( .I(n6351), .Z(n6350) );
  BUFFD0 U6345 ( .I(n6352), .Z(n6351) );
  BUFFD0 U6346 ( .I(n6353), .Z(n6352) );
  BUFFD0 U6347 ( .I(n6354), .Z(n6353) );
  BUFFD0 U6348 ( .I(n6355), .Z(n6354) );
  BUFFD0 U6349 ( .I(n6356), .Z(n6355) );
  BUFFD0 U6350 ( .I(n6357), .Z(n6356) );
  BUFFD0 U6351 ( .I(n6358), .Z(n6357) );
  BUFFD0 U6352 ( .I(n6359), .Z(n6358) );
  BUFFD0 U6353 ( .I(n6360), .Z(n6359) );
  BUFFD0 U6354 ( .I(n6361), .Z(n6360) );
  BUFFD0 U6355 ( .I(n6362), .Z(n6361) );
  BUFFD0 U6356 ( .I(n6363), .Z(n6362) );
  BUFFD0 U6357 ( .I(n6364), .Z(n6363) );
  BUFFD0 U6358 ( .I(n6365), .Z(n6364) );
  BUFFD0 U6359 ( .I(n6367), .Z(n6365) );
  BUFFD0 U6360 ( .I(n2217), .Z(n6366) );
  BUFFD0 U6361 ( .I(n6368), .Z(n6367) );
  BUFFD0 U6362 ( .I(n6369), .Z(n6368) );
  BUFFD0 U6363 ( .I(n6370), .Z(n6369) );
  BUFFD0 U6364 ( .I(n6371), .Z(n6370) );
  BUFFD0 U6365 ( .I(n6372), .Z(n6371) );
  BUFFD0 U6366 ( .I(n6373), .Z(n6372) );
  BUFFD0 U6367 ( .I(n6374), .Z(n6373) );
  BUFFD0 U6368 ( .I(n6375), .Z(n6374) );
  BUFFD0 U6369 ( .I(n6376), .Z(n6375) );
  BUFFD0 U6370 ( .I(n6377), .Z(n6376) );
  BUFFD0 U6371 ( .I(n6378), .Z(n6377) );
  BUFFD0 U6372 ( .I(n6379), .Z(n6378) );
  BUFFD0 U6373 ( .I(n6380), .Z(n6379) );
  BUFFD0 U6374 ( .I(n6381), .Z(n6380) );
  BUFFD0 U6375 ( .I(n6382), .Z(n6381) );
  BUFFD0 U6376 ( .I(n6383), .Z(n6382) );
  BUFFD0 U6377 ( .I(n6384), .Z(n6383) );
  BUFFD0 U6378 ( .I(n6385), .Z(n6384) );
  BUFFD0 U6379 ( .I(n6386), .Z(n6385) );
  BUFFD0 U6380 ( .I(n6387), .Z(n6386) );
  BUFFD0 U6381 ( .I(n6388), .Z(n6387) );
  BUFFD0 U6382 ( .I(n6389), .Z(n6388) );
  BUFFD0 U6383 ( .I(n6390), .Z(n6389) );
  BUFFD0 U6384 ( .I(n6391), .Z(n6390) );
  BUFFD0 U6385 ( .I(n6392), .Z(n6391) );
  BUFFD0 U6386 ( .I(n6393), .Z(n6392) );
  BUFFD0 U6387 ( .I(n6394), .Z(n6393) );
  BUFFD0 U6388 ( .I(n6395), .Z(n6394) );
  BUFFD0 U6389 ( .I(n6396), .Z(n6395) );
  BUFFD0 U6390 ( .I(n6397), .Z(n6396) );
  BUFFD0 U6391 ( .I(n6398), .Z(n6397) );
  BUFFD0 U6392 ( .I(n6399), .Z(n6398) );
  BUFFD0 U6393 ( .I(n8699), .Z(n6399) );
  BUFFD0 U6394 ( .I(n8696), .Z(n6400) );
  BUFFD0 U6395 ( .I(n6402), .Z(n6401) );
  BUFFD0 U6396 ( .I(n6403), .Z(n6402) );
  BUFFD0 U6397 ( .I(n6404), .Z(n6403) );
  BUFFD0 U6398 ( .I(n6405), .Z(n6404) );
  BUFFD0 U6399 ( .I(n6406), .Z(n6405) );
  BUFFD0 U6400 ( .I(n6407), .Z(n6406) );
  BUFFD0 U6401 ( .I(n6408), .Z(n6407) );
  BUFFD0 U6402 ( .I(n6409), .Z(n6408) );
  BUFFD0 U6403 ( .I(n6410), .Z(n6409) );
  BUFFD0 U6404 ( .I(n6411), .Z(n6410) );
  BUFFD0 U6405 ( .I(n6412), .Z(n6411) );
  BUFFD0 U6406 ( .I(n6413), .Z(n6412) );
  BUFFD0 U6407 ( .I(n6414), .Z(n6413) );
  BUFFD0 U6408 ( .I(n6415), .Z(n6414) );
  BUFFD0 U6409 ( .I(n6416), .Z(n6415) );
  BUFFD0 U6410 ( .I(n6417), .Z(n6416) );
  BUFFD0 U6411 ( .I(n6418), .Z(n6417) );
  BUFFD0 U6412 ( .I(n6419), .Z(n6418) );
  BUFFD0 U6413 ( .I(n6420), .Z(n6419) );
  BUFFD0 U6414 ( .I(n6421), .Z(n6420) );
  BUFFD0 U6415 ( .I(n6422), .Z(n6421) );
  BUFFD0 U6416 ( .I(n6423), .Z(n6422) );
  BUFFD0 U6417 ( .I(n6424), .Z(n6423) );
  BUFFD0 U6418 ( .I(n6425), .Z(n6424) );
  BUFFD0 U6419 ( .I(n6426), .Z(n6425) );
  BUFFD0 U6420 ( .I(n6427), .Z(n6426) );
  BUFFD0 U6421 ( .I(n6428), .Z(n6427) );
  BUFFD0 U6422 ( .I(n6429), .Z(n6428) );
  BUFFD0 U6423 ( .I(n6430), .Z(n6429) );
  BUFFD0 U6424 ( .I(n6431), .Z(n6430) );
  BUFFD0 U6425 ( .I(n6432), .Z(n6431) );
  BUFFD0 U6426 ( .I(n6433), .Z(n6432) );
  BUFFD0 U6427 ( .I(n6434), .Z(n6433) );
  BUFFD0 U6428 ( .I(n6435), .Z(n6434) );
  BUFFD0 U6429 ( .I(n6436), .Z(n6435) );
  BUFFD0 U6430 ( .I(n6437), .Z(n6436) );
  BUFFD0 U6431 ( .I(n6438), .Z(n6437) );
  BUFFD0 U6432 ( .I(n6439), .Z(n6438) );
  BUFFD0 U6433 ( .I(n6440), .Z(n6439) );
  BUFFD0 U6434 ( .I(n6441), .Z(n6440) );
  BUFFD0 U6435 ( .I(n6442), .Z(n6441) );
  BUFFD0 U6436 ( .I(n6443), .Z(n6442) );
  BUFFD0 U6437 ( .I(n6444), .Z(n6443) );
  BUFFD0 U6438 ( .I(n6445), .Z(n6444) );
  BUFFD0 U6439 ( .I(n6446), .Z(n6445) );
  BUFFD0 U6440 ( .I(n6447), .Z(n6446) );
  BUFFD0 U6441 ( .I(n6448), .Z(n6447) );
  BUFFD0 U6442 ( .I(n6449), .Z(n6448) );
  BUFFD0 U6443 ( .I(n6450), .Z(n6449) );
  BUFFD0 U6444 ( .I(n6451), .Z(n6450) );
  BUFFD0 U6445 ( .I(n6452), .Z(n6451) );
  BUFFD0 U6446 ( .I(n6453), .Z(n6452) );
  BUFFD0 U6447 ( .I(n6454), .Z(n6453) );
  BUFFD0 U6448 ( .I(n6455), .Z(n6454) );
  BUFFD0 U6449 ( .I(n6456), .Z(n6455) );
  BUFFD0 U6450 ( .I(n6457), .Z(n6456) );
  BUFFD0 U6451 ( .I(n6458), .Z(n6457) );
  BUFFD0 U6452 ( .I(n6459), .Z(n6458) );
  BUFFD0 U6453 ( .I(n6460), .Z(n6459) );
  BUFFD0 U6454 ( .I(n6461), .Z(n6460) );
  BUFFD0 U6455 ( .I(n6462), .Z(n6461) );
  BUFFD0 U6456 ( .I(n6463), .Z(n6462) );
  BUFFD0 U6457 ( .I(n6464), .Z(n6463) );
  BUFFD0 U6458 ( .I(n6465), .Z(n6464) );
  BUFFD0 U6459 ( .I(n6466), .Z(n6465) );
  BUFFD0 U6460 ( .I(n6467), .Z(n6466) );
  BUFFD0 U6461 ( .I(n6468), .Z(n6467) );
  BUFFD0 U6462 ( .I(n6469), .Z(n6468) );
  BUFFD0 U6463 ( .I(n6470), .Z(n6469) );
  BUFFD0 U6464 ( .I(n6471), .Z(n6470) );
  BUFFD0 U6465 ( .I(n6472), .Z(n6471) );
  BUFFD0 U6466 ( .I(n6473), .Z(n6472) );
  BUFFD0 U6467 ( .I(n6474), .Z(n6473) );
  BUFFD0 U6468 ( .I(n6475), .Z(n6474) );
  BUFFD0 U6469 ( .I(n6476), .Z(n6475) );
  BUFFD0 U6470 ( .I(n6477), .Z(n6476) );
  BUFFD0 U6471 ( .I(n6478), .Z(n6477) );
  BUFFD0 U6472 ( .I(n6479), .Z(n6478) );
  BUFFD0 U6473 ( .I(n6480), .Z(n6479) );
  BUFFD0 U6474 ( .I(n6481), .Z(n6480) );
  BUFFD0 U6475 ( .I(n6482), .Z(n6481) );
  BUFFD0 U6476 ( .I(n6483), .Z(n6482) );
  BUFFD0 U6477 ( .I(n6484), .Z(n6483) );
  BUFFD0 U6478 ( .I(n6485), .Z(n6484) );
  BUFFD0 U6479 ( .I(n6486), .Z(n6485) );
  BUFFD0 U6480 ( .I(n6487), .Z(n6486) );
  BUFFD0 U6481 ( .I(n6488), .Z(n6487) );
  BUFFD0 U6482 ( .I(n6489), .Z(n6488) );
  BUFFD0 U6483 ( .I(n6490), .Z(n6489) );
  BUFFD0 U6484 ( .I(n6491), .Z(n6490) );
  BUFFD0 U6485 ( .I(n6492), .Z(n6491) );
  BUFFD0 U6486 ( .I(n6493), .Z(n6492) );
  BUFFD0 U6487 ( .I(n6494), .Z(n6493) );
  BUFFD0 U6488 ( .I(n6495), .Z(n6494) );
  BUFFD0 U6489 ( .I(n6496), .Z(n6495) );
  BUFFD0 U6490 ( .I(n6497), .Z(n6496) );
  BUFFD0 U6491 ( .I(n6498), .Z(n6497) );
  BUFFD0 U6492 ( .I(n6499), .Z(n6498) );
  BUFFD0 U6493 ( .I(n6500), .Z(n6499) );
  BUFFD0 U6494 ( .I(n6501), .Z(n6500) );
  BUFFD0 U6495 ( .I(n6502), .Z(n6501) );
  BUFFD0 U6496 ( .I(n6503), .Z(n6502) );
  BUFFD0 U6497 ( .I(n6504), .Z(n6503) );
  BUFFD0 U6498 ( .I(n6505), .Z(n6504) );
  BUFFD0 U6499 ( .I(n6506), .Z(n6505) );
  BUFFD0 U6500 ( .I(n6507), .Z(n6506) );
  BUFFD0 U6501 ( .I(n6508), .Z(n6507) );
  BUFFD0 U6502 ( .I(n6509), .Z(n6508) );
  BUFFD0 U6503 ( .I(n6510), .Z(n6509) );
  BUFFD0 U6504 ( .I(n6511), .Z(n6510) );
  BUFFD0 U6505 ( .I(n6512), .Z(n6511) );
  BUFFD0 U6506 ( .I(n6513), .Z(n6512) );
  BUFFD0 U6507 ( .I(n6514), .Z(n6513) );
  BUFFD0 U6508 ( .I(n6515), .Z(n6514) );
  BUFFD0 U6509 ( .I(n6516), .Z(n6515) );
  BUFFD0 U6510 ( .I(n6517), .Z(n6516) );
  BUFFD0 U6511 ( .I(n6518), .Z(n6517) );
  BUFFD0 U6512 ( .I(n6519), .Z(n6518) );
  BUFFD0 U6513 ( .I(n6520), .Z(n6519) );
  BUFFD0 U6514 ( .I(n6521), .Z(n6520) );
  BUFFD0 U6515 ( .I(n6522), .Z(n6521) );
  BUFFD0 U6516 ( .I(n6523), .Z(n6522) );
  BUFFD0 U6517 ( .I(n6524), .Z(n6523) );
  BUFFD0 U6518 ( .I(n6525), .Z(n6524) );
  BUFFD0 U6519 ( .I(n6526), .Z(n6525) );
  BUFFD0 U6520 ( .I(n6527), .Z(n6526) );
  BUFFD0 U6521 ( .I(n6528), .Z(n6527) );
  BUFFD0 U6522 ( .I(n6529), .Z(n6528) );
  BUFFD0 U6523 ( .I(n6530), .Z(n6529) );
  BUFFD0 U6524 ( .I(n6531), .Z(n6530) );
  BUFFD0 U6525 ( .I(n6532), .Z(n6531) );
  BUFFD0 U6526 ( .I(n6533), .Z(n6532) );
  BUFFD0 U6527 ( .I(n6534), .Z(n6533) );
  BUFFD0 U6528 ( .I(n6535), .Z(n6534) );
  BUFFD0 U6529 ( .I(n6536), .Z(n6535) );
  BUFFD0 U6530 ( .I(n6537), .Z(n6536) );
  BUFFD0 U6531 ( .I(n6538), .Z(n6537) );
  BUFFD0 U6532 ( .I(n6539), .Z(n6538) );
  BUFFD0 U6533 ( .I(n6540), .Z(n6539) );
  BUFFD0 U6534 ( .I(n6541), .Z(n6540) );
  BUFFD0 U6535 ( .I(n6542), .Z(n6541) );
  BUFFD0 U6536 ( .I(n6543), .Z(n6542) );
  BUFFD0 U6537 ( .I(n6544), .Z(n6543) );
  BUFFD0 U6538 ( .I(n6545), .Z(n6544) );
  BUFFD0 U6539 ( .I(n6546), .Z(n6545) );
  BUFFD0 U6540 ( .I(n6547), .Z(n6546) );
  BUFFD0 U6541 ( .I(n6548), .Z(n6547) );
  BUFFD0 U6542 ( .I(n6549), .Z(n6548) );
  BUFFD0 U6543 ( .I(n6550), .Z(n6549) );
  BUFFD0 U6544 ( .I(n6551), .Z(n6550) );
  BUFFD0 U6545 ( .I(n6552), .Z(n6551) );
  BUFFD0 U6546 ( .I(n6553), .Z(n6552) );
  BUFFD0 U6547 ( .I(n6554), .Z(n6553) );
  BUFFD0 U6548 ( .I(n6555), .Z(n6554) );
  BUFFD0 U6549 ( .I(n6556), .Z(n6555) );
  BUFFD0 U6550 ( .I(n6557), .Z(n6556) );
  BUFFD0 U6551 ( .I(n6558), .Z(n6557) );
  BUFFD0 U6552 ( .I(n6559), .Z(n6558) );
  BUFFD0 U6553 ( .I(n6560), .Z(n6559) );
  BUFFD0 U6554 ( .I(n6561), .Z(n6560) );
  BUFFD0 U6555 ( .I(n6562), .Z(n6561) );
  BUFFD0 U6556 ( .I(n6563), .Z(n6562) );
  BUFFD0 U6557 ( .I(n6564), .Z(n6563) );
  BUFFD0 U6558 ( .I(n6565), .Z(n6564) );
  BUFFD0 U6559 ( .I(n6566), .Z(n6565) );
  BUFFD0 U6560 ( .I(n6567), .Z(n6566) );
  BUFFD0 U6561 ( .I(n6568), .Z(n6567) );
  BUFFD0 U6562 ( .I(n6569), .Z(n6568) );
  BUFFD0 U6563 ( .I(n6570), .Z(n6569) );
  BUFFD0 U6564 ( .I(n6571), .Z(n6570) );
  BUFFD0 U6565 ( .I(n6572), .Z(n6571) );
  BUFFD0 U6566 ( .I(n6573), .Z(n6572) );
  BUFFD0 U6567 ( .I(n6574), .Z(n6573) );
  BUFFD0 U6568 ( .I(n6575), .Z(n6574) );
  BUFFD0 U6569 ( .I(n6576), .Z(n6575) );
  BUFFD0 U6570 ( .I(n6577), .Z(n6576) );
  BUFFD0 U6571 ( .I(n6578), .Z(n6577) );
  BUFFD0 U6572 ( .I(n8697), .Z(n6578) );
  BUFFD0 U6573 ( .I(n8694), .Z(n6579) );
  BUFFD0 U6574 ( .I(n6581), .Z(n6580) );
  BUFFD0 U6575 ( .I(n6582), .Z(n6581) );
  BUFFD0 U6576 ( .I(n6583), .Z(n6582) );
  BUFFD0 U6577 ( .I(n6584), .Z(n6583) );
  BUFFD0 U6578 ( .I(n6585), .Z(n6584) );
  BUFFD0 U6579 ( .I(n6586), .Z(n6585) );
  BUFFD0 U6580 ( .I(n6587), .Z(n6586) );
  BUFFD0 U6581 ( .I(n6588), .Z(n6587) );
  BUFFD0 U6582 ( .I(n6589), .Z(n6588) );
  BUFFD0 U6583 ( .I(n6590), .Z(n6589) );
  BUFFD0 U6584 ( .I(n6591), .Z(n6590) );
  BUFFD0 U6585 ( .I(n6592), .Z(n6591) );
  BUFFD0 U6586 ( .I(n6593), .Z(n6592) );
  BUFFD0 U6587 ( .I(n6594), .Z(n6593) );
  BUFFD0 U6588 ( .I(n6595), .Z(n6594) );
  BUFFD0 U6589 ( .I(n6596), .Z(n6595) );
  BUFFD0 U6590 ( .I(n6597), .Z(n6596) );
  BUFFD0 U6591 ( .I(n6598), .Z(n6597) );
  BUFFD0 U6592 ( .I(n6599), .Z(n6598) );
  BUFFD0 U6593 ( .I(n6600), .Z(n6599) );
  BUFFD0 U6594 ( .I(n6601), .Z(n6600) );
  BUFFD0 U6595 ( .I(n6602), .Z(n6601) );
  BUFFD0 U6596 ( .I(n6603), .Z(n6602) );
  BUFFD0 U6597 ( .I(n6604), .Z(n6603) );
  BUFFD0 U6598 ( .I(n6605), .Z(n6604) );
  BUFFD0 U6599 ( .I(n6606), .Z(n6605) );
  BUFFD0 U6600 ( .I(n6607), .Z(n6606) );
  BUFFD0 U6601 ( .I(n6608), .Z(n6607) );
  BUFFD0 U6602 ( .I(n6609), .Z(n6608) );
  BUFFD0 U6603 ( .I(n6610), .Z(n6609) );
  BUFFD0 U6604 ( .I(n6611), .Z(n6610) );
  BUFFD0 U6605 ( .I(n6612), .Z(n6611) );
  BUFFD0 U6606 ( .I(n6613), .Z(n6612) );
  BUFFD0 U6607 ( .I(n6614), .Z(n6613) );
  BUFFD0 U6608 ( .I(n6615), .Z(n6614) );
  BUFFD0 U6609 ( .I(n6616), .Z(n6615) );
  BUFFD0 U6610 ( .I(n6617), .Z(n6616) );
  BUFFD0 U6611 ( .I(n6618), .Z(n6617) );
  BUFFD0 U6612 ( .I(n6619), .Z(n6618) );
  BUFFD0 U6613 ( .I(n6620), .Z(n6619) );
  BUFFD0 U6614 ( .I(n6621), .Z(n6620) );
  BUFFD0 U6615 ( .I(n6622), .Z(n6621) );
  BUFFD0 U6616 ( .I(n6623), .Z(n6622) );
  BUFFD0 U6617 ( .I(n6624), .Z(n6623) );
  BUFFD0 U6618 ( .I(n6625), .Z(n6624) );
  BUFFD0 U6619 ( .I(n6626), .Z(n6625) );
  BUFFD0 U6620 ( .I(n6627), .Z(n6626) );
  BUFFD0 U6621 ( .I(n6628), .Z(n6627) );
  BUFFD0 U6622 ( .I(n6629), .Z(n6628) );
  BUFFD0 U6623 ( .I(n6630), .Z(n6629) );
  BUFFD0 U6624 ( .I(n6631), .Z(n6630) );
  BUFFD0 U6625 ( .I(n6632), .Z(n6631) );
  BUFFD0 U6626 ( .I(n6633), .Z(n6632) );
  BUFFD0 U6627 ( .I(n6634), .Z(n6633) );
  BUFFD0 U6628 ( .I(n6635), .Z(n6634) );
  BUFFD0 U6629 ( .I(n6636), .Z(n6635) );
  BUFFD0 U6630 ( .I(n6637), .Z(n6636) );
  BUFFD0 U6631 ( .I(n6638), .Z(n6637) );
  BUFFD0 U6632 ( .I(n6639), .Z(n6638) );
  BUFFD0 U6633 ( .I(n6640), .Z(n6639) );
  BUFFD0 U6634 ( .I(n6641), .Z(n6640) );
  BUFFD0 U6635 ( .I(n6642), .Z(n6641) );
  BUFFD0 U6636 ( .I(n6643), .Z(n6642) );
  BUFFD0 U6637 ( .I(n6644), .Z(n6643) );
  BUFFD0 U6638 ( .I(n6645), .Z(n6644) );
  BUFFD0 U6639 ( .I(n6646), .Z(n6645) );
  BUFFD0 U6640 ( .I(n6647), .Z(n6646) );
  BUFFD0 U6641 ( .I(n6648), .Z(n6647) );
  BUFFD0 U6642 ( .I(n6649), .Z(n6648) );
  BUFFD0 U6643 ( .I(n6650), .Z(n6649) );
  BUFFD0 U6644 ( .I(n6651), .Z(n6650) );
  BUFFD0 U6645 ( .I(n6652), .Z(n6651) );
  BUFFD0 U6646 ( .I(n6653), .Z(n6652) );
  BUFFD0 U6647 ( .I(n6654), .Z(n6653) );
  BUFFD0 U6648 ( .I(n6655), .Z(n6654) );
  BUFFD0 U6649 ( .I(n6656), .Z(n6655) );
  BUFFD0 U6650 ( .I(n6657), .Z(n6656) );
  BUFFD0 U6651 ( .I(n6658), .Z(n6657) );
  BUFFD0 U6652 ( .I(n6659), .Z(n6658) );
  BUFFD0 U6653 ( .I(n6660), .Z(n6659) );
  BUFFD0 U6654 ( .I(n6661), .Z(n6660) );
  BUFFD0 U6655 ( .I(n6662), .Z(n6661) );
  BUFFD0 U6656 ( .I(n6663), .Z(n6662) );
  BUFFD0 U6657 ( .I(n6664), .Z(n6663) );
  BUFFD0 U6658 ( .I(n6665), .Z(n6664) );
  BUFFD0 U6659 ( .I(n6666), .Z(n6665) );
  BUFFD0 U6660 ( .I(n6667), .Z(n6666) );
  BUFFD0 U6661 ( .I(n6668), .Z(n6667) );
  BUFFD0 U6662 ( .I(n6669), .Z(n6668) );
  BUFFD0 U6663 ( .I(n6670), .Z(n6669) );
  BUFFD0 U6664 ( .I(n6671), .Z(n6670) );
  BUFFD0 U6665 ( .I(n6672), .Z(n6671) );
  BUFFD0 U6666 ( .I(n6673), .Z(n6672) );
  BUFFD0 U6667 ( .I(n6674), .Z(n6673) );
  BUFFD0 U6668 ( .I(n6675), .Z(n6674) );
  BUFFD0 U6669 ( .I(n6676), .Z(n6675) );
  BUFFD0 U6670 ( .I(n6677), .Z(n6676) );
  BUFFD0 U6671 ( .I(n6678), .Z(n6677) );
  BUFFD0 U6672 ( .I(n6679), .Z(n6678) );
  BUFFD0 U6673 ( .I(n6680), .Z(n6679) );
  BUFFD0 U6674 ( .I(n6681), .Z(n6680) );
  BUFFD0 U6675 ( .I(n6682), .Z(n6681) );
  BUFFD0 U6676 ( .I(n6683), .Z(n6682) );
  BUFFD0 U6677 ( .I(n6684), .Z(n6683) );
  BUFFD0 U6678 ( .I(n6685), .Z(n6684) );
  BUFFD0 U6679 ( .I(n6686), .Z(n6685) );
  BUFFD0 U6680 ( .I(n6687), .Z(n6686) );
  BUFFD0 U6681 ( .I(n6688), .Z(n6687) );
  BUFFD0 U6682 ( .I(n6689), .Z(n6688) );
  BUFFD0 U6683 ( .I(n6690), .Z(n6689) );
  BUFFD0 U6684 ( .I(n6691), .Z(n6690) );
  BUFFD0 U6685 ( .I(n6692), .Z(n6691) );
  BUFFD0 U6686 ( .I(n6693), .Z(n6692) );
  BUFFD0 U6687 ( .I(n6694), .Z(n6693) );
  BUFFD0 U6688 ( .I(n6695), .Z(n6694) );
  BUFFD0 U6689 ( .I(n6696), .Z(n6695) );
  BUFFD0 U6690 ( .I(n6697), .Z(n6696) );
  BUFFD0 U6691 ( .I(n6698), .Z(n6697) );
  BUFFD0 U6692 ( .I(n6699), .Z(n6698) );
  BUFFD0 U6693 ( .I(n6700), .Z(n6699) );
  BUFFD0 U6694 ( .I(n6701), .Z(n6700) );
  BUFFD0 U6695 ( .I(n6702), .Z(n6701) );
  BUFFD0 U6696 ( .I(n6703), .Z(n6702) );
  BUFFD0 U6697 ( .I(n6704), .Z(n6703) );
  BUFFD0 U6698 ( .I(n6705), .Z(n6704) );
  BUFFD0 U6699 ( .I(n6706), .Z(n6705) );
  BUFFD0 U6700 ( .I(n6707), .Z(n6706) );
  BUFFD0 U6701 ( .I(n6708), .Z(n6707) );
  BUFFD0 U6702 ( .I(n6709), .Z(n6708) );
  BUFFD0 U6703 ( .I(n6710), .Z(n6709) );
  BUFFD0 U6704 ( .I(n6711), .Z(n6710) );
  BUFFD0 U6705 ( .I(n6712), .Z(n6711) );
  BUFFD0 U6706 ( .I(n6713), .Z(n6712) );
  BUFFD0 U6707 ( .I(n6714), .Z(n6713) );
  BUFFD0 U6708 ( .I(n6715), .Z(n6714) );
  BUFFD0 U6709 ( .I(n6716), .Z(n6715) );
  BUFFD0 U6710 ( .I(n6717), .Z(n6716) );
  BUFFD0 U6711 ( .I(n6718), .Z(n6717) );
  BUFFD0 U6712 ( .I(n6719), .Z(n6718) );
  BUFFD0 U6713 ( .I(n6720), .Z(n6719) );
  BUFFD0 U6714 ( .I(n6721), .Z(n6720) );
  BUFFD0 U6715 ( .I(n6722), .Z(n6721) );
  BUFFD0 U6716 ( .I(n6723), .Z(n6722) );
  BUFFD0 U6717 ( .I(n6724), .Z(n6723) );
  BUFFD0 U6718 ( .I(n6725), .Z(n6724) );
  BUFFD0 U6719 ( .I(n6726), .Z(n6725) );
  BUFFD0 U6720 ( .I(n6727), .Z(n6726) );
  BUFFD0 U6721 ( .I(n6728), .Z(n6727) );
  BUFFD0 U6722 ( .I(n6729), .Z(n6728) );
  BUFFD0 U6723 ( .I(n6730), .Z(n6729) );
  BUFFD0 U6724 ( .I(n6731), .Z(n6730) );
  BUFFD0 U6725 ( .I(n6732), .Z(n6731) );
  BUFFD0 U6726 ( .I(n6733), .Z(n6732) );
  BUFFD0 U6727 ( .I(n6734), .Z(n6733) );
  BUFFD0 U6728 ( .I(n6735), .Z(n6734) );
  BUFFD0 U6729 ( .I(n6736), .Z(n6735) );
  BUFFD0 U6730 ( .I(n6737), .Z(n6736) );
  BUFFD0 U6731 ( .I(n6738), .Z(n6737) );
  BUFFD0 U6732 ( .I(n6739), .Z(n6738) );
  BUFFD0 U6733 ( .I(n6740), .Z(n6739) );
  BUFFD0 U6734 ( .I(n6741), .Z(n6740) );
  BUFFD0 U6735 ( .I(n6742), .Z(n6741) );
  BUFFD0 U6736 ( .I(n6743), .Z(n6742) );
  BUFFD0 U6737 ( .I(n6744), .Z(n6743) );
  BUFFD0 U6738 ( .I(n6745), .Z(n6744) );
  BUFFD0 U6739 ( .I(n6746), .Z(n6745) );
  BUFFD0 U6740 ( .I(n6747), .Z(n6746) );
  BUFFD0 U6741 ( .I(n6748), .Z(n6747) );
  BUFFD0 U6742 ( .I(n6749), .Z(n6748) );
  BUFFD0 U6743 ( .I(n6750), .Z(n6749) );
  BUFFD0 U6744 ( .I(n6751), .Z(n6750) );
  BUFFD0 U6745 ( .I(n6752), .Z(n6751) );
  BUFFD0 U6746 ( .I(n6753), .Z(n6752) );
  BUFFD0 U6747 ( .I(n6754), .Z(n6753) );
  BUFFD0 U6748 ( .I(n6755), .Z(n6754) );
  BUFFD0 U6749 ( .I(n6756), .Z(n6755) );
  BUFFD0 U6750 ( .I(n6757), .Z(n6756) );
  BUFFD0 U6751 ( .I(n8695), .Z(n6757) );
  BUFFD0 U6752 ( .I(n6759), .Z(n6758) );
  BUFFD0 U6753 ( .I(n6760), .Z(n6759) );
  BUFFD0 U6754 ( .I(n6761), .Z(n6760) );
  BUFFD0 U6755 ( .I(n6762), .Z(n6761) );
  BUFFD0 U6756 ( .I(n6763), .Z(n6762) );
  BUFFD0 U6757 ( .I(n6764), .Z(n6763) );
  BUFFD0 U6758 ( .I(n6765), .Z(n6764) );
  BUFFD0 U6759 ( .I(n6766), .Z(n6765) );
  BUFFD0 U6760 ( .I(n6767), .Z(n6766) );
  BUFFD0 U6761 ( .I(n6768), .Z(n6767) );
  BUFFD0 U6762 ( .I(n6769), .Z(n6768) );
  BUFFD0 U6763 ( .I(n6770), .Z(n6769) );
  BUFFD0 U6764 ( .I(n6771), .Z(n6770) );
  BUFFD0 U6765 ( .I(n6772), .Z(n6771) );
  BUFFD0 U6766 ( .I(n6773), .Z(n6772) );
  BUFFD0 U6767 ( .I(n6774), .Z(n6773) );
  BUFFD0 U6768 ( .I(n6775), .Z(n6774) );
  BUFFD0 U6769 ( .I(n6776), .Z(n6775) );
  BUFFD0 U6770 ( .I(n6777), .Z(n6776) );
  BUFFD0 U6771 ( .I(n6778), .Z(n6777) );
  BUFFD0 U6772 ( .I(n6779), .Z(n6778) );
  BUFFD0 U6773 ( .I(n6780), .Z(n6779) );
  BUFFD0 U6774 ( .I(n6781), .Z(n6780) );
  BUFFD0 U6775 ( .I(n6782), .Z(n6781) );
  BUFFD0 U6776 ( .I(n6783), .Z(n6782) );
  BUFFD0 U6777 ( .I(n6784), .Z(n6783) );
  BUFFD0 U6778 ( .I(n6785), .Z(n6784) );
  BUFFD0 U6779 ( .I(n6786), .Z(n6785) );
  BUFFD0 U6780 ( .I(n6787), .Z(n6786) );
  BUFFD0 U6781 ( .I(n6788), .Z(n6787) );
  BUFFD0 U6782 ( .I(n6789), .Z(n6788) );
  BUFFD0 U6783 ( .I(n6790), .Z(n6789) );
  BUFFD0 U6784 ( .I(n6791), .Z(n6790) );
  BUFFD0 U6785 ( .I(n6792), .Z(n6791) );
  BUFFD0 U6786 ( .I(n6793), .Z(n6792) );
  BUFFD0 U6787 ( .I(n6794), .Z(n6793) );
  BUFFD0 U6788 ( .I(n6795), .Z(n6794) );
  BUFFD0 U6789 ( .I(n6796), .Z(n6795) );
  BUFFD0 U6790 ( .I(n6797), .Z(n6796) );
  BUFFD0 U6791 ( .I(n6798), .Z(n6797) );
  BUFFD0 U6792 ( .I(n6799), .Z(n6798) );
  BUFFD0 U6793 ( .I(n6800), .Z(n6799) );
  BUFFD0 U6794 ( .I(n6801), .Z(n6800) );
  BUFFD0 U6795 ( .I(n6802), .Z(n6801) );
  BUFFD0 U6796 ( .I(n6803), .Z(n6802) );
  BUFFD0 U6797 ( .I(n6804), .Z(n6803) );
  BUFFD0 U6798 ( .I(n6805), .Z(n6804) );
  BUFFD0 U6799 ( .I(n6806), .Z(n6805) );
  BUFFD0 U6800 ( .I(n6807), .Z(n6806) );
  BUFFD0 U6801 ( .I(n6808), .Z(n6807) );
  BUFFD0 U6802 ( .I(n6809), .Z(n6808) );
  BUFFD0 U6803 ( .I(n6810), .Z(n6809) );
  BUFFD0 U6804 ( .I(n6811), .Z(n6810) );
  BUFFD0 U6805 ( .I(n6812), .Z(n6811) );
  BUFFD0 U6806 ( .I(n6813), .Z(n6812) );
  BUFFD0 U6807 ( .I(n6814), .Z(n6813) );
  BUFFD0 U6808 ( .I(n6815), .Z(n6814) );
  BUFFD0 U6809 ( .I(n6816), .Z(n6815) );
  BUFFD0 U6810 ( .I(n6817), .Z(n6816) );
  BUFFD0 U6811 ( .I(n6818), .Z(n6817) );
  BUFFD0 U6812 ( .I(n6819), .Z(n6818) );
  BUFFD0 U6813 ( .I(n6820), .Z(n6819) );
  BUFFD0 U6814 ( .I(n6821), .Z(n6820) );
  BUFFD0 U6815 ( .I(n6822), .Z(n6821) );
  BUFFD0 U6816 ( .I(n6823), .Z(n6822) );
  BUFFD0 U6817 ( .I(n6824), .Z(n6823) );
  BUFFD0 U6818 ( .I(n6825), .Z(n6824) );
  BUFFD0 U6819 ( .I(n6826), .Z(n6825) );
  BUFFD0 U6820 ( .I(n6827), .Z(n6826) );
  BUFFD0 U6821 ( .I(n6828), .Z(n6827) );
  BUFFD0 U6822 ( .I(n6829), .Z(n6828) );
  BUFFD0 U6823 ( .I(n6830), .Z(n6829) );
  BUFFD0 U6824 ( .I(n6831), .Z(n6830) );
  BUFFD0 U6825 ( .I(n6832), .Z(n6831) );
  BUFFD0 U6826 ( .I(n6833), .Z(n6832) );
  BUFFD0 U6827 ( .I(n6834), .Z(n6833) );
  BUFFD0 U6828 ( .I(n6835), .Z(n6834) );
  BUFFD0 U6829 ( .I(n6836), .Z(n6835) );
  BUFFD0 U6830 ( .I(n6837), .Z(n6836) );
  BUFFD0 U6831 ( .I(n6838), .Z(n6837) );
  BUFFD0 U6832 ( .I(n6839), .Z(n6838) );
  BUFFD0 U6833 ( .I(n6840), .Z(n6839) );
  BUFFD0 U6834 ( .I(n6841), .Z(n6840) );
  BUFFD0 U6835 ( .I(n6842), .Z(n6841) );
  BUFFD0 U6836 ( .I(n6843), .Z(n6842) );
  BUFFD0 U6837 ( .I(n6844), .Z(n6843) );
  BUFFD0 U6838 ( .I(n6845), .Z(n6844) );
  BUFFD0 U6839 ( .I(n6846), .Z(n6845) );
  BUFFD0 U6840 ( .I(n6847), .Z(n6846) );
  BUFFD0 U6841 ( .I(n6848), .Z(n6847) );
  BUFFD0 U6842 ( .I(n6849), .Z(n6848) );
  BUFFD0 U6843 ( .I(n6850), .Z(n6849) );
  BUFFD0 U6844 ( .I(n6851), .Z(n6850) );
  BUFFD0 U6845 ( .I(n6852), .Z(n6851) );
  BUFFD0 U6846 ( .I(n6853), .Z(n6852) );
  BUFFD0 U6847 ( .I(n6854), .Z(n6853) );
  BUFFD0 U6848 ( .I(n6855), .Z(n6854) );
  BUFFD0 U6849 ( .I(n6856), .Z(n6855) );
  BUFFD0 U6850 ( .I(n6857), .Z(n6856) );
  BUFFD0 U6851 ( .I(n6858), .Z(n6857) );
  BUFFD0 U6852 ( .I(n6859), .Z(n6858) );
  BUFFD0 U6853 ( .I(n6860), .Z(n6859) );
  BUFFD0 U6854 ( .I(n6861), .Z(n6860) );
  BUFFD0 U6855 ( .I(n6862), .Z(n6861) );
  BUFFD0 U6856 ( .I(n6863), .Z(n6862) );
  BUFFD0 U6857 ( .I(n6864), .Z(n6863) );
  BUFFD0 U6858 ( .I(n6865), .Z(n6864) );
  BUFFD0 U6859 ( .I(n6866), .Z(n6865) );
  BUFFD0 U6860 ( .I(n6867), .Z(n6866) );
  BUFFD0 U6861 ( .I(n6868), .Z(n6867) );
  BUFFD0 U6862 ( .I(n6869), .Z(n6868) );
  BUFFD0 U6863 ( .I(n6870), .Z(n6869) );
  BUFFD0 U6864 ( .I(n6871), .Z(n6870) );
  BUFFD0 U6865 ( .I(n6872), .Z(n6871) );
  BUFFD0 U6866 ( .I(n6873), .Z(n6872) );
  BUFFD0 U6867 ( .I(n6874), .Z(n6873) );
  BUFFD0 U6868 ( .I(n6875), .Z(n6874) );
  BUFFD0 U6869 ( .I(n6876), .Z(n6875) );
  BUFFD0 U6870 ( .I(n6877), .Z(n6876) );
  BUFFD0 U6871 ( .I(n6878), .Z(n6877) );
  BUFFD0 U6872 ( .I(n6879), .Z(n6878) );
  BUFFD0 U6873 ( .I(n6880), .Z(n6879) );
  BUFFD0 U6874 ( .I(n6881), .Z(n6880) );
  BUFFD0 U6875 ( .I(n6882), .Z(n6881) );
  BUFFD0 U6876 ( .I(n6883), .Z(n6882) );
  BUFFD0 U6877 ( .I(n6884), .Z(n6883) );
  BUFFD0 U6878 ( .I(n6885), .Z(n6884) );
  BUFFD0 U6879 ( .I(n6886), .Z(n6885) );
  BUFFD0 U6880 ( .I(n6887), .Z(n6886) );
  BUFFD0 U6881 ( .I(n6888), .Z(n6887) );
  BUFFD0 U6882 ( .I(n6889), .Z(n6888) );
  BUFFD0 U6883 ( .I(n6890), .Z(n6889) );
  BUFFD0 U6884 ( .I(n6891), .Z(n6890) );
  BUFFD0 U6885 ( .I(n6892), .Z(n6891) );
  BUFFD0 U6886 ( .I(n6893), .Z(n6892) );
  BUFFD0 U6887 ( .I(n6894), .Z(n6893) );
  BUFFD0 U6888 ( .I(n6895), .Z(n6894) );
  BUFFD0 U6889 ( .I(n6896), .Z(n6895) );
  BUFFD0 U6890 ( .I(n6897), .Z(n6896) );
  BUFFD0 U6891 ( .I(n6898), .Z(n6897) );
  BUFFD0 U6892 ( .I(n6899), .Z(n6898) );
  BUFFD0 U6893 ( .I(n6901), .Z(n6899) );
  BUFFD0 U6894 ( .I(n8692), .Z(n6900) );
  BUFFD0 U6895 ( .I(n6902), .Z(n6901) );
  BUFFD0 U6896 ( .I(n6903), .Z(n6902) );
  BUFFD0 U6897 ( .I(n6904), .Z(n6903) );
  BUFFD0 U6898 ( .I(n6905), .Z(n6904) );
  BUFFD0 U6899 ( .I(n6906), .Z(n6905) );
  BUFFD0 U6900 ( .I(n6907), .Z(n6906) );
  BUFFD0 U6901 ( .I(n6908), .Z(n6907) );
  BUFFD0 U6902 ( .I(n6909), .Z(n6908) );
  BUFFD0 U6903 ( .I(n6910), .Z(n6909) );
  BUFFD0 U6904 ( .I(n6911), .Z(n6910) );
  BUFFD0 U6905 ( .I(n6912), .Z(n6911) );
  BUFFD0 U6906 ( .I(n6913), .Z(n6912) );
  BUFFD0 U6907 ( .I(n6914), .Z(n6913) );
  BUFFD0 U6908 ( .I(n6915), .Z(n6914) );
  BUFFD0 U6909 ( .I(n6916), .Z(n6915) );
  BUFFD0 U6910 ( .I(n6917), .Z(n6916) );
  BUFFD0 U6911 ( .I(n6918), .Z(n6917) );
  BUFFD0 U6912 ( .I(n6919), .Z(n6918) );
  BUFFD0 U6913 ( .I(n6920), .Z(n6919) );
  BUFFD0 U6914 ( .I(n6921), .Z(n6920) );
  BUFFD0 U6915 ( .I(n6922), .Z(n6921) );
  BUFFD0 U6916 ( .I(n6923), .Z(n6922) );
  BUFFD0 U6917 ( .I(n6924), .Z(n6923) );
  BUFFD0 U6918 ( .I(n6925), .Z(n6924) );
  BUFFD0 U6919 ( .I(n6926), .Z(n6925) );
  BUFFD0 U6920 ( .I(n6927), .Z(n6926) );
  BUFFD0 U6921 ( .I(n6928), .Z(n6927) );
  BUFFD0 U6922 ( .I(n6929), .Z(n6928) );
  BUFFD0 U6923 ( .I(n6930), .Z(n6929) );
  BUFFD0 U6924 ( .I(n6931), .Z(n6930) );
  BUFFD0 U6925 ( .I(n6932), .Z(n6931) );
  BUFFD0 U6926 ( .I(n6933), .Z(n6932) );
  BUFFD0 U6927 ( .I(n8689), .Z(n6934) );
  BUFFD0 U6928 ( .I(n6936), .Z(n6935) );
  BUFFD0 U6929 ( .I(n6937), .Z(n6936) );
  BUFFD0 U6930 ( .I(n6938), .Z(n6937) );
  BUFFD0 U6931 ( .I(n6939), .Z(n6938) );
  BUFFD0 U6932 ( .I(n6940), .Z(n6939) );
  BUFFD0 U6933 ( .I(n6941), .Z(n6940) );
  BUFFD0 U6934 ( .I(n6942), .Z(n6941) );
  BUFFD0 U6935 ( .I(n6943), .Z(n6942) );
  BUFFD0 U6936 ( .I(n6944), .Z(n6943) );
  BUFFD0 U6937 ( .I(n6945), .Z(n6944) );
  BUFFD0 U6938 ( .I(n6946), .Z(n6945) );
  BUFFD0 U6939 ( .I(n6947), .Z(n6946) );
  BUFFD0 U6940 ( .I(n6948), .Z(n6947) );
  BUFFD0 U6941 ( .I(n6949), .Z(n6948) );
  BUFFD0 U6942 ( .I(n6950), .Z(n6949) );
  BUFFD0 U6943 ( .I(n6951), .Z(n6950) );
  BUFFD0 U6944 ( .I(n6952), .Z(n6951) );
  BUFFD0 U6945 ( .I(n6953), .Z(n6952) );
  BUFFD0 U6946 ( .I(n6954), .Z(n6953) );
  BUFFD0 U6947 ( .I(n6955), .Z(n6954) );
  BUFFD0 U6948 ( .I(n6956), .Z(n6955) );
  BUFFD0 U6949 ( .I(n6957), .Z(n6956) );
  BUFFD0 U6950 ( .I(n6958), .Z(n6957) );
  BUFFD0 U6951 ( .I(n6959), .Z(n6958) );
  BUFFD0 U6952 ( .I(n6960), .Z(n6959) );
  BUFFD0 U6953 ( .I(n6961), .Z(n6960) );
  BUFFD0 U6954 ( .I(n6962), .Z(n6961) );
  BUFFD0 U6955 ( .I(n6963), .Z(n6962) );
  BUFFD0 U6956 ( .I(n6964), .Z(n6963) );
  BUFFD0 U6957 ( .I(n6965), .Z(n6964) );
  BUFFD0 U6958 ( .I(n6966), .Z(n6965) );
  BUFFD0 U6959 ( .I(n6967), .Z(n6966) );
  BUFFD0 U6960 ( .I(n6968), .Z(n6967) );
  BUFFD0 U6961 ( .I(n6969), .Z(n6968) );
  BUFFD0 U6962 ( .I(n6970), .Z(n6969) );
  BUFFD0 U6963 ( .I(n6971), .Z(n6970) );
  BUFFD0 U6964 ( .I(n6972), .Z(n6971) );
  BUFFD0 U6965 ( .I(n6973), .Z(n6972) );
  BUFFD0 U6966 ( .I(n6974), .Z(n6973) );
  BUFFD0 U6967 ( .I(n6975), .Z(n6974) );
  BUFFD0 U6968 ( .I(n6976), .Z(n6975) );
  BUFFD0 U6969 ( .I(n6977), .Z(n6976) );
  BUFFD0 U6970 ( .I(n6978), .Z(n6977) );
  BUFFD0 U6971 ( .I(n6979), .Z(n6978) );
  BUFFD0 U6972 ( .I(n6980), .Z(n6979) );
  BUFFD0 U6973 ( .I(n6981), .Z(n6980) );
  BUFFD0 U6974 ( .I(n6982), .Z(n6981) );
  BUFFD0 U6975 ( .I(n6983), .Z(n6982) );
  BUFFD0 U6976 ( .I(n6984), .Z(n6983) );
  BUFFD0 U6977 ( .I(n6985), .Z(n6984) );
  BUFFD0 U6978 ( .I(n6986), .Z(n6985) );
  BUFFD0 U6979 ( .I(n6987), .Z(n6986) );
  BUFFD0 U6980 ( .I(n6988), .Z(n6987) );
  BUFFD0 U6981 ( .I(n6989), .Z(n6988) );
  BUFFD0 U6982 ( .I(n6990), .Z(n6989) );
  BUFFD0 U6983 ( .I(n6991), .Z(n6990) );
  BUFFD0 U6984 ( .I(n6992), .Z(n6991) );
  BUFFD0 U6985 ( .I(n6993), .Z(n6992) );
  BUFFD0 U6986 ( .I(n6994), .Z(n6993) );
  BUFFD0 U6987 ( .I(n6995), .Z(n6994) );
  BUFFD0 U6988 ( .I(n6996), .Z(n6995) );
  BUFFD0 U6989 ( .I(n6997), .Z(n6996) );
  BUFFD0 U6990 ( .I(n6998), .Z(n6997) );
  BUFFD0 U6991 ( .I(n6999), .Z(n6998) );
  BUFFD0 U6992 ( .I(n7000), .Z(n6999) );
  BUFFD0 U6993 ( .I(n7001), .Z(n7000) );
  BUFFD0 U6994 ( .I(n7002), .Z(n7001) );
  BUFFD0 U6995 ( .I(n7003), .Z(n7002) );
  BUFFD0 U6996 ( .I(n7004), .Z(n7003) );
  BUFFD0 U6997 ( .I(n7005), .Z(n7004) );
  BUFFD0 U6998 ( .I(n7006), .Z(n7005) );
  BUFFD0 U6999 ( .I(n7007), .Z(n7006) );
  BUFFD0 U7000 ( .I(n7008), .Z(n7007) );
  BUFFD0 U7001 ( .I(n7009), .Z(n7008) );
  BUFFD0 U7002 ( .I(n7010), .Z(n7009) );
  BUFFD0 U7003 ( .I(n7011), .Z(n7010) );
  BUFFD0 U7004 ( .I(n7012), .Z(n7011) );
  BUFFD0 U7005 ( .I(n7013), .Z(n7012) );
  BUFFD0 U7006 ( .I(n7014), .Z(n7013) );
  BUFFD0 U7007 ( .I(n7015), .Z(n7014) );
  BUFFD0 U7008 ( .I(n7016), .Z(n7015) );
  BUFFD0 U7009 ( .I(n7017), .Z(n7016) );
  BUFFD0 U7010 ( .I(n7018), .Z(n7017) );
  BUFFD0 U7011 ( .I(n7019), .Z(n7018) );
  BUFFD0 U7012 ( .I(n7020), .Z(n7019) );
  BUFFD0 U7013 ( .I(n7021), .Z(n7020) );
  BUFFD0 U7014 ( .I(n7022), .Z(n7021) );
  BUFFD0 U7015 ( .I(n7023), .Z(n7022) );
  BUFFD0 U7016 ( .I(n7024), .Z(n7023) );
  BUFFD0 U7017 ( .I(n7025), .Z(n7024) );
  BUFFD0 U7018 ( .I(n7026), .Z(n7025) );
  BUFFD0 U7019 ( .I(n7027), .Z(n7026) );
  BUFFD0 U7020 ( .I(n7028), .Z(n7027) );
  BUFFD0 U7021 ( .I(n7029), .Z(n7028) );
  BUFFD0 U7022 ( .I(n7030), .Z(n7029) );
  BUFFD0 U7023 ( .I(n7031), .Z(n7030) );
  BUFFD0 U7024 ( .I(n7032), .Z(n7031) );
  BUFFD0 U7025 ( .I(n7033), .Z(n7032) );
  BUFFD0 U7026 ( .I(n7034), .Z(n7033) );
  BUFFD0 U7027 ( .I(n7035), .Z(n7034) );
  BUFFD0 U7028 ( .I(n7036), .Z(n7035) );
  BUFFD0 U7029 ( .I(n7037), .Z(n7036) );
  BUFFD0 U7030 ( .I(n7038), .Z(n7037) );
  BUFFD0 U7031 ( .I(n7039), .Z(n7038) );
  BUFFD0 U7032 ( .I(n7040), .Z(n7039) );
  BUFFD0 U7033 ( .I(n7041), .Z(n7040) );
  BUFFD0 U7034 ( .I(n7042), .Z(n7041) );
  BUFFD0 U7035 ( .I(n7043), .Z(n7042) );
  BUFFD0 U7036 ( .I(n7044), .Z(n7043) );
  BUFFD0 U7037 ( .I(n7045), .Z(n7044) );
  BUFFD0 U7038 ( .I(n7046), .Z(n7045) );
  BUFFD0 U7039 ( .I(n7047), .Z(n7046) );
  BUFFD0 U7040 ( .I(n7048), .Z(n7047) );
  BUFFD0 U7041 ( .I(n7049), .Z(n7048) );
  BUFFD0 U7042 ( .I(n7050), .Z(n7049) );
  BUFFD0 U7043 ( .I(n7051), .Z(n7050) );
  BUFFD0 U7044 ( .I(n7052), .Z(n7051) );
  BUFFD0 U7045 ( .I(n7053), .Z(n7052) );
  BUFFD0 U7046 ( .I(n7054), .Z(n7053) );
  BUFFD0 U7047 ( .I(n7055), .Z(n7054) );
  BUFFD0 U7048 ( .I(n7056), .Z(n7055) );
  BUFFD0 U7049 ( .I(n7057), .Z(n7056) );
  BUFFD0 U7050 ( .I(n7058), .Z(n7057) );
  BUFFD0 U7051 ( .I(n7059), .Z(n7058) );
  BUFFD0 U7052 ( .I(n7060), .Z(n7059) );
  BUFFD0 U7053 ( .I(n7061), .Z(n7060) );
  BUFFD0 U7054 ( .I(n7062), .Z(n7061) );
  BUFFD0 U7055 ( .I(n7063), .Z(n7062) );
  BUFFD0 U7056 ( .I(n7064), .Z(n7063) );
  BUFFD0 U7057 ( .I(n7065), .Z(n7064) );
  BUFFD0 U7058 ( .I(n7066), .Z(n7065) );
  BUFFD0 U7059 ( .I(n7067), .Z(n7066) );
  BUFFD0 U7060 ( .I(n7068), .Z(n7067) );
  BUFFD0 U7061 ( .I(n7069), .Z(n7068) );
  BUFFD0 U7062 ( .I(n7070), .Z(n7069) );
  BUFFD0 U7063 ( .I(n7071), .Z(n7070) );
  BUFFD0 U7064 ( .I(n7072), .Z(n7071) );
  BUFFD0 U7065 ( .I(n7073), .Z(n7072) );
  BUFFD0 U7066 ( .I(n7074), .Z(n7073) );
  BUFFD0 U7067 ( .I(n7075), .Z(n7074) );
  BUFFD0 U7068 ( .I(n7076), .Z(n7075) );
  BUFFD0 U7069 ( .I(n7077), .Z(n7076) );
  BUFFD0 U7070 ( .I(n7078), .Z(n7077) );
  BUFFD0 U7071 ( .I(n7079), .Z(n7078) );
  BUFFD0 U7072 ( .I(n7080), .Z(n7079) );
  BUFFD0 U7073 ( .I(n7081), .Z(n7080) );
  BUFFD0 U7074 ( .I(n7082), .Z(n7081) );
  BUFFD0 U7075 ( .I(n7083), .Z(n7082) );
  BUFFD0 U7076 ( .I(n7084), .Z(n7083) );
  BUFFD0 U7077 ( .I(n7085), .Z(n7084) );
  BUFFD0 U7078 ( .I(n7086), .Z(n7085) );
  BUFFD0 U7079 ( .I(n7087), .Z(n7086) );
  BUFFD0 U7080 ( .I(n7088), .Z(n7087) );
  BUFFD0 U7081 ( .I(n7089), .Z(n7088) );
  BUFFD0 U7082 ( .I(n7090), .Z(n7089) );
  BUFFD0 U7083 ( .I(n7091), .Z(n7090) );
  BUFFD0 U7084 ( .I(n7092), .Z(n7091) );
  BUFFD0 U7085 ( .I(n7093), .Z(n7092) );
  BUFFD0 U7086 ( .I(n7094), .Z(n7093) );
  BUFFD0 U7087 ( .I(n7095), .Z(n7094) );
  BUFFD0 U7088 ( .I(n7096), .Z(n7095) );
  BUFFD0 U7089 ( .I(n7097), .Z(n7096) );
  BUFFD0 U7090 ( .I(n7098), .Z(n7097) );
  BUFFD0 U7091 ( .I(n7099), .Z(n7098) );
  BUFFD0 U7092 ( .I(n7100), .Z(n7099) );
  BUFFD0 U7093 ( .I(n7101), .Z(n7100) );
  BUFFD0 U7094 ( .I(n7102), .Z(n7101) );
  BUFFD0 U7095 ( .I(n7103), .Z(n7102) );
  BUFFD0 U7096 ( .I(n7104), .Z(n7103) );
  BUFFD0 U7097 ( .I(n7105), .Z(n7104) );
  BUFFD0 U7098 ( .I(n7106), .Z(n7105) );
  BUFFD0 U7099 ( .I(n7107), .Z(n7106) );
  BUFFD0 U7100 ( .I(n7108), .Z(n7107) );
  BUFFD0 U7101 ( .I(n7109), .Z(n7108) );
  BUFFD0 U7102 ( .I(n7110), .Z(n7109) );
  BUFFD0 U7103 ( .I(n7111), .Z(n7110) );
  BUFFD0 U7104 ( .I(n7112), .Z(n7111) );
  BUFFD0 U7105 ( .I(n8690), .Z(n7112) );
  BUFFD0 U7106 ( .I(n7114), .Z(n7113) );
  BUFFD0 U7107 ( .I(n7115), .Z(n7114) );
  BUFFD0 U7108 ( .I(n7116), .Z(n7115) );
  BUFFD0 U7109 ( .I(n7117), .Z(n7116) );
  BUFFD0 U7110 ( .I(n7118), .Z(n7117) );
  BUFFD0 U7111 ( .I(n7119), .Z(n7118) );
  BUFFD0 U7112 ( .I(n7120), .Z(n7119) );
  BUFFD0 U7113 ( .I(n7121), .Z(n7120) );
  BUFFD0 U7114 ( .I(n7122), .Z(n7121) );
  BUFFD0 U7115 ( .I(n7123), .Z(n7122) );
  BUFFD0 U7116 ( .I(n7124), .Z(n7123) );
  BUFFD0 U7117 ( .I(n7125), .Z(n7124) );
  BUFFD0 U7118 ( .I(n7126), .Z(n7125) );
  BUFFD0 U7119 ( .I(n7127), .Z(n7126) );
  BUFFD0 U7120 ( .I(n7128), .Z(n7127) );
  BUFFD0 U7121 ( .I(n7129), .Z(n7128) );
  BUFFD0 U7122 ( .I(n7130), .Z(n7129) );
  BUFFD0 U7123 ( .I(n7131), .Z(n7130) );
  BUFFD0 U7124 ( .I(n7132), .Z(n7131) );
  BUFFD0 U7125 ( .I(n7133), .Z(n7132) );
  BUFFD0 U7126 ( .I(n7134), .Z(n7133) );
  BUFFD0 U7127 ( .I(n7135), .Z(n7134) );
  BUFFD0 U7128 ( .I(n7136), .Z(n7135) );
  BUFFD0 U7129 ( .I(n7137), .Z(n7136) );
  BUFFD0 U7130 ( .I(n7138), .Z(n7137) );
  BUFFD0 U7131 ( .I(n7139), .Z(n7138) );
  BUFFD0 U7132 ( .I(n7140), .Z(n7139) );
  BUFFD0 U7133 ( .I(n7141), .Z(n7140) );
  BUFFD0 U7134 ( .I(n7142), .Z(n7141) );
  BUFFD0 U7135 ( .I(n7143), .Z(n7142) );
  BUFFD0 U7136 ( .I(n7144), .Z(n7143) );
  BUFFD0 U7137 ( .I(n7145), .Z(n7144) );
  BUFFD0 U7138 ( .I(n7146), .Z(n7145) );
  BUFFD0 U7139 ( .I(n7147), .Z(n7146) );
  BUFFD0 U7140 ( .I(n7148), .Z(n7147) );
  BUFFD0 U7141 ( .I(n7149), .Z(n7148) );
  BUFFD0 U7142 ( .I(n7150), .Z(n7149) );
  BUFFD0 U7143 ( .I(n7151), .Z(n7150) );
  BUFFD0 U7144 ( .I(n7152), .Z(n7151) );
  BUFFD0 U7145 ( .I(n7153), .Z(n7152) );
  BUFFD0 U7146 ( .I(n7154), .Z(n7153) );
  BUFFD0 U7147 ( .I(n7155), .Z(n7154) );
  BUFFD0 U7148 ( .I(n7156), .Z(n7155) );
  BUFFD0 U7149 ( .I(n7157), .Z(n7156) );
  BUFFD0 U7150 ( .I(n7158), .Z(n7157) );
  BUFFD0 U7151 ( .I(n7159), .Z(n7158) );
  BUFFD0 U7152 ( .I(n7160), .Z(n7159) );
  BUFFD0 U7153 ( .I(n7161), .Z(n7160) );
  BUFFD0 U7154 ( .I(n7162), .Z(n7161) );
  BUFFD0 U7155 ( .I(n7163), .Z(n7162) );
  BUFFD0 U7156 ( .I(n7164), .Z(n7163) );
  BUFFD0 U7157 ( .I(n7165), .Z(n7164) );
  BUFFD0 U7158 ( .I(n7166), .Z(n7165) );
  BUFFD0 U7159 ( .I(n7167), .Z(n7166) );
  BUFFD0 U7160 ( .I(n7168), .Z(n7167) );
  BUFFD0 U7161 ( .I(n7169), .Z(n7168) );
  BUFFD0 U7162 ( .I(n7170), .Z(n7169) );
  BUFFD0 U7163 ( .I(n7171), .Z(n7170) );
  BUFFD0 U7164 ( .I(n7172), .Z(n7171) );
  BUFFD0 U7165 ( .I(n7173), .Z(n7172) );
  BUFFD0 U7166 ( .I(n7174), .Z(n7173) );
  BUFFD0 U7167 ( .I(n7175), .Z(n7174) );
  BUFFD0 U7168 ( .I(n7176), .Z(n7175) );
  BUFFD0 U7169 ( .I(n7177), .Z(n7176) );
  BUFFD0 U7170 ( .I(n7178), .Z(n7177) );
  BUFFD0 U7171 ( .I(n7179), .Z(n7178) );
  BUFFD0 U7172 ( .I(n7180), .Z(n7179) );
  BUFFD0 U7173 ( .I(n7181), .Z(n7180) );
  BUFFD0 U7174 ( .I(n7182), .Z(n7181) );
  BUFFD0 U7175 ( .I(n7183), .Z(n7182) );
  BUFFD0 U7176 ( .I(n7184), .Z(n7183) );
  BUFFD0 U7177 ( .I(n7185), .Z(n7184) );
  BUFFD0 U7178 ( .I(n7186), .Z(n7185) );
  BUFFD0 U7179 ( .I(n7187), .Z(n7186) );
  BUFFD0 U7180 ( .I(n7188), .Z(n7187) );
  BUFFD0 U7181 ( .I(n7189), .Z(n7188) );
  BUFFD0 U7182 ( .I(n7190), .Z(n7189) );
  BUFFD0 U7183 ( .I(n7191), .Z(n7190) );
  BUFFD0 U7184 ( .I(n7192), .Z(n7191) );
  BUFFD0 U7185 ( .I(n7193), .Z(n7192) );
  BUFFD0 U7186 ( .I(n7194), .Z(n7193) );
  BUFFD0 U7187 ( .I(n7195), .Z(n7194) );
  BUFFD0 U7188 ( .I(n7196), .Z(n7195) );
  BUFFD0 U7189 ( .I(n7197), .Z(n7196) );
  BUFFD0 U7190 ( .I(n7198), .Z(n7197) );
  BUFFD0 U7191 ( .I(n7199), .Z(n7198) );
  BUFFD0 U7192 ( .I(n7200), .Z(n7199) );
  BUFFD0 U7193 ( .I(n7201), .Z(n7200) );
  BUFFD0 U7194 ( .I(n7202), .Z(n7201) );
  BUFFD0 U7195 ( .I(n7203), .Z(n7202) );
  BUFFD0 U7196 ( .I(n7204), .Z(n7203) );
  BUFFD0 U7197 ( .I(n7205), .Z(n7204) );
  BUFFD0 U7198 ( .I(n7206), .Z(n7205) );
  BUFFD0 U7199 ( .I(n7207), .Z(n7206) );
  BUFFD0 U7200 ( .I(n7208), .Z(n7207) );
  BUFFD0 U7201 ( .I(n7209), .Z(n7208) );
  BUFFD0 U7202 ( .I(n7210), .Z(n7209) );
  BUFFD0 U7203 ( .I(n7211), .Z(n7210) );
  BUFFD0 U7204 ( .I(n7212), .Z(n7211) );
  BUFFD0 U7205 ( .I(n7213), .Z(n7212) );
  BUFFD0 U7206 ( .I(n7214), .Z(n7213) );
  BUFFD0 U7207 ( .I(n7215), .Z(n7214) );
  BUFFD0 U7208 ( .I(n7216), .Z(n7215) );
  BUFFD0 U7209 ( .I(n7217), .Z(n7216) );
  BUFFD0 U7210 ( .I(n7218), .Z(n7217) );
  BUFFD0 U7211 ( .I(n7219), .Z(n7218) );
  BUFFD0 U7212 ( .I(n7220), .Z(n7219) );
  BUFFD0 U7213 ( .I(n7221), .Z(n7220) );
  BUFFD0 U7214 ( .I(n7222), .Z(n7221) );
  BUFFD0 U7215 ( .I(n7223), .Z(n7222) );
  BUFFD0 U7216 ( .I(n7224), .Z(n7223) );
  BUFFD0 U7217 ( .I(n7225), .Z(n7224) );
  BUFFD0 U7218 ( .I(n7226), .Z(n7225) );
  BUFFD0 U7219 ( .I(n7227), .Z(n7226) );
  BUFFD0 U7220 ( .I(n7228), .Z(n7227) );
  BUFFD0 U7221 ( .I(n7229), .Z(n7228) );
  BUFFD0 U7222 ( .I(n7230), .Z(n7229) );
  BUFFD0 U7223 ( .I(n7231), .Z(n7230) );
  BUFFD0 U7224 ( .I(n7232), .Z(n7231) );
  BUFFD0 U7225 ( .I(n7233), .Z(n7232) );
  BUFFD0 U7226 ( .I(n7234), .Z(n7233) );
  BUFFD0 U7227 ( .I(n7235), .Z(n7234) );
  BUFFD0 U7228 ( .I(n7236), .Z(n7235) );
  BUFFD0 U7229 ( .I(n7237), .Z(n7236) );
  BUFFD0 U7230 ( .I(n7238), .Z(n7237) );
  BUFFD0 U7231 ( .I(n7239), .Z(n7238) );
  BUFFD0 U7232 ( .I(n7240), .Z(n7239) );
  BUFFD0 U7233 ( .I(n7241), .Z(n7240) );
  BUFFD0 U7234 ( .I(n7242), .Z(n7241) );
  BUFFD0 U7235 ( .I(n7243), .Z(n7242) );
  BUFFD0 U7236 ( .I(n7244), .Z(n7243) );
  BUFFD0 U7237 ( .I(n7245), .Z(n7244) );
  BUFFD0 U7238 ( .I(n7246), .Z(n7245) );
  BUFFD0 U7239 ( .I(n7247), .Z(n7246) );
  BUFFD0 U7240 ( .I(n7248), .Z(n7247) );
  BUFFD0 U7241 ( .I(n7249), .Z(n7248) );
  BUFFD0 U7242 ( .I(n7250), .Z(n7249) );
  BUFFD0 U7243 ( .I(n7251), .Z(n7250) );
  BUFFD0 U7244 ( .I(n7252), .Z(n7251) );
  BUFFD0 U7245 ( .I(n7253), .Z(n7252) );
  BUFFD0 U7246 ( .I(n7254), .Z(n7253) );
  BUFFD0 U7247 ( .I(n7256), .Z(n7254) );
  BUFFD0 U7248 ( .I(n2219), .Z(n7255) );
  BUFFD0 U7249 ( .I(n7257), .Z(n7256) );
  BUFFD0 U7250 ( .I(n7258), .Z(n7257) );
  BUFFD0 U7251 ( .I(n7259), .Z(n7258) );
  BUFFD0 U7252 ( .I(n7260), .Z(n7259) );
  BUFFD0 U7253 ( .I(n7261), .Z(n7260) );
  BUFFD0 U7254 ( .I(n7262), .Z(n7261) );
  BUFFD0 U7255 ( .I(n7263), .Z(n7262) );
  BUFFD0 U7256 ( .I(n7264), .Z(n7263) );
  BUFFD0 U7257 ( .I(n7265), .Z(n7264) );
  BUFFD0 U7258 ( .I(n7266), .Z(n7265) );
  BUFFD0 U7259 ( .I(n7267), .Z(n7266) );
  BUFFD0 U7260 ( .I(n7268), .Z(n7267) );
  BUFFD0 U7261 ( .I(n7269), .Z(n7268) );
  BUFFD0 U7262 ( .I(n7270), .Z(n7269) );
  BUFFD0 U7263 ( .I(n7271), .Z(n7270) );
  BUFFD0 U7264 ( .I(n7272), .Z(n7271) );
  BUFFD0 U7265 ( .I(n7273), .Z(n7272) );
  BUFFD0 U7266 ( .I(n7274), .Z(n7273) );
  BUFFD0 U7267 ( .I(n7275), .Z(n7274) );
  BUFFD0 U7268 ( .I(n7276), .Z(n7275) );
  BUFFD0 U7269 ( .I(n7277), .Z(n7276) );
  BUFFD0 U7270 ( .I(n7278), .Z(n7277) );
  BUFFD0 U7271 ( .I(n7279), .Z(n7278) );
  BUFFD0 U7272 ( .I(n7280), .Z(n7279) );
  BUFFD0 U7273 ( .I(n7281), .Z(n7280) );
  BUFFD0 U7274 ( .I(n7282), .Z(n7281) );
  BUFFD0 U7275 ( .I(n7283), .Z(n7282) );
  BUFFD0 U7276 ( .I(n7284), .Z(n7283) );
  BUFFD0 U7277 ( .I(n7285), .Z(n7284) );
  BUFFD0 U7278 ( .I(n7286), .Z(n7285) );
  BUFFD0 U7279 ( .I(n7287), .Z(n7286) );
  BUFFD0 U7280 ( .I(n7288), .Z(n7287) );
  BUFFD0 U7281 ( .I(n8688), .Z(n7288) );
  BUFFD0 U7282 ( .I(n8750), .Z(n7289) );
  BUFFD0 U7283 ( .I(n7291), .Z(n7290) );
  BUFFD0 U7284 ( .I(n7292), .Z(n7291) );
  BUFFD0 U7285 ( .I(n7293), .Z(n7292) );
  BUFFD0 U7286 ( .I(n7294), .Z(n7293) );
  BUFFD0 U7287 ( .I(n7295), .Z(n7294) );
  BUFFD0 U7288 ( .I(n7296), .Z(n7295) );
  BUFFD0 U7289 ( .I(n7297), .Z(n7296) );
  BUFFD0 U7290 ( .I(n7298), .Z(n7297) );
  BUFFD0 U7291 ( .I(n7299), .Z(n7298) );
  BUFFD0 U7292 ( .I(n7300), .Z(n7299) );
  BUFFD0 U7293 ( .I(n7301), .Z(n7300) );
  BUFFD0 U7294 ( .I(n7302), .Z(n7301) );
  BUFFD0 U7295 ( .I(n7303), .Z(n7302) );
  BUFFD0 U7296 ( .I(n7304), .Z(n7303) );
  BUFFD0 U7297 ( .I(n7305), .Z(n7304) );
  BUFFD0 U7298 ( .I(n7306), .Z(n7305) );
  BUFFD0 U7299 ( .I(n7307), .Z(n7306) );
  BUFFD0 U7300 ( .I(n7308), .Z(n7307) );
  BUFFD0 U7301 ( .I(n7309), .Z(n7308) );
  BUFFD0 U7302 ( .I(n7310), .Z(n7309) );
  BUFFD0 U7303 ( .I(n7311), .Z(n7310) );
  BUFFD0 U7304 ( .I(n7312), .Z(n7311) );
  BUFFD0 U7305 ( .I(n7313), .Z(n7312) );
  BUFFD0 U7306 ( .I(n7314), .Z(n7313) );
  BUFFD0 U7307 ( .I(n7315), .Z(n7314) );
  BUFFD0 U7308 ( .I(n7316), .Z(n7315) );
  BUFFD0 U7309 ( .I(n7317), .Z(n7316) );
  BUFFD0 U7310 ( .I(n7318), .Z(n7317) );
  BUFFD0 U7311 ( .I(n7319), .Z(n7318) );
  BUFFD0 U7312 ( .I(n7320), .Z(n7319) );
  BUFFD0 U7313 ( .I(n7321), .Z(n7320) );
  BUFFD0 U7314 ( .I(n7322), .Z(n7321) );
  BUFFD0 U7315 ( .I(n7323), .Z(n7322) );
  BUFFD0 U7316 ( .I(n7324), .Z(n7323) );
  BUFFD0 U7317 ( .I(n7325), .Z(n7324) );
  BUFFD0 U7318 ( .I(n7326), .Z(n7325) );
  BUFFD0 U7319 ( .I(n7327), .Z(n7326) );
  BUFFD0 U7320 ( .I(n7328), .Z(n7327) );
  BUFFD0 U7321 ( .I(n7329), .Z(n7328) );
  BUFFD0 U7322 ( .I(n7330), .Z(n7329) );
  BUFFD0 U7323 ( .I(n7331), .Z(n7330) );
  BUFFD0 U7324 ( .I(n7332), .Z(n7331) );
  BUFFD0 U7325 ( .I(n7333), .Z(n7332) );
  BUFFD0 U7326 ( .I(n7334), .Z(n7333) );
  BUFFD0 U7327 ( .I(n7335), .Z(n7334) );
  BUFFD0 U7328 ( .I(n7336), .Z(n7335) );
  BUFFD0 U7329 ( .I(n7337), .Z(n7336) );
  BUFFD0 U7330 ( .I(n7338), .Z(n7337) );
  BUFFD0 U7331 ( .I(n7339), .Z(n7338) );
  BUFFD0 U7332 ( .I(n7340), .Z(n7339) );
  BUFFD0 U7333 ( .I(n7341), .Z(n7340) );
  BUFFD0 U7334 ( .I(n7342), .Z(n7341) );
  BUFFD0 U7335 ( .I(n7343), .Z(n7342) );
  BUFFD0 U7336 ( .I(n7344), .Z(n7343) );
  BUFFD0 U7337 ( .I(n7345), .Z(n7344) );
  BUFFD0 U7338 ( .I(n7346), .Z(n7345) );
  BUFFD0 U7339 ( .I(n7347), .Z(n7346) );
  BUFFD0 U7340 ( .I(n7348), .Z(n7347) );
  BUFFD0 U7341 ( .I(n7349), .Z(n7348) );
  BUFFD0 U7342 ( .I(n7350), .Z(n7349) );
  BUFFD0 U7343 ( .I(n7351), .Z(n7350) );
  BUFFD0 U7344 ( .I(n7352), .Z(n7351) );
  BUFFD0 U7345 ( .I(n7353), .Z(n7352) );
  BUFFD0 U7346 ( .I(n7354), .Z(n7353) );
  BUFFD0 U7347 ( .I(n7355), .Z(n7354) );
  BUFFD0 U7348 ( .I(n7356), .Z(n7355) );
  BUFFD0 U7349 ( .I(n7357), .Z(n7356) );
  BUFFD0 U7350 ( .I(n7358), .Z(n7357) );
  BUFFD0 U7351 ( .I(n7359), .Z(n7358) );
  BUFFD0 U7352 ( .I(n7360), .Z(n7359) );
  BUFFD0 U7353 ( .I(n7361), .Z(n7360) );
  BUFFD0 U7354 ( .I(n7362), .Z(n7361) );
  BUFFD0 U7355 ( .I(n7363), .Z(n7362) );
  BUFFD0 U7356 ( .I(n7364), .Z(n7363) );
  BUFFD0 U7357 ( .I(n7365), .Z(n7364) );
  BUFFD0 U7358 ( .I(n7366), .Z(n7365) );
  BUFFD0 U7359 ( .I(n7367), .Z(n7366) );
  BUFFD0 U7360 ( .I(n7368), .Z(n7367) );
  BUFFD0 U7361 ( .I(n7369), .Z(n7368) );
  BUFFD0 U7362 ( .I(n7370), .Z(n7369) );
  BUFFD0 U7363 ( .I(n7371), .Z(n7370) );
  BUFFD0 U7364 ( .I(n7372), .Z(n7371) );
  BUFFD0 U7365 ( .I(n7373), .Z(n7372) );
  BUFFD0 U7366 ( .I(n7374), .Z(n7373) );
  BUFFD0 U7367 ( .I(n7375), .Z(n7374) );
  BUFFD0 U7368 ( .I(n7376), .Z(n7375) );
  BUFFD0 U7369 ( .I(n7377), .Z(n7376) );
  BUFFD0 U7370 ( .I(n7378), .Z(n7377) );
  BUFFD0 U7371 ( .I(n7379), .Z(n7378) );
  BUFFD0 U7372 ( .I(n7380), .Z(n7379) );
  BUFFD0 U7373 ( .I(n7381), .Z(n7380) );
  BUFFD0 U7374 ( .I(n7382), .Z(n7381) );
  BUFFD0 U7375 ( .I(n7383), .Z(n7382) );
  BUFFD0 U7376 ( .I(n7384), .Z(n7383) );
  BUFFD0 U7377 ( .I(n7385), .Z(n7384) );
  BUFFD0 U7378 ( .I(n7386), .Z(n7385) );
  BUFFD0 U7379 ( .I(n7387), .Z(n7386) );
  BUFFD0 U7380 ( .I(n7388), .Z(n7387) );
  BUFFD0 U7381 ( .I(n7389), .Z(n7388) );
  BUFFD0 U7382 ( .I(n7390), .Z(n7389) );
  BUFFD0 U7383 ( .I(n7391), .Z(n7390) );
  BUFFD0 U7384 ( .I(n7392), .Z(n7391) );
  BUFFD0 U7385 ( .I(n7393), .Z(n7392) );
  BUFFD0 U7386 ( .I(n7394), .Z(n7393) );
  BUFFD0 U7387 ( .I(n7395), .Z(n7394) );
  BUFFD0 U7388 ( .I(n7396), .Z(n7395) );
  BUFFD0 U7389 ( .I(n7397), .Z(n7396) );
  BUFFD0 U7390 ( .I(n7398), .Z(n7397) );
  BUFFD0 U7391 ( .I(n7399), .Z(n7398) );
  BUFFD0 U7392 ( .I(n7400), .Z(n7399) );
  BUFFD0 U7393 ( .I(n7401), .Z(n7400) );
  BUFFD0 U7394 ( .I(n7402), .Z(n7401) );
  BUFFD0 U7395 ( .I(n7403), .Z(n7402) );
  BUFFD0 U7396 ( .I(n7404), .Z(n7403) );
  BUFFD0 U7397 ( .I(n7405), .Z(n7404) );
  BUFFD0 U7398 ( .I(n7406), .Z(n7405) );
  BUFFD0 U7399 ( .I(n7407), .Z(n7406) );
  BUFFD0 U7400 ( .I(n7408), .Z(n7407) );
  BUFFD0 U7401 ( .I(n7409), .Z(n7408) );
  BUFFD0 U7402 ( .I(n7410), .Z(n7409) );
  BUFFD0 U7403 ( .I(n7411), .Z(n7410) );
  BUFFD0 U7404 ( .I(n7412), .Z(n7411) );
  BUFFD0 U7405 ( .I(n7413), .Z(n7412) );
  BUFFD0 U7406 ( .I(n7414), .Z(n7413) );
  BUFFD0 U7407 ( .I(n7415), .Z(n7414) );
  BUFFD0 U7408 ( .I(n7416), .Z(n7415) );
  BUFFD0 U7409 ( .I(n7417), .Z(n7416) );
  BUFFD0 U7410 ( .I(n7418), .Z(n7417) );
  BUFFD0 U7411 ( .I(n7419), .Z(n7418) );
  BUFFD0 U7412 ( .I(n7420), .Z(n7419) );
  BUFFD0 U7413 ( .I(n7421), .Z(n7420) );
  BUFFD0 U7414 ( .I(n7422), .Z(n7421) );
  BUFFD0 U7415 ( .I(n7423), .Z(n7422) );
  BUFFD0 U7416 ( .I(n7424), .Z(n7423) );
  BUFFD0 U7417 ( .I(n7425), .Z(n7424) );
  BUFFD0 U7418 ( .I(n7426), .Z(n7425) );
  BUFFD0 U7419 ( .I(n7427), .Z(n7426) );
  BUFFD0 U7420 ( .I(n7428), .Z(n7427) );
  BUFFD0 U7421 ( .I(n7429), .Z(n7428) );
  BUFFD0 U7422 ( .I(n7430), .Z(n7429) );
  BUFFD0 U7423 ( .I(n7431), .Z(n7430) );
  BUFFD0 U7424 ( .I(n7432), .Z(n7431) );
  BUFFD0 U7425 ( .I(n7433), .Z(n7432) );
  BUFFD0 U7426 ( .I(n7434), .Z(n7433) );
  BUFFD0 U7427 ( .I(n7435), .Z(n7434) );
  BUFFD0 U7428 ( .I(n7436), .Z(n7435) );
  BUFFD0 U7429 ( .I(n7437), .Z(n7436) );
  BUFFD0 U7430 ( .I(n7438), .Z(n7437) );
  BUFFD0 U7431 ( .I(n7439), .Z(n7438) );
  BUFFD0 U7432 ( .I(n7440), .Z(n7439) );
  BUFFD0 U7433 ( .I(n7441), .Z(n7440) );
  BUFFD0 U7434 ( .I(n7442), .Z(n7441) );
  BUFFD0 U7435 ( .I(n7443), .Z(n7442) );
  BUFFD0 U7436 ( .I(n7444), .Z(n7443) );
  BUFFD0 U7437 ( .I(n7445), .Z(n7444) );
  BUFFD0 U7438 ( .I(n7446), .Z(n7445) );
  BUFFD0 U7439 ( .I(n7447), .Z(n7446) );
  BUFFD0 U7440 ( .I(n7448), .Z(n7447) );
  BUFFD0 U7441 ( .I(n7449), .Z(n7448) );
  BUFFD0 U7442 ( .I(n7450), .Z(n7449) );
  BUFFD0 U7443 ( .I(n7451), .Z(n7450) );
  BUFFD0 U7444 ( .I(n7452), .Z(n7451) );
  BUFFD0 U7445 ( .I(n7453), .Z(n7452) );
  BUFFD0 U7446 ( .I(n7454), .Z(n7453) );
  BUFFD0 U7447 ( .I(n7455), .Z(n7454) );
  BUFFD0 U7448 ( .I(n7456), .Z(n7455) );
  BUFFD0 U7449 ( .I(n7457), .Z(n7456) );
  BUFFD0 U7450 ( .I(n7458), .Z(n7457) );
  BUFFD0 U7451 ( .I(n7459), .Z(n7458) );
  BUFFD0 U7452 ( .I(n7460), .Z(n7459) );
  BUFFD0 U7453 ( .I(n7461), .Z(n7460) );
  BUFFD0 U7454 ( .I(n7462), .Z(n7461) );
  BUFFD0 U7455 ( .I(n7463), .Z(n7462) );
  BUFFD0 U7456 ( .I(n7464), .Z(n7463) );
  BUFFD0 U7457 ( .I(n7465), .Z(n7464) );
  BUFFD0 U7458 ( .I(n8751), .Z(n7465) );
  BUFFD0 U7459 ( .I(n8745), .Z(n7466) );
  BUFFD0 U7460 ( .I(n7468), .Z(n7467) );
  BUFFD0 U7461 ( .I(n7469), .Z(n7468) );
  BUFFD0 U7462 ( .I(n7470), .Z(n7469) );
  BUFFD0 U7463 ( .I(n7471), .Z(n7470) );
  BUFFD0 U7464 ( .I(n7472), .Z(n7471) );
  BUFFD0 U7465 ( .I(n7473), .Z(n7472) );
  BUFFD0 U7466 ( .I(n7474), .Z(n7473) );
  BUFFD0 U7467 ( .I(n7475), .Z(n7474) );
  BUFFD0 U7468 ( .I(n7476), .Z(n7475) );
  BUFFD0 U7469 ( .I(n7477), .Z(n7476) );
  BUFFD0 U7470 ( .I(n7478), .Z(n7477) );
  BUFFD0 U7471 ( .I(n7479), .Z(n7478) );
  BUFFD0 U7472 ( .I(n7480), .Z(n7479) );
  BUFFD0 U7473 ( .I(n7481), .Z(n7480) );
  BUFFD0 U7474 ( .I(n7482), .Z(n7481) );
  BUFFD0 U7475 ( .I(n7483), .Z(n7482) );
  BUFFD0 U7476 ( .I(n7484), .Z(n7483) );
  BUFFD0 U7477 ( .I(n7485), .Z(n7484) );
  BUFFD0 U7478 ( .I(n7486), .Z(n7485) );
  BUFFD0 U7479 ( .I(n7487), .Z(n7486) );
  BUFFD0 U7480 ( .I(n7488), .Z(n7487) );
  BUFFD0 U7481 ( .I(n7489), .Z(n7488) );
  BUFFD0 U7482 ( .I(n7490), .Z(n7489) );
  BUFFD0 U7483 ( .I(n7491), .Z(n7490) );
  BUFFD0 U7484 ( .I(n7492), .Z(n7491) );
  BUFFD0 U7485 ( .I(n7493), .Z(n7492) );
  BUFFD0 U7486 ( .I(n7494), .Z(n7493) );
  BUFFD0 U7487 ( .I(n7495), .Z(n7494) );
  BUFFD0 U7488 ( .I(n7496), .Z(n7495) );
  BUFFD0 U7489 ( .I(n7497), .Z(n7496) );
  BUFFD0 U7490 ( .I(n7498), .Z(n7497) );
  BUFFD0 U7491 ( .I(n7499), .Z(n7498) );
  BUFFD0 U7492 ( .I(n7500), .Z(n7499) );
  BUFFD0 U7493 ( .I(n7501), .Z(n7500) );
  BUFFD0 U7494 ( .I(n7502), .Z(n7501) );
  BUFFD0 U7495 ( .I(n7503), .Z(n7502) );
  BUFFD0 U7496 ( .I(n7504), .Z(n7503) );
  BUFFD0 U7497 ( .I(n7505), .Z(n7504) );
  BUFFD0 U7498 ( .I(n7506), .Z(n7505) );
  BUFFD0 U7499 ( .I(n7507), .Z(n7506) );
  BUFFD0 U7500 ( .I(n7508), .Z(n7507) );
  BUFFD0 U7501 ( .I(n7509), .Z(n7508) );
  BUFFD0 U7502 ( .I(n7510), .Z(n7509) );
  BUFFD0 U7503 ( .I(n7511), .Z(n7510) );
  BUFFD0 U7504 ( .I(n7512), .Z(n7511) );
  BUFFD0 U7505 ( .I(n7513), .Z(n7512) );
  BUFFD0 U7506 ( .I(n7514), .Z(n7513) );
  BUFFD0 U7507 ( .I(n7515), .Z(n7514) );
  BUFFD0 U7508 ( .I(n7516), .Z(n7515) );
  BUFFD0 U7509 ( .I(n7517), .Z(n7516) );
  BUFFD0 U7510 ( .I(n7518), .Z(n7517) );
  BUFFD0 U7511 ( .I(n7519), .Z(n7518) );
  BUFFD0 U7512 ( .I(n7520), .Z(n7519) );
  BUFFD0 U7513 ( .I(n7521), .Z(n7520) );
  BUFFD0 U7514 ( .I(n7522), .Z(n7521) );
  BUFFD0 U7515 ( .I(n7523), .Z(n7522) );
  BUFFD0 U7516 ( .I(n7524), .Z(n7523) );
  BUFFD0 U7517 ( .I(n7525), .Z(n7524) );
  BUFFD0 U7518 ( .I(n7526), .Z(n7525) );
  BUFFD0 U7519 ( .I(n7527), .Z(n7526) );
  BUFFD0 U7520 ( .I(n7528), .Z(n7527) );
  BUFFD0 U7521 ( .I(n7529), .Z(n7528) );
  BUFFD0 U7522 ( .I(n7530), .Z(n7529) );
  BUFFD0 U7523 ( .I(n7531), .Z(n7530) );
  BUFFD0 U7524 ( .I(n7532), .Z(n7531) );
  BUFFD0 U7525 ( .I(n7533), .Z(n7532) );
  BUFFD0 U7526 ( .I(n7534), .Z(n7533) );
  BUFFD0 U7527 ( .I(n7535), .Z(n7534) );
  BUFFD0 U7528 ( .I(n7536), .Z(n7535) );
  BUFFD0 U7529 ( .I(n7537), .Z(n7536) );
  BUFFD0 U7530 ( .I(n7538), .Z(n7537) );
  BUFFD0 U7531 ( .I(n7539), .Z(n7538) );
  BUFFD0 U7532 ( .I(n7540), .Z(n7539) );
  BUFFD0 U7533 ( .I(n7541), .Z(n7540) );
  BUFFD0 U7534 ( .I(n7542), .Z(n7541) );
  BUFFD0 U7535 ( .I(n7543), .Z(n7542) );
  BUFFD0 U7536 ( .I(n7544), .Z(n7543) );
  BUFFD0 U7537 ( .I(n7545), .Z(n7544) );
  BUFFD0 U7538 ( .I(n7546), .Z(n7545) );
  BUFFD0 U7539 ( .I(n7547), .Z(n7546) );
  BUFFD0 U7540 ( .I(n7548), .Z(n7547) );
  BUFFD0 U7541 ( .I(n7549), .Z(n7548) );
  BUFFD0 U7542 ( .I(n7550), .Z(n7549) );
  BUFFD0 U7543 ( .I(n7551), .Z(n7550) );
  BUFFD0 U7544 ( .I(n7552), .Z(n7551) );
  BUFFD0 U7545 ( .I(n7553), .Z(n7552) );
  BUFFD0 U7546 ( .I(n7554), .Z(n7553) );
  BUFFD0 U7547 ( .I(n7555), .Z(n7554) );
  BUFFD0 U7548 ( .I(n7556), .Z(n7555) );
  BUFFD0 U7549 ( .I(n7557), .Z(n7556) );
  BUFFD0 U7550 ( .I(n7558), .Z(n7557) );
  BUFFD0 U7551 ( .I(n7559), .Z(n7558) );
  BUFFD0 U7552 ( .I(n7560), .Z(n7559) );
  BUFFD0 U7553 ( .I(n7561), .Z(n7560) );
  BUFFD0 U7554 ( .I(n7562), .Z(n7561) );
  BUFFD0 U7555 ( .I(n7563), .Z(n7562) );
  BUFFD0 U7556 ( .I(n7564), .Z(n7563) );
  BUFFD0 U7557 ( .I(n7565), .Z(n7564) );
  BUFFD0 U7558 ( .I(n7566), .Z(n7565) );
  BUFFD0 U7559 ( .I(n7567), .Z(n7566) );
  BUFFD0 U7560 ( .I(n7568), .Z(n7567) );
  BUFFD0 U7561 ( .I(n7569), .Z(n7568) );
  BUFFD0 U7562 ( .I(n7570), .Z(n7569) );
  BUFFD0 U7563 ( .I(n7571), .Z(n7570) );
  BUFFD0 U7564 ( .I(n7572), .Z(n7571) );
  BUFFD0 U7565 ( .I(n7573), .Z(n7572) );
  BUFFD0 U7566 ( .I(n7574), .Z(n7573) );
  BUFFD0 U7567 ( .I(n7575), .Z(n7574) );
  BUFFD0 U7568 ( .I(n7576), .Z(n7575) );
  BUFFD0 U7569 ( .I(n7577), .Z(n7576) );
  BUFFD0 U7570 ( .I(n7578), .Z(n7577) );
  BUFFD0 U7571 ( .I(n7579), .Z(n7578) );
  BUFFD0 U7572 ( .I(n7580), .Z(n7579) );
  BUFFD0 U7573 ( .I(n7581), .Z(n7580) );
  BUFFD0 U7574 ( .I(n7582), .Z(n7581) );
  BUFFD0 U7575 ( .I(n7583), .Z(n7582) );
  BUFFD0 U7576 ( .I(n7584), .Z(n7583) );
  BUFFD0 U7577 ( .I(n7585), .Z(n7584) );
  BUFFD0 U7578 ( .I(n7586), .Z(n7585) );
  BUFFD0 U7579 ( .I(n7587), .Z(n7586) );
  BUFFD0 U7580 ( .I(n7588), .Z(n7587) );
  BUFFD0 U7581 ( .I(n7589), .Z(n7588) );
  BUFFD0 U7582 ( .I(n7590), .Z(n7589) );
  BUFFD0 U7583 ( .I(n7591), .Z(n7590) );
  BUFFD0 U7584 ( .I(n7592), .Z(n7591) );
  BUFFD0 U7585 ( .I(n7593), .Z(n7592) );
  BUFFD0 U7586 ( .I(n7594), .Z(n7593) );
  BUFFD0 U7587 ( .I(n7595), .Z(n7594) );
  BUFFD0 U7588 ( .I(n7596), .Z(n7595) );
  BUFFD0 U7589 ( .I(n7597), .Z(n7596) );
  BUFFD0 U7590 ( .I(n7598), .Z(n7597) );
  BUFFD0 U7591 ( .I(n7599), .Z(n7598) );
  BUFFD0 U7592 ( .I(n7600), .Z(n7599) );
  BUFFD0 U7593 ( .I(n7601), .Z(n7600) );
  BUFFD0 U7594 ( .I(n7602), .Z(n7601) );
  BUFFD0 U7595 ( .I(n7603), .Z(n7602) );
  BUFFD0 U7596 ( .I(n7604), .Z(n7603) );
  BUFFD0 U7597 ( .I(n7605), .Z(n7604) );
  BUFFD0 U7598 ( .I(n7606), .Z(n7605) );
  BUFFD0 U7599 ( .I(n7607), .Z(n7606) );
  BUFFD0 U7600 ( .I(n7608), .Z(n7607) );
  BUFFD0 U7601 ( .I(n7609), .Z(n7608) );
  BUFFD0 U7602 ( .I(n7610), .Z(n7609) );
  BUFFD0 U7603 ( .I(n7611), .Z(n7610) );
  BUFFD0 U7604 ( .I(n7612), .Z(n7611) );
  BUFFD0 U7605 ( .I(n7613), .Z(n7612) );
  BUFFD0 U7606 ( .I(n7614), .Z(n7613) );
  BUFFD0 U7607 ( .I(n7615), .Z(n7614) );
  BUFFD0 U7608 ( .I(n7616), .Z(n7615) );
  BUFFD0 U7609 ( .I(n7617), .Z(n7616) );
  BUFFD0 U7610 ( .I(n7618), .Z(n7617) );
  BUFFD0 U7611 ( .I(n7619), .Z(n7618) );
  BUFFD0 U7612 ( .I(n7620), .Z(n7619) );
  BUFFD0 U7613 ( .I(n7621), .Z(n7620) );
  BUFFD0 U7614 ( .I(n7622), .Z(n7621) );
  BUFFD0 U7615 ( .I(n7623), .Z(n7622) );
  BUFFD0 U7616 ( .I(n7624), .Z(n7623) );
  BUFFD0 U7617 ( .I(n7625), .Z(n7624) );
  BUFFD0 U7618 ( .I(n7626), .Z(n7625) );
  BUFFD0 U7619 ( .I(n7627), .Z(n7626) );
  BUFFD0 U7620 ( .I(n7628), .Z(n7627) );
  BUFFD0 U7621 ( .I(n7629), .Z(n7628) );
  BUFFD0 U7622 ( .I(n7630), .Z(n7629) );
  BUFFD0 U7623 ( .I(n7631), .Z(n7630) );
  BUFFD0 U7624 ( .I(n7632), .Z(n7631) );
  BUFFD0 U7625 ( .I(n7633), .Z(n7632) );
  BUFFD0 U7626 ( .I(n7634), .Z(n7633) );
  BUFFD0 U7627 ( .I(n7635), .Z(n7634) );
  BUFFD0 U7628 ( .I(n7636), .Z(n7635) );
  BUFFD0 U7629 ( .I(n7637), .Z(n7636) );
  BUFFD0 U7630 ( .I(n7638), .Z(n7637) );
  BUFFD0 U7631 ( .I(n7639), .Z(n7638) );
  BUFFD0 U7632 ( .I(n7640), .Z(n7639) );
  BUFFD0 U7633 ( .I(n7641), .Z(n7640) );
  BUFFD0 U7634 ( .I(n7642), .Z(n7641) );
  BUFFD0 U7635 ( .I(n7643), .Z(n7642) );
  BUFFD0 U7636 ( .I(n7644), .Z(n7643) );
  BUFFD0 U7637 ( .I(n8746), .Z(n7644) );
  BUFFD0 U7638 ( .I(n8747), .Z(n7645) );
  BUFFD0 U7639 ( .I(n7647), .Z(n7646) );
  BUFFD0 U7640 ( .I(n7648), .Z(n7647) );
  BUFFD0 U7641 ( .I(n7649), .Z(n7648) );
  BUFFD0 U7642 ( .I(n7650), .Z(n7649) );
  BUFFD0 U7643 ( .I(n7651), .Z(n7650) );
  BUFFD0 U7644 ( .I(n7652), .Z(n7651) );
  BUFFD0 U7645 ( .I(n7653), .Z(n7652) );
  BUFFD0 U7646 ( .I(n7654), .Z(n7653) );
  BUFFD0 U7647 ( .I(n7655), .Z(n7654) );
  BUFFD0 U7648 ( .I(n7656), .Z(n7655) );
  BUFFD0 U7649 ( .I(n7657), .Z(n7656) );
  BUFFD0 U7650 ( .I(n7658), .Z(n7657) );
  BUFFD0 U7651 ( .I(n7659), .Z(n7658) );
  BUFFD0 U7652 ( .I(n7660), .Z(n7659) );
  BUFFD0 U7653 ( .I(n7661), .Z(n7660) );
  BUFFD0 U7654 ( .I(n7662), .Z(n7661) );
  BUFFD0 U7655 ( .I(n7663), .Z(n7662) );
  BUFFD0 U7656 ( .I(n7664), .Z(n7663) );
  BUFFD0 U7657 ( .I(n7665), .Z(n7664) );
  BUFFD0 U7658 ( .I(n7666), .Z(n7665) );
  BUFFD0 U7659 ( .I(n7667), .Z(n7666) );
  BUFFD0 U7660 ( .I(n7668), .Z(n7667) );
  BUFFD0 U7661 ( .I(n7669), .Z(n7668) );
  BUFFD0 U7662 ( .I(n7670), .Z(n7669) );
  BUFFD0 U7663 ( .I(n7671), .Z(n7670) );
  BUFFD0 U7664 ( .I(n7672), .Z(n7671) );
  BUFFD0 U7665 ( .I(n7673), .Z(n7672) );
  BUFFD0 U7666 ( .I(n7674), .Z(n7673) );
  BUFFD0 U7667 ( .I(n7675), .Z(n7674) );
  BUFFD0 U7668 ( .I(n7676), .Z(n7675) );
  BUFFD0 U7669 ( .I(n7677), .Z(n7676) );
  BUFFD0 U7670 ( .I(n7678), .Z(n7677) );
  BUFFD0 U7671 ( .I(n7679), .Z(n7678) );
  BUFFD0 U7672 ( .I(n7680), .Z(n7679) );
  BUFFD0 U7673 ( .I(n7681), .Z(n7680) );
  BUFFD0 U7674 ( .I(n7682), .Z(n7681) );
  BUFFD0 U7675 ( .I(n7683), .Z(n7682) );
  BUFFD0 U7676 ( .I(n7684), .Z(n7683) );
  BUFFD0 U7677 ( .I(n7685), .Z(n7684) );
  BUFFD0 U7678 ( .I(n7686), .Z(n7685) );
  BUFFD0 U7679 ( .I(n7687), .Z(n7686) );
  BUFFD0 U7680 ( .I(n7688), .Z(n7687) );
  BUFFD0 U7681 ( .I(n7689), .Z(n7688) );
  BUFFD0 U7682 ( .I(n7690), .Z(n7689) );
  BUFFD0 U7683 ( .I(n7691), .Z(n7690) );
  BUFFD0 U7684 ( .I(n7692), .Z(n7691) );
  BUFFD0 U7685 ( .I(n7693), .Z(n7692) );
  BUFFD0 U7686 ( .I(n7694), .Z(n7693) );
  BUFFD0 U7687 ( .I(n7695), .Z(n7694) );
  BUFFD0 U7688 ( .I(n7696), .Z(n7695) );
  BUFFD0 U7689 ( .I(n7697), .Z(n7696) );
  BUFFD0 U7690 ( .I(n7698), .Z(n7697) );
  BUFFD0 U7691 ( .I(n7699), .Z(n7698) );
  BUFFD0 U7692 ( .I(n7700), .Z(n7699) );
  BUFFD0 U7693 ( .I(n7701), .Z(n7700) );
  BUFFD0 U7694 ( .I(n7702), .Z(n7701) );
  BUFFD0 U7695 ( .I(n7703), .Z(n7702) );
  BUFFD0 U7696 ( .I(n7704), .Z(n7703) );
  BUFFD0 U7697 ( .I(n7705), .Z(n7704) );
  BUFFD0 U7698 ( .I(n7706), .Z(n7705) );
  BUFFD0 U7699 ( .I(n7707), .Z(n7706) );
  BUFFD0 U7700 ( .I(n7708), .Z(n7707) );
  BUFFD0 U7701 ( .I(n7709), .Z(n7708) );
  BUFFD0 U7702 ( .I(n7710), .Z(n7709) );
  BUFFD0 U7703 ( .I(n7711), .Z(n7710) );
  BUFFD0 U7704 ( .I(n7712), .Z(n7711) );
  BUFFD0 U7705 ( .I(n7713), .Z(n7712) );
  BUFFD0 U7706 ( .I(n7714), .Z(n7713) );
  BUFFD0 U7707 ( .I(n7715), .Z(n7714) );
  BUFFD0 U7708 ( .I(n7716), .Z(n7715) );
  BUFFD0 U7709 ( .I(n7717), .Z(n7716) );
  BUFFD0 U7710 ( .I(n7718), .Z(n7717) );
  BUFFD0 U7711 ( .I(n7719), .Z(n7718) );
  BUFFD0 U7712 ( .I(n7720), .Z(n7719) );
  BUFFD0 U7713 ( .I(n7721), .Z(n7720) );
  BUFFD0 U7714 ( .I(n7722), .Z(n7721) );
  BUFFD0 U7715 ( .I(n7723), .Z(n7722) );
  BUFFD0 U7716 ( .I(n7724), .Z(n7723) );
  BUFFD0 U7717 ( .I(n7725), .Z(n7724) );
  BUFFD0 U7718 ( .I(n7726), .Z(n7725) );
  BUFFD0 U7719 ( .I(n7727), .Z(n7726) );
  BUFFD0 U7720 ( .I(n7728), .Z(n7727) );
  BUFFD0 U7721 ( .I(n7729), .Z(n7728) );
  BUFFD0 U7722 ( .I(n7730), .Z(n7729) );
  BUFFD0 U7723 ( .I(n7731), .Z(n7730) );
  BUFFD0 U7724 ( .I(n7732), .Z(n7731) );
  BUFFD0 U7725 ( .I(n7733), .Z(n7732) );
  BUFFD0 U7726 ( .I(n7734), .Z(n7733) );
  BUFFD0 U7727 ( .I(n7735), .Z(n7734) );
  BUFFD0 U7728 ( .I(n7736), .Z(n7735) );
  BUFFD0 U7729 ( .I(n7737), .Z(n7736) );
  BUFFD0 U7730 ( .I(n7738), .Z(n7737) );
  BUFFD0 U7731 ( .I(n7739), .Z(n7738) );
  BUFFD0 U7732 ( .I(n7740), .Z(n7739) );
  BUFFD0 U7733 ( .I(n7741), .Z(n7740) );
  BUFFD0 U7734 ( .I(n7742), .Z(n7741) );
  BUFFD0 U7735 ( .I(n7743), .Z(n7742) );
  BUFFD0 U7736 ( .I(n7744), .Z(n7743) );
  BUFFD0 U7737 ( .I(n7745), .Z(n7744) );
  BUFFD0 U7738 ( .I(n7746), .Z(n7745) );
  BUFFD0 U7739 ( .I(n7747), .Z(n7746) );
  BUFFD0 U7740 ( .I(n7748), .Z(n7747) );
  BUFFD0 U7741 ( .I(n7749), .Z(n7748) );
  BUFFD0 U7742 ( .I(n7750), .Z(n7749) );
  BUFFD0 U7743 ( .I(n7751), .Z(n7750) );
  BUFFD0 U7744 ( .I(n7752), .Z(n7751) );
  BUFFD0 U7745 ( .I(n7753), .Z(n7752) );
  BUFFD0 U7746 ( .I(n7754), .Z(n7753) );
  BUFFD0 U7747 ( .I(n7755), .Z(n7754) );
  BUFFD0 U7748 ( .I(n7756), .Z(n7755) );
  BUFFD0 U7749 ( .I(n7757), .Z(n7756) );
  BUFFD0 U7750 ( .I(n7758), .Z(n7757) );
  BUFFD0 U7751 ( .I(n7759), .Z(n7758) );
  BUFFD0 U7752 ( .I(n7760), .Z(n7759) );
  BUFFD0 U7753 ( .I(n7761), .Z(n7760) );
  BUFFD0 U7754 ( .I(n7762), .Z(n7761) );
  BUFFD0 U7755 ( .I(n7763), .Z(n7762) );
  BUFFD0 U7756 ( .I(n7764), .Z(n7763) );
  BUFFD0 U7757 ( .I(n7765), .Z(n7764) );
  BUFFD0 U7758 ( .I(n7766), .Z(n7765) );
  BUFFD0 U7759 ( .I(n7767), .Z(n7766) );
  BUFFD0 U7760 ( .I(n7768), .Z(n7767) );
  BUFFD0 U7761 ( .I(n7769), .Z(n7768) );
  BUFFD0 U7762 ( .I(n7770), .Z(n7769) );
  BUFFD0 U7763 ( .I(n7771), .Z(n7770) );
  BUFFD0 U7764 ( .I(n7772), .Z(n7771) );
  BUFFD0 U7765 ( .I(n7773), .Z(n7772) );
  BUFFD0 U7766 ( .I(n7774), .Z(n7773) );
  BUFFD0 U7767 ( .I(n7775), .Z(n7774) );
  BUFFD0 U7768 ( .I(n7776), .Z(n7775) );
  BUFFD0 U7769 ( .I(n7777), .Z(n7776) );
  BUFFD0 U7770 ( .I(n7778), .Z(n7777) );
  BUFFD0 U7771 ( .I(n7779), .Z(n7778) );
  BUFFD0 U7772 ( .I(n7780), .Z(n7779) );
  BUFFD0 U7773 ( .I(n7781), .Z(n7780) );
  BUFFD0 U7774 ( .I(n7782), .Z(n7781) );
  BUFFD0 U7775 ( .I(n7783), .Z(n7782) );
  BUFFD0 U7776 ( .I(n7784), .Z(n7783) );
  BUFFD0 U7777 ( .I(n7785), .Z(n7784) );
  BUFFD0 U7778 ( .I(n7786), .Z(n7785) );
  BUFFD0 U7779 ( .I(n7787), .Z(n7786) );
  BUFFD0 U7780 ( .I(n7788), .Z(n7787) );
  BUFFD0 U7781 ( .I(n7789), .Z(n7788) );
  BUFFD0 U7782 ( .I(n7790), .Z(n7789) );
  BUFFD0 U7783 ( .I(n7791), .Z(n7790) );
  BUFFD0 U7784 ( .I(n7792), .Z(n7791) );
  BUFFD0 U7785 ( .I(n7793), .Z(n7792) );
  BUFFD0 U7786 ( .I(n7794), .Z(n7793) );
  BUFFD0 U7787 ( .I(n7795), .Z(n7794) );
  BUFFD0 U7788 ( .I(n7796), .Z(n7795) );
  BUFFD0 U7789 ( .I(n7797), .Z(n7796) );
  BUFFD0 U7790 ( .I(n7798), .Z(n7797) );
  BUFFD0 U7791 ( .I(n7799), .Z(n7798) );
  BUFFD0 U7792 ( .I(n7800), .Z(n7799) );
  BUFFD0 U7793 ( .I(n7801), .Z(n7800) );
  BUFFD0 U7794 ( .I(n7802), .Z(n7801) );
  BUFFD0 U7795 ( .I(n7803), .Z(n7802) );
  BUFFD0 U7796 ( .I(n7804), .Z(n7803) );
  BUFFD0 U7797 ( .I(n7805), .Z(n7804) );
  BUFFD0 U7798 ( .I(n7806), .Z(n7805) );
  BUFFD0 U7799 ( .I(n7807), .Z(n7806) );
  BUFFD0 U7800 ( .I(n7808), .Z(n7807) );
  BUFFD0 U7801 ( .I(n7809), .Z(n7808) );
  BUFFD0 U7802 ( .I(n7810), .Z(n7809) );
  BUFFD0 U7803 ( .I(n7811), .Z(n7810) );
  BUFFD0 U7804 ( .I(n7812), .Z(n7811) );
  BUFFD0 U7805 ( .I(n7813), .Z(n7812) );
  BUFFD0 U7806 ( .I(n7814), .Z(n7813) );
  BUFFD0 U7807 ( .I(n7815), .Z(n7814) );
  BUFFD0 U7808 ( .I(n7816), .Z(n7815) );
  BUFFD0 U7809 ( .I(n7817), .Z(n7816) );
  BUFFD0 U7810 ( .I(n7818), .Z(n7817) );
  BUFFD0 U7811 ( .I(n7819), .Z(n7818) );
  BUFFD0 U7812 ( .I(n7820), .Z(n7819) );
  BUFFD0 U7813 ( .I(n7821), .Z(n7820) );
  BUFFD0 U7814 ( .I(n7822), .Z(n7821) );
  BUFFD0 U7815 ( .I(n7823), .Z(n7822) );
  BUFFD0 U7816 ( .I(n8748), .Z(n7823) );
  BUFFD0 U7817 ( .I(n7825), .Z(n7824) );
  BUFFD0 U7818 ( .I(n7826), .Z(n7825) );
  BUFFD0 U7819 ( .I(n8681), .Z(n7826) );
  CKAN2D0 U7820 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U7821 ( .I(N48), .ZN(n8289) );
  INVD1 U7822 ( .I(DataI[17]), .ZN(n8727) );
  INVD1 U7823 ( .I(DataI[21]), .ZN(n8736) );
  INVD1 U7824 ( .I(DataI[22]), .ZN(n8738) );
  INVD1 U7825 ( .I(DataI[24]), .ZN(n8744) );
  INVD1 U7826 ( .I(DataI[25]), .ZN(n8746) );
  INVD1 U7827 ( .I(DataI[26]), .ZN(n8748) );
  INVD1 U7828 ( .I(DataI[27]), .ZN(n8751) );
  INVD1 U7829 ( .I(DataI[28]), .ZN(n8754) );
  INVD1 U7830 ( .I(DataI[29]), .ZN(n8756) );
  INVD1 U7831 ( .I(DataI[30]), .ZN(n8758) );
  INVD1 U7832 ( .I(DataI[31]), .ZN(n8761) );
  INVD1 U7833 ( .I(DataI[0]), .ZN(n8688) );
  INVD1 U7834 ( .I(DataI[1]), .ZN(n8690) );
  INVD1 U7835 ( .I(DataI[3]), .ZN(n8695) );
  INVD1 U7836 ( .I(DataI[4]), .ZN(n8697) );
  INVD1 U7837 ( .I(DataI[5]), .ZN(n8699) );
  INVD1 U7838 ( .I(DataI[6]), .ZN(n8702) );
  INVD1 U7839 ( .I(DataI[7]), .ZN(n8704) );
  INVD1 U7840 ( .I(DataI[8]), .ZN(n8706) );
  INVD1 U7841 ( .I(DataI[9]), .ZN(n8709) );
  INVD1 U7842 ( .I(DataI[10]), .ZN(n8711) );
  INVD1 U7843 ( .I(DataI[11]), .ZN(n8713) );
  INVD1 U7844 ( .I(DataI[12]), .ZN(n8715) );
  INVD1 U7845 ( .I(DataI[13]), .ZN(n8718) );
  INVD1 U7846 ( .I(DataI[14]), .ZN(n8720) );
  INVD1 U7847 ( .I(DataI[15]), .ZN(n8722) );
  INVD1 U7848 ( .I(DataI[16]), .ZN(n8725) );
  INVD1 U7849 ( .I(DataI[18]), .ZN(n8729) );
  INVD1 U7850 ( .I(DataI[19]), .ZN(n8731) );
  INVD1 U7851 ( .I(DataI[20]), .ZN(n8734) );
  INVD1 U7852 ( .I(DataI[23]), .ZN(n8741) );
  BUFFD1 U7853 ( .I(n8447), .Z(n8358) );
  BUFFD1 U7854 ( .I(n8447), .Z(n8359) );
  BUFFD1 U7855 ( .I(n8447), .Z(n8360) );
  BUFFD1 U7856 ( .I(n8447), .Z(n8361) );
  BUFFD1 U7857 ( .I(n8446), .Z(n8362) );
  BUFFD1 U7858 ( .I(n8446), .Z(n8363) );
  BUFFD1 U7859 ( .I(n8446), .Z(n8364) );
  BUFFD1 U7860 ( .I(n8446), .Z(n8365) );
  BUFFD1 U7861 ( .I(n8445), .Z(n8366) );
  BUFFD1 U7862 ( .I(n8445), .Z(n8367) );
  BUFFD1 U7863 ( .I(n8445), .Z(n8368) );
  BUFFD1 U7864 ( .I(n8445), .Z(n8369) );
  BUFFD1 U7865 ( .I(n8444), .Z(n8370) );
  BUFFD1 U7866 ( .I(n8444), .Z(n8371) );
  BUFFD1 U7867 ( .I(n8444), .Z(n8372) );
  BUFFD1 U7868 ( .I(n8444), .Z(n8373) );
  BUFFD1 U7869 ( .I(n8443), .Z(n8374) );
  BUFFD1 U7870 ( .I(n8443), .Z(n8375) );
  BUFFD1 U7871 ( .I(n8443), .Z(n8376) );
  BUFFD1 U7872 ( .I(n8443), .Z(n8377) );
  BUFFD1 U7873 ( .I(n8442), .Z(n8378) );
  BUFFD1 U7874 ( .I(n8442), .Z(n8379) );
  BUFFD1 U7875 ( .I(n8442), .Z(n8380) );
  BUFFD1 U7876 ( .I(n8442), .Z(n8381) );
  BUFFD1 U7877 ( .I(n8441), .Z(n8382) );
  BUFFD1 U7878 ( .I(n8441), .Z(n8383) );
  BUFFD1 U7879 ( .I(n8441), .Z(n8384) );
  BUFFD1 U7880 ( .I(n8441), .Z(n8385) );
  BUFFD1 U7881 ( .I(n8440), .Z(n8386) );
  BUFFD1 U7882 ( .I(n8440), .Z(n8387) );
  BUFFD1 U7883 ( .I(n8440), .Z(n8388) );
  BUFFD1 U7884 ( .I(n8440), .Z(n8389) );
  BUFFD1 U7885 ( .I(n8439), .Z(n8390) );
  BUFFD1 U7886 ( .I(n8439), .Z(n8391) );
  BUFFD1 U7887 ( .I(n8439), .Z(n8392) );
  BUFFD1 U7888 ( .I(n8439), .Z(n8393) );
  BUFFD1 U7889 ( .I(n8438), .Z(n8394) );
  BUFFD1 U7890 ( .I(n8438), .Z(n8395) );
  BUFFD1 U7891 ( .I(n8438), .Z(n8396) );
  BUFFD1 U7892 ( .I(n8438), .Z(n8397) );
  BUFFD1 U7893 ( .I(n8437), .Z(n8398) );
  BUFFD1 U7894 ( .I(n8437), .Z(n8399) );
  BUFFD1 U7895 ( .I(n8437), .Z(n8400) );
  BUFFD1 U7896 ( .I(n8437), .Z(n8401) );
  BUFFD1 U7897 ( .I(n8436), .Z(n8402) );
  BUFFD1 U7898 ( .I(n8436), .Z(n8403) );
  BUFFD1 U7899 ( .I(n8436), .Z(n8404) );
  BUFFD1 U7900 ( .I(n8436), .Z(n8405) );
  BUFFD1 U7901 ( .I(n8435), .Z(n8406) );
  BUFFD1 U7902 ( .I(n8435), .Z(n8407) );
  BUFFD1 U7903 ( .I(n8435), .Z(n8408) );
  BUFFD1 U7904 ( .I(n8435), .Z(n8409) );
  BUFFD1 U7905 ( .I(n8434), .Z(n8410) );
  BUFFD1 U7906 ( .I(n8434), .Z(n8411) );
  BUFFD1 U7907 ( .I(n8434), .Z(n8412) );
  BUFFD1 U7908 ( .I(n8434), .Z(n8413) );
  BUFFD1 U7909 ( .I(n8433), .Z(n8414) );
  BUFFD1 U7910 ( .I(n8433), .Z(n8415) );
  BUFFD1 U7911 ( .I(n8433), .Z(n8416) );
  BUFFD1 U7912 ( .I(n8433), .Z(n8417) );
  BUFFD1 U7913 ( .I(n8432), .Z(n8418) );
  BUFFD1 U7914 ( .I(n8432), .Z(n8419) );
  BUFFD1 U7915 ( .I(n8432), .Z(n8420) );
  BUFFD1 U7916 ( .I(n8432), .Z(n8421) );
  BUFFD1 U7917 ( .I(n8431), .Z(n8422) );
  BUFFD1 U7918 ( .I(n8431), .Z(n8423) );
  BUFFD1 U7919 ( .I(n8431), .Z(n8424) );
  BUFFD1 U7920 ( .I(n8431), .Z(n8425) );
  BUFFD1 U7921 ( .I(n8430), .Z(n8426) );
  BUFFD1 U7922 ( .I(n8430), .Z(n8427) );
  BUFFD1 U7923 ( .I(n8430), .Z(n8428) );
  BUFFD1 U7924 ( .I(n8430), .Z(n8429) );
  BUFFD1 U7925 ( .I(n8452), .Z(n8334) );
  BUFFD1 U7926 ( .I(n8452), .Z(n8335) );
  BUFFD1 U7927 ( .I(n8452), .Z(n8336) );
  BUFFD1 U7928 ( .I(n8452), .Z(n8337) );
  BUFFD1 U7929 ( .I(n8451), .Z(n8338) );
  BUFFD1 U7930 ( .I(n8451), .Z(n8339) );
  BUFFD1 U7931 ( .I(n8451), .Z(n8340) );
  BUFFD1 U7932 ( .I(n8451), .Z(n8341) );
  BUFFD1 U7933 ( .I(n8450), .Z(n8342) );
  BUFFD1 U7934 ( .I(n8450), .Z(n8343) );
  BUFFD1 U7935 ( .I(n8450), .Z(n8344) );
  BUFFD1 U7936 ( .I(n8450), .Z(n8345) );
  BUFFD1 U7937 ( .I(n8450), .Z(n8346) );
  BUFFD1 U7938 ( .I(n8450), .Z(n8347) );
  BUFFD1 U7939 ( .I(n8450), .Z(n8348) );
  BUFFD1 U7940 ( .I(n8450), .Z(n8349) );
  BUFFD1 U7941 ( .I(n8449), .Z(n8350) );
  BUFFD1 U7942 ( .I(n8449), .Z(n8351) );
  BUFFD1 U7943 ( .I(n8449), .Z(n8352) );
  BUFFD1 U7944 ( .I(n8449), .Z(n8353) );
  BUFFD1 U7945 ( .I(n8448), .Z(n8354) );
  BUFFD1 U7946 ( .I(n8448), .Z(n8355) );
  BUFFD1 U7947 ( .I(n8448), .Z(n8356) );
  BUFFD1 U7948 ( .I(n8448), .Z(n8357) );
  BUFFD1 U7949 ( .I(n8455), .Z(n8447) );
  BUFFD1 U7950 ( .I(n8455), .Z(n8446) );
  BUFFD1 U7951 ( .I(n8456), .Z(n8445) );
  BUFFD1 U7952 ( .I(n8456), .Z(n8444) );
  BUFFD1 U7953 ( .I(n8457), .Z(n8443) );
  BUFFD1 U7954 ( .I(n8457), .Z(n8442) );
  BUFFD1 U7955 ( .I(n8458), .Z(n8441) );
  BUFFD1 U7956 ( .I(n8458), .Z(n8440) );
  BUFFD1 U7957 ( .I(n8459), .Z(n8439) );
  BUFFD1 U7958 ( .I(n8459), .Z(n8438) );
  BUFFD1 U7959 ( .I(n8460), .Z(n8437) );
  BUFFD1 U7960 ( .I(n8460), .Z(n8436) );
  BUFFD1 U7961 ( .I(n8461), .Z(n8435) );
  BUFFD1 U7962 ( .I(n8461), .Z(n8434) );
  BUFFD1 U7963 ( .I(n8461), .Z(n8433) );
  BUFFD1 U7964 ( .I(n8462), .Z(n8432) );
  BUFFD1 U7965 ( .I(n8462), .Z(n8431) );
  BUFFD1 U7966 ( .I(n8462), .Z(n8430) );
  BUFFD1 U7967 ( .I(n8317), .Z(n8319) );
  BUFFD1 U7968 ( .I(n8314), .Z(n8321) );
  BUFFD1 U7969 ( .I(n8317), .Z(n8320) );
  BUFFD1 U7970 ( .I(n8321), .Z(n8322) );
  BUFFD1 U7971 ( .I(n8315), .Z(n8323) );
  BUFFD1 U7972 ( .I(n8316), .Z(n8324) );
  BUFFD1 U7973 ( .I(n8316), .Z(n8325) );
  BUFFD1 U7974 ( .I(n8316), .Z(n8326) );
  BUFFD1 U7975 ( .I(n8315), .Z(n8327) );
  BUFFD1 U7976 ( .I(n8315), .Z(n8328) );
  BUFFD1 U7977 ( .I(n8301), .Z(n8313) );
  BUFFD1 U7978 ( .I(n8301), .Z(n8312) );
  BUFFD1 U7979 ( .I(n8301), .Z(n8311) );
  BUFFD1 U7980 ( .I(n8303), .Z(n8305) );
  BUFFD1 U7981 ( .I(n8303), .Z(n8306) );
  BUFFD1 U7982 ( .I(n8302), .Z(n8309) );
  BUFFD1 U7983 ( .I(n8303), .Z(n8307) );
  BUFFD1 U7984 ( .I(n8302), .Z(n8310) );
  BUFFD1 U7985 ( .I(n8302), .Z(n8308) );
  BUFFD1 U7986 ( .I(n8317), .Z(n8318) );
  BUFFD1 U7987 ( .I(n8622), .Z(n8620) );
  BUFFD1 U7988 ( .I(n8623), .Z(n8619) );
  BUFFD1 U7989 ( .I(n8623), .Z(n8618) );
  BUFFD1 U7990 ( .I(n8636), .Z(n8617) );
  BUFFD1 U7991 ( .I(n8529), .Z(n8616) );
  BUFFD1 U7992 ( .I(n8624), .Z(n8615) );
  BUFFD1 U7993 ( .I(n8624), .Z(n8614) );
  BUFFD1 U7994 ( .I(n8625), .Z(n8613) );
  BUFFD1 U7995 ( .I(n8625), .Z(n8612) );
  BUFFD1 U7996 ( .I(n8626), .Z(n8611) );
  BUFFD1 U7997 ( .I(n8626), .Z(n8610) );
  BUFFD1 U7998 ( .I(n8627), .Z(n8609) );
  BUFFD1 U7999 ( .I(n8627), .Z(n8608) );
  BUFFD1 U8000 ( .I(n8628), .Z(n8607) );
  BUFFD1 U8001 ( .I(n8628), .Z(n8606) );
  BUFFD1 U8002 ( .I(n8629), .Z(n8605) );
  BUFFD1 U8003 ( .I(n8629), .Z(n8604) );
  BUFFD1 U8004 ( .I(n8677), .Z(n8603) );
  BUFFD1 U8005 ( .I(n8630), .Z(n8602) );
  BUFFD1 U8006 ( .I(n8630), .Z(n8601) );
  BUFFD1 U8007 ( .I(n8631), .Z(n8600) );
  BUFFD1 U8008 ( .I(n8631), .Z(n8599) );
  BUFFD1 U8009 ( .I(n8632), .Z(n8598) );
  BUFFD1 U8010 ( .I(n8632), .Z(n8597) );
  BUFFD1 U8011 ( .I(n8633), .Z(n8596) );
  BUFFD1 U8012 ( .I(n8633), .Z(n8595) );
  BUFFD1 U8013 ( .I(n8634), .Z(n8594) );
  BUFFD1 U8014 ( .I(n8634), .Z(n8593) );
  BUFFD1 U8015 ( .I(n8635), .Z(n8592) );
  BUFFD1 U8016 ( .I(n8635), .Z(n8591) );
  BUFFD1 U8017 ( .I(n8636), .Z(n8590) );
  BUFFD1 U8018 ( .I(n8636), .Z(n8589) );
  BUFFD1 U8019 ( .I(n8637), .Z(n8588) );
  BUFFD1 U8020 ( .I(n8637), .Z(n8587) );
  BUFFD1 U8021 ( .I(n8638), .Z(n8586) );
  BUFFD1 U8022 ( .I(n8638), .Z(n8585) );
  BUFFD1 U8023 ( .I(n8639), .Z(n8584) );
  BUFFD1 U8024 ( .I(n8639), .Z(n8583) );
  BUFFD1 U8025 ( .I(n8640), .Z(n8582) );
  BUFFD1 U8026 ( .I(n8670), .Z(n8581) );
  BUFFD1 U8027 ( .I(n8675), .Z(n8580) );
  BUFFD1 U8028 ( .I(n8641), .Z(n8579) );
  BUFFD1 U8029 ( .I(n8641), .Z(n8578) );
  BUFFD1 U8030 ( .I(n8642), .Z(n8577) );
  BUFFD1 U8031 ( .I(n8642), .Z(n8576) );
  BUFFD1 U8032 ( .I(n8643), .Z(n8575) );
  BUFFD1 U8033 ( .I(n8643), .Z(n8574) );
  BUFFD1 U8034 ( .I(n8644), .Z(n8573) );
  BUFFD1 U8035 ( .I(n8644), .Z(n8572) );
  BUFFD1 U8036 ( .I(n8645), .Z(n8571) );
  BUFFD1 U8037 ( .I(n8645), .Z(n8570) );
  BUFFD1 U8038 ( .I(n8646), .Z(n8569) );
  BUFFD1 U8039 ( .I(n8646), .Z(n8568) );
  BUFFD1 U8040 ( .I(n8647), .Z(n8567) );
  BUFFD1 U8041 ( .I(n8647), .Z(n8566) );
  BUFFD1 U8042 ( .I(n8648), .Z(n8565) );
  BUFFD1 U8043 ( .I(n8648), .Z(n8564) );
  BUFFD1 U8044 ( .I(n8649), .Z(n8563) );
  BUFFD1 U8045 ( .I(n8649), .Z(n8562) );
  BUFFD1 U8046 ( .I(n8650), .Z(n8561) );
  BUFFD1 U8047 ( .I(n8650), .Z(n8560) );
  BUFFD1 U8048 ( .I(n8651), .Z(n8559) );
  BUFFD1 U8049 ( .I(n8651), .Z(n8558) );
  BUFFD1 U8050 ( .I(n8652), .Z(n8557) );
  BUFFD1 U8051 ( .I(n8652), .Z(n8556) );
  BUFFD1 U8052 ( .I(n8653), .Z(n8555) );
  BUFFD1 U8053 ( .I(n8653), .Z(n8554) );
  BUFFD1 U8054 ( .I(n8654), .Z(n8553) );
  BUFFD1 U8055 ( .I(n8654), .Z(n8552) );
  BUFFD1 U8056 ( .I(n8655), .Z(n8551) );
  BUFFD1 U8057 ( .I(n8655), .Z(n8550) );
  BUFFD1 U8058 ( .I(n8656), .Z(n8549) );
  BUFFD1 U8059 ( .I(n8656), .Z(n8548) );
  BUFFD1 U8060 ( .I(n8657), .Z(n8547) );
  BUFFD1 U8061 ( .I(n8657), .Z(n8546) );
  BUFFD1 U8062 ( .I(n8658), .Z(n8545) );
  BUFFD1 U8063 ( .I(n8658), .Z(n8544) );
  BUFFD1 U8064 ( .I(n8659), .Z(n8543) );
  BUFFD1 U8065 ( .I(n8659), .Z(n8542) );
  BUFFD1 U8066 ( .I(n8660), .Z(n8541) );
  BUFFD1 U8067 ( .I(n8660), .Z(n8540) );
  BUFFD1 U8068 ( .I(n8661), .Z(n8539) );
  BUFFD1 U8069 ( .I(n8661), .Z(n8538) );
  BUFFD1 U8070 ( .I(n8662), .Z(n8537) );
  BUFFD1 U8071 ( .I(n8662), .Z(n8536) );
  BUFFD1 U8072 ( .I(n8622), .Z(n8621) );
  BUFFD1 U8073 ( .I(n8453), .Z(n8451) );
  BUFFD1 U8074 ( .I(n8333), .Z(n8450) );
  BUFFD1 U8075 ( .I(n8454), .Z(n8449) );
  BUFFD1 U8076 ( .I(n8454), .Z(n8448) );
  BUFFD1 U8077 ( .I(n8453), .Z(n8452) );
  BUFFD1 U8078 ( .I(n8329), .Z(n8455) );
  BUFFD1 U8079 ( .I(n8329), .Z(n8456) );
  BUFFD1 U8080 ( .I(n8329), .Z(n8457) );
  BUFFD1 U8081 ( .I(n8330), .Z(n8458) );
  BUFFD1 U8082 ( .I(n8330), .Z(n8459) );
  BUFFD1 U8083 ( .I(n8330), .Z(n8460) );
  BUFFD1 U8084 ( .I(n8331), .Z(n8461) );
  BUFFD1 U8085 ( .I(n8331), .Z(n8462) );
  BUFFD1 U8086 ( .I(N44), .Z(n8317) );
  BUFFD1 U8087 ( .I(n8686), .Z(n8293) );
  BUFFD1 U8088 ( .I(n8686), .Z(n8292) );
  BUFFD1 U8089 ( .I(n8300), .Z(n8303) );
  BUFFD1 U8090 ( .I(n8300), .Z(n8302) );
  BUFFD1 U8091 ( .I(n8314), .Z(n8316) );
  BUFFD1 U8092 ( .I(n8300), .Z(n8301) );
  BUFFD1 U8093 ( .I(n8314), .Z(n8315) );
  BUFFD1 U8094 ( .I(n8300), .Z(n8304) );
  BUFFD1 U8095 ( .I(n8676), .Z(n8624) );
  BUFFD1 U8096 ( .I(n8676), .Z(n8625) );
  BUFFD1 U8097 ( .I(n8676), .Z(n8626) );
  BUFFD1 U8098 ( .I(n8675), .Z(n8627) );
  BUFFD1 U8099 ( .I(n8675), .Z(n8628) );
  BUFFD1 U8100 ( .I(n8675), .Z(n8629) );
  BUFFD1 U8101 ( .I(n8674), .Z(n8630) );
  BUFFD1 U8102 ( .I(n8674), .Z(n8631) );
  BUFFD1 U8103 ( .I(n8674), .Z(n8632) );
  BUFFD1 U8104 ( .I(n8672), .Z(n8633) );
  BUFFD1 U8105 ( .I(n8672), .Z(n8634) );
  BUFFD1 U8106 ( .I(n8672), .Z(n8635) );
  BUFFD1 U8107 ( .I(n8671), .Z(n8636) );
  BUFFD1 U8108 ( .I(n8671), .Z(n8637) );
  BUFFD1 U8109 ( .I(n8671), .Z(n8638) );
  BUFFD1 U8110 ( .I(n8670), .Z(n8639) );
  BUFFD1 U8111 ( .I(n8670), .Z(n8640) );
  BUFFD1 U8112 ( .I(n8671), .Z(n8641) );
  BUFFD1 U8113 ( .I(n8669), .Z(n8642) );
  BUFFD1 U8114 ( .I(n8669), .Z(n8643) );
  BUFFD1 U8115 ( .I(n8669), .Z(n8644) );
  BUFFD1 U8116 ( .I(n8668), .Z(n8645) );
  BUFFD1 U8117 ( .I(n8668), .Z(n8646) );
  BUFFD1 U8118 ( .I(n8668), .Z(n8647) );
  BUFFD1 U8119 ( .I(n8667), .Z(n8648) );
  BUFFD1 U8120 ( .I(n8667), .Z(n8649) );
  BUFFD1 U8121 ( .I(n8667), .Z(n8650) );
  BUFFD1 U8122 ( .I(n8666), .Z(n8651) );
  BUFFD1 U8123 ( .I(n8666), .Z(n8652) );
  BUFFD1 U8124 ( .I(n8666), .Z(n8653) );
  BUFFD1 U8125 ( .I(n8665), .Z(n8654) );
  BUFFD1 U8126 ( .I(n8665), .Z(n8655) );
  BUFFD1 U8127 ( .I(n8665), .Z(n8656) );
  BUFFD1 U8128 ( .I(n8664), .Z(n8657) );
  BUFFD1 U8129 ( .I(n8664), .Z(n8658) );
  BUFFD1 U8130 ( .I(n8664), .Z(n8659) );
  BUFFD1 U8131 ( .I(n8663), .Z(n8660) );
  BUFFD1 U8132 ( .I(n8663), .Z(n8661) );
  BUFFD1 U8133 ( .I(n8663), .Z(n8662) );
  BUFFD1 U8134 ( .I(n8677), .Z(n8622) );
  BUFFD1 U8135 ( .I(n8677), .Z(n8623) );
  BUFFD1 U8136 ( .I(n8333), .Z(n8454) );
  BUFFD1 U8137 ( .I(n8333), .Z(n8453) );
  BUFFD1 U8138 ( .I(n8332), .Z(n8329) );
  BUFFD1 U8139 ( .I(n8332), .Z(n8330) );
  INVD1 U8140 ( .I(N85), .ZN(n8528) );
  BUFFD1 U8141 ( .I(n8294), .Z(n8299) );
  BUFFD1 U8142 ( .I(n8295), .Z(n8297) );
  BUFFD1 U8143 ( .I(n8295), .Z(n8298) );
  BUFFD1 U8144 ( .I(N44), .Z(n8314) );
  BUFFD1 U8145 ( .I(N45), .Z(n8300) );
  BUFFD1 U8146 ( .I(n8295), .Z(n8296) );
  BUFFD1 U8147 ( .I(n8664), .Z(n8676) );
  BUFFD1 U8148 ( .I(n8529), .Z(n8675) );
  BUFFD1 U8149 ( .I(n8640), .Z(n8674) );
  BUFFD1 U8150 ( .I(n8533), .Z(n8673) );
  BUFFD1 U8151 ( .I(n8533), .Z(n8672) );
  BUFFD1 U8152 ( .I(n8532), .Z(n8671) );
  BUFFD1 U8153 ( .I(n8532), .Z(n8670) );
  BUFFD1 U8154 ( .I(n8636), .Z(n8669) );
  BUFFD1 U8155 ( .I(n8531), .Z(n8668) );
  BUFFD1 U8156 ( .I(n8531), .Z(n8667) );
  BUFFD1 U8157 ( .I(n8530), .Z(n8666) );
  BUFFD1 U8158 ( .I(n8530), .Z(n8665) );
  BUFFD1 U8159 ( .I(n8529), .Z(n8664) );
  BUFFD1 U8160 ( .I(n8529), .Z(n8663) );
  BUFFD1 U8161 ( .I(ClockW), .Z(n8677) );
  BUFFD1 U8162 ( .I(n108), .Z(n8332) );
  BUFFD1 U8163 ( .I(n108), .Z(n8331) );
  BUFFD1 U8164 ( .I(n108), .Z(n8333) );
  XOR3D1 U8165 ( .A1(n80), .A2(n8710), .A3(n81), .Z(n79) );
  XOR3D1 U8166 ( .A1(n8730), .A2(n8728), .A3(n82), .Z(n81) );
  XOR3D1 U8167 ( .A1(n83), .A2(n8726), .A3(n84), .Z(n82) );
  XOR3D1 U8168 ( .A1(n8698), .A2(n8696), .A3(n76), .Z(n75) );
  XOR3D1 U8169 ( .A1(n77), .A2(n8694), .A3(n78), .Z(n76) );
  XOR3D1 U8170 ( .A1(n8714), .A2(n8712), .A3(n79), .Z(n78) );
  XOR3D1 U8171 ( .A1(n8687), .A2(n74), .A3(n75), .Z(n73) );
  XOR3D1 U8172 ( .A1(n2090), .A2(n2083), .A3(n92), .Z(n90) );
  XOR3D1 U8173 ( .A1(N65), .A2(n93), .A3(n94), .Z(n92) );
  XOR3D1 U8174 ( .A1(N60), .A2(N59), .A3(n95), .Z(n94) );
  XOR3D1 U8175 ( .A1(n96), .A2(N58), .A3(n97), .Z(n95) );
  XOR3D1 U8176 ( .A1(n2091), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D1 U8177 ( .A1(n2084), .A2(n2098), .A3(n89), .Z(n88) );
  BUFFD1 U8178 ( .I(n8685), .Z(n8295) );
  BUFFD1 U8179 ( .I(n8685), .Z(n8294) );
  INVD1 U8180 ( .I(n8289), .ZN(n8290) );
  INVD1 U8181 ( .I(n8289), .ZN(n8291) );
  BUFFD1 U8182 ( .I(N47), .Z(n8686) );
  INVD1 U8183 ( .I(n7836), .ZN(n8488) );
  INVD1 U8184 ( .I(n7836), .ZN(n8487) );
  INVD1 U8185 ( .I(n7837), .ZN(n8486) );
  INVD1 U8186 ( .I(n7837), .ZN(n8485) );
  INVD1 U8187 ( .I(n7838), .ZN(n8484) );
  INVD1 U8188 ( .I(n7838), .ZN(n8483) );
  INVD1 U8189 ( .I(n7839), .ZN(n8482) );
  INVD1 U8190 ( .I(n7839), .ZN(n8481) );
  INVD1 U8191 ( .I(n7840), .ZN(n8480) );
  INVD1 U8192 ( .I(n7840), .ZN(n8479) );
  INVD1 U8193 ( .I(n7841), .ZN(n8478) );
  INVD1 U8194 ( .I(n7841), .ZN(n8477) );
  INVD1 U8195 ( .I(n7842), .ZN(n8476) );
  INVD1 U8196 ( .I(n7842), .ZN(n8475) );
  INVD1 U8197 ( .I(n7843), .ZN(n8474) );
  INVD1 U8198 ( .I(n7843), .ZN(n8473) );
  INVD1 U8199 ( .I(n7844), .ZN(n8472) );
  INVD1 U8200 ( .I(n7844), .ZN(n8471) );
  INVD1 U8201 ( .I(n7845), .ZN(n8470) );
  INVD1 U8202 ( .I(n7845), .ZN(n8469) );
  INVD1 U8203 ( .I(n7846), .ZN(n8468) );
  INVD1 U8204 ( .I(n7846), .ZN(n8467) );
  INVD1 U8205 ( .I(n7847), .ZN(n8466) );
  INVD1 U8206 ( .I(n7847), .ZN(n8465) );
  INVD1 U8207 ( .I(n7848), .ZN(n8464) );
  INVD1 U8208 ( .I(n7848), .ZN(n8463) );
  INVD1 U8209 ( .I(n7849), .ZN(n8526) );
  INVD1 U8210 ( .I(n7849), .ZN(n8525) );
  INVD1 U8211 ( .I(n7850), .ZN(n8524) );
  INVD1 U8212 ( .I(n7850), .ZN(n8523) );
  INVD1 U8213 ( .I(n7851), .ZN(n8522) );
  INVD1 U8214 ( .I(n7851), .ZN(n8521) );
  INVD1 U8215 ( .I(n7852), .ZN(n8520) );
  INVD1 U8216 ( .I(n7852), .ZN(n8519) );
  INVD1 U8217 ( .I(n7853), .ZN(n8518) );
  INVD1 U8218 ( .I(n7853), .ZN(n8517) );
  INVD1 U8219 ( .I(n7854), .ZN(n8516) );
  INVD1 U8220 ( .I(n7854), .ZN(n8515) );
  INVD1 U8221 ( .I(n7855), .ZN(n8514) );
  INVD1 U8222 ( .I(n7855), .ZN(n8513) );
  INVD1 U8223 ( .I(n7856), .ZN(n8512) );
  INVD1 U8224 ( .I(n7856), .ZN(n8511) );
  INVD1 U8225 ( .I(n7828), .ZN(n8510) );
  INVD1 U8226 ( .I(n7828), .ZN(n8509) );
  INVD1 U8227 ( .I(n7829), .ZN(n8508) );
  INVD1 U8228 ( .I(n7829), .ZN(n8507) );
  INVD1 U8229 ( .I(n7830), .ZN(n8506) );
  INVD1 U8230 ( .I(n7830), .ZN(n8505) );
  INVD1 U8231 ( .I(n7831), .ZN(n8504) );
  INVD1 U8232 ( .I(n7831), .ZN(n8503) );
  INVD1 U8233 ( .I(n7832), .ZN(n8502) );
  INVD1 U8234 ( .I(n7832), .ZN(n8501) );
  INVD1 U8235 ( .I(n7833), .ZN(n8500) );
  INVD1 U8236 ( .I(n7833), .ZN(n8499) );
  INVD1 U8237 ( .I(n7834), .ZN(n8498) );
  INVD1 U8238 ( .I(n7834), .ZN(n8497) );
  INVD1 U8239 ( .I(n7835), .ZN(n8496) );
  INVD1 U8240 ( .I(n7835), .ZN(n8495) );
  INVD1 U8241 ( .I(n7857), .ZN(n8494) );
  INVD1 U8242 ( .I(n7857), .ZN(n8493) );
  INVD1 U8243 ( .I(n7858), .ZN(n8492) );
  INVD1 U8244 ( .I(n7858), .ZN(n8491) );
  INVD1 U8245 ( .I(n7859), .ZN(n8490) );
  INVD1 U8246 ( .I(n7859), .ZN(n8489) );
  BUFFD1 U8247 ( .I(n8680), .Z(n8683) );
  BUFFD1 U8248 ( .I(n8680), .Z(n8682) );
  BUFFD1 U8249 ( .I(n8681), .Z(n8684) );
  BUFFD1 U8250 ( .I(n8534), .Z(n8533) );
  BUFFD1 U8251 ( .I(n8534), .Z(n8532) );
  BUFFD1 U8252 ( .I(n8535), .Z(n8531) );
  BUFFD1 U8253 ( .I(n8535), .Z(n8530) );
  BUFFD1 U8254 ( .I(n8535), .Z(n8529) );
  INVD1 U8255 ( .I(n8679), .ZN(n8678) );
  INVD1 U8256 ( .I(Reset), .ZN(n108) );
  INVD1 U8257 ( .I(n7113), .ZN(n8687) );
  INVD1 U8258 ( .I(n6224), .ZN(n8698) );
  INVD1 U8259 ( .I(n4980), .ZN(n8714) );
  INVD1 U8260 ( .I(n3738), .ZN(n8730) );
  INVD1 U8261 ( .I(n5869), .ZN(n8703) );
  INVD1 U8262 ( .I(n5690), .ZN(n8705) );
  INVD1 U8263 ( .I(n4625), .ZN(n8719) );
  INVD1 U8264 ( .I(n4446), .ZN(n8721) );
  INVD1 U8265 ( .I(n3383), .ZN(n8735) );
  INVD1 U8266 ( .I(n3204), .ZN(n8737) );
  INVD1 U8267 ( .I(n7467), .ZN(n8745) );
  INVD1 U8268 ( .I(n7646), .ZN(n8747) );
  INVD1 U8269 ( .I(n2494), .ZN(n8755) );
  INVD1 U8270 ( .I(n2315), .ZN(n8757) );
  INVD1 U8271 ( .I(n6935), .ZN(n8689) );
  INVD1 U8272 ( .I(n6580), .ZN(n8694) );
  INVD1 U8273 ( .I(n6401), .ZN(n8696) );
  INVD1 U8274 ( .I(n5334), .ZN(n8710) );
  INVD1 U8275 ( .I(n5155), .ZN(n8712) );
  INVD1 U8276 ( .I(n4090), .ZN(n8726) );
  INVD1 U8277 ( .I(n3911), .ZN(n8728) );
  INVD1 U8278 ( .I(n6048), .ZN(n8700) );
  INVD1 U8279 ( .I(n5513), .ZN(n8707) );
  INVD1 U8280 ( .I(n4804), .ZN(n8716) );
  INVD1 U8281 ( .I(n4269), .ZN(n8723) );
  INVD1 U8282 ( .I(n3562), .ZN(n8732) );
  INVD1 U8283 ( .I(n3027), .ZN(n8739) );
  INVD1 U8284 ( .I(n2850), .ZN(n8742) );
  INVD1 U8285 ( .I(n7290), .ZN(n8749) );
  INVD1 U8286 ( .I(n2673), .ZN(n8752) );
  INVD1 U8287 ( .I(n2221), .ZN(n8759) );
  INVD1 U8288 ( .I(n6048), .ZN(n8701) );
  INVD1 U8289 ( .I(n5513), .ZN(n8708) );
  INVD1 U8290 ( .I(n4804), .ZN(n8717) );
  INVD1 U8291 ( .I(n4269), .ZN(n8724) );
  INVD1 U8292 ( .I(n3562), .ZN(n8733) );
  INVD1 U8293 ( .I(n3027), .ZN(n8740) );
  INVD1 U8294 ( .I(n2850), .ZN(n8743) );
  INVD1 U8295 ( .I(n7290), .ZN(n8750) );
  INVD1 U8296 ( .I(n2673), .ZN(n8753) );
  INVD1 U8297 ( .I(n2221), .ZN(n8760) );
  BUFFD1 U8298 ( .I(N46), .Z(n8685) );
  OR2D1 U8299 ( .A1(n69), .A2(n101), .Z(n7828) );
  OR2D1 U8300 ( .A1(n68), .A2(n101), .Z(n7829) );
  OR2D1 U8301 ( .A1(n67), .A2(n101), .Z(n7830) );
  OR2D1 U8302 ( .A1(n99), .A2(n101), .Z(n7831) );
  OR2D1 U8303 ( .A1(n98), .A2(n101), .Z(n7832) );
  OR2D1 U8304 ( .A1(n85), .A2(n101), .Z(n7833) );
  OR2D1 U8305 ( .A1(n72), .A2(n101), .Z(n7834) );
  OR2D1 U8306 ( .A1(n71), .A2(n101), .Z(n7835) );
  ND3D1 U8307 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U8308 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  INVD1 U8309 ( .I(AddrW[2]), .ZN(n105) );
  OR2D1 U8310 ( .A1(n70), .A2(n99), .Z(n7836) );
  OR2D1 U8311 ( .A1(n70), .A2(n98), .Z(n7837) );
  OR2D1 U8312 ( .A1(n70), .A2(n85), .Z(n7838) );
  OR2D1 U8313 ( .A1(n70), .A2(n72), .Z(n7839) );
  OR2D1 U8314 ( .A1(n70), .A2(n71), .Z(n7840) );
  OR2D1 U8315 ( .A1(n66), .A2(n69), .Z(n7841) );
  OR2D1 U8316 ( .A1(n66), .A2(n68), .Z(n7842) );
  OR2D1 U8317 ( .A1(n66), .A2(n67), .Z(n7843) );
  OR2D1 U8318 ( .A1(n66), .A2(n99), .Z(n7844) );
  OR2D1 U8319 ( .A1(n66), .A2(n98), .Z(n7845) );
  OR2D1 U8320 ( .A1(n66), .A2(n85), .Z(n7846) );
  OR2D1 U8321 ( .A1(n66), .A2(n72), .Z(n7847) );
  OR2D1 U8322 ( .A1(n66), .A2(n71), .Z(n7848) );
  OR2D1 U8323 ( .A1(n69), .A2(n103), .Z(n7849) );
  OR2D1 U8324 ( .A1(n68), .A2(n103), .Z(n7850) );
  OR2D1 U8325 ( .A1(n67), .A2(n103), .Z(n7851) );
  OR2D1 U8326 ( .A1(n99), .A2(n103), .Z(n7852) );
  OR2D1 U8327 ( .A1(n98), .A2(n103), .Z(n7853) );
  OR2D1 U8328 ( .A1(n85), .A2(n103), .Z(n7854) );
  OR2D1 U8329 ( .A1(n72), .A2(n103), .Z(n7855) );
  OR2D1 U8330 ( .A1(n71), .A2(n103), .Z(n7856) );
  OR2D1 U8331 ( .A1(n69), .A2(n70), .Z(n7857) );
  OR2D1 U8332 ( .A1(n68), .A2(n70), .Z(n7858) );
  OR2D1 U8333 ( .A1(n67), .A2(n70), .Z(n7859) );
  BUFFD1 U8334 ( .I(Read), .Z(n8680) );
  BUFFD1 U8335 ( .I(Read), .Z(n8681) );
  INVD1 U8336 ( .I(ClockR), .ZN(n8679) );
  BUFFD1 U8337 ( .I(ClockW), .Z(n8534) );
  BUFFD1 U8338 ( .I(ClockW), .Z(n8535) );
  MUX4ND0 U8339 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n8321), .S1(n8301), 
        .ZN(n8188) );
  MUX4ND0 U8340 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n8321), .S1(n8303), 
        .ZN(n8201) );
  MUX4D0 U8341 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n8315), .S1(n8302), 
        .Z(n8189) );
  MUX4D0 U8342 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n8318), .S1(N45), .Z(
        n8202) );
  MUX4D0 U8343 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n8321), .S1(n8302), 
        .Z(n8215) );
  MUX4D0 U8344 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n8315), .S1(n8302), 
        .Z(n8228) );
  MUX4D0 U8345 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n8318), .S1(n8303), .Z(
        n8193) );
  MUX4D0 U8346 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n8318), .S1(n8302), 
        .Z(n8191) );
  MUX4D0 U8347 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n8316), .S1(n8303), .Z(
        n8206) );
  MUX4D0 U8348 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n8315), .S1(n8300), 
        .Z(n8204) );
  MUX4D0 U8349 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n8315), .S1(n8303), .Z(
        n8219) );
  MUX4D0 U8350 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n8318), .S1(n8304), 
        .Z(n8217) );
  MUX4D0 U8351 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n8316), .S1(n8303), .Z(
        n8232) );
  MUX4D0 U8352 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n8314), .S1(n8302), 
        .Z(n8230) );
  MUX4D0 U8353 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n8315), .S1(n8300), .Z(
        n8258) );
  MUX4D0 U8354 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n8314), .S1(n8303), 
        .Z(n8190) );
  MUX4D0 U8355 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n8316), .S1(n8304), 
        .Z(n8203) );
  MUX4D0 U8356 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n8316), .S1(n8304), 
        .Z(n8216) );
  MUX4D0 U8357 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n8316), .S1(n8304), 
        .Z(n8229) );
  MUX4D0 U8358 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n8318), .S1(n8301), .Z(
        n8194) );
  MUX4D0 U8359 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n8316), .S1(n8304), 
        .Z(n8192) );
  MUX4D0 U8360 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n8316), .S1(n8302), .Z(
        n8207) );
  MUX4D0 U8361 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n8318), .S1(n8302), 
        .Z(n8205) );
  MUX4D0 U8362 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n8315), .S1(n8304), .Z(
        n8220) );
  MUX4D0 U8363 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n8314), .S1(n8304), 
        .Z(n8218) );
  MUX4D0 U8364 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n8315), .S1(n8302), .Z(
        n8233) );
  MUX4D0 U8365 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n8314), .S1(n8304), 
        .Z(n8231) );
  MUX4D0 U8366 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n8316), .S1(n8304), .Z(
        n8259) );
  MUX4D0 U8367 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n8318), .S1(n8304), .Z(
        n8272) );
  MUX4ND0 U8368 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(N44), .S1(n8304), .ZN(
        n8279) );
  MUX4ND0 U8369 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n8321), .S1(n8301), 
        .ZN(n8214) );
  MUX4ND0 U8370 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n8317), .S1(n8302), 
        .ZN(n8227) );
  MUX4ND0 U8371 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(N44), .S1(n8304), .ZN(
        n8240) );
  MUX4ND0 U8372 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n8315), .S1(n8304), 
        .ZN(n8253) );
  MUX4ND0 U8373 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n8314), .S1(n8304), 
        .ZN(n8266) );
  MUX4ND0 U8374 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n8321), .S1(n8310), 
        .ZN(n8032) );
  MUX4ND0 U8375 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n8321), .S1(n8301), 
        .ZN(n8045) );
  MUX4ND0 U8376 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n8321), .S1(n8306), 
        .ZN(n8058) );
  MUX4ND0 U8377 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n8321), .S1(N45), .ZN(
        n8071) );
  MUX4ND0 U8378 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n8321), .S1(N45), .ZN(
        n8084) );
  MUX4ND0 U8379 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n8321), .S1(N45), .ZN(
        n8097) );
  MUX4ND0 U8380 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n8321), .S1(n8300), 
        .ZN(n8110) );
  MUX4ND0 U8381 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n8321), .S1(n8300), 
        .ZN(n8123) );
  MUX4ND0 U8382 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n8321), .S1(n8303), 
        .ZN(n8136) );
  MUX4ND0 U8383 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n8321), .S1(N45), .ZN(
        n8149) );
  MUX4ND0 U8384 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n8321), .S1(N45), .ZN(
        n8162) );
  MUX4ND0 U8385 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n8321), .S1(n8300), 
        .ZN(n8175) );
  MUX4D0 U8386 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n8314), .S1(n8300), 
        .Z(n8280) );
  MUX4D0 U8387 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n8322), .S1(n8311), .Z(
        n7864) );
  MUX4D0 U8388 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n8323), .S1(n8308), .Z(
        n7877) );
  MUX4D0 U8389 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n8322), .S1(n8310), .Z(
        n7890) );
  MUX4D0 U8390 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n8316), .S1(n8301), .Z(
        n7903) );
  MUX4D0 U8391 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n8328), .S1(n8305), .Z(
        n7916) );
  MUX4D0 U8392 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n8323), .S1(n8305), .Z(
        n7929) );
  MUX4D0 U8393 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n8323), .S1(n8306), .Z(
        n7942) );
  MUX4D0 U8394 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n8324), .S1(n8306), .Z(
        n7955) );
  MUX4D0 U8395 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n8322), .S1(n8306), .Z(
        n7968) );
  MUX4D0 U8396 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n8317), .S1(n8307), .Z(
        n7981) );
  MUX4D0 U8397 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n8317), .S1(n8307), 
        .Z(n7994) );
  MUX4D0 U8398 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n8322), .S1(n8308), 
        .Z(n8007) );
  MUX4D0 U8399 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n8322), .S1(n8309), 
        .Z(n8020) );
  MUX4D0 U8400 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n8323), .S1(n8309), 
        .Z(n8033) );
  MUX4D0 U8401 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n8323), .S1(n8309), 
        .Z(n8046) );
  MUX4D0 U8402 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n8324), .S1(n8310), 
        .Z(n8059) );
  MUX4D0 U8403 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n8324), .S1(n8310), 
        .Z(n8072) );
  MUX4D0 U8404 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n8325), .S1(n8310), 
        .Z(n8085) );
  MUX4D0 U8405 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n8325), .S1(n8310), 
        .Z(n8098) );
  MUX4D0 U8406 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n8326), .S1(n8300), 
        .Z(n8111) );
  MUX4D0 U8407 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n8326), .S1(n8303), 
        .Z(n8124) );
  MUX4D0 U8408 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n8327), .S1(n8303), 
        .Z(n8137) );
  MUX4D0 U8409 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n8327), .S1(n8310), 
        .Z(n8150) );
  MUX4D0 U8410 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n8328), .S1(n8306), 
        .Z(n8163) );
  MUX4D0 U8411 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n8328), .S1(n8313), 
        .Z(n8176) );
  MUX4D0 U8412 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n8314), .S1(n8304), 
        .Z(n8241) );
  MUX4D0 U8413 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n8318), .S1(n8302), 
        .Z(n8254) );
  MUX4D0 U8414 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n8316), .S1(n8304), 
        .Z(n8267) );
  MUX4D0 U8415 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(N44), .S1(N45), .Z(n8284) );
  MUX4D0 U8416 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(N44), .S1(n8300), .Z(
        n8282) );
  MUX4D0 U8417 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n8324), .S1(n8301), .Z(
        n7868) );
  MUX4D0 U8418 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n8317), .S1(n8308), .Z(
        n7866) );
  MUX4D0 U8419 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n8316), .S1(n8301), .Z(
        n7879) );
  MUX4D0 U8420 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n8325), .S1(n8310), .Z(
        n7881) );
  MUX4D0 U8421 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n8318), .S1(N45), .Z(
        n7892) );
  MUX4D0 U8422 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n8325), .S1(n8306), .Z(
        n7894) );
  MUX4D0 U8423 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n8315), .S1(n8309), .Z(
        n7907) );
  MUX4D0 U8424 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n8327), .S1(N45), .Z(
        n7905) );
  MUX4D0 U8425 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n8315), .S1(n8305), .Z(
        n7920) );
  MUX4D0 U8426 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n8326), .S1(n8305), .Z(
        n7918) );
  MUX4D0 U8427 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(N44), .S1(n8305), .Z(n7933) );
  MUX4D0 U8428 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n8325), .S1(n8305), .Z(
        n7931) );
  MUX4D0 U8429 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n8328), .S1(n8306), .Z(
        n7944) );
  MUX4D0 U8430 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n8315), .S1(n8306), .Z(
        n7946) );
  MUX4D0 U8431 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n8324), .S1(n8306), .Z(
        n7957) );
  MUX4D0 U8432 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n8322), .S1(n8306), .Z(
        n7959) );
  MUX4D0 U8433 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n8324), .S1(n8307), .Z(
        n7970) );
  MUX4D0 U8434 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n8316), .S1(n8307), .Z(
        n7972) );
  MUX4D0 U8435 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n8317), .S1(n8307), .Z(
        n7985) );
  MUX4D0 U8436 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n8318), .S1(n8305), .Z(
        n7983) );
  MUX4D0 U8437 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n8327), .S1(n8308), .Z(
        n7998) );
  MUX4D0 U8438 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n8314), .S1(n8308), 
        .Z(n7996) );
  MUX4D0 U8439 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n8322), .S1(n8308), .Z(
        n8011) );
  MUX4D0 U8440 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n8322), .S1(n8308), 
        .Z(n8009) );
  MUX4D0 U8441 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n8322), .S1(n8309), 
        .Z(n8022) );
  MUX4D0 U8442 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n8322), .S1(n8309), .Z(
        n8024) );
  MUX4D0 U8443 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n8323), .S1(n8309), 
        .Z(n8035) );
  MUX4D0 U8444 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n8323), .S1(n8310), .Z(
        n8037) );
  MUX4D0 U8445 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n8323), .S1(n8309), .Z(
        n8050) );
  MUX4D0 U8446 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n8323), .S1(n8309), 
        .Z(n8048) );
  MUX4D0 U8447 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n8324), .S1(n8310), .Z(
        n8063) );
  MUX4D0 U8448 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n8324), .S1(n8310), 
        .Z(n8061) );
  MUX4D0 U8449 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n8324), .S1(n8311), .Z(
        n8076) );
  MUX4D0 U8450 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n8324), .S1(n8311), 
        .Z(n8074) );
  MUX4D0 U8451 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n8325), .S1(n8307), .Z(
        n8089) );
  MUX4D0 U8452 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n8325), .S1(n8310), 
        .Z(n8087) );
  MUX4D0 U8453 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n8325), .S1(n8310), .Z(
        n8102) );
  MUX4D0 U8454 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n8325), .S1(n8308), 
        .Z(n8100) );
  MUX4D0 U8455 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n8326), .S1(n8303), .Z(
        n8115) );
  MUX4D0 U8456 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n8326), .S1(n8307), 
        .Z(n8113) );
  MUX4D0 U8457 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n8326), .S1(n8302), 
        .Z(n8126) );
  MUX4D0 U8458 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n8326), .S1(n8303), .Z(
        n8128) );
  MUX4D0 U8459 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n8327), .S1(n8306), .Z(
        n8141) );
  MUX4D0 U8460 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n8327), .S1(n8302), 
        .Z(n8139) );
  MUX4D0 U8461 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n8327), .S1(n8309), .Z(
        n8154) );
  MUX4D0 U8462 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n8327), .S1(n8301), 
        .Z(n8152) );
  MUX4D0 U8463 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n8328), .S1(n8301), .Z(
        n8167) );
  MUX4D0 U8464 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n8328), .S1(n8301), 
        .Z(n8165) );
  MUX4D0 U8465 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n8327), .S1(n8313), .Z(
        n8180) );
  MUX4D0 U8466 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n8328), .S1(n8313), 
        .Z(n8178) );
  MUX4D0 U8467 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(N44), .S1(n8303), .Z(
        n8245) );
  MUX4D0 U8468 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(N44), .S1(N45), .Z(
        n8243) );
  MUX4D0 U8469 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(N44), .S1(n8302), .Z(
        n8256) );
  MUX4D0 U8470 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n8317), .S1(n8300), .Z(
        n8271) );
  MUX4D0 U8471 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n8316), .S1(n8301), 
        .Z(n8269) );
  MUX4D0 U8472 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n8317), .S1(n8300), 
        .Z(n8281) );
  MUX4D0 U8473 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n8328), .S1(n8310), .Z(
        n7865) );
  MUX4D0 U8474 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n8322), .S1(n8300), .Z(
        n7878) );
  MUX4D0 U8475 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n8327), .S1(n8309), .Z(
        n7891) );
  MUX4D0 U8476 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n8327), .S1(N45), .Z(
        n7904) );
  MUX4D0 U8477 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n8325), .S1(n8305), .Z(
        n7917) );
  MUX4D0 U8478 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n8318), .S1(n8305), .Z(
        n7930) );
  MUX4D0 U8479 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n8322), .S1(n8306), .Z(
        n7943) );
  MUX4D0 U8480 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n8324), .S1(n8306), .Z(
        n7956) );
  MUX4D0 U8481 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n8321), .S1(n8307), .Z(
        n7969) );
  MUX4D0 U8482 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n8314), .S1(n8307), .Z(
        n7982) );
  MUX4D0 U8483 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n8326), .S1(n8307), 
        .Z(n7995) );
  MUX4D0 U8484 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n8322), .S1(n8308), 
        .Z(n8008) );
  MUX4D0 U8485 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n8322), .S1(n8308), 
        .Z(n8021) );
  MUX4D0 U8486 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n8323), .S1(n8309), 
        .Z(n8034) );
  MUX4D0 U8487 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n8323), .S1(n8308), 
        .Z(n8047) );
  MUX4D0 U8488 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n8324), .S1(n8309), 
        .Z(n8060) );
  MUX4D0 U8489 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n8324), .S1(n8311), 
        .Z(n8073) );
  MUX4D0 U8490 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n8325), .S1(n8311), 
        .Z(n8086) );
  MUX4D0 U8491 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n8325), .S1(n8309), 
        .Z(n8099) );
  MUX4D0 U8492 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n8326), .S1(n8301), 
        .Z(n8112) );
  MUX4D0 U8493 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n8326), .S1(n8303), 
        .Z(n8125) );
  MUX4D0 U8494 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n8327), .S1(n8303), 
        .Z(n8138) );
  MUX4D0 U8495 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n8327), .S1(n8307), 
        .Z(n8151) );
  MUX4D0 U8496 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n8328), .S1(n8308), 
        .Z(n8164) );
  MUX4D0 U8497 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n8328), .S1(n8313), 
        .Z(n8177) );
  MUX4D0 U8498 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n8317), .S1(n8303), 
        .Z(n8242) );
  MUX4D0 U8499 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n8318), .S1(n8304), 
        .Z(n8255) );
  MUX4D0 U8500 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n8318), .S1(n8304), 
        .Z(n8268) );
  MUX4D0 U8501 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(N44), .S1(N45), .Z(n8285) );
  MUX4D0 U8502 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(N44), .S1(n8300), .Z(
        n8283) );
  MUX4D0 U8503 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n8324), .S1(n8307), .Z(
        n7869) );
  MUX4D0 U8504 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n8324), .S1(n8309), .Z(
        n7867) );
  MUX4D0 U8505 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n8318), .S1(n8306), .Z(
        n7880) );
  MUX4D0 U8506 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n8314), .S1(n8301), .Z(
        n7882) );
  MUX4D0 U8507 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n8316), .S1(N45), .Z(
        n7893) );
  MUX4D0 U8508 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n8317), .S1(n8308), .Z(
        n7895) );
  MUX4D0 U8509 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n8326), .S1(n8305), .Z(
        n7908) );
  MUX4D0 U8510 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n8318), .S1(n8307), .Z(
        n7906) );
  MUX4D0 U8511 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n8323), .S1(n8305), .Z(
        n7921) );
  MUX4D0 U8512 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n8318), .S1(n8305), .Z(
        n7919) );
  MUX4D0 U8513 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n8324), .S1(n8305), .Z(
        n7934) );
  MUX4D0 U8514 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n8317), .S1(n8305), .Z(
        n7932) );
  MUX4D0 U8515 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n8318), .S1(n8306), .Z(
        n7945) );
  MUX4D0 U8516 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n8316), .S1(n8306), .Z(
        n7947) );
  MUX4D0 U8517 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n8323), .S1(n8306), .Z(
        n7958) );
  MUX4D0 U8518 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n8325), .S1(n8306), .Z(
        n7960) );
  MUX4D0 U8519 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n8328), .S1(n8307), .Z(
        n7971) );
  MUX4D0 U8520 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n8323), .S1(n8307), .Z(
        n7973) );
  MUX4D0 U8521 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n8314), .S1(n8307), .Z(
        n7986) );
  MUX4D0 U8522 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n8314), .S1(n8307), .Z(
        n7984) );
  MUX4D0 U8523 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n8328), .S1(n8308), .Z(
        n7999) );
  MUX4D0 U8524 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n8315), .S1(n8308), 
        .Z(n7997) );
  MUX4D0 U8525 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n8322), .S1(n8308), .Z(
        n8012) );
  MUX4D0 U8526 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n8322), .S1(n8308), 
        .Z(n8010) );
  MUX4D0 U8527 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n8322), .S1(n8309), 
        .Z(n8023) );
  MUX4D0 U8528 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n8323), .S1(n8309), .Z(
        n8025) );
  MUX4D0 U8529 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n8323), .S1(n8310), 
        .Z(n8036) );
  MUX4D0 U8530 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n8323), .S1(n8309), .Z(
        n8038) );
  MUX4D0 U8531 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n8324), .S1(n8310), .Z(
        n8051) );
  MUX4D0 U8532 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n8323), .S1(n8310), 
        .Z(n8049) );
  MUX4D0 U8533 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n8324), .S1(n8310), .Z(
        n8064) );
  MUX4D0 U8534 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n8324), .S1(n8310), 
        .Z(n8062) );
  MUX4D0 U8535 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n8325), .S1(n8311), .Z(
        n8077) );
  MUX4D0 U8536 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n8324), .S1(n8310), 
        .Z(n8075) );
  MUX4D0 U8537 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n8325), .S1(n8305), .Z(
        n8090) );
  MUX4D0 U8538 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n8325), .S1(n8308), 
        .Z(n8088) );
  MUX4D0 U8539 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n8326), .S1(n8309), .Z(
        n8103) );
  MUX4D0 U8540 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n8325), .S1(n8306), 
        .Z(n8101) );
  MUX4D0 U8541 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n8326), .S1(n8302), .Z(
        n8116) );
  MUX4D0 U8542 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n8326), .S1(n8303), 
        .Z(n8114) );
  MUX4D0 U8543 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n8326), .S1(n8302), 
        .Z(n8127) );
  MUX4D0 U8544 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n8327), .S1(n8302), .Z(
        n8129) );
  MUX4D0 U8545 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n8327), .S1(n8307), .Z(
        n8142) );
  MUX4D0 U8546 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n8327), .S1(n8303), 
        .Z(n8140) );
  MUX4D0 U8547 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n8328), .S1(n8302), .Z(
        n8155) );
  MUX4D0 U8548 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n8327), .S1(n8301), 
        .Z(n8153) );
  MUX4D0 U8549 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n8328), .S1(n8308), .Z(
        n8168) );
  MUX4D0 U8550 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n8328), .S1(n8301), 
        .Z(n8166) );
  MUX4D0 U8551 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n8328), .S1(n8300), .Z(
        n8181) );
  MUX4D0 U8552 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n8328), .S1(n8300), 
        .Z(n8179) );
  MUX4D0 U8553 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(N44), .S1(n8304), .Z(
        n8246) );
  MUX4D0 U8554 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(N44), .S1(n8300), .Z(
        n8244) );
  MUX4D0 U8555 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n8316), .S1(n8301), 
        .Z(n8257) );
  MUX4D0 U8556 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n8317), .S1(n8300), 
        .Z(n8270) );
  MUX4ND0 U8557 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n8328), .S1(n8305), .ZN(
        n7863) );
  MUX4ND0 U8558 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n8326), .S1(n8305), .ZN(
        n7876) );
  MUX4ND0 U8559 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n8315), .S1(n8305), .ZN(
        n7889) );
  MUX4ND0 U8560 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n8326), .S1(n8307), .ZN(
        n7902) );
  MUX4ND0 U8561 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n8322), .S1(n8309), .ZN(
        n7915) );
  MUX4ND0 U8562 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n8322), .S1(n8304), .ZN(
        n7928) );
  MUX4ND0 U8563 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n8326), .S1(n8311), .ZN(
        n7941) );
  MUX4ND0 U8564 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n8322), .S1(n8307), .ZN(
        n7954) );
  MUX4ND0 U8565 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n8315), .S1(n8308), .ZN(
        n7967) );
  MUX4ND0 U8566 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n8315), .S1(n8306), .ZN(
        n7980) );
  MUX4ND0 U8567 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n8325), .S1(n8311), 
        .ZN(n7993) );
  MUX4ND0 U8568 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n8323), .S1(n8305), 
        .ZN(n8006) );
  MUX4ND0 U8569 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n8323), .S1(n8305), 
        .ZN(n8019) );
  ND3D1 U8570 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U8571 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U8572 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U8573 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U8574 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U8575 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U8576 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U8577 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  ND3D1 U8578 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U8579 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U8580 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U8581 ( .I(AddrW[1]), .ZN(n106) );
  INVD1 U8582 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U8583 ( .I(AddrW[4]), .ZN(n102) );
  CKAN2D0 U8584 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  CKAN2D0 U8585 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U8586 ( .I0(n7861), .I1(n7862), .I2(n7863), .S0(n8311), .S1(n8296), 
        .ZN(n7860) );
  MUX3ND0 U8587 ( .I0(n7870), .I1(n7871), .I2(n2198), .S0(N47), .S1(n8290), 
        .ZN(N82) );
  MUX3ND0 U8588 ( .I0(n7874), .I1(n7875), .I2(n7876), .S0(n8313), .S1(n8296), 
        .ZN(n7873) );
  MUX3ND0 U8589 ( .I0(n7883), .I1(n7884), .I2(n2196), .S0(N47), .S1(n8290), 
        .ZN(N81) );
  MUX3ND0 U8590 ( .I0(n7887), .I1(n7888), .I2(n7889), .S0(n8313), .S1(n8297), 
        .ZN(n7886) );
  MUX3ND0 U8591 ( .I0(n7896), .I1(n7897), .I2(n2194), .S0(N47), .S1(n8290), 
        .ZN(N80) );
  MUX3ND0 U8592 ( .I0(n7900), .I1(n7901), .I2(n7902), .S0(n8312), .S1(n8297), 
        .ZN(n7899) );
  MUX3ND0 U8593 ( .I0(n7909), .I1(n7910), .I2(n2213), .S0(n8686), .S1(n8290), 
        .ZN(N79) );
  MUX3ND0 U8594 ( .I0(n7913), .I1(n7914), .I2(n7915), .S0(n8313), .S1(n8297), 
        .ZN(n7912) );
  MUX3ND0 U8595 ( .I0(n7922), .I1(n7923), .I2(n2200), .S0(N47), .S1(n8290), 
        .ZN(N78) );
  MUX3ND0 U8596 ( .I0(n7926), .I1(n7927), .I2(n7928), .S0(n8312), .S1(n8297), 
        .ZN(n7925) );
  MUX3ND0 U8597 ( .I0(n7935), .I1(n7936), .I2(n2204), .S0(N47), .S1(n8290), 
        .ZN(N77) );
  MUX3ND0 U8598 ( .I0(n7939), .I1(n7940), .I2(n7941), .S0(n8312), .S1(n8297), 
        .ZN(n7938) );
  MUX3ND0 U8599 ( .I0(n7948), .I1(n7949), .I2(n2202), .S0(N47), .S1(n8290), 
        .ZN(N76) );
  MUX3ND0 U8600 ( .I0(n7952), .I1(n7953), .I2(n7954), .S0(n8312), .S1(n8297), 
        .ZN(n7951) );
  MUX3ND0 U8601 ( .I0(n7961), .I1(n7962), .I2(n2191), .S0(N47), .S1(n8290), 
        .ZN(N75) );
  MUX3ND0 U8602 ( .I0(n7965), .I1(n7966), .I2(n7967), .S0(n8311), .S1(n8297), 
        .ZN(n7964) );
  MUX3ND0 U8603 ( .I0(n7974), .I1(n7975), .I2(n2212), .S0(n8686), .S1(n8290), 
        .ZN(N74) );
  MUX3ND0 U8604 ( .I0(n7978), .I1(n7979), .I2(n7980), .S0(n8311), .S1(n8297), 
        .ZN(n7977) );
  MUX3ND0 U8605 ( .I0(n7987), .I1(n7988), .I2(n2209), .S0(n8686), .S1(n8290), 
        .ZN(N73) );
  MUX3ND0 U8606 ( .I0(n7991), .I1(n7992), .I2(n7993), .S0(n8312), .S1(n8297), 
        .ZN(n7990) );
  MUX3ND0 U8607 ( .I0(n8000), .I1(n8001), .I2(n2195), .S0(N47), .S1(n8290), 
        .ZN(N72) );
  MUX3ND0 U8608 ( .I0(n8004), .I1(n8005), .I2(n8006), .S0(n8312), .S1(n8297), 
        .ZN(n8003) );
  MUX3ND0 U8609 ( .I0(n8013), .I1(n8014), .I2(n2160), .S0(N47), .S1(n8290), 
        .ZN(N71) );
  MUX3ND0 U8610 ( .I0(n8017), .I1(n8018), .I2(n8019), .S0(n8312), .S1(n8297), 
        .ZN(n8016) );
  MUX3ND0 U8611 ( .I0(n8030), .I1(n8031), .I2(n8032), .S0(n8313), .S1(n8297), 
        .ZN(n8029) );
  MUX3ND0 U8612 ( .I0(n8039), .I1(n8040), .I2(n2161), .S0(n8686), .S1(n8290), 
        .ZN(N69) );
  MUX3ND0 U8613 ( .I0(n8043), .I1(n8044), .I2(n8045), .S0(n8312), .S1(n8297), 
        .ZN(n8042) );
  MUX3ND0 U8614 ( .I0(n8052), .I1(n8053), .I2(n2166), .S0(N47), .S1(n8290), 
        .ZN(N68) );
  MUX3ND0 U8615 ( .I0(n8056), .I1(n8057), .I2(n8058), .S0(n8312), .S1(n8298), 
        .ZN(n8055) );
  MUX3ND0 U8616 ( .I0(n8065), .I1(n8066), .I2(n2155), .S0(n8686), .S1(n8290), 
        .ZN(N67) );
  MUX3ND0 U8617 ( .I0(n8069), .I1(n8070), .I2(n8071), .S0(n8313), .S1(n8298), 
        .ZN(n8068) );
  MUX3ND0 U8618 ( .I0(n8082), .I1(n8083), .I2(n8084), .S0(n8313), .S1(n8298), 
        .ZN(n8081) );
  MUX3ND0 U8619 ( .I0(n8095), .I1(n8096), .I2(n8097), .S0(n8313), .S1(n8298), 
        .ZN(n8094) );
  MUX3ND0 U8620 ( .I0(n8108), .I1(n8109), .I2(n8110), .S0(n8313), .S1(n8298), 
        .ZN(n8107) );
  MUX3ND0 U8621 ( .I0(n8117), .I1(n8118), .I2(n903), .S0(n8293), .S1(n8290), 
        .ZN(N63) );
  MUX3ND0 U8622 ( .I0(n8121), .I1(n8122), .I2(n8123), .S0(n8313), .S1(n8298), 
        .ZN(n8120) );
  MUX3ND0 U8623 ( .I0(n8134), .I1(n8135), .I2(n8136), .S0(n8313), .S1(n8298), 
        .ZN(n8133) );
  MUX3ND0 U8624 ( .I0(n8147), .I1(n8148), .I2(n8149), .S0(n8313), .S1(n8298), 
        .ZN(n8146) );
  MUX3ND0 U8625 ( .I0(n8160), .I1(n8161), .I2(n8162), .S0(n8312), .S1(n8298), 
        .ZN(n8159) );
  MUX3ND0 U8626 ( .I0(n8173), .I1(n8174), .I2(n8175), .S0(n8311), .S1(n8298), 
        .ZN(n8172) );
  MUX3ND0 U8627 ( .I0(n8186), .I1(n8187), .I2(n8188), .S0(n8312), .S1(n8298), 
        .ZN(n8185) );
  MUX3ND0 U8628 ( .I0(n8199), .I1(n8200), .I2(n8201), .S0(n8311), .S1(n8298), 
        .ZN(n8198) );
  MUX3ND0 U8629 ( .I0(n8212), .I1(n8213), .I2(n8214), .S0(n8311), .S1(n8298), 
        .ZN(n8211) );
  MUX3ND0 U8630 ( .I0(n8225), .I1(n8226), .I2(n8227), .S0(n8312), .S1(n8296), 
        .ZN(n8224) );
  MUX3ND0 U8631 ( .I0(n8238), .I1(n8239), .I2(n8240), .S0(n8311), .S1(n8294), 
        .ZN(n8237) );
  MUX3ND0 U8632 ( .I0(n8251), .I1(n8252), .I2(n8253), .S0(n8313), .S1(n8296), 
        .ZN(n8250) );
  MUX3ND0 U8633 ( .I0(n8264), .I1(n8265), .I2(n8266), .S0(n8312), .S1(n8295), 
        .ZN(n8263) );
  MUX3ND0 U8634 ( .I0(n8273), .I1(n8274), .I2(n111), .S0(n8293), .S1(n8291), 
        .ZN(N51) );
  MUX3ND0 U8635 ( .I0(n8277), .I1(n8278), .I2(n8279), .S0(n8313), .S1(n8295), 
        .ZN(n8276) );
  MUX3ND0 U8636 ( .I0(n8286), .I1(n8287), .I2(n8288), .S0(n8293), .S1(n8291), 
        .ZN(N50) );
  MUX2ND0 U8637 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n8318), 
        .ZN(n7862) );
  MUX2ND0 U8638 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n8318), 
        .ZN(n7861) );
  MUX3ND0 U8639 ( .I0(n7865), .I1(n7864), .I2(n7860), .S0(n8295), .S1(n8293), 
        .ZN(n7872) );
  MUX2ND0 U8640 ( .I0(n7867), .I1(n7866), .S(n8294), .ZN(n7871) );
  MUX2ND0 U8641 ( .I0(n7869), .I1(n7868), .S(n8294), .ZN(n7870) );
  MUX2ND0 U8642 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n8319), 
        .ZN(n7875) );
  MUX2ND0 U8643 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n8319), 
        .ZN(n7874) );
  MUX3ND0 U8644 ( .I0(n7878), .I1(n7877), .I2(n7873), .S0(n8296), .S1(n8293), 
        .ZN(n7885) );
  MUX2ND0 U8645 ( .I0(n7880), .I1(n7879), .S(n8294), .ZN(n7884) );
  MUX2ND0 U8646 ( .I0(n7882), .I1(n7881), .S(n8298), .ZN(n7883) );
  MUX2ND0 U8647 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n8319), 
        .ZN(n7888) );
  MUX2ND0 U8648 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n8319), 
        .ZN(n7887) );
  MUX3ND0 U8649 ( .I0(n7891), .I1(n7890), .I2(n7886), .S0(n8298), .S1(n8293), 
        .ZN(n7898) );
  MUX2ND0 U8650 ( .I0(n7893), .I1(n7892), .S(n8685), .ZN(n7897) );
  MUX2ND0 U8651 ( .I0(n7895), .I1(n7894), .S(N46), .ZN(n7896) );
  MUX2ND0 U8652 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n8319), 
        .ZN(n7901) );
  MUX2ND0 U8653 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n8320), 
        .ZN(n7900) );
  MUX3ND0 U8654 ( .I0(n7904), .I1(n7903), .I2(n7899), .S0(n8299), .S1(n8293), 
        .ZN(n7911) );
  MUX2ND0 U8655 ( .I0(n7906), .I1(n7905), .S(n8685), .ZN(n7910) );
  MUX2ND0 U8656 ( .I0(n7908), .I1(n7907), .S(n8685), .ZN(n7909) );
  MUX2ND0 U8657 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n8320), 
        .ZN(n7914) );
  MUX2ND0 U8658 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n8320), 
        .ZN(n7913) );
  MUX3ND0 U8659 ( .I0(n7917), .I1(n7916), .I2(n7912), .S0(n8298), .S1(n8293), 
        .ZN(n7924) );
  MUX2ND0 U8660 ( .I0(n7919), .I1(n7918), .S(n8295), .ZN(n7923) );
  MUX2ND0 U8661 ( .I0(n7921), .I1(n7920), .S(n8294), .ZN(n7922) );
  MUX2ND0 U8662 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n8320), 
        .ZN(n7927) );
  MUX2ND0 U8663 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n8314), 
        .ZN(n7926) );
  MUX3ND0 U8664 ( .I0(n7930), .I1(n7929), .I2(n7925), .S0(n8299), .S1(n8293), 
        .ZN(n7937) );
  MUX2ND0 U8665 ( .I0(n7932), .I1(n7931), .S(n8685), .ZN(n7936) );
  MUX2ND0 U8666 ( .I0(n7934), .I1(n7933), .S(n8294), .ZN(n7935) );
  MUX2ND0 U8667 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n8314), 
        .ZN(n7940) );
  MUX2ND0 U8668 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n8317), 
        .ZN(n7939) );
  MUX3ND0 U8669 ( .I0(n7943), .I1(n7942), .I2(n7938), .S0(n8299), .S1(n8686), 
        .ZN(n7950) );
  MUX2ND0 U8670 ( .I0(n7945), .I1(n7944), .S(N46), .ZN(n7949) );
  MUX2ND0 U8671 ( .I0(n7947), .I1(n7946), .S(N46), .ZN(n7948) );
  MUX2ND0 U8672 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n8317), 
        .ZN(n7953) );
  MUX2ND0 U8673 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n8317), 
        .ZN(n7952) );
  MUX3ND0 U8674 ( .I0(n7956), .I1(n7955), .I2(n7951), .S0(n8295), .S1(n8686), 
        .ZN(n7963) );
  MUX2ND0 U8675 ( .I0(n7958), .I1(n7957), .S(n8295), .ZN(n7962) );
  MUX2ND0 U8676 ( .I0(n7960), .I1(n7959), .S(n8297), .ZN(n7961) );
  MUX2ND0 U8677 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n8327), 
        .ZN(n7966) );
  MUX2ND0 U8678 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n8314), 
        .ZN(n7965) );
  MUX3ND0 U8679 ( .I0(n7969), .I1(n7968), .I2(n7964), .S0(n8296), .S1(n8686), 
        .ZN(n7976) );
  MUX2ND0 U8680 ( .I0(n7971), .I1(n7970), .S(n8685), .ZN(n7975) );
  MUX2ND0 U8681 ( .I0(n7973), .I1(n7972), .S(N46), .ZN(n7974) );
  MUX2ND0 U8682 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n8317), 
        .ZN(n7979) );
  MUX2ND0 U8683 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n8325), 
        .ZN(n7978) );
  MUX3ND0 U8684 ( .I0(n7982), .I1(n7981), .I2(n7977), .S0(n8299), .S1(n8686), 
        .ZN(n7989) );
  MUX2ND0 U8685 ( .I0(n7984), .I1(n7983), .S(N46), .ZN(n7988) );
  MUX2ND0 U8686 ( .I0(n7986), .I1(n7985), .S(n8296), .ZN(n7987) );
  MUX2ND0 U8687 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n8326), 
        .ZN(n7992) );
  MUX2ND0 U8688 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n8314), 
        .ZN(n7991) );
  MUX3ND0 U8689 ( .I0(n7995), .I1(n7994), .I2(n7990), .S0(n8299), .S1(n8686), 
        .ZN(n8002) );
  MUX2ND0 U8690 ( .I0(n7997), .I1(n7996), .S(n8297), .ZN(n8001) );
  MUX2ND0 U8691 ( .I0(n7999), .I1(n7998), .S(n8299), .ZN(n8000) );
  MUX2ND0 U8692 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n8315), 
        .ZN(n8005) );
  MUX2ND0 U8693 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n8327), 
        .ZN(n8004) );
  MUX3ND0 U8694 ( .I0(n8008), .I1(n8007), .I2(n8003), .S0(n8295), .S1(n8686), 
        .ZN(n8015) );
  MUX2ND0 U8695 ( .I0(n8010), .I1(n8009), .S(n8296), .ZN(n8014) );
  MUX2ND0 U8696 ( .I0(n8012), .I1(n8011), .S(n8297), .ZN(n8013) );
  MUX2ND0 U8697 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n8316), 
        .ZN(n8018) );
  MUX2ND0 U8698 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n8326), 
        .ZN(n8017) );
  MUX3ND0 U8699 ( .I0(n8021), .I1(n8020), .I2(n8016), .S0(n8299), .S1(N47), 
        .ZN(n8028) );
  MUX2ND0 U8700 ( .I0(n8023), .I1(n8022), .S(n8297), .ZN(n8027) );
  MUX2ND0 U8701 ( .I0(n8025), .I1(n8024), .S(n8295), .ZN(n8026) );
  MUX2ND0 U8702 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n8321), 
        .ZN(n8031) );
  MUX2ND0 U8703 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n8315), 
        .ZN(n8030) );
  MUX3ND0 U8704 ( .I0(n8034), .I1(n8033), .I2(n8029), .S0(n8299), .S1(N47), 
        .ZN(n8041) );
  MUX2ND0 U8705 ( .I0(n8036), .I1(n8035), .S(n8299), .ZN(n8040) );
  MUX2ND0 U8706 ( .I0(n8038), .I1(n8037), .S(n8296), .ZN(n8039) );
  MUX2ND0 U8707 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n8317), 
        .ZN(n8044) );
  MUX2ND0 U8708 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n8327), 
        .ZN(n8043) );
  MUX3ND0 U8709 ( .I0(n8047), .I1(n8046), .I2(n8042), .S0(n8294), .S1(n8686), 
        .ZN(n8054) );
  MUX2ND0 U8710 ( .I0(n8049), .I1(n8048), .S(n8294), .ZN(n8053) );
  MUX2ND0 U8711 ( .I0(n8051), .I1(n8050), .S(n8295), .ZN(n8052) );
  MUX2ND0 U8712 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n8321), 
        .ZN(n8057) );
  MUX2ND0 U8713 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n8325), 
        .ZN(n8056) );
  MUX3ND0 U8714 ( .I0(n8060), .I1(n8059), .I2(n8055), .S0(n8296), .S1(N47), 
        .ZN(n8067) );
  MUX2ND0 U8715 ( .I0(n8062), .I1(n8061), .S(n8297), .ZN(n8066) );
  MUX2ND0 U8716 ( .I0(n8064), .I1(n8063), .S(n8294), .ZN(n8065) );
  MUX2ND0 U8717 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n8314), 
        .ZN(n8070) );
  MUX2ND0 U8718 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n8320), 
        .ZN(n8069) );
  MUX3ND0 U8719 ( .I0(n8073), .I1(n8072), .I2(n8068), .S0(n8299), .S1(N47), 
        .ZN(n8080) );
  MUX2ND0 U8720 ( .I0(n8075), .I1(n8074), .S(n8294), .ZN(n8079) );
  MUX2ND0 U8721 ( .I0(n8077), .I1(n8076), .S(n8295), .ZN(n8078) );
  MUX2ND0 U8722 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n8320), 
        .ZN(n8083) );
  MUX2ND0 U8723 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n8320), 
        .ZN(n8082) );
  MUX3ND0 U8724 ( .I0(n8086), .I1(n8085), .I2(n8081), .S0(n8299), .S1(N47), 
        .ZN(n8093) );
  MUX2ND0 U8725 ( .I0(n8088), .I1(n8087), .S(n8295), .ZN(n8092) );
  MUX2ND0 U8726 ( .I0(n8090), .I1(n8089), .S(n8685), .ZN(n8091) );
  MUX2ND0 U8727 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n8320), 
        .ZN(n8096) );
  MUX2ND0 U8728 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n8320), 
        .ZN(n8095) );
  MUX3ND0 U8729 ( .I0(n8099), .I1(n8098), .I2(n8094), .S0(n8299), .S1(n8293), 
        .ZN(n8106) );
  MUX2ND0 U8730 ( .I0(n8101), .I1(n8100), .S(n8685), .ZN(n8105) );
  MUX2ND0 U8731 ( .I0(n8103), .I1(n8102), .S(n8685), .ZN(n8104) );
  MUX2ND0 U8732 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n8320), 
        .ZN(n8109) );
  MUX2ND0 U8733 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n8320), 
        .ZN(n8108) );
  MUX3ND0 U8734 ( .I0(n8112), .I1(n8111), .I2(n8107), .S0(n8295), .S1(n8292), 
        .ZN(n8119) );
  MUX2ND0 U8735 ( .I0(n8114), .I1(n8113), .S(n8685), .ZN(n8118) );
  MUX2ND0 U8736 ( .I0(n8116), .I1(n8115), .S(n8685), .ZN(n8117) );
  MUX2ND0 U8737 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n8320), 
        .ZN(n8122) );
  MUX2ND0 U8738 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n8320), 
        .ZN(n8121) );
  MUX3ND0 U8739 ( .I0(n8125), .I1(n8124), .I2(n8120), .S0(n8299), .S1(n8292), 
        .ZN(n8132) );
  MUX2ND0 U8740 ( .I0(n8127), .I1(n8126), .S(n8685), .ZN(n8131) );
  MUX2ND0 U8741 ( .I0(n8129), .I1(n8128), .S(n8685), .ZN(n8130) );
  MUX2ND0 U8742 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n8320), 
        .ZN(n8135) );
  MUX2ND0 U8743 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n8320), 
        .ZN(n8134) );
  MUX3ND0 U8744 ( .I0(n8138), .I1(n8137), .I2(n8133), .S0(n8294), .S1(n8292), 
        .ZN(n8145) );
  MUX2ND0 U8745 ( .I0(n8140), .I1(n8139), .S(n8685), .ZN(n8144) );
  MUX2ND0 U8746 ( .I0(n8142), .I1(n8141), .S(n8685), .ZN(n8143) );
  MUX2ND0 U8747 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n8320), 
        .ZN(n8148) );
  MUX2ND0 U8748 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n8320), 
        .ZN(n8147) );
  MUX3ND0 U8749 ( .I0(n8151), .I1(n8150), .I2(n8146), .S0(n8294), .S1(n8292), 
        .ZN(n8158) );
  MUX2ND0 U8750 ( .I0(n8153), .I1(n8152), .S(n8294), .ZN(n8157) );
  MUX2ND0 U8751 ( .I0(n8155), .I1(n8154), .S(n8685), .ZN(n8156) );
  MUX2ND0 U8752 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n8320), 
        .ZN(n8161) );
  MUX2ND0 U8753 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n8320), 
        .ZN(n8160) );
  MUX3ND0 U8754 ( .I0(n8164), .I1(n8163), .I2(n8159), .S0(n8299), .S1(n8292), 
        .ZN(n8171) );
  MUX2ND0 U8755 ( .I0(n8166), .I1(n8165), .S(n8297), .ZN(n8170) );
  MUX2ND0 U8756 ( .I0(n8168), .I1(n8167), .S(n8295), .ZN(n8169) );
  MUX2ND0 U8757 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n8320), 
        .ZN(n8174) );
  MUX2ND0 U8758 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n8319), 
        .ZN(n8173) );
  MUX3ND0 U8759 ( .I0(n8177), .I1(n8176), .I2(n8172), .S0(n8299), .S1(n8292), 
        .ZN(n8184) );
  MUX2ND0 U8760 ( .I0(n8179), .I1(n8178), .S(n8294), .ZN(n8183) );
  MUX2ND0 U8761 ( .I0(n8181), .I1(n8180), .S(n8295), .ZN(n8182) );
  MUX2ND0 U8762 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n8319), 
        .ZN(n8187) );
  MUX2ND0 U8763 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n8319), 
        .ZN(n8186) );
  MUX3ND0 U8764 ( .I0(n8190), .I1(n8189), .I2(n8185), .S0(n8299), .S1(n8292), 
        .ZN(n8197) );
  MUX2ND0 U8765 ( .I0(n8192), .I1(n8191), .S(n8294), .ZN(n8196) );
  MUX2ND0 U8766 ( .I0(n8194), .I1(n8193), .S(n8294), .ZN(n8195) );
  MUX2ND0 U8767 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n8319), 
        .ZN(n8200) );
  MUX2ND0 U8768 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n8319), 
        .ZN(n8199) );
  MUX3ND0 U8769 ( .I0(n8203), .I1(n8202), .I2(n8198), .S0(n8298), .S1(n8292), 
        .ZN(n8210) );
  MUX2ND0 U8770 ( .I0(n8205), .I1(n8204), .S(n8295), .ZN(n8209) );
  MUX2ND0 U8771 ( .I0(n8207), .I1(n8206), .S(n8296), .ZN(n8208) );
  MUX2ND0 U8772 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n8319), 
        .ZN(n8213) );
  MUX2ND0 U8773 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n8319), 
        .ZN(n8212) );
  MUX3ND0 U8774 ( .I0(n8216), .I1(n8215), .I2(n8211), .S0(n8299), .S1(n8292), 
        .ZN(n8223) );
  MUX2ND0 U8775 ( .I0(n8218), .I1(n8217), .S(n8296), .ZN(n8222) );
  MUX2ND0 U8776 ( .I0(n8220), .I1(n8219), .S(n8296), .ZN(n8221) );
  MUX2ND0 U8777 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n8319), 
        .ZN(n8226) );
  MUX2ND0 U8778 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n8319), 
        .ZN(n8225) );
  MUX3ND0 U8779 ( .I0(n8229), .I1(n8228), .I2(n8224), .S0(n8296), .S1(n8292), 
        .ZN(n8236) );
  MUX2ND0 U8780 ( .I0(n8231), .I1(n8230), .S(n8294), .ZN(n8235) );
  MUX2ND0 U8781 ( .I0(n8233), .I1(n8232), .S(n8296), .ZN(n8234) );
  MUX2ND0 U8782 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n8319), 
        .ZN(n8239) );
  MUX2ND0 U8783 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n8319), 
        .ZN(n8238) );
  MUX3ND0 U8784 ( .I0(n8242), .I1(n8241), .I2(n8237), .S0(n8294), .S1(n8292), 
        .ZN(n8249) );
  MUX2ND0 U8785 ( .I0(n8244), .I1(n8243), .S(n8685), .ZN(n8248) );
  MUX2ND0 U8786 ( .I0(n8246), .I1(n8245), .S(n8685), .ZN(n8247) );
  MUX2ND0 U8787 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n8319), 
        .ZN(n8252) );
  MUX2ND0 U8788 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n8319), 
        .ZN(n8251) );
  MUX3ND0 U8789 ( .I0(n8255), .I1(n8254), .I2(n8250), .S0(n8295), .S1(n8292), 
        .ZN(n8262) );
  MUX2ND0 U8790 ( .I0(n8257), .I1(n8256), .S(n8297), .ZN(n8261) );
  MUX2ND0 U8791 ( .I0(n8259), .I1(n8258), .S(n8685), .ZN(n8260) );
  MUX2ND0 U8792 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n8319), 
        .ZN(n8265) );
  MUX2ND0 U8793 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n8319), 
        .ZN(n8264) );
  MUX3ND0 U8794 ( .I0(n8268), .I1(n8267), .I2(n8263), .S0(n8299), .S1(n8292), 
        .ZN(n8275) );
  MUX2ND0 U8795 ( .I0(n8270), .I1(n8269), .S(n8296), .ZN(n8274) );
  MUX2ND0 U8796 ( .I0(n8272), .I1(n8271), .S(n8296), .ZN(n8273) );
  MUX2ND0 U8797 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n8318), 
        .ZN(n8278) );
  MUX2ND0 U8798 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n8317), 
        .ZN(n8277) );
  MUX3ND0 U8799 ( .I0(n8281), .I1(n8280), .I2(n8276), .S0(n8295), .S1(n8293), 
        .ZN(n8288) );
  MUX2ND0 U8800 ( .I0(n8283), .I1(n8282), .S(n8296), .ZN(n8287) );
  MUX2ND0 U8801 ( .I0(n8285), .I1(n8284), .S(n8294), .ZN(n8286) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n2, \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  BUFFD0 U1 ( .I(n2), .Z(SUM[0]) );
  CKXOR2D0 U2 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U3 ( .CLK(A[0]), .CN(n2) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n7, \carry[4] , \carry[3] , \carry[2] , n1, n2, n4, n5;

  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(n4), .CO(\carry[2] ), .S(n7) );
  INVD8 U1 ( .I(n7), .ZN(n1) );
  INVD1 U2 ( .I(n1), .ZN(n2) );
  CKBD0 U3 ( .CLK(n2), .C(SUM[1]) );
  CKNXD16 U4 ( .I(n4), .ZN(SUM[0]) );
  INVD0 U5 ( .I(n5), .ZN(n4) );
  CKNXD16 U6 ( .I(A[0]), .ZN(n5) );
  CKXOR2D0 U7 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
endmodule

