
module Deserializer ( ParOut, ParValid, DecoderParClk, FIFOEmpty, FIFOFull, 
        ParOutClk, SerialIn, FIFOReadCmd, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, FIFOReadCmd, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n2, n4;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFO_Top_AWid5_DWid32 FIFO_U1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(FIFOReadCmd), .WriteIn(
        ParValidDecode), .Clocker(DecoderParClk), .Reseter(Reset) );
  DesDecoder_DWid32 DesDecoder_U1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(Reset) );
  SerialRx SerialRx_U1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(Reset) );
  DFCNQD1 ParValidReg_reg ( .D(N35), .CP(ParOutClk), .CDN(n2), .Q(ParValid) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n2), .Q(ParOut[31])
         );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n2), .Q(ParOut[30])
         );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n2), .Q(ParOut[29])
         );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n2), .Q(ParOut[28])
         );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n2), .Q(ParOut[27])
         );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n2), .Q(ParOut[26])
         );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n2), .Q(ParOut[25])
         );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n2), .Q(ParOut[24])
         );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n2), .Q(ParOut[23])
         );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n2), .Q(ParOut[22])
         );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n2), .Q(ParOut[21])
         );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n2), .Q(ParOut[20])
         );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n2), .Q(ParOut[19])
         );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n2), .Q(ParOut[18])
         );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n2), .Q(ParOut[17])
         );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n2), .Q(ParOut[16])
         );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n2), .Q(ParOut[15])
         );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n2), .Q(ParOut[14])
         );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n2), .Q(ParOut[13])
         );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n2), .Q(ParOut[12])
         );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n2), .Q(ParOut[11])
         );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n2), .Q(ParOut[10])
         );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n2), .Q(ParOut[9])
         );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n2), .Q(ParOut[8])
         );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n2), .Q(ParOut[7])
         );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n2), .Q(ParOut[6]) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n2), .Q(ParOut[5]) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n2), .Q(ParOut[4]) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n2), .Q(ParOut[3]) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n2), .Q(ParOut[2]) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n2), .Q(ParOut[1]) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n2), .Q(ParOut[0]) );
  INVD2 U38 ( .I(Reset), .ZN(n2) );
  AN2D0 U39 ( .A1(FIFO_Out[6]), .A2(FIFOReadCmd), .Z(N9) );
  AN2D0 U40 ( .A1(FIFO_Out[5]), .A2(FIFOReadCmd), .Z(N8) );
  AN2D0 U41 ( .A1(FIFO_Out[4]), .A2(FIFOReadCmd), .Z(N7) );
  AN2D0 U42 ( .A1(FIFO_Out[3]), .A2(FIFOReadCmd), .Z(N6) );
  AN2D0 U43 ( .A1(FIFO_Out[2]), .A2(FIFOReadCmd), .Z(N5) );
  AN2D0 U44 ( .A1(FIFO_Out[1]), .A2(FIFOReadCmd), .Z(N4) );
  NR2D0 U45 ( .A1(FIFOEmpty), .A2(n4), .ZN(N35) );
  CKND0 U46 ( .CLK(FIFOReadCmd), .CN(n4) );
  AN2D0 U47 ( .A1(FIFO_Out[31]), .A2(FIFOReadCmd), .Z(N34) );
  AN2D0 U48 ( .A1(FIFO_Out[30]), .A2(FIFOReadCmd), .Z(N33) );
  AN2D0 U49 ( .A1(FIFO_Out[29]), .A2(FIFOReadCmd), .Z(N32) );
  AN2D0 U50 ( .A1(FIFO_Out[28]), .A2(FIFOReadCmd), .Z(N31) );
  AN2D0 U51 ( .A1(FIFO_Out[27]), .A2(FIFOReadCmd), .Z(N30) );
  AN2D0 U52 ( .A1(FIFO_Out[0]), .A2(FIFOReadCmd), .Z(N3) );
  AN2D0 U53 ( .A1(FIFO_Out[26]), .A2(FIFOReadCmd), .Z(N29) );
  AN2D0 U54 ( .A1(FIFO_Out[25]), .A2(FIFOReadCmd), .Z(N28) );
  AN2D0 U55 ( .A1(FIFO_Out[24]), .A2(FIFOReadCmd), .Z(N27) );
  AN2D0 U56 ( .A1(FIFO_Out[23]), .A2(FIFOReadCmd), .Z(N26) );
  AN2D0 U57 ( .A1(FIFO_Out[22]), .A2(FIFOReadCmd), .Z(N25) );
  AN2D0 U58 ( .A1(FIFO_Out[21]), .A2(FIFOReadCmd), .Z(N24) );
  AN2D0 U59 ( .A1(FIFO_Out[20]), .A2(FIFOReadCmd), .Z(N23) );
  AN2D0 U60 ( .A1(FIFO_Out[19]), .A2(FIFOReadCmd), .Z(N22) );
  AN2D0 U61 ( .A1(FIFO_Out[18]), .A2(FIFOReadCmd), .Z(N21) );
  AN2D0 U62 ( .A1(FIFO_Out[17]), .A2(FIFOReadCmd), .Z(N20) );
  AN2D0 U63 ( .A1(FIFO_Out[16]), .A2(FIFOReadCmd), .Z(N19) );
  AN2D0 U64 ( .A1(FIFO_Out[15]), .A2(FIFOReadCmd), .Z(N18) );
  AN2D0 U65 ( .A1(FIFO_Out[14]), .A2(FIFOReadCmd), .Z(N17) );
  AN2D0 U66 ( .A1(FIFO_Out[13]), .A2(FIFOReadCmd), .Z(N16) );
  AN2D0 U67 ( .A1(FIFO_Out[12]), .A2(FIFOReadCmd), .Z(N15) );
  AN2D0 U68 ( .A1(FIFO_Out[11]), .A2(FIFOReadCmd), .Z(N14) );
  AN2D0 U69 ( .A1(FIFO_Out[10]), .A2(FIFOReadCmd), .Z(N13) );
  AN2D0 U70 ( .A1(FIFO_Out[9]), .A2(FIFOReadCmd), .Z(N12) );
  AN2D0 U71 ( .A1(FIFO_Out[8]), .A2(FIFOReadCmd), .Z(N11) );
  AN2D0 U72 ( .A1(FIFO_Out[7]), .A2(FIFOReadCmd), .Z(N10) );
endmodule


module FIFO_Top_AWid5_DWid32 ( Dout, Din, Full, Empty, ReadIn, WriteIn, 
        Clocker, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, Clocker, Reseter;
  output Full, Empty;
  wire   SM_MemReadCmd, SM_MemWriteCmd, Mem_Enable, n1;
  wire   [4:0] SM_MemAddr;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), .WriteReq(WriteIn), .Clk(
        Clocker), .Reset(Reseter) );
  Mem1kx32_AWid5_DWid32 RegFile1 ( .DataO(Dout), .DataI(Din), .Addr(SM_MemAddr), .ClockIn(Clocker), .ChipEna(Mem_Enable), .Read(SM_MemReadCmd), .Write(
        SM_MemWriteCmd), .Reset(Reseter) );
  AOI211XD4 U1 ( .A1(SM_MemWriteCmd), .A2(SM_MemReadCmd), .B(Full), .C(Empty), 
        .ZN(Mem_Enable) );
  MUX2D2 U2 ( .I0(SM_WriteAddr[4]), .I1(SM_ReadAddr[4]), .S(n1), .Z(
        SM_MemAddr[4]) );
  MUX2D4 U3 ( .I0(SM_WriteAddr[3]), .I1(SM_ReadAddr[3]), .S(n1), .Z(
        SM_MemAddr[3]) );
  MUX2D0 U4 ( .I0(SM_WriteAddr[2]), .I1(SM_ReadAddr[2]), .S(n1), .Z(
        SM_MemAddr[2]) );
  MUX2D0 U5 ( .I0(SM_WriteAddr[1]), .I1(SM_ReadAddr[1]), .S(n1), .Z(
        SM_MemAddr[1]) );
  MUX2D0 U6 ( .I0(SM_WriteAddr[0]), .I1(SM_ReadAddr[0]), .S(n1), .Z(
        SM_MemAddr[0]) );
  INR2D0 U7 ( .A1(SM_MemReadCmd), .B1(SM_MemWriteCmd), .ZN(n1) );
endmodule


module DesDecoder_DWid32 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   N12, N44, N49, N50, N51, N52, N53, N62, N63, N65, N66, N67, N68, N69,
         N70, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n123, n124, n125, n126, n127, n128,
         n129, n130, n133, n134, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n155, n156, n157, n158, n159, n160, n161, n162,
         n164, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n131, n132,
         n135, n136, n137, n138, n149, n150, n151, n152, n153, n154, n163,
         n165, n166, n167, n168, n179, n180, n181, n182, n183, n184, n185,
         n186, n254, n255, n256, n257, n258, n259;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  DFNCND2 UnLoad_reg ( .D(N44), .CPN(n96), .CDN(n253), .QN(n117) );
  LHQD1 \Count32_reg[0]  ( .E(N69), .D(N65), .Q(Count32[0]) );
  LHQD1 \Count32_reg[1]  ( .E(N69), .D(N66), .Q(Count32[1]) );
  LHQD1 \Count32_reg[2]  ( .E(N69), .D(N67), .Q(Count32[2]) );
  LHQD1 \Count32_reg[3]  ( .E(N69), .D(N68), .Q(Count32[3]) );
  LHQD1 \Count32_reg[4]  ( .E(N69), .D(N70), .Q(Count32[4]) );
  LHQD1 ParClkReg_reg ( .E(N62), .D(N63), .Q(ParClk) );
  DesDecoder_DWid32_DW01_inc_0 \SerClockGen/add_170_C252_S2  ( .A(Count32), 
        .SUM({N53, N52, N51, N50, N49}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(FrameSR[62]), .CPN(n95), .CDN(n253), .QN(n123) );
  DFNCND1 \DecodeReg_reg[31]  ( .D(n251), .CPN(n96), .CDN(n91), .QN(n255) );
  DFNCND1 \DecodeReg_reg[30]  ( .D(n250), .CPN(n95), .CDN(n93), .QN(n254) );
  DFNCND1 \DecodeReg_reg[29]  ( .D(n249), .CPN(n97), .CDN(n94), .QN(n186) );
  DFNCND1 \DecodeReg_reg[28]  ( .D(n248), .CPN(n96), .CDN(n92), .QN(n185) );
  DFNCND1 \DecodeReg_reg[27]  ( .D(n247), .CPN(n95), .CDN(n253), .QN(n184) );
  DFNCND1 \DecodeReg_reg[26]  ( .D(n246), .CPN(n97), .CDN(n91), .QN(n183) );
  DFNCND1 \DecodeReg_reg[25]  ( .D(n245), .CPN(n252), .CDN(n93), .QN(n182) );
  DFNCND1 \DecodeReg_reg[24]  ( .D(n244), .CPN(n97), .CDN(n94), .QN(n181) );
  DFNCND1 \DecodeReg_reg[23]  ( .D(n243), .CPN(n252), .CDN(n92), .QN(n180) );
  DFNCND1 \DecodeReg_reg[22]  ( .D(n242), .CPN(n96), .CDN(n253), .QN(n179) );
  DFNCND1 \DecodeReg_reg[21]  ( .D(n241), .CPN(n252), .CDN(n91), .QN(n168) );
  DFNCND1 \DecodeReg_reg[20]  ( .D(n240), .CPN(n97), .CDN(n253), .QN(n167) );
  DFNCND1 \DecodeReg_reg[19]  ( .D(n239), .CPN(n95), .CDN(n94), .QN(n166) );
  DFNCND1 \DecodeReg_reg[18]  ( .D(n238), .CPN(n97), .CDN(n93), .QN(n165) );
  DFNCND1 \DecodeReg_reg[17]  ( .D(n237), .CPN(n95), .CDN(n94), .QN(n163) );
  DFNCND1 \DecodeReg_reg[16]  ( .D(n236), .CPN(n252), .CDN(n92), .QN(n154) );
  DFNCND1 \DecodeReg_reg[15]  ( .D(n235), .CPN(n252), .CDN(n94), .QN(n153) );
  DFNCND1 \DecodeReg_reg[14]  ( .D(n234), .CPN(n96), .CDN(n93), .QN(n152) );
  DFNCND1 \DecodeReg_reg[13]  ( .D(n233), .CPN(n97), .CDN(n253), .QN(n151) );
  DFNCND1 \DecodeReg_reg[12]  ( .D(n232), .CPN(n95), .CDN(n93), .QN(n150) );
  DFNCND1 \DecodeReg_reg[11]  ( .D(n231), .CPN(n95), .CDN(n94), .QN(n149) );
  DFNCND1 \DecodeReg_reg[10]  ( .D(n230), .CPN(n96), .CDN(n92), .QN(n138) );
  DFNCND1 \DecodeReg_reg[9]  ( .D(n229), .CPN(n95), .CDN(n253), .QN(n137) );
  DFNCND1 \DecodeReg_reg[8]  ( .D(n228), .CPN(n97), .CDN(n92), .QN(n136) );
  DFNCND1 \DecodeReg_reg[7]  ( .D(n227), .CPN(n97), .CDN(n94), .QN(n135) );
  DFNCND1 \DecodeReg_reg[6]  ( .D(n226), .CPN(n97), .CDN(n91), .QN(n132) );
  DFNCND1 \DecodeReg_reg[5]  ( .D(n225), .CPN(n96), .CDN(n93), .QN(n131) );
  DFNCND1 \DecodeReg_reg[4]  ( .D(n224), .CPN(n252), .CDN(n92), .QN(n122) );
  DFNCND1 \DecodeReg_reg[3]  ( .D(n223), .CPN(n96), .CDN(n93), .QN(n121) );
  DFNCND1 \DecodeReg_reg[2]  ( .D(n222), .CPN(n97), .CDN(n94), .QN(n120) );
  DFNCND1 \DecodeReg_reg[1]  ( .D(n221), .CPN(n96), .CDN(n93), .QN(n119) );
  DFNCND1 \DecodeReg_reg[0]  ( .D(n220), .CPN(n252), .CDN(n91), .QN(n118) );
  DFNCND1 \FrameSR_reg[8]  ( .D(FrameSR[7]), .CPN(n96), .CDN(n93), .Q(
        FrameSR[8]), .QN(n178) );
  DFNCND1 \FrameSR_reg[9]  ( .D(FrameSR[8]), .CPN(n252), .CDN(n93), .Q(
        FrameSR[9]), .QN(n177) );
  DFNCND1 \FrameSR_reg[10]  ( .D(FrameSR[9]), .CPN(n252), .CDN(n91), .Q(
        FrameSR[10]), .QN(n176) );
  DFNCND1 \FrameSR_reg[11]  ( .D(FrameSR[10]), .CPN(n96), .CDN(n91), .Q(
        FrameSR[11]), .QN(n175) );
  DFNCND1 \FrameSR_reg[12]  ( .D(FrameSR[11]), .CPN(n97), .CDN(n91), .Q(
        FrameSR[12]), .QN(n174) );
  DFNCND1 \FrameSR_reg[13]  ( .D(FrameSR[12]), .CPN(n97), .CDN(n91), .Q(
        FrameSR[13]), .QN(n173) );
  DFNCND1 \FrameSR_reg[14]  ( .D(FrameSR[13]), .CPN(n95), .CDN(n91), .Q(
        FrameSR[14]), .QN(n172) );
  DFNCND1 \FrameSR_reg[15]  ( .D(FrameSR[14]), .CPN(n252), .CDN(n91), .Q(
        FrameSR[15]), .QN(n171) );
  DFNCND1 \FrameSR_reg[16]  ( .D(FrameSR[15]), .CPN(n96), .CDN(n91), .Q(
        FrameSR[16]), .QN(n170) );
  DFNCND1 \FrameSR_reg[17]  ( .D(FrameSR[16]), .CPN(n97), .CDN(n91), .Q(
        FrameSR[17]), .QN(n169) );
  DFNCND1 \FrameSR_reg[22]  ( .D(FrameSR[21]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[22]), .QN(n164) );
  DFNCND1 \FrameSR_reg[24]  ( .D(FrameSR[23]), .CPN(n252), .CDN(n94), .Q(
        FrameSR[24]), .QN(n162) );
  DFNCND1 \FrameSR_reg[25]  ( .D(FrameSR[24]), .CPN(n95), .CDN(n93), .Q(
        FrameSR[25]), .QN(n161) );
  DFNCND1 \FrameSR_reg[26]  ( .D(FrameSR[25]), .CPN(n97), .CDN(n253), .Q(
        FrameSR[26]), .QN(n160) );
  DFNCND1 \FrameSR_reg[27]  ( .D(FrameSR[26]), .CPN(n96), .CDN(n92), .Q(
        FrameSR[27]), .QN(n159) );
  DFNCND1 \FrameSR_reg[28]  ( .D(FrameSR[27]), .CPN(n252), .CDN(n93), .Q(
        FrameSR[28]), .QN(n158) );
  DFNCND1 \FrameSR_reg[29]  ( .D(FrameSR[28]), .CPN(n95), .CDN(n94), .Q(
        FrameSR[29]), .QN(n157) );
  DFNCND1 \FrameSR_reg[30]  ( .D(FrameSR[29]), .CPN(n97), .CDN(n94), .Q(
        FrameSR[30]), .QN(n156) );
  DFNCND1 \FrameSR_reg[31]  ( .D(FrameSR[30]), .CPN(n97), .CDN(n93), .Q(
        FrameSR[31]), .QN(n155) );
  DFNCND1 \FrameSR_reg[33]  ( .D(FrameSR[32]), .CPN(n97), .CDN(n93), .Q(
        FrameSR[33]), .QN(n259) );
  DFNCND1 \FrameSR_reg[34]  ( .D(FrameSR[33]), .CPN(n97), .CDN(n94), .Q(
        FrameSR[34]), .QN(n257) );
  DFNCND1 \FrameSR_reg[35]  ( .D(FrameSR[34]), .CPN(n97), .CDN(n93), .Q(
        FrameSR[35]), .QN(n258) );
  DFNCND1 \FrameSR_reg[38]  ( .D(FrameSR[37]), .CPN(n97), .CDN(n94), .Q(
        FrameSR[38]), .QN(n148) );
  DFNCND1 \FrameSR_reg[39]  ( .D(FrameSR[38]), .CPN(n97), .CDN(n93), .Q(
        FrameSR[39]), .QN(n147) );
  DFNCND1 \FrameSR_reg[40]  ( .D(FrameSR[39]), .CPN(n97), .CDN(n91), .Q(
        FrameSR[40]), .QN(n146) );
  DFNCND1 \FrameSR_reg[41]  ( .D(FrameSR[40]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[41]), .QN(n145) );
  DFNCND1 \FrameSR_reg[42]  ( .D(FrameSR[41]), .CPN(n96), .CDN(n92), .Q(
        FrameSR[42]), .QN(n144) );
  DFNCND1 \FrameSR_reg[43]  ( .D(FrameSR[42]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[43]), .QN(n143) );
  DFNCND1 \FrameSR_reg[44]  ( .D(FrameSR[43]), .CPN(n96), .CDN(n93), .Q(
        FrameSR[44]), .QN(n142) );
  DFNCND1 \FrameSR_reg[45]  ( .D(FrameSR[44]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[45]), .QN(n141) );
  DFNCND1 \FrameSR_reg[46]  ( .D(FrameSR[45]), .CPN(n96), .CDN(n91), .Q(
        FrameSR[46]), .QN(n140) );
  DFNCND1 \FrameSR_reg[47]  ( .D(FrameSR[46]), .CPN(n96), .CDN(n92), .Q(
        FrameSR[47]), .QN(n139) );
  DFNCND1 \FrameSR_reg[52]  ( .D(FrameSR[51]), .CPN(n95), .CDN(n253), .Q(
        FrameSR[52]), .QN(n134) );
  DFNCND1 \FrameSR_reg[53]  ( .D(FrameSR[52]), .CPN(n95), .CDN(n253), .Q(
        FrameSR[53]), .QN(n133) );
  DFNCND1 \FrameSR_reg[56]  ( .D(FrameSR[55]), .CPN(n95), .CDN(n91), .Q(
        FrameSR[56]), .QN(n130) );
  DFNCND1 \FrameSR_reg[57]  ( .D(FrameSR[56]), .CPN(n95), .CDN(n93), .Q(
        FrameSR[57]), .QN(n129) );
  DFNCND1 \FrameSR_reg[58]  ( .D(FrameSR[57]), .CPN(n95), .CDN(n93), .Q(
        FrameSR[58]), .QN(n128) );
  DFNCND1 \FrameSR_reg[59]  ( .D(FrameSR[58]), .CPN(n95), .CDN(n94), .Q(
        FrameSR[59]), .QN(n127) );
  DFNCND1 \FrameSR_reg[60]  ( .D(FrameSR[59]), .CPN(n95), .CDN(n92), .Q(
        FrameSR[60]), .QN(n126) );
  DFNCND1 \FrameSR_reg[61]  ( .D(FrameSR[60]), .CPN(n252), .CDN(n92), .Q(
        FrameSR[61]), .QN(n125) );
  DFNCND1 \FrameSR_reg[62]  ( .D(FrameSR[61]), .CPN(n97), .CDN(n253), .Q(
        FrameSR[62]), .QN(n124) );
  DFNCND1 doParSync_reg ( .D(N12), .CPN(n252), .CDN(n94), .Q(n256) );
  DFNCND1 \FrameSR_reg[19]  ( .D(FrameSR[18]), .CPN(n252), .CDN(n91), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(FrameSR[50]), .CPN(n95), .CDN(n94), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(FrameSR[35]), .CPN(n97), .CDN(n92), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n252), .CDN(n94), .Q(FrameSR[0])
         );
  DFNCND1 \FrameSR_reg[1]  ( .D(FrameSR[0]), .CPN(n252), .CDN(n92), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(FrameSR[1]), .CPN(n95), .CDN(n253), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(FrameSR[3]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(FrameSR[4]), .CPN(n97), .CDN(n94), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(FrameSR[5]), .CPN(n96), .CDN(n91), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(FrameSR[17]), .CPN(n95), .CDN(n91), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(FrameSR[19]), .CPN(n252), .CDN(n91), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(FrameSR[20]), .CPN(n96), .CDN(n92), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(FrameSR[22]), .CPN(n252), .CDN(n91), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(FrameSR[31]), .CPN(n97), .CDN(n92), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(FrameSR[36]), .CPN(n97), .CDN(n94), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(FrameSR[47]), .CPN(n96), .CDN(n253), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(FrameSR[48]), .CPN(n96), .CDN(n91), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(FrameSR[49]), .CPN(n96), .CDN(n92), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(FrameSR[53]), .CPN(n95), .CDN(n92), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(FrameSR[54]), .CPN(n95), .CDN(n91), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(FrameSR[2]), .CPN(n95), .CDN(n94), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(FrameSR[6]), .CPN(n252), .CDN(n93), .Q(
        FrameSR[7]) );
  DFNCND1 ParValidReg_reg ( .D(n187), .CPN(n95), .CDN(n93), .Q(ParValid), .QN(
        n57) );
  DFNCND1 \ParOutReg_reg[0]  ( .D(n219), .CPN(n95), .CDN(n94), .Q(ParOut[0]), 
        .QN(n89) );
  DFNCND1 \ParOutReg_reg[2]  ( .D(n217), .CPN(n252), .CDN(n94), .Q(ParOut[2]), 
        .QN(n87) );
  DFNCND1 \ParOutReg_reg[5]  ( .D(n214), .CPN(n95), .CDN(n91), .Q(ParOut[5]), 
        .QN(n84) );
  DFNCND1 \ParOutReg_reg[6]  ( .D(n213), .CPN(n97), .CDN(n253), .Q(ParOut[6]), 
        .QN(n83) );
  DFNCND1 \ParOutReg_reg[9]  ( .D(n210), .CPN(n96), .CDN(n94), .Q(ParOut[9]), 
        .QN(n80) );
  DFNCND1 \ParOutReg_reg[12]  ( .D(n207), .CPN(n252), .CDN(n91), .Q(ParOut[12]), .QN(n77) );
  DFNCND1 \ParOutReg_reg[13]  ( .D(n206), .CPN(n252), .CDN(n93), .Q(ParOut[13]), .QN(n76) );
  DFNCND1 \ParOutReg_reg[16]  ( .D(n203), .CPN(n95), .CDN(n94), .Q(ParOut[16]), 
        .QN(n73) );
  DFNCND1 \ParOutReg_reg[19]  ( .D(n200), .CPN(n96), .CDN(n253), .Q(ParOut[19]), .QN(n70) );
  DFNCND1 \ParOutReg_reg[20]  ( .D(n199), .CPN(n252), .CDN(n93), .Q(ParOut[20]), .QN(n69) );
  DFNCND1 \ParOutReg_reg[23]  ( .D(n196), .CPN(n95), .CDN(n253), .Q(ParOut[23]), .QN(n66) );
  DFNCND1 \ParOutReg_reg[24]  ( .D(n195), .CPN(n97), .CDN(n92), .Q(ParOut[24]), 
        .QN(n65) );
  DFNCND1 \ParOutReg_reg[27]  ( .D(n192), .CPN(n95), .CDN(n94), .Q(ParOut[27]), 
        .QN(n62) );
  DFNCND1 \ParOutReg_reg[28]  ( .D(n191), .CPN(n97), .CDN(n93), .Q(ParOut[28]), 
        .QN(n61) );
  DFNCND1 \ParOutReg_reg[31]  ( .D(n188), .CPN(n252), .CDN(n92), .Q(ParOut[31]), .QN(n58) );
  DFNCND1 \ParOutReg_reg[1]  ( .D(n218), .CPN(n95), .CDN(n93), .Q(ParOut[1]), 
        .QN(n88) );
  DFNCND1 \ParOutReg_reg[3]  ( .D(n216), .CPN(n252), .CDN(n92), .Q(ParOut[3]), 
        .QN(n86) );
  DFNCND1 \ParOutReg_reg[4]  ( .D(n215), .CPN(n96), .CDN(n91), .Q(ParOut[4]), 
        .QN(n85) );
  DFNCND1 \ParOutReg_reg[10]  ( .D(n209), .CPN(n252), .CDN(n93), .Q(ParOut[10]), .QN(n79) );
  DFNCND1 \ParOutReg_reg[11]  ( .D(n208), .CPN(n95), .CDN(n91), .Q(ParOut[11]), 
        .QN(n78) );
  DFNCND1 \ParOutReg_reg[17]  ( .D(n202), .CPN(n97), .CDN(n92), .Q(ParOut[17]), 
        .QN(n72) );
  DFNCND1 \ParOutReg_reg[18]  ( .D(n201), .CPN(n95), .CDN(n92), .Q(ParOut[18]), 
        .QN(n71) );
  DFNCND1 \ParOutReg_reg[7]  ( .D(n212), .CPN(n96), .CDN(n253), .Q(ParOut[7]), 
        .QN(n82) );
  DFNCND1 \ParOutReg_reg[8]  ( .D(n211), .CPN(n95), .CDN(n93), .Q(ParOut[8]), 
        .QN(n81) );
  DFNCND1 \ParOutReg_reg[14]  ( .D(n205), .CPN(n97), .CDN(n92), .Q(ParOut[14]), 
        .QN(n75) );
  DFNCND1 \ParOutReg_reg[15]  ( .D(n204), .CPN(n96), .CDN(n92), .Q(ParOut[15]), 
        .QN(n74) );
  DFNCND1 \ParOutReg_reg[21]  ( .D(n198), .CPN(n97), .CDN(n92), .Q(ParOut[21]), 
        .QN(n68) );
  DFNCND1 \ParOutReg_reg[22]  ( .D(n197), .CPN(n96), .CDN(n94), .Q(ParOut[22]), 
        .QN(n67) );
  DFNCND1 \ParOutReg_reg[25]  ( .D(n194), .CPN(n252), .CDN(n91), .Q(ParOut[25]), .QN(n64) );
  DFNCND1 \ParOutReg_reg[26]  ( .D(n193), .CPN(n97), .CDN(n253), .Q(ParOut[26]), .QN(n63) );
  DFNCND1 \ParOutReg_reg[29]  ( .D(n190), .CPN(n252), .CDN(n253), .Q(
        ParOut[29]), .QN(n60) );
  DFNCND1 \ParOutReg_reg[30]  ( .D(n189), .CPN(n252), .CDN(n94), .Q(ParOut[30]), .QN(n59) );
  LHCND1 SerClock_reg ( .E(SerValid), .D(SerClk), .CDN(n253), .Q(n252) );
  INVD1 U3 ( .I(Reset), .ZN(n253) );
  INR2XD2 U4 ( .A1(n105), .B1(n106), .ZN(N44) );
  AN4D1 U5 ( .A1(n109), .A2(n110), .A3(n111), .A4(n112), .Z(n105) );
  BUFFD1 U6 ( .I(n92), .Z(n91) );
  BUFFD1 U7 ( .I(n93), .Z(n92) );
  BUFFD1 U8 ( .I(n94), .Z(n93) );
  BUFFD1 U9 ( .I(n253), .Z(n94) );
  BUFFD1 U10 ( .I(n252), .Z(n95) );
  BUFFD1 U11 ( .I(n252), .Z(n96) );
  BUFFD1 U12 ( .I(n252), .Z(n97) );
  MUX2ND0 U13 ( .I0(n255), .I1(n123), .S(N44), .ZN(n251) );
  MUX2ND0 U14 ( .I0(n254), .I1(n124), .S(N44), .ZN(n250) );
  MUX2ND0 U15 ( .I0(n186), .I1(n125), .S(N44), .ZN(n249) );
  MUX2ND0 U16 ( .I0(n185), .I1(n126), .S(N44), .ZN(n248) );
  MUX2ND0 U17 ( .I0(n184), .I1(n127), .S(N44), .ZN(n247) );
  MUX2ND0 U18 ( .I0(n183), .I1(n128), .S(N44), .ZN(n246) );
  MUX2ND0 U19 ( .I0(n182), .I1(n129), .S(N44), .ZN(n245) );
  MUX2ND0 U20 ( .I0(n181), .I1(n130), .S(N44), .ZN(n244) );
  MUX2ND0 U21 ( .I0(n180), .I1(n139), .S(N44), .ZN(n243) );
  MUX2ND0 U22 ( .I0(n179), .I1(n140), .S(N44), .ZN(n242) );
  MUX2ND0 U23 ( .I0(n168), .I1(n141), .S(N44), .ZN(n241) );
  MUX2ND0 U24 ( .I0(n167), .I1(n142), .S(N44), .ZN(n240) );
  MUX2ND0 U25 ( .I0(n166), .I1(n143), .S(N44), .ZN(n239) );
  MUX2ND0 U26 ( .I0(n165), .I1(n144), .S(N44), .ZN(n238) );
  MUX2ND0 U27 ( .I0(n163), .I1(n145), .S(N44), .ZN(n237) );
  MUX2ND0 U28 ( .I0(n154), .I1(n146), .S(N44), .ZN(n236) );
  MUX2ND0 U29 ( .I0(n153), .I1(n155), .S(N44), .ZN(n235) );
  MUX2ND0 U30 ( .I0(n152), .I1(n156), .S(N44), .ZN(n234) );
  MUX2ND0 U31 ( .I0(n151), .I1(n157), .S(N44), .ZN(n233) );
  MUX2ND0 U32 ( .I0(n150), .I1(n158), .S(N44), .ZN(n232) );
  MUX2ND0 U33 ( .I0(n149), .I1(n159), .S(N44), .ZN(n231) );
  MUX2ND0 U34 ( .I0(n138), .I1(n160), .S(N44), .ZN(n230) );
  MUX2ND0 U35 ( .I0(n137), .I1(n161), .S(N44), .ZN(n229) );
  MUX2ND0 U36 ( .I0(n136), .I1(n162), .S(N44), .ZN(n228) );
  MUX2ND0 U37 ( .I0(n135), .I1(n171), .S(N44), .ZN(n227) );
  MUX2ND0 U38 ( .I0(n132), .I1(n172), .S(N44), .ZN(n226) );
  MUX2ND0 U39 ( .I0(n131), .I1(n173), .S(N44), .ZN(n225) );
  MUX2ND0 U40 ( .I0(n122), .I1(n174), .S(N44), .ZN(n224) );
  MUX2ND0 U41 ( .I0(n121), .I1(n175), .S(N44), .ZN(n223) );
  MUX2ND0 U42 ( .I0(n120), .I1(n176), .S(N44), .ZN(n222) );
  MUX2ND0 U43 ( .I0(n119), .I1(n177), .S(N44), .ZN(n221) );
  MUX2ND0 U44 ( .I0(n118), .I1(n178), .S(N44), .ZN(n220) );
  MUX2ND0 U45 ( .I0(n118), .I1(n89), .S(n117), .ZN(n219) );
  MUX2ND0 U46 ( .I0(n119), .I1(n88), .S(n117), .ZN(n218) );
  MUX2ND0 U47 ( .I0(n120), .I1(n87), .S(n117), .ZN(n217) );
  MUX2ND0 U48 ( .I0(n121), .I1(n86), .S(n117), .ZN(n216) );
  MUX2ND0 U49 ( .I0(n122), .I1(n85), .S(n117), .ZN(n215) );
  MUX2ND0 U50 ( .I0(n131), .I1(n84), .S(n117), .ZN(n214) );
  MUX2ND0 U51 ( .I0(n132), .I1(n83), .S(n117), .ZN(n213) );
  MUX2ND0 U52 ( .I0(n135), .I1(n82), .S(n117), .ZN(n212) );
  MUX2ND0 U53 ( .I0(n136), .I1(n81), .S(n117), .ZN(n211) );
  MUX2ND0 U54 ( .I0(n137), .I1(n80), .S(n117), .ZN(n210) );
  MUX2ND0 U55 ( .I0(n138), .I1(n79), .S(n117), .ZN(n209) );
  MUX2ND0 U56 ( .I0(n149), .I1(n78), .S(n117), .ZN(n208) );
  MUX2ND0 U57 ( .I0(n150), .I1(n77), .S(n117), .ZN(n207) );
  MUX2ND0 U58 ( .I0(n151), .I1(n76), .S(n117), .ZN(n206) );
  MUX2ND0 U59 ( .I0(n152), .I1(n75), .S(n117), .ZN(n205) );
  MUX2ND0 U60 ( .I0(n153), .I1(n74), .S(n117), .ZN(n204) );
  MUX2ND0 U61 ( .I0(n154), .I1(n73), .S(n117), .ZN(n203) );
  MUX2ND0 U62 ( .I0(n163), .I1(n72), .S(n117), .ZN(n202) );
  MUX2ND0 U63 ( .I0(n165), .I1(n71), .S(n117), .ZN(n201) );
  MUX2ND0 U64 ( .I0(n166), .I1(n70), .S(n117), .ZN(n200) );
  MUX2ND0 U65 ( .I0(n167), .I1(n69), .S(n117), .ZN(n199) );
  MUX2ND0 U66 ( .I0(n168), .I1(n68), .S(n117), .ZN(n198) );
  MUX2ND0 U67 ( .I0(n179), .I1(n67), .S(n117), .ZN(n197) );
  MUX2ND0 U68 ( .I0(n180), .I1(n66), .S(n117), .ZN(n196) );
  MUX2ND0 U69 ( .I0(n181), .I1(n65), .S(n117), .ZN(n195) );
  MUX2ND0 U70 ( .I0(n182), .I1(n64), .S(n117), .ZN(n194) );
  MUX2ND0 U71 ( .I0(n183), .I1(n63), .S(n117), .ZN(n193) );
  MUX2ND0 U72 ( .I0(n184), .I1(n62), .S(n117), .ZN(n192) );
  MUX2ND0 U73 ( .I0(n185), .I1(n61), .S(n117), .ZN(n191) );
  MUX2ND0 U74 ( .I0(n186), .I1(n60), .S(n117), .ZN(n190) );
  MUX2ND0 U75 ( .I0(n254), .I1(n59), .S(n117), .ZN(n189) );
  MUX2ND0 U76 ( .I0(n255), .I1(n58), .S(n117), .ZN(n188) );
  OAI21D0 U77 ( .A1(n57), .A2(n98), .B(n117), .ZN(n187) );
  CKND0 U78 ( .CLK(ParClk), .CN(n98) );
  INR2D0 U79 ( .A1(N53), .B1(n99), .ZN(N70) );
  CKND2D0 U80 ( .A1(n100), .A2(n92), .ZN(N69) );
  INR2D0 U81 ( .A1(N52), .B1(n99), .ZN(N68) );
  INR2D0 U82 ( .A1(N51), .B1(n99), .ZN(N67) );
  NR2D0 U83 ( .A1(n99), .A2(n101), .ZN(N66) );
  NR2D0 U84 ( .A1(n99), .A2(n102), .ZN(N65) );
  NR2D0 U85 ( .A1(ParClk), .A2(n99), .ZN(N63) );
  IND3D0 U86 ( .A1(n256), .B1(n92), .B2(SerValid), .ZN(n99) );
  OAI21D0 U87 ( .A1(n103), .A2(n100), .B(n92), .ZN(N62) );
  CKND0 U88 ( .CLK(SerValid), .CN(n100) );
  AOI31D0 U89 ( .A1(n102), .A2(n101), .A3(n104), .B(n256), .ZN(n103) );
  NR3D0 U90 ( .A1(N51), .A2(N53), .A3(N52), .ZN(n104) );
  CKND0 U91 ( .CLK(N50), .CN(n101) );
  CKND0 U92 ( .CLK(N49), .CN(n102) );
  NR2D0 U93 ( .A1(n105), .A2(n106), .ZN(N12) );
  CKND2D0 U94 ( .A1(n107), .A2(n108), .ZN(n106) );
  NR4D0 U95 ( .A1(FrameSR[3]), .A2(FrameSR[2]), .A3(FrameSR[1]), .A4(
        FrameSR[0]), .ZN(n108) );
  NR4D0 U96 ( .A1(FrameSR[7]), .A2(FrameSR[6]), .A3(FrameSR[5]), .A4(
        FrameSR[4]), .ZN(n107) );
  NR4D0 U97 ( .A1(n113), .A2(FrameSR[54]), .A3(n134), .A4(FrameSR[55]), .ZN(
        n112) );
  ND3D0 U98 ( .A1(FrameSR[36]), .A2(FrameSR[19]), .A3(FrameSR[51]), .ZN(n113)
         );
  NR4D0 U99 ( .A1(n114), .A2(FrameSR[23]), .A3(FrameSR[37]), .A4(FrameSR[32]), 
        .ZN(n111) );
  ND3D0 U100 ( .A1(n147), .A2(n133), .A3(n148), .ZN(n114) );
  NR4D0 U101 ( .A1(n115), .A2(FrameSR[20]), .A3(FrameSR[18]), .A4(FrameSR[21]), 
        .ZN(n110) );
  ND3D0 U102 ( .A1(n169), .A2(n164), .A3(n170), .ZN(n115) );
  NR4D0 U103 ( .A1(n116), .A2(FrameSR[49]), .A3(FrameSR[48]), .A4(FrameSR[50]), 
        .ZN(n109) );
  ND3D0 U104 ( .A1(n258), .A2(n259), .A3(n257), .ZN(n116) );
endmodule


module SerialRx ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;


  PLLTop PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(Reset) );
  BUFFD0 U1 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, Clk, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, Clk, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, \CurState[1] , N72, N73, N74,
         N75, N76, N88, N89, N90, N91, N92, N105, N106, N107, N108, N109, N122,
         N123, N124, N125, N126, N142, N144, N146, N148, N150, N153, N156,
         N159, N162, N165, N167, N170, N173, N176, N179, N182, N184, N185,
         N188, N189, N198, N199, N200, N209, N210, N211, N212, N215, N218,
         N221, N224, N227, N230, N233, N236, N239, \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71;
  wire   [2:0] NextState;

  LHQD1 \WriteCount_tri_enable_reg[0]  ( .E(N198), .D(N199), .Q(N9) );
  LHQD1 \ReadCount_reg[0]  ( .E(N209), .D(N167), .Q(N224) );
  LHQD1 \WriteCount_reg[4]  ( .E(N198), .D(N162), .Q(N227) );
  LHQD1 \ReadCount_reg[4]  ( .E(N209), .D(N179), .Q(N212) );
  LHQD1 \NextState_reg[1]  ( .E(N188), .D(N144), .Q(NextState[1]) );
  LHQD1 \NextState_reg[0]  ( .E(N188), .D(N142), .Q(NextState[0]) );
  LHQD1 \NextState_reg[2]  ( .E(N188), .D(N146), .Q(NextState[2]) );
  LHQD1 EmptyFIFOReg_reg ( .E(N211), .D(N182), .Q(EmptyFIFO) );
  LHQD1 \ReadCount_tri_enable_reg[4]  ( .E(N209), .D(N210), .Q(N0) );
  LHQD1 \ReadCount_tri_enable_reg[2]  ( .E(N209), .D(N210), .Q(N2) );
  LHQD1 \ReadCount_tri_enable_reg[0]  ( .E(N209), .D(N210), .Q(N4) );
  LHQD1 \ReadCount_tri_enable_reg[1]  ( .E(N209), .D(N210), .Q(N3) );
  LHQD1 \ReadCount_tri_enable_reg[3]  ( .E(N209), .D(N210), .Q(N1) );
  LHQD1 \WriteCount_tri_enable_reg[4]  ( .E(N198), .D(N199), .Q(N5) );
  LHQD1 \WriteCount_tri_enable_reg[2]  ( .E(N198), .D(N199), .Q(N7) );
  LHQD1 \WriteCount_tri_enable_reg[1]  ( .E(N198), .D(N199), .Q(N8) );
  LHQD1 \WriteCount_tri_enable_reg[3]  ( .E(N198), .D(N199), .Q(N6) );
  LHQD1 FullFIFOReg_reg ( .E(N189), .D(N148), .Q(FullFIFO) );
  LHQD1 ReadCmdReg_reg ( .E(N185), .D(N184), .Q(ReadCmd) );
  LHQD1 WriteCmdReg_reg ( .E(N200), .D(N165), .Q(WriteCmd) );
  LHQD1 \ReadCount_reg[1]  ( .E(N209), .D(N170), .Q(N221) );
  LHQD1 \WriteCount_reg[1]  ( .E(N198), .D(N153), .Q(N236) );
  LHQD1 \WriteCount_reg[2]  ( .E(N198), .D(N156), .Q(N233) );
  LHQD1 \ReadCount_reg[2]  ( .E(N209), .D(N173), .Q(N218) );
  LHQD1 \WriteCount_reg[3]  ( .E(N198), .D(N159), .Q(N230) );
  LHQD1 \ReadCount_reg[3]  ( .E(N209), .D(N176), .Q(N215) );
  LHQD1 \WriteCount_reg[0]  ( .E(N198), .D(N150), .Q(N239) );
  BUFTD1 \WriteCount_tri[0]  ( .I(N239), .OE(n92), .Z(WriteAddr[0]) );
  BUFTD1 \WriteCount_tri[1]  ( .I(N236), .OE(n91), .Z(WriteAddr[1]) );
  BUFTD1 \WriteCount_tri[2]  ( .I(N233), .OE(n90), .Z(WriteAddr[2]) );
  BUFTD1 \WriteCount_tri[3]  ( .I(N230), .OE(n89), .Z(WriteAddr[3]) );
  BUFTD1 \WriteCount_tri[4]  ( .I(N227), .OE(n88), .Z(WriteAddr[4]) );
  BUFTD1 \ReadCount_tri[0]  ( .I(N224), .OE(n87), .Z(ReadAddr[0]) );
  BUFTD1 \ReadCount_tri[1]  ( .I(N221), .OE(n86), .Z(ReadAddr[1]) );
  BUFTD1 \ReadCount_tri[2]  ( .I(N218), .OE(n85), .Z(ReadAddr[2]) );
  BUFTD1 \ReadCount_tri[3]  ( .I(N215), .OE(n84), .Z(ReadAddr[3]) );
  BUFTD1 \ReadCount_tri[4]  ( .I(N212), .OE(n83), .Z(ReadAddr[4]) );
  FIFOStateM_AWid5_DW01_inc_0 add_183 ( .A({N76, N75, N74, N73, N72}), .SUM({
        N92, N91, N90, N89, N88}) );
  FIFOStateM_AWid5_DW01_inc_1 r147 ( .A(WriteAddr), .SUM({N76, N75, N74, N73, 
        N72}) );
  FIFOStateM_AWid5_DW01_inc_2 add_196 ( .A({N126, N125, N124, N123, N122}), 
        .SUM({N109, N108, N107, N106, N105}) );
  FIFOStateM_AWid5_DW01_inc_3 r133 ( .A({\U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , 
        \U3/U1/Z_1 , \U3/U1/Z_0 }), .SUM({N126, N125, N124, N123, N122}) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(Clk), .CDN(n93), .Q(
        \CurState[1] ) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(Clk), .CDN(n93), .Q(n70) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(Clk), .CDN(n93), .Q(n71) );
  AOI21D1 U3 ( .A1(n16), .A2(n19), .B(Clk), .ZN(N198) );
  AOI21D1 U4 ( .A1(n12), .A2(n22), .B(Clk), .ZN(N209) );
  CKND0 U5 ( .CLK(N9), .CN(n92) );
  CKND0 U6 ( .CLK(N8), .CN(n91) );
  CKND0 U7 ( .CLK(N7), .CN(n90) );
  CKND0 U8 ( .CLK(N6), .CN(n89) );
  CKND0 U9 ( .CLK(N5), .CN(n88) );
  CKND0 U10 ( .CLK(N4), .CN(n87) );
  CKND0 U11 ( .CLK(N3), .CN(n86) );
  CKND0 U12 ( .CLK(N2), .CN(n85) );
  CKND0 U13 ( .CLK(N1), .CN(n84) );
  CKND0 U14 ( .CLK(N0), .CN(n83) );
  IOA22D0 U15 ( .B1(n3), .B2(n4), .A1(n5), .A2(ReadAddr[4]), .ZN(\U3/U1/Z_4 )
         );
  IOA22D0 U16 ( .B1(n3), .B2(n6), .A1(n5), .A2(ReadAddr[3]), .ZN(\U3/U1/Z_3 )
         );
  IOA22D0 U17 ( .B1(n3), .B2(n7), .A1(n5), .A2(ReadAddr[2]), .ZN(\U3/U1/Z_2 )
         );
  IOA22D0 U18 ( .B1(n3), .B2(n8), .A1(n5), .A2(ReadAddr[1]), .ZN(\U3/U1/Z_1 )
         );
  IOA22D0 U19 ( .B1(n3), .B2(n9), .A1(n5), .A2(ReadAddr[0]), .ZN(\U3/U1/Z_0 )
         );
  CKND2D0 U20 ( .A1(n10), .A2(n93), .ZN(n3) );
  AOI21D0 U21 ( .A1(n11), .A2(n12), .B(Clk), .ZN(N211) );
  AN2D0 U22 ( .A1(N182), .A2(n13), .Z(N210) );
  AOI31D0 U23 ( .A1(n14), .A2(n15), .A3(n16), .B(Clk), .ZN(N200) );
  CKND0 U24 ( .CLK(N184), .CN(n15) );
  CKND2D0 U25 ( .A1(n17), .A2(n18), .ZN(n14) );
  AN2D0 U26 ( .A1(N148), .A2(n13), .Z(N199) );
  AOI21D0 U27 ( .A1(n20), .A2(n21), .B(Clk), .ZN(N189) );
  AOI31D0 U28 ( .A1(n16), .A2(n22), .A3(n23), .B(Clk), .ZN(N188) );
  NR2D0 U29 ( .A1(n24), .A2(n25), .ZN(n23) );
  MUX2ND0 U30 ( .I0(n26), .I1(n71), .S(n70), .ZN(n25) );
  CKND2D0 U31 ( .A1(n71), .A2(n27), .ZN(n26) );
  INR3D0 U32 ( .A1(n21), .B1(n28), .B2(n10), .ZN(n16) );
  CKND2D0 U33 ( .A1(n29), .A2(Reset), .ZN(n21) );
  IND2D0 U34 ( .A1(N209), .B1(n30), .ZN(N185) );
  OAI21D0 U35 ( .A1(n28), .A2(n24), .B(n13), .ZN(n30) );
  CKND0 U36 ( .CLK(Clk), .CN(n13) );
  OAI22D0 U37 ( .A1(n31), .A2(n11), .B1(n32), .B2(n33), .ZN(n24) );
  NR2D0 U38 ( .A1(n32), .A2(n34), .ZN(n28) );
  CKND0 U39 ( .CLK(n5), .CN(n22) );
  OAI211D0 U40 ( .A1(n31), .A2(n19), .B(n35), .C(n36), .ZN(n5) );
  ND3D0 U41 ( .A1(n36), .A2(n19), .A3(n37), .ZN(N184) );
  OA21D0 U42 ( .A1(n11), .A2(n31), .B(n35), .Z(n37) );
  CKND2D0 U43 ( .A1(n17), .A2(n38), .ZN(n35) );
  CKND0 U44 ( .CLK(n39), .CN(n11) );
  NR2D0 U45 ( .A1(n12), .A2(n18), .ZN(N182) );
  CKND0 U46 ( .CLK(n32), .CN(n18) );
  OAI22D0 U47 ( .A1(n40), .A2(n41), .B1(n4), .B2(n42), .ZN(N179) );
  CKND0 U48 ( .CLK(N126), .CN(n41) );
  OAI22D0 U49 ( .A1(n40), .A2(n43), .B1(n6), .B2(n42), .ZN(N176) );
  CKND0 U50 ( .CLK(N125), .CN(n43) );
  OAI22D0 U51 ( .A1(n40), .A2(n44), .B1(n7), .B2(n42), .ZN(N173) );
  CKND0 U52 ( .CLK(WriteAddr[2]), .CN(n7) );
  CKND0 U53 ( .CLK(N124), .CN(n44) );
  OAI22D0 U54 ( .A1(n40), .A2(n45), .B1(n8), .B2(n42), .ZN(N170) );
  CKND0 U55 ( .CLK(WriteAddr[1]), .CN(n8) );
  CKND0 U56 ( .CLK(N123), .CN(n45) );
  OAI22D0 U57 ( .A1(n40), .A2(n46), .B1(n9), .B2(n42), .ZN(N167) );
  CKND2D0 U58 ( .A1(n29), .A2(n93), .ZN(n42) );
  CKND0 U59 ( .CLK(Reset), .CN(n93) );
  CKND0 U60 ( .CLK(WriteAddr[0]), .CN(n9) );
  CKND0 U61 ( .CLK(N122), .CN(n46) );
  INR2D0 U62 ( .A1(n20), .B1(n47), .ZN(n40) );
  OAI21D0 U63 ( .A1(n38), .A2(n48), .B(n49), .ZN(N165) );
  NR2D0 U64 ( .A1(n17), .A2(n50), .ZN(n48) );
  AO222D0 U65 ( .A1(ReadAddr[4]), .A2(n51), .B1(N126), .B2(n10), .C1(N76), 
        .C2(n50), .Z(N162) );
  AO222D0 U66 ( .A1(ReadAddr[3]), .A2(n51), .B1(N125), .B2(n10), .C1(N75), 
        .C2(n50), .Z(N159) );
  AO222D0 U67 ( .A1(ReadAddr[2]), .A2(n51), .B1(N124), .B2(n10), .C1(N74), 
        .C2(n50), .Z(N156) );
  AO222D0 U68 ( .A1(ReadAddr[1]), .A2(n51), .B1(N123), .B2(n10), .C1(N73), 
        .C2(n50), .Z(N153) );
  AO222D0 U69 ( .A1(ReadAddr[0]), .A2(n51), .B1(N122), .B2(n10), .C1(N72), 
        .C2(n50), .Z(N150) );
  CKND0 U70 ( .CLK(n34), .CN(n50) );
  NR2D0 U71 ( .A1(n19), .A2(n38), .ZN(N148) );
  OAI21D0 U72 ( .A1(n38), .A2(n52), .B(n19), .ZN(N146) );
  AOI21D0 U73 ( .A1(n53), .A2(n47), .B(n17), .ZN(n52) );
  CKND0 U74 ( .CLK(n54), .CN(n53) );
  ND4D0 U75 ( .A1(n36), .A2(n33), .A3(n49), .A4(n55), .ZN(N144) );
  AOI22D0 U76 ( .A1(n47), .A2(n54), .B1(n39), .B2(n31), .ZN(n55) );
  CKND0 U77 ( .CLK(n38), .CN(n31) );
  ND3D0 U78 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n54) );
  NR3D0 U79 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n58) );
  CKXOR2D0 U80 ( .A1(ReadAddr[3]), .A2(N91), .Z(n61) );
  CKXOR2D0 U81 ( .A1(ReadAddr[1]), .A2(N89), .Z(n60) );
  CKXOR2D0 U82 ( .A1(ReadAddr[0]), .A2(N88), .Z(n59) );
  XNR2D0 U83 ( .A1(N90), .A2(ReadAddr[2]), .ZN(n57) );
  XNR2D0 U84 ( .A1(N92), .A2(ReadAddr[4]), .ZN(n56) );
  CKND0 U85 ( .CLK(n10), .CN(n49) );
  NR2D0 U86 ( .A1(n32), .A2(n12), .ZN(n10) );
  CKND0 U87 ( .CLK(n29), .CN(n12) );
  NR3D0 U88 ( .A1(n71), .A2(n70), .A3(\CurState[1] ), .ZN(n29) );
  CKND2D0 U89 ( .A1(WriteReq), .A2(n62), .ZN(n32) );
  CKND2D0 U90 ( .A1(n38), .A2(n47), .ZN(n36) );
  OAI211D0 U91 ( .A1(n38), .A2(n34), .B(n63), .C(n20), .ZN(N142) );
  NR2D0 U92 ( .A1(n51), .A2(n17), .ZN(n20) );
  CKND0 U93 ( .CLK(n33), .CN(n17) );
  ND3D0 U94 ( .A1(n71), .A2(n27), .A3(n70), .ZN(n33) );
  CKND0 U95 ( .CLK(n19), .CN(n51) );
  ND3D0 U96 ( .A1(n71), .A2(\CurState[1] ), .A3(n70), .ZN(n19) );
  OAI31D0 U97 ( .A1(n64), .A2(n65), .A3(n66), .B(n47), .ZN(n63) );
  XNR2D0 U98 ( .A1(n4), .A2(N109), .ZN(n66) );
  CKND0 U99 ( .CLK(WriteAddr[4]), .CN(n4) );
  XNR2D0 U100 ( .A1(n6), .A2(N108), .ZN(n65) );
  CKND0 U101 ( .CLK(WriteAddr[3]), .CN(n6) );
  ND3D0 U102 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n64) );
  XNR2D0 U103 ( .A1(N106), .A2(WriteAddr[1]), .ZN(n69) );
  XNR2D0 U104 ( .A1(N107), .A2(WriteAddr[2]), .ZN(n68) );
  XNR2D0 U105 ( .A1(N105), .A2(WriteAddr[0]), .ZN(n67) );
  NR2D0 U106 ( .A1(n39), .A2(n47), .ZN(n34) );
  INR3D0 U107 ( .A1(n71), .B1(n27), .B2(n70), .ZN(n47) );
  NR3D0 U108 ( .A1(n71), .A2(n70), .A3(n27), .ZN(n39) );
  CKND0 U109 ( .CLK(\CurState[1] ), .CN(n27) );
  NR2D0 U110 ( .A1(n62), .A2(WriteReq), .ZN(n38) );
  CKND0 U111 ( .CLK(ReadReq), .CN(n62) );
endmodule


module Mem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, Addr, ClockIn, 
        ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] Addr;
  input ClockIn, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N75, N76, N77, N78, N79, ChipClock, DreadyReg,
         \Storage[31][32] , \Storage[31][31] , \Storage[31][30] ,
         \Storage[31][29] , \Storage[31][28] , \Storage[31][27] ,
         \Storage[31][26] , \Storage[31][25] , \Storage[31][24] ,
         \Storage[31][23] , \Storage[31][22] , \Storage[31][21] ,
         \Storage[31][20] , \Storage[31][19] , \Storage[31][18] ,
         \Storage[31][17] , \Storage[31][16] , \Storage[31][15] ,
         \Storage[31][14] , \Storage[31][13] , \Storage[31][12] ,
         \Storage[31][11] , \Storage[31][10] , \Storage[31][9] ,
         \Storage[31][8] , \Storage[31][7] , \Storage[31][6] ,
         \Storage[31][5] , \Storage[31][4] , \Storage[31][3] ,
         \Storage[31][2] , \Storage[31][1] , \Storage[31][0] ,
         \Storage[30][32] , \Storage[30][31] , \Storage[30][30] ,
         \Storage[30][29] , \Storage[30][28] , \Storage[30][27] ,
         \Storage[30][26] , \Storage[30][25] , \Storage[30][24] ,
         \Storage[30][23] , \Storage[30][22] , \Storage[30][21] ,
         \Storage[30][20] , \Storage[30][19] , \Storage[30][18] ,
         \Storage[30][17] , \Storage[30][16] , \Storage[30][15] ,
         \Storage[30][14] , \Storage[30][13] , \Storage[30][12] ,
         \Storage[30][11] , \Storage[30][10] , \Storage[30][9] ,
         \Storage[30][8] , \Storage[30][7] , \Storage[30][6] ,
         \Storage[30][5] , \Storage[30][4] , \Storage[30][3] ,
         \Storage[30][2] , \Storage[30][1] , \Storage[30][0] ,
         \Storage[29][32] , \Storage[29][31] , \Storage[29][30] ,
         \Storage[29][29] , \Storage[29][28] , \Storage[29][27] ,
         \Storage[29][26] , \Storage[29][25] , \Storage[29][24] ,
         \Storage[29][23] , \Storage[29][22] , \Storage[29][21] ,
         \Storage[29][20] , \Storage[29][19] , \Storage[29][18] ,
         \Storage[29][17] , \Storage[29][16] , \Storage[29][15] ,
         \Storage[29][14] , \Storage[29][13] , \Storage[29][12] ,
         \Storage[29][11] , \Storage[29][10] , \Storage[29][9] ,
         \Storage[29][8] , \Storage[29][7] , \Storage[29][6] ,
         \Storage[29][5] , \Storage[29][4] , \Storage[29][3] ,
         \Storage[29][2] , \Storage[29][1] , \Storage[29][0] ,
         \Storage[28][32] , \Storage[28][31] , \Storage[28][30] ,
         \Storage[28][29] , \Storage[28][28] , \Storage[28][27] ,
         \Storage[28][26] , \Storage[28][25] , \Storage[28][24] ,
         \Storage[28][23] , \Storage[28][22] , \Storage[28][21] ,
         \Storage[28][20] , \Storage[28][19] , \Storage[28][18] ,
         \Storage[28][17] , \Storage[28][16] , \Storage[28][15] ,
         \Storage[28][14] , \Storage[28][13] , \Storage[28][12] ,
         \Storage[28][11] , \Storage[28][10] , \Storage[28][9] ,
         \Storage[28][8] , \Storage[28][7] , \Storage[28][6] ,
         \Storage[28][5] , \Storage[28][4] , \Storage[28][3] ,
         \Storage[28][2] , \Storage[28][1] , \Storage[28][0] ,
         \Storage[27][32] , \Storage[27][31] , \Storage[27][30] ,
         \Storage[27][29] , \Storage[27][28] , \Storage[27][27] ,
         \Storage[27][26] , \Storage[27][25] , \Storage[27][24] ,
         \Storage[27][23] , \Storage[27][22] , \Storage[27][21] ,
         \Storage[27][20] , \Storage[27][19] , \Storage[27][18] ,
         \Storage[27][17] , \Storage[27][16] , \Storage[27][15] ,
         \Storage[27][14] , \Storage[27][13] , \Storage[27][12] ,
         \Storage[27][11] , \Storage[27][10] , \Storage[27][9] ,
         \Storage[27][8] , \Storage[27][7] , \Storage[27][6] ,
         \Storage[27][5] , \Storage[27][4] , \Storage[27][3] ,
         \Storage[27][2] , \Storage[27][1] , \Storage[27][0] ,
         \Storage[26][32] , \Storage[26][31] , \Storage[26][30] ,
         \Storage[26][29] , \Storage[26][28] , \Storage[26][27] ,
         \Storage[26][26] , \Storage[26][25] , \Storage[26][24] ,
         \Storage[26][23] , \Storage[26][22] , \Storage[26][21] ,
         \Storage[26][20] , \Storage[26][19] , \Storage[26][18] ,
         \Storage[26][17] , \Storage[26][16] , \Storage[26][15] ,
         \Storage[26][14] , \Storage[26][13] , \Storage[26][12] ,
         \Storage[26][11] , \Storage[26][10] , \Storage[26][9] ,
         \Storage[26][8] , \Storage[26][7] , \Storage[26][6] ,
         \Storage[26][5] , \Storage[26][4] , \Storage[26][3] ,
         \Storage[26][2] , \Storage[26][1] , \Storage[26][0] ,
         \Storage[25][32] , \Storage[25][31] , \Storage[25][30] ,
         \Storage[25][29] , \Storage[25][28] , \Storage[25][27] ,
         \Storage[25][26] , \Storage[25][25] , \Storage[25][24] ,
         \Storage[25][23] , \Storage[25][22] , \Storage[25][21] ,
         \Storage[25][20] , \Storage[25][19] , \Storage[25][18] ,
         \Storage[25][17] , \Storage[25][16] , \Storage[25][15] ,
         \Storage[25][14] , \Storage[25][13] , \Storage[25][12] ,
         \Storage[25][11] , \Storage[25][10] , \Storage[25][9] ,
         \Storage[25][8] , \Storage[25][7] , \Storage[25][6] ,
         \Storage[25][5] , \Storage[25][4] , \Storage[25][3] ,
         \Storage[25][2] , \Storage[25][1] , \Storage[25][0] ,
         \Storage[24][32] , \Storage[24][31] , \Storage[24][30] ,
         \Storage[24][29] , \Storage[24][28] , \Storage[24][27] ,
         \Storage[24][26] , \Storage[24][25] , \Storage[24][24] ,
         \Storage[24][23] , \Storage[24][22] , \Storage[24][21] ,
         \Storage[24][20] , \Storage[24][19] , \Storage[24][18] ,
         \Storage[24][17] , \Storage[24][16] , \Storage[24][15] ,
         \Storage[24][14] , \Storage[24][13] , \Storage[24][12] ,
         \Storage[24][11] , \Storage[24][10] , \Storage[24][9] ,
         \Storage[24][8] , \Storage[24][7] , \Storage[24][6] ,
         \Storage[24][5] , \Storage[24][4] , \Storage[24][3] ,
         \Storage[24][2] , \Storage[24][1] , \Storage[24][0] ,
         \Storage[23][32] , \Storage[23][31] , \Storage[23][30] ,
         \Storage[23][29] , \Storage[23][28] , \Storage[23][27] ,
         \Storage[23][26] , \Storage[23][25] , \Storage[23][24] ,
         \Storage[23][23] , \Storage[23][22] , \Storage[23][21] ,
         \Storage[23][20] , \Storage[23][19] , \Storage[23][18] ,
         \Storage[23][17] , \Storage[23][16] , \Storage[23][15] ,
         \Storage[23][14] , \Storage[23][13] , \Storage[23][12] ,
         \Storage[23][11] , \Storage[23][10] , \Storage[23][9] ,
         \Storage[23][8] , \Storage[23][7] , \Storage[23][6] ,
         \Storage[23][5] , \Storage[23][4] , \Storage[23][3] ,
         \Storage[23][2] , \Storage[23][1] , \Storage[23][0] ,
         \Storage[22][32] , \Storage[22][31] , \Storage[22][30] ,
         \Storage[22][29] , \Storage[22][28] , \Storage[22][27] ,
         \Storage[22][26] , \Storage[22][25] , \Storage[22][24] ,
         \Storage[22][23] , \Storage[22][22] , \Storage[22][21] ,
         \Storage[22][20] , \Storage[22][19] , \Storage[22][18] ,
         \Storage[22][17] , \Storage[22][16] , \Storage[22][15] ,
         \Storage[22][14] , \Storage[22][13] , \Storage[22][12] ,
         \Storage[22][11] , \Storage[22][10] , \Storage[22][9] ,
         \Storage[22][8] , \Storage[22][7] , \Storage[22][6] ,
         \Storage[22][5] , \Storage[22][4] , \Storage[22][3] ,
         \Storage[22][2] , \Storage[22][1] , \Storage[22][0] ,
         \Storage[21][32] , \Storage[21][31] , \Storage[21][30] ,
         \Storage[21][29] , \Storage[21][28] , \Storage[21][27] ,
         \Storage[21][26] , \Storage[21][25] , \Storage[21][24] ,
         \Storage[21][23] , \Storage[21][22] , \Storage[21][21] ,
         \Storage[21][20] , \Storage[21][19] , \Storage[21][18] ,
         \Storage[21][17] , \Storage[21][16] , \Storage[21][15] ,
         \Storage[21][14] , \Storage[21][13] , \Storage[21][12] ,
         \Storage[21][11] , \Storage[21][10] , \Storage[21][9] ,
         \Storage[21][8] , \Storage[21][7] , \Storage[21][6] ,
         \Storage[21][5] , \Storage[21][4] , \Storage[21][3] ,
         \Storage[21][2] , \Storage[21][1] , \Storage[21][0] ,
         \Storage[20][32] , \Storage[20][31] , \Storage[20][30] ,
         \Storage[20][29] , \Storage[20][28] , \Storage[20][27] ,
         \Storage[20][26] , \Storage[20][25] , \Storage[20][24] ,
         \Storage[20][23] , \Storage[20][22] , \Storage[20][21] ,
         \Storage[20][20] , \Storage[20][19] , \Storage[20][18] ,
         \Storage[20][17] , \Storage[20][16] , \Storage[20][15] ,
         \Storage[20][14] , \Storage[20][13] , \Storage[20][12] ,
         \Storage[20][11] , \Storage[20][10] , \Storage[20][9] ,
         \Storage[20][8] , \Storage[20][7] , \Storage[20][6] ,
         \Storage[20][5] , \Storage[20][4] , \Storage[20][3] ,
         \Storage[20][2] , \Storage[20][1] , \Storage[20][0] ,
         \Storage[19][32] , \Storage[19][31] , \Storage[19][30] ,
         \Storage[19][29] , \Storage[19][28] , \Storage[19][27] ,
         \Storage[19][26] , \Storage[19][25] , \Storage[19][24] ,
         \Storage[19][23] , \Storage[19][22] , \Storage[19][21] ,
         \Storage[19][20] , \Storage[19][19] , \Storage[19][18] ,
         \Storage[19][17] , \Storage[19][16] , \Storage[19][15] ,
         \Storage[19][14] , \Storage[19][13] , \Storage[19][12] ,
         \Storage[19][11] , \Storage[19][10] , \Storage[19][9] ,
         \Storage[19][8] , \Storage[19][7] , \Storage[19][6] ,
         \Storage[19][5] , \Storage[19][4] , \Storage[19][3] ,
         \Storage[19][2] , \Storage[19][1] , \Storage[19][0] ,
         \Storage[18][32] , \Storage[18][31] , \Storage[18][30] ,
         \Storage[18][29] , \Storage[18][28] , \Storage[18][27] ,
         \Storage[18][26] , \Storage[18][25] , \Storage[18][24] ,
         \Storage[18][23] , \Storage[18][22] , \Storage[18][21] ,
         \Storage[18][20] , \Storage[18][19] , \Storage[18][18] ,
         \Storage[18][17] , \Storage[18][16] , \Storage[18][15] ,
         \Storage[18][14] , \Storage[18][13] , \Storage[18][12] ,
         \Storage[18][11] , \Storage[18][10] , \Storage[18][9] ,
         \Storage[18][8] , \Storage[18][7] , \Storage[18][6] ,
         \Storage[18][5] , \Storage[18][4] , \Storage[18][3] ,
         \Storage[18][2] , \Storage[18][1] , \Storage[18][0] ,
         \Storage[17][32] , \Storage[17][31] , \Storage[17][30] ,
         \Storage[17][29] , \Storage[17][28] , \Storage[17][27] ,
         \Storage[17][26] , \Storage[17][25] , \Storage[17][24] ,
         \Storage[17][23] , \Storage[17][22] , \Storage[17][21] ,
         \Storage[17][20] , \Storage[17][19] , \Storage[17][18] ,
         \Storage[17][17] , \Storage[17][16] , \Storage[17][15] ,
         \Storage[17][14] , \Storage[17][13] , \Storage[17][12] ,
         \Storage[17][11] , \Storage[17][10] , \Storage[17][9] ,
         \Storage[17][8] , \Storage[17][7] , \Storage[17][6] ,
         \Storage[17][5] , \Storage[17][4] , \Storage[17][3] ,
         \Storage[17][2] , \Storage[17][1] , \Storage[17][0] ,
         \Storage[16][32] , \Storage[16][31] , \Storage[16][30] ,
         \Storage[16][29] , \Storage[16][28] , \Storage[16][27] ,
         \Storage[16][26] , \Storage[16][25] , \Storage[16][24] ,
         \Storage[16][23] , \Storage[16][22] , \Storage[16][21] ,
         \Storage[16][20] , \Storage[16][19] , \Storage[16][18] ,
         \Storage[16][17] , \Storage[16][16] , \Storage[16][15] ,
         \Storage[16][14] , \Storage[16][13] , \Storage[16][12] ,
         \Storage[16][11] , \Storage[16][10] , \Storage[16][9] ,
         \Storage[16][8] , \Storage[16][7] , \Storage[16][6] ,
         \Storage[16][5] , \Storage[16][4] , \Storage[16][3] ,
         \Storage[16][2] , \Storage[16][1] , \Storage[16][0] ,
         \Storage[15][32] , \Storage[15][31] , \Storage[15][30] ,
         \Storage[15][29] , \Storage[15][28] , \Storage[15][27] ,
         \Storage[15][26] , \Storage[15][25] , \Storage[15][24] ,
         \Storage[15][23] , \Storage[15][22] , \Storage[15][21] ,
         \Storage[15][20] , \Storage[15][19] , \Storage[15][18] ,
         \Storage[15][17] , \Storage[15][16] , \Storage[15][15] ,
         \Storage[15][14] , \Storage[15][13] , \Storage[15][12] ,
         \Storage[15][11] , \Storage[15][10] , \Storage[15][9] ,
         \Storage[15][8] , \Storage[15][7] , \Storage[15][6] ,
         \Storage[15][5] , \Storage[15][4] , \Storage[15][3] ,
         \Storage[15][2] , \Storage[15][1] , \Storage[15][0] ,
         \Storage[14][32] , \Storage[14][31] , \Storage[14][30] ,
         \Storage[14][29] , \Storage[14][28] , \Storage[14][27] ,
         \Storage[14][26] , \Storage[14][25] , \Storage[14][24] ,
         \Storage[14][23] , \Storage[14][22] , \Storage[14][21] ,
         \Storage[14][20] , \Storage[14][19] , \Storage[14][18] ,
         \Storage[14][17] , \Storage[14][16] , \Storage[14][15] ,
         \Storage[14][14] , \Storage[14][13] , \Storage[14][12] ,
         \Storage[14][11] , \Storage[14][10] , \Storage[14][9] ,
         \Storage[14][8] , \Storage[14][7] , \Storage[14][6] ,
         \Storage[14][5] , \Storage[14][4] , \Storage[14][3] ,
         \Storage[14][2] , \Storage[14][1] , \Storage[14][0] ,
         \Storage[13][32] , \Storage[13][31] , \Storage[13][30] ,
         \Storage[13][29] , \Storage[13][28] , \Storage[13][27] ,
         \Storage[13][26] , \Storage[13][25] , \Storage[13][24] ,
         \Storage[13][23] , \Storage[13][22] , \Storage[13][21] ,
         \Storage[13][20] , \Storage[13][19] , \Storage[13][18] ,
         \Storage[13][17] , \Storage[13][16] , \Storage[13][15] ,
         \Storage[13][14] , \Storage[13][13] , \Storage[13][12] ,
         \Storage[13][11] , \Storage[13][10] , \Storage[13][9] ,
         \Storage[13][8] , \Storage[13][7] , \Storage[13][6] ,
         \Storage[13][5] , \Storage[13][4] , \Storage[13][3] ,
         \Storage[13][2] , \Storage[13][1] , \Storage[13][0] ,
         \Storage[12][32] , \Storage[12][31] , \Storage[12][30] ,
         \Storage[12][29] , \Storage[12][28] , \Storage[12][27] ,
         \Storage[12][26] , \Storage[12][25] , \Storage[12][24] ,
         \Storage[12][23] , \Storage[12][22] , \Storage[12][21] ,
         \Storage[12][20] , \Storage[12][19] , \Storage[12][18] ,
         \Storage[12][17] , \Storage[12][16] , \Storage[12][15] ,
         \Storage[12][14] , \Storage[12][13] , \Storage[12][12] ,
         \Storage[12][11] , \Storage[12][10] , \Storage[12][9] ,
         \Storage[12][8] , \Storage[12][7] , \Storage[12][6] ,
         \Storage[12][5] , \Storage[12][4] , \Storage[12][3] ,
         \Storage[12][2] , \Storage[12][1] , \Storage[12][0] ,
         \Storage[11][32] , \Storage[11][31] , \Storage[11][30] ,
         \Storage[11][29] , \Storage[11][28] , \Storage[11][27] ,
         \Storage[11][26] , \Storage[11][25] , \Storage[11][24] ,
         \Storage[11][23] , \Storage[11][22] , \Storage[11][21] ,
         \Storage[11][20] , \Storage[11][19] , \Storage[11][18] ,
         \Storage[11][17] , \Storage[11][16] , \Storage[11][15] ,
         \Storage[11][14] , \Storage[11][13] , \Storage[11][12] ,
         \Storage[11][11] , \Storage[11][10] , \Storage[11][9] ,
         \Storage[11][8] , \Storage[11][7] , \Storage[11][6] ,
         \Storage[11][5] , \Storage[11][4] , \Storage[11][3] ,
         \Storage[11][2] , \Storage[11][1] , \Storage[11][0] ,
         \Storage[10][32] , \Storage[10][31] , \Storage[10][30] ,
         \Storage[10][29] , \Storage[10][28] , \Storage[10][27] ,
         \Storage[10][26] , \Storage[10][25] , \Storage[10][24] ,
         \Storage[10][23] , \Storage[10][22] , \Storage[10][21] ,
         \Storage[10][20] , \Storage[10][19] , \Storage[10][18] ,
         \Storage[10][17] , \Storage[10][16] , \Storage[10][15] ,
         \Storage[10][14] , \Storage[10][13] , \Storage[10][12] ,
         \Storage[10][11] , \Storage[10][10] , \Storage[10][9] ,
         \Storage[10][8] , \Storage[10][7] , \Storage[10][6] ,
         \Storage[10][5] , \Storage[10][4] , \Storage[10][3] ,
         \Storage[10][2] , \Storage[10][1] , \Storage[10][0] ,
         \Storage[9][32] , \Storage[9][31] , \Storage[9][30] ,
         \Storage[9][29] , \Storage[9][28] , \Storage[9][27] ,
         \Storage[9][26] , \Storage[9][25] , \Storage[9][24] ,
         \Storage[9][23] , \Storage[9][22] , \Storage[9][21] ,
         \Storage[9][20] , \Storage[9][19] , \Storage[9][18] ,
         \Storage[9][17] , \Storage[9][16] , \Storage[9][15] ,
         \Storage[9][14] , \Storage[9][13] , \Storage[9][12] ,
         \Storage[9][11] , \Storage[9][10] , \Storage[9][9] , \Storage[9][8] ,
         \Storage[9][7] , \Storage[9][6] , \Storage[9][5] , \Storage[9][4] ,
         \Storage[9][3] , \Storage[9][2] , \Storage[9][1] , \Storage[9][0] ,
         \Storage[8][32] , \Storage[8][31] , \Storage[8][30] ,
         \Storage[8][29] , \Storage[8][28] , \Storage[8][27] ,
         \Storage[8][26] , \Storage[8][25] , \Storage[8][24] ,
         \Storage[8][23] , \Storage[8][22] , \Storage[8][21] ,
         \Storage[8][20] , \Storage[8][19] , \Storage[8][18] ,
         \Storage[8][17] , \Storage[8][16] , \Storage[8][15] ,
         \Storage[8][14] , \Storage[8][13] , \Storage[8][12] ,
         \Storage[8][11] , \Storage[8][10] , \Storage[8][9] , \Storage[8][8] ,
         \Storage[8][7] , \Storage[8][6] , \Storage[8][5] , \Storage[8][4] ,
         \Storage[8][3] , \Storage[8][2] , \Storage[8][1] , \Storage[8][0] ,
         \Storage[7][32] , \Storage[7][31] , \Storage[7][30] ,
         \Storage[7][29] , \Storage[7][28] , \Storage[7][27] ,
         \Storage[7][26] , \Storage[7][25] , \Storage[7][24] ,
         \Storage[7][23] , \Storage[7][22] , \Storage[7][21] ,
         \Storage[7][20] , \Storage[7][19] , \Storage[7][18] ,
         \Storage[7][17] , \Storage[7][16] , \Storage[7][15] ,
         \Storage[7][14] , \Storage[7][13] , \Storage[7][12] ,
         \Storage[7][11] , \Storage[7][10] , \Storage[7][9] , \Storage[7][8] ,
         \Storage[7][7] , \Storage[7][6] , \Storage[7][5] , \Storage[7][4] ,
         \Storage[7][3] , \Storage[7][2] , \Storage[7][1] , \Storage[7][0] ,
         \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N116, N117, N1240, N1273,
         N1306, N1339, N1372, N1405, N1438, N1471, N1504, N1537, N1570, N1603,
         N1636, N1669, N1702, N1735, N1768, N1801, N1834, N1867, N1900, N1933,
         N1966, N1999, N2032, N2065, N2098, N2131, N2164, N2197, N2230, N2263,
         N2264, N2327, N2328, N2330, N2333, N2336, N2339, N2342, N2345, N2348,
         N2351, N2354, N2357, N2360, N2363, N2366, N2369, N2372, N2375, N2378,
         N2381, N2384, N2387, N2390, N2393, N2396, N2399, N2402, N2405, N2408,
         N2411, N2414, N2417, N2420, N2423, \DataOreg[9] , \DataOreg[8] ,
         \DataOreg[7] , \DataOreg[6] , \DataOreg[5] , \DataOreg[4] ,
         \DataOreg[3] , \DataOreg[31] , \DataOreg[30] , \DataOreg[2] ,
         \DataOreg[29] , \DataOreg[28] , \DataOreg[27] , \DataOreg[26] ,
         \DataOreg[25] , \DataOreg[24] , \DataOreg[23] , \DataOreg[22] ,
         \DataOreg[21] , \DataOreg[20] , \DataOreg[1] , \DataOreg[19] ,
         \DataOreg[18] , \DataOreg[17] , \DataOreg[16] , \DataOreg[15] ,
         \DataOreg[14] , \DataOreg[13] , \DataOreg[12] , \DataOreg[11] ,
         \DataOreg[10] , \DataOreg[0] , n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608;
  assign N75 = Addr[0];
  assign N76 = Addr[1];
  assign N77 = Addr[2];
  assign N78 = Addr[3];
  assign N79 = Addr[4];

  BUFTD1 \DataOreg_tri[0]  ( .I(N2423), .OE(n173), .Z(\DataOreg[0] ) );
  BUFTD1 \DataOreg_tri[1]  ( .I(N2420), .OE(n172), .Z(\DataOreg[1] ) );
  BUFTD1 \DataOreg_tri[2]  ( .I(N2417), .OE(n171), .Z(\DataOreg[2] ) );
  BUFTD1 \DataOreg_tri[3]  ( .I(N2414), .OE(n170), .Z(\DataOreg[3] ) );
  BUFTD1 \DataOreg_tri[4]  ( .I(N2411), .OE(n169), .Z(\DataOreg[4] ) );
  BUFTD1 \DataOreg_tri[5]  ( .I(N2408), .OE(n168), .Z(\DataOreg[5] ) );
  BUFTD1 \DataOreg_tri[6]  ( .I(N2405), .OE(n167), .Z(\DataOreg[6] ) );
  BUFTD1 \DataOreg_tri[7]  ( .I(N2402), .OE(n166), .Z(\DataOreg[7] ) );
  BUFTD1 \DataOreg_tri[8]  ( .I(N2399), .OE(n165), .Z(\DataOreg[8] ) );
  BUFTD1 \DataOreg_tri[9]  ( .I(N2396), .OE(n164), .Z(\DataOreg[9] ) );
  BUFTD1 \DataOreg_tri[10]  ( .I(N2393), .OE(n163), .Z(\DataOreg[10] ) );
  BUFTD1 \DataOreg_tri[11]  ( .I(N2390), .OE(n162), .Z(\DataOreg[11] ) );
  BUFTD1 \DataOreg_tri[12]  ( .I(N2387), .OE(n161), .Z(\DataOreg[12] ) );
  BUFTD1 \DataOreg_tri[13]  ( .I(N2384), .OE(n160), .Z(\DataOreg[13] ) );
  BUFTD1 \DataOreg_tri[14]  ( .I(N2381), .OE(n159), .Z(\DataOreg[14] ) );
  BUFTD1 \DataOreg_tri[15]  ( .I(N2378), .OE(n158), .Z(\DataOreg[15] ) );
  BUFTD1 \DataOreg_tri[16]  ( .I(N2375), .OE(n157), .Z(\DataOreg[16] ) );
  BUFTD1 \DataOreg_tri[17]  ( .I(N2372), .OE(n156), .Z(\DataOreg[17] ) );
  BUFTD1 \DataOreg_tri[18]  ( .I(N2369), .OE(n155), .Z(\DataOreg[18] ) );
  BUFTD1 \DataOreg_tri[19]  ( .I(N2366), .OE(n154), .Z(\DataOreg[19] ) );
  BUFTD1 \DataOreg_tri[20]  ( .I(N2363), .OE(n153), .Z(\DataOreg[20] ) );
  BUFTD1 \DataOreg_tri[21]  ( .I(N2360), .OE(n152), .Z(\DataOreg[21] ) );
  BUFTD1 \DataOreg_tri[22]  ( .I(N2357), .OE(n151), .Z(\DataOreg[22] ) );
  BUFTD1 \DataOreg_tri[23]  ( .I(N2354), .OE(n150), .Z(\DataOreg[23] ) );
  BUFTD1 \DataOreg_tri[24]  ( .I(N2351), .OE(n149), .Z(\DataOreg[24] ) );
  BUFTD1 \DataOreg_tri[25]  ( .I(N2348), .OE(n148), .Z(\DataOreg[25] ) );
  BUFTD1 \DataOreg_tri[26]  ( .I(N2345), .OE(n147), .Z(\DataOreg[26] ) );
  BUFTD1 \DataOreg_tri[27]  ( .I(N2342), .OE(n146), .Z(\DataOreg[27] ) );
  BUFTD1 \DataOreg_tri[28]  ( .I(N2339), .OE(n145), .Z(\DataOreg[28] ) );
  BUFTD1 \DataOreg_tri[29]  ( .I(N2336), .OE(n144), .Z(\DataOreg[29] ) );
  BUFTD1 \DataOreg_tri[30]  ( .I(N2333), .OE(n143), .Z(\DataOreg[30] ) );
  BUFTD1 \DataOreg_tri[31]  ( .I(N2330), .OE(n142), .Z(\DataOreg[31] ) );
  BUFTD1 \DataO_tri[0]  ( .I(\DataOreg[0] ), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD1 \DataO_tri[1]  ( .I(\DataOreg[1] ), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD1 \DataO_tri[2]  ( .I(\DataOreg[2] ), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD1 \DataO_tri[3]  ( .I(\DataOreg[3] ), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD1 \DataO_tri[4]  ( .I(\DataOreg[4] ), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD1 \DataO_tri[5]  ( .I(\DataOreg[5] ), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD1 \DataO_tri[6]  ( .I(\DataOreg[6] ), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD1 \DataO_tri[7]  ( .I(\DataOreg[7] ), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD1 \DataO_tri[8]  ( .I(\DataOreg[8] ), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD1 \DataO_tri[9]  ( .I(\DataOreg[9] ), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD1 \DataO_tri[10]  ( .I(\DataOreg[10] ), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD1 \DataO_tri[11]  ( .I(\DataOreg[11] ), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD1 \DataO_tri[12]  ( .I(\DataOreg[12] ), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD1 \DataO_tri[13]  ( .I(\DataOreg[13] ), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD1 \DataO_tri[14]  ( .I(\DataOreg[14] ), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD1 \DataO_tri[15]  ( .I(\DataOreg[15] ), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD1 \DataO_tri[16]  ( .I(\DataOreg[16] ), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD1 \DataO_tri[17]  ( .I(\DataOreg[17] ), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD1 \DataO_tri[18]  ( .I(\DataOreg[18] ), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD1 \DataO_tri[19]  ( .I(\DataOreg[19] ), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD1 \DataO_tri[20]  ( .I(\DataOreg[20] ), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD1 \DataO_tri[21]  ( .I(\DataOreg[21] ), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD1 \DataO_tri[22]  ( .I(\DataOreg[22] ), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD1 \DataO_tri[23]  ( .I(\DataOreg[23] ), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD1 \DataO_tri[24]  ( .I(\DataOreg[24] ), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD1 \DataO_tri[25]  ( .I(\DataOreg[25] ), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD1 \DataO_tri[26]  ( .I(\DataOreg[26] ), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD1 \DataO_tri[27]  ( .I(\DataOreg[27] ), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD1 \DataO_tri[28]  ( .I(\DataOreg[28] ), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD1 \DataO_tri[29]  ( .I(\DataOreg[29] ), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD1 \DataO_tri[30]  ( .I(\DataOreg[30] ), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD1 \DataO_tri[31]  ( .I(\DataOreg[31] ), .OE(ChipEna), .Z(DataO[31]) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(DataI[31]), .E(N2032), .CP(n59), .CDN(
        n29), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(DataI[30]), .E(N2032), .CP(n69), .CDN(
        n29), .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(N117), .E(N2098), .CP(n48), .CDN(n7), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(N2098), .CP(n68), .CDN(
        n27), .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(DataI[30]), .E(N2098), .CP(n58), .CDN(
        n27), .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(DataI[29]), .E(N2098), .CP(n64), .CDN(
        n27), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(N2098), .CP(n43), .CDN(
        n27), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(N2098), .CP(n42), .CDN(
        n27), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(DataI[26]), .E(N2098), .CP(n65), .CDN(
        n27), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(DataI[25]), .E(N2098), .CP(n44), .CDN(
        n27), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(N2098), .CP(n62), .CDN(
        n26), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(N2098), .CP(n62), .CDN(
        n26), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(DataI[22]), .E(N2098), .CP(n70), .CDN(
        n26), .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(DataI[21]), .E(N2098), .CP(n66), .CDN(
        n26), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(N2098), .CP(n45), .CDN(
        n26), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(N2098), .CP(n49), .CDN(
        n26), .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(DataI[18]), .E(N2098), .CP(n64), .CDN(
        n26), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(DataI[17]), .E(N2098), .CP(n56), .CDN(
        n26), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(N2098), .CP(n71), .CDN(
        n26), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(DataI[15]), .E(N2098), .CP(n55), .CDN(
        n26), .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(DataI[14]), .E(N2098), .CP(n73), .CDN(
        n26), .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(N2098), .CP(n72), .CDN(
        n25), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(DataI[12]), .E(N2098), .CP(n67), .CDN(
        n25), .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(DataI[11]), .E(N2098), .CP(n60), .CDN(
        n25), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(DataI[10]), .E(N2098), .CP(n67), .CDN(
        n25), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(DataI[9]), .E(N2098), .CP(n71), .CDN(n25), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(DataI[8]), .E(N2098), .CP(n50), .CDN(n25), 
        .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(DataI[7]), .E(N2098), .CP(n58), .CDN(n28), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(DataI[6]), .E(N2098), .CP(n58), .CDN(n30), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(DataI[5]), .E(N2098), .CP(n49), .CDN(n30), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(DataI[4]), .E(N2098), .CP(n45), .CDN(n35), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(DataI[3]), .E(N2098), .CP(n56), .CDN(n34), 
        .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(DataI[2]), .E(N2098), .CP(n54), .CDN(n37), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(N2098), .CP(n51), .CDN(n2), 
        .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(DataI[0]), .E(N2098), .CP(n44), .CDN(n4), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(N117), .E(N2032), .CP(n47), .CDN(n7), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(DataI[29]), .E(N2032), .CP(n59), .CDN(
        n29), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(DataI[28]), .E(N2032), .CP(n45), .CDN(
        n29), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(DataI[27]), .E(N2032), .CP(n61), .CDN(
        n29), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(DataI[26]), .E(N2032), .CP(n60), .CDN(
        n29), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(DataI[25]), .E(N2032), .CP(n73), .CDN(
        n29), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(DataI[24]), .E(N2032), .CP(n72), .CDN(
        n29), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(DataI[23]), .E(N2032), .CP(n48), .CDN(
        n29), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(DataI[22]), .E(N2032), .CP(n50), .CDN(
        n29), .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(DataI[21]), .E(N2032), .CP(n70), .CDN(
        n29), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(DataI[20]), .E(N2032), .CP(n65), .CDN(
        n23), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(DataI[19]), .E(N2032), .CP(n64), .CDN(
        n41), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(DataI[18]), .E(N2032), .CP(n63), .CDN(
        n40), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(DataI[17]), .E(N2032), .CP(n72), .CDN(
        n38), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(DataI[16]), .E(N2032), .CP(n58), .CDN(
        n10), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(DataI[15]), .E(N2032), .CP(n47), .CDN(
        n14), .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(DataI[14]), .E(N2032), .CP(n70), .CDN(
        n37), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(DataI[13]), .E(N2032), .CP(n66), .CDN(
        n36), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(DataI[12]), .E(N2032), .CP(n62), .CDN(
        n39), .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(DataI[11]), .E(N2032), .CP(n57), .CDN(
        n41), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(DataI[10]), .E(N2032), .CP(n71), .CDN(
        n27), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(DataI[9]), .E(N2032), .CP(n66), .CDN(n20), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(DataI[8]), .E(N2032), .CP(n68), .CDN(n24), 
        .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(DataI[7]), .E(N2032), .CP(n70), .CDN(n29), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(DataI[6]), .E(N2032), .CP(n63), .CDN(n6), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(DataI[5]), .E(N2032), .CP(n67), .CDN(n10), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(DataI[4]), .E(N2032), .CP(n42), .CDN(n14), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(DataI[3]), .E(N2032), .CP(n56), .CDN(n33), 
        .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(DataI[2]), .E(N2032), .CP(n54), .CDN(n16), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(DataI[1]), .E(N2032), .CP(n51), .CDN(n7), 
        .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(DataI[0]), .E(N2032), .CP(n44), .CDN(n4), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(N117), .E(N2230), .CP(n48), .CDN(n7), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(N2230), .CP(n55), .CDN(
        n18), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(N2230), .CP(n64), .CDN(
        n18), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(N2230), .CP(n63), .CDN(
        n18), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(N2230), .CP(n62), .CDN(
        n18), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(N2230), .CP(n64), .CDN(
        n18), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(N2230), .CP(n61), .CDN(
        n18), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(N2230), .CP(n60), .CDN(
        n18), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(N2230), .CP(n66), .CDN(
        n18), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(N2230), .CP(n61), .CDN(
        n18), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(N2230), .CP(n66), .CDN(
        n18), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(N2230), .CP(n72), .CDN(
        n17), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(N2230), .CP(n67), .CDN(
        n17), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(N2230), .CP(n68), .CDN(
        n17), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(N2230), .CP(n53), .CDN(
        n17), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(N2230), .CP(n73), .CDN(
        n17), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(N2230), .CP(n74), .CDN(
        n17), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(N2230), .CP(n46), .CDN(
        n17), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(N2230), .CP(n46), .CDN(
        n17), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(N2230), .CP(n43), .CDN(
        n17), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(DataI[12]), .E(N2230), .CP(n48), .CDN(
        n17), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(N2230), .CP(n50), .CDN(
        n17), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(N2230), .CP(n52), .CDN(
        n16), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(DataI[9]), .E(N2230), .CP(n64), .CDN(n16), 
        .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(N2230), .CP(n62), .CDN(n16), 
        .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(N2230), .CP(n44), .CDN(n16), 
        .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(DataI[6]), .E(N2230), .CP(n62), .CDN(n5), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(DataI[5]), .E(N2230), .CP(n62), .CDN(n14), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(N2230), .CP(n60), .CDN(n12), 
        .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(N2230), .CP(n57), .CDN(n34), 
        .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(DataI[2]), .E(N2230), .CP(n55), .CDN(n18), 
        .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(N2230), .CP(n51), .CDN(n38), 
        .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(DataI[0]), .E(N2230), .CP(n45), .CDN(n4), 
        .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(N117), .E(N2197), .CP(n48), .CDN(n7), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(N2197), .CP(n59), .CDN(
        n21), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(N2197), .CP(n44), .CDN(
        n20), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(N2197), .CP(n63), .CDN(
        n20), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(N2197), .CP(n48), .CDN(
        n20), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(DataI[27]), .E(N2197), .CP(n51), .CDN(
        n20), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(N2197), .CP(n42), .CDN(
        n20), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(N2197), .CP(n74), .CDN(
        n20), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(N2197), .CP(n65), .CDN(
        n20), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(DataI[23]), .E(N2197), .CP(n66), .CDN(
        n20), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(N2197), .CP(n71), .CDN(
        n20), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(N2197), .CP(n64), .CDN(
        n20), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(N2197), .CP(n62), .CDN(
        n20), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(N2197), .CP(n60), .CDN(
        n19), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(N2197), .CP(n53), .CDN(
        n19), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(N2197), .CP(n42), .CDN(
        n19), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(N2197), .CP(n49), .CDN(
        n19), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(N2197), .CP(n71), .CDN(
        n19), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(N2197), .CP(n69), .CDN(
        n19), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(DataI[13]), .E(N2197), .CP(n58), .CDN(
        n19), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(N2197), .CP(n47), .CDN(
        n19), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(N2197), .CP(n67), .CDN(
        n19), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(N2197), .CP(n72), .CDN(
        n19), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(N2197), .CP(n65), .CDN(n19), 
        .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(N2197), .CP(n58), .CDN(n18), 
        .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(N2197), .CP(n66), .CDN(n30), 
        .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(DataI[6]), .E(N2197), .CP(n63), .CDN(n7), 
        .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(DataI[5]), .E(N2197), .CP(n63), .CDN(n3), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(N2197), .CP(n46), .CDN(n13), 
        .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(N2197), .CP(n57), .CDN(n30), 
        .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(N2197), .CP(n54), .CDN(n17), 
        .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(N2197), .CP(n51), .CDN(n36), 
        .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(DataI[0]), .E(N2197), .CP(n45), .CDN(n4), 
        .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(N117), .E(N2164), .CP(n48), .CDN(n7), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(N2164), .CP(n69), .CDN(
        n23), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(DataI[30]), .E(N2164), .CP(n71), .CDN(
        n23), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(DataI[29]), .E(N2164), .CP(n53), .CDN(
        n23), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(N2164), .CP(n42), .CDN(
        n22), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(N2164), .CP(n66), .CDN(
        n22), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(DataI[26]), .E(N2164), .CP(n45), .CDN(
        n22), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(DataI[25]), .E(N2164), .CP(n64), .CDN(
        n22), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(N2164), .CP(n67), .CDN(
        n22), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(N2164), .CP(n63), .CDN(
        n22), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(DataI[22]), .E(N2164), .CP(n53), .CDN(
        n22), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(DataI[21]), .E(N2164), .CP(n73), .CDN(
        n22), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(N2164), .CP(n63), .CDN(
        n22), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(N2164), .CP(n43), .CDN(
        n22), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(DataI[18]), .E(N2164), .CP(n73), .CDN(
        n22), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(DataI[17]), .E(N2164), .CP(n57), .CDN(
        n21), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(N2164), .CP(n72), .CDN(
        n21), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(DataI[15]), .E(N2164), .CP(n43), .CDN(
        n21), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(DataI[14]), .E(N2164), .CP(n45), .CDN(
        n21), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(N2164), .CP(n46), .CDN(
        n21), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(DataI[12]), .E(N2164), .CP(n42), .CDN(
        n21), .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(DataI[11]), .E(N2164), .CP(n63), .CDN(
        n21), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(DataI[10]), .E(N2164), .CP(n71), .CDN(
        n21), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(DataI[9]), .E(N2164), .CP(n52), .CDN(n21), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(DataI[8]), .E(N2164), .CP(n70), .CDN(n21), 
        .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(DataI[7]), .E(N2164), .CP(n61), .CDN(n39), 
        .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(DataI[6]), .E(N2164), .CP(n59), .CDN(n4), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(DataI[5]), .E(N2164), .CP(n61), .CDN(n27), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(DataI[4]), .E(N2164), .CP(n67), .CDN(n11), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(DataI[3]), .E(N2164), .CP(n57), .CDN(n27), 
        .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(DataI[2]), .E(N2164), .CP(n54), .CDN(n19), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(DataI[1]), .E(N2164), .CP(n51), .CDN(n39), 
        .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(DataI[0]), .E(N2164), .CP(n45), .CDN(n4), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \DataOreg_tri_enable_reg[31]  ( .D(N2328), .E(N2327), .CP(n42), 
        .CDN(n32), .Q(N32) );
  EDFCNQD1 \DataOreg_tri_enable_reg[30]  ( .D(N2328), .E(N2327), .CP(n50), 
        .CDN(n33), .Q(N33) );
  EDFCNQD1 \DataOreg_tri_enable_reg[29]  ( .D(N2328), .E(N2327), .CP(n63), 
        .CDN(n33), .Q(N34) );
  EDFCNQD1 \DataOreg_tri_enable_reg[28]  ( .D(N2328), .E(N2327), .CP(n46), 
        .CDN(n174), .Q(N35) );
  EDFCNQD1 \DataOreg_tri_enable_reg[27]  ( .D(N2328), .E(N2327), .CP(n73), 
        .CDN(n35), .Q(N36) );
  EDFCNQD1 \DataOreg_tri_enable_reg[26]  ( .D(N2328), .E(N2327), .CP(n52), 
        .CDN(n25), .Q(N37) );
  EDFCNQD1 \DataOreg_tri_enable_reg[25]  ( .D(N2328), .E(N2327), .CP(n54), 
        .CDN(n40), .Q(N38) );
  EDFCNQD1 \DataOreg_tri_enable_reg[24]  ( .D(N2328), .E(N2327), .CP(n59), 
        .CDN(n13), .Q(N39) );
  EDFCNQD1 \DataOreg_tri_enable_reg[23]  ( .D(N2328), .E(N2327), .CP(n63), 
        .CDN(n7), .Q(N40) );
  EDFCNQD1 \DataOreg_tri_enable_reg[22]  ( .D(N2328), .E(N2327), .CP(n62), 
        .CDN(n7), .Q(N41) );
  EDFCNQD1 \DataOreg_tri_enable_reg[21]  ( .D(N2328), .E(N2327), .CP(n64), 
        .CDN(n2), .Q(N42) );
  EDFCNQD1 \DataOreg_tri_enable_reg[20]  ( .D(N2328), .E(N2327), .CP(n71), 
        .CDN(n7), .Q(N43) );
  EDFCNQD1 \DataOreg_tri_enable_reg[19]  ( .D(N2328), .E(N2327), .CP(n54), 
        .CDN(n36), .Q(N44) );
  EDFCNQD1 \DataOreg_tri_enable_reg[18]  ( .D(N2328), .E(N2327), .CP(n58), 
        .CDN(n28), .Q(N45) );
  EDFCNQD1 \DataOreg_tri_enable_reg[17]  ( .D(N2328), .E(N2327), .CP(n53), 
        .CDN(n29), .Q(N46) );
  EDFCNQD1 \DataOreg_tri_enable_reg[16]  ( .D(N2328), .E(N2327), .CP(n66), 
        .CDN(n17), .Q(N47) );
  EDFCNQD1 \DataOreg_tri_enable_reg[15]  ( .D(N2328), .E(N2327), .CP(n58), 
        .CDN(n4), .Q(N48) );
  EDFCNQD1 \DataOreg_tri_enable_reg[14]  ( .D(N2328), .E(N2327), .CP(n47), 
        .CDN(n30), .Q(N49) );
  EDFCNQD1 \DataOreg_tri_enable_reg[13]  ( .D(N2328), .E(N2327), .CP(n73), 
        .CDN(n35), .Q(N50) );
  EDFCNQD1 \DataOreg_tri_enable_reg[12]  ( .D(N2328), .E(N2327), .CP(n43), 
        .CDN(n32), .Q(N51) );
  EDFCNQD1 \DataOreg_tri_enable_reg[11]  ( .D(N2328), .E(N2327), .CP(n47), 
        .CDN(n38), .Q(N52) );
  EDFCNQD1 \DataOreg_tri_enable_reg[10]  ( .D(N2328), .E(N2327), .CP(n59), 
        .CDN(n40), .Q(N53) );
  EDFCNQD1 \DataOreg_tri_enable_reg[9]  ( .D(N2328), .E(N2327), .CP(n48), 
        .CDN(n37), .Q(N54) );
  EDFCNQD1 \DataOreg_tri_enable_reg[8]  ( .D(N2328), .E(N2327), .CP(n70), 
        .CDN(n2), .Q(N55) );
  EDFCNQD1 \DataOreg_tri_enable_reg[7]  ( .D(N2328), .E(N2327), .CP(n51), 
        .CDN(n7), .Q(N56) );
  EDFCNQD1 \DataOreg_tri_enable_reg[6]  ( .D(N2328), .E(N2327), .CP(n60), 
        .CDN(n5), .Q(N57) );
  EDFCNQD1 \DataOreg_tri_enable_reg[5]  ( .D(N2328), .E(N2327), .CP(n53), 
        .CDN(n6), .Q(N58) );
  EDFCNQD1 \DataOreg_tri_enable_reg[4]  ( .D(N2328), .E(N2327), .CP(n64), 
        .CDN(n25), .Q(N59) );
  EDFCNQD1 \DataOreg_tri_enable_reg[3]  ( .D(N2328), .E(N2327), .CP(n43), 
        .CDN(n24), .Q(N60) );
  EDFCNQD1 \DataOreg_tri_enable_reg[2]  ( .D(N2328), .E(N2327), .CP(n61), 
        .CDN(n25), .Q(N61) );
  EDFCNQD1 \DataOreg_tri_enable_reg[1]  ( .D(N2328), .E(N2327), .CP(n63), 
        .CDN(n26), .Q(N62) );
  EDFCNQD1 \DataOreg_tri_enable_reg[0]  ( .D(N2328), .E(N2327), .CP(n62), 
        .CDN(n23), .Q(N63) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(N117), .E(N2131), .CP(n48), .CDN(n7), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(N2131), .CP(n48), .CDN(
        n25), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(N2131), .CP(n61), .CDN(
        n25), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(DataI[29]), .E(N2131), .CP(n68), .CDN(
        n25), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(N2131), .CP(n57), .CDN(
        n25), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(N2131), .CP(n68), .CDN(
        n25), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(N2131), .CP(n50), .CDN(
        n24), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(N2131), .CP(n51), .CDN(
        n24), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(N2131), .CP(n66), .CDN(
        n24), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(N2131), .CP(n64), .CDN(
        n24), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(DataI[22]), .E(N2131), .CP(n47), .CDN(
        n24), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(N2131), .CP(n65), .CDN(
        n24), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(N2131), .CP(n58), .CDN(
        n24), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(N2131), .CP(n57), .CDN(
        n24), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(N2131), .CP(n55), .CDN(
        n24), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(DataI[17]), .E(N2131), .CP(n44), .CDN(
        n24), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(N2131), .CP(n58), .CDN(
        n24), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(DataI[15]), .E(N2131), .CP(n51), .CDN(
        n23), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(DataI[14]), .E(N2131), .CP(n60), .CDN(
        n23), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(N2131), .CP(n49), .CDN(
        n23), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(N2131), .CP(n57), .CDN(
        n23), .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(N2131), .CP(n54), .CDN(
        n23), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(DataI[10]), .E(N2131), .CP(n62), .CDN(
        n23), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(N2131), .CP(n67), .CDN(n23), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(N2131), .CP(n50), .CDN(n23), 
        .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(DataI[7]), .E(N2131), .CP(n70), .CDN(n38), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(DataI[6]), .E(N2131), .CP(n61), .CDN(n2), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(N2131), .CP(n49), .CDN(n20), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(DataI[4]), .E(N2131), .CP(n72), .CDN(n19), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(DataI[3]), .E(N2131), .CP(n57), .CDN(n32), 
        .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(DataI[2]), .E(N2131), .CP(n54), .CDN(n18), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(DataI[1]), .E(N2131), .CP(n51), .CDN(n23), 
        .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(N2131), .CP(n44), .CDN(n4), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(N117), .E(N2065), .CP(n47), .CDN(n7), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(N2065), .CP(n72), .CDN(
        n27), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(DataI[30]), .E(N2065), .CP(n67), .CDN(
        n26), .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(N2065), .CP(n62), .CDN(
        n35), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(N2065), .CP(n64), .CDN(
        n32), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(N2065), .CP(n50), .CDN(
        n30), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(DataI[26]), .E(N2065), .CP(ChipClock), 
        .CDN(n33), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(DataI[25]), .E(N2065), .CP(n74), .CDN(
        n38), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(N2065), .CP(n65), .CDN(
        n40), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(N2065), .CP(n50), .CDN(
        n37), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(DataI[22]), .E(N2065), .CP(ChipClock), 
        .CDN(n28), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(DataI[21]), .E(N2065), .CP(n53), .CDN(
        n28), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(N2065), .CP(n59), .CDN(
        n28), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(N2065), .CP(n65), .CDN(
        n28), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(DataI[18]), .E(N2065), .CP(n69), .CDN(
        n28), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(N2065), .CP(n50), .CDN(
        n28), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(N2065), .CP(n74), .CDN(
        n28), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(N2065), .CP(n59), .CDN(
        n28), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(DataI[14]), .E(N2065), .CP(n48), .CDN(
        n28), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(N2065), .CP(n54), .CDN(
        n28), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(DataI[12]), .E(N2065), .CP(n73), .CDN(
        n28), .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(DataI[11]), .E(N2065), .CP(n71), .CDN(
        n27), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(N2065), .CP(n42), .CDN(
        n27), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(DataI[9]), .E(N2065), .CP(n69), .CDN(n27), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(DataI[8]), .E(N2065), .CP(n70), .CDN(n27), 
        .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(N2065), .CP(n65), .CDN(n40), 
        .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(DataI[6]), .E(N2065), .CP(n59), .CDN(n15), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(DataI[5]), .E(N2065), .CP(n66), .CDN(n37), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(DataI[4]), .E(N2065), .CP(n59), .CDN(n7), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(N2065), .CP(n56), .CDN(n28), 
        .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(N2065), .CP(n54), .CDN(n29), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(N2065), .CP(n51), .CDN(n5), 
        .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(DataI[0]), .E(N2065), .CP(n44), .CDN(n4), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(N117), .E(N1966), .CP(n47), .CDN(n7), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(DataI[31]), .E(N1966), .CP(n70), .CDN(
        n13), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(DataI[30]), .E(N1966), .CP(n46), .CDN(
        n10), .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(DataI[29]), .E(N1966), .CP(n68), .CDN(
        n16), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(DataI[28]), .E(N1966), .CP(n62), .CDN(
        n12), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(DataI[27]), .E(N1966), .CP(n44), .CDN(
        n26), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(DataI[26]), .E(N1966), .CP(n64), .CDN(
        n20), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(DataI[25]), .E(N1966), .CP(n70), .CDN(n3), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(DataI[24]), .E(N1966), .CP(n74), .CDN(
        n32), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(DataI[23]), .E(N1966), .CP(n70), .CDN(
        n33), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(DataI[22]), .E(N1966), .CP(n57), .CDN(
        n34), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(DataI[21]), .E(N1966), .CP(n68), .CDN(
        n30), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(DataI[20]), .E(N1966), .CP(n56), .CDN(
        n15), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(DataI[19]), .E(N1966), .CP(n74), .CDN(n4), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(DataI[18]), .E(N1966), .CP(n73), .CDN(
        n174), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(DataI[17]), .E(N1966), .CP(n68), .CDN(
        n40), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(DataI[16]), .E(N1966), .CP(n69), .CDN(
        n174), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(DataI[15]), .E(N1966), .CP(n42), .CDN(
        n38), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(DataI[14]), .E(N1966), .CP(n74), .CDN(
        n16), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(DataI[13]), .E(N1966), .CP(n64), .CDN(
        n18), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(DataI[12]), .E(N1966), .CP(n74), .CDN(
        n17), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(DataI[11]), .E(N1966), .CP(n57), .CDN(
        n19), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(DataI[10]), .E(N1966), .CP(n48), .CDN(
        n21), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(DataI[9]), .E(N1966), .CP(n73), .CDN(n9), 
        .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(DataI[8]), .E(N1966), .CP(n68), .CDN(n8), 
        .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(DataI[7]), .E(N1966), .CP(n53), .CDN(n37), 
        .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(DataI[6]), .E(N1966), .CP(n60), .CDN(n14), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(DataI[5]), .E(N1966), .CP(n70), .CDN(n39), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(DataI[4]), .E(N1966), .CP(n69), .CDN(n22), 
        .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(DataI[3]), .E(N1966), .CP(n56), .CDN(n11), 
        .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(DataI[2]), .E(N1966), .CP(n54), .CDN(n34), 
        .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(DataI[1]), .E(N1966), .CP(n50), .CDN(n3), 
        .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(DataI[0]), .E(N1966), .CP(n44), .CDN(n4), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(N117), .E(N1933), .CP(n47), .CDN(n7), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(DataI[31]), .E(N1933), .CP(n47), .CDN(
        n35), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(DataI[30]), .E(N1933), .CP(n60), .CDN(
        n37), .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(DataI[29]), .E(N1933), .CP(n53), .CDN(
        n39), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(DataI[28]), .E(N1933), .CP(n51), .CDN(
        n38), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(N1933), .CP(n59), .CDN(
        n35), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(DataI[26]), .E(N1933), .CP(n68), .CDN(
        n36), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(DataI[25]), .E(N1933), .CP(n69), .CDN(
        n12), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(DataI[24]), .E(N1933), .CP(n64), .CDN(n8), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(N1933), .CP(n63), .CDN(
        n35), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(DataI[22]), .E(N1933), .CP(n73), .CDN(
        n12), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(DataI[21]), .E(N1933), .CP(n50), .CDN(
        n19), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(DataI[20]), .E(N1933), .CP(n50), .CDN(
        n17), .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(DataI[19]), .E(N1933), .CP(n60), .CDN(
        n18), .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(N1933), .CP(n71), .CDN(
        n16), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(DataI[17]), .E(N1933), .CP(n69), .CDN(
        n21), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(DataI[16]), .E(N1933), .CP(n64), .CDN(
        n20), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(DataI[15]), .E(N1933), .CP(n57), .CDN(
        n23), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(DataI[14]), .E(N1933), .CP(n65), .CDN(
        n22), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(DataI[13]), .E(N1933), .CP(n74), .CDN(
        n40), .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(DataI[12]), .E(N1933), .CP(n68), .CDN(
        n12), .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(DataI[11]), .E(N1933), .CP(ChipClock), 
        .CDN(n18), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(DataI[10]), .E(N1933), .CP(n72), .CDN(
        n16), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(DataI[9]), .E(N1933), .CP(n67), .CDN(n3), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(DataI[8]), .E(N1933), .CP(n62), .CDN(n25), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(DataI[7]), .E(N1933), .CP(n54), .CDN(n36), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(DataI[6]), .E(N1933), .CP(n66), .CDN(n12), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(DataI[5]), .E(N1933), .CP(n72), .CDN(n20), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(DataI[4]), .E(N1933), .CP(n46), .CDN(n3), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(DataI[3]), .E(N1933), .CP(n56), .CDN(n30), 
        .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(DataI[2]), .E(N1933), .CP(n54), .CDN(n5), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(DataI[1]), .E(N1933), .CP(n50), .CDN(n41), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(DataI[0]), .E(N1933), .CP(n44), .CDN(n4), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N117), .E(N1834), .CP(n47), .CDN(n6), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(DataI[31]), .E(N1834), .CP(n58), .CDN(
        n10), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(DataI[30]), .E(N1834), .CP(n63), .CDN(
        n10), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(N1834), .CP(n52), .CDN(n9), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(DataI[28]), .E(N1834), .CP(n62), .CDN(n9), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(DataI[27]), .E(N1834), .CP(n51), .CDN(n9), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(DataI[26]), .E(N1834), .CP(n69), .CDN(n9), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(DataI[25]), .E(N1834), .CP(n73), .CDN(n9), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(DataI[24]), .E(N1834), .CP(n63), .CDN(n9), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(DataI[23]), .E(N1834), .CP(n72), .CDN(n9), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(DataI[22]), .E(N1834), .CP(n67), .CDN(n9), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(DataI[21]), .E(N1834), .CP(n42), .CDN(n9), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(N1834), .CP(n70), .CDN(n9), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(DataI[19]), .E(N1834), .CP(n44), .CDN(n9), .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(DataI[18]), .E(N1834), .CP(n65), .CDN(n8), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(N1834), .CP(n65), .CDN(n8), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(DataI[16]), .E(N1834), .CP(n46), .CDN(n8), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(N1834), .CP(n72), .CDN(n8), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(DataI[14]), .E(N1834), .CP(n58), .CDN(n8), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(DataI[13]), .E(N1834), .CP(n46), .CDN(n8), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(DataI[12]), .E(N1834), .CP(n68), .CDN(n8), .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(DataI[11]), .E(N1834), .CP(n59), .CDN(n8), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(N1834), .CP(n70), .CDN(n8), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(DataI[9]), .E(N1834), .CP(n58), .CDN(n8), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(DataI[8]), .E(N1834), .CP(n66), .CDN(n8), 
        .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(N1834), .CP(n49), .CDN(n17), 
        .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(DataI[6]), .E(N1834), .CP(n46), .CDN(n30), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(DataI[5]), .E(N1834), .CP(n69), .CDN(n21), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(DataI[4]), .E(N1834), .CP(n44), .CDN(n15), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(N1834), .CP(n56), .CDN(n8), 
        .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(DataI[2]), .E(N1834), .CP(n53), .CDN(n40), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(N1834), .CP(n50), .CDN(n14), 
        .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(DataI[0]), .E(N1834), .CP(n44), .CDN(n3), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(N117), .E(N1801), .CP(n47), .CDN(n6), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(DataI[31]), .E(N1801), .CP(n69), .CDN(
        n12), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(DataI[30]), .E(N1801), .CP(n58), .CDN(
        n12), .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(DataI[29]), .E(N1801), .CP(n46), .CDN(
        n12), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(DataI[28]), .E(N1801), .CP(n59), .CDN(
        n12), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(DataI[27]), .E(N1801), .CP(n57), .CDN(
        n11), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(DataI[26]), .E(N1801), .CP(n51), .CDN(
        n11), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(DataI[25]), .E(N1801), .CP(n45), .CDN(
        n11), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(DataI[24]), .E(N1801), .CP(n61), .CDN(
        n11), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(DataI[23]), .E(N1801), .CP(n74), .CDN(
        n11), .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(DataI[22]), .E(N1801), .CP(n69), .CDN(
        n11), .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(DataI[21]), .E(N1801), .CP(n48), .CDN(
        n11), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(DataI[20]), .E(N1801), .CP(n47), .CDN(
        n11), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(DataI[19]), .E(N1801), .CP(n49), .CDN(
        n11), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(DataI[18]), .E(N1801), .CP(n70), .CDN(
        n11), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(DataI[17]), .E(N1801), .CP(n66), .CDN(
        n11), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(DataI[16]), .E(N1801), .CP(n50), .CDN(
        n10), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(DataI[15]), .E(N1801), .CP(n71), .CDN(
        n10), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(DataI[14]), .E(N1801), .CP(n64), .CDN(
        n10), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(DataI[13]), .E(N1801), .CP(n62), .CDN(
        n10), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(DataI[12]), .E(N1801), .CP(n63), .CDN(
        n10), .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(DataI[11]), .E(N1801), .CP(n59), .CDN(
        n10), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(DataI[10]), .E(N1801), .CP(n60), .CDN(
        n10), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(DataI[9]), .E(N1801), .CP(n61), .CDN(n10), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(DataI[8]), .E(N1801), .CP(n44), .CDN(n10), 
        .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(DataI[7]), .E(N1801), .CP(n50), .CDN(n17), 
        .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(DataI[6]), .E(N1801), .CP(n60), .CDN(n19), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(DataI[5]), .E(N1801), .CP(n45), .CDN(n35), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(DataI[4]), .E(N1801), .CP(n43), .CDN(n26), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(DataI[3]), .E(N1801), .CP(n56), .CDN(n21), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(DataI[2]), .E(N1801), .CP(n53), .CDN(n20), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(DataI[1]), .E(N1801), .CP(n50), .CDN(n18), 
        .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(DataI[0]), .E(N1801), .CP(n43), .CDN(n3), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N117), .E(N1702), .CP(n46), .CDN(n6), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(N1702), .CP(n60), .CDN(
        n31), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(N1702), .CP(n49), .CDN(n6), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(N1702), .CP(n49), .CDN(
        n38), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(N1702), .CP(n66), .CDN(n3), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(N1702), .CP(n64), .CDN(n4), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(N1702), .CP(n54), .CDN(
        n37), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(N1702), .CP(n56), .CDN(
        n41), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(N1702), .CP(n43), .CDN(
        n39), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(N1702), .CP(n44), .CDN(
        n37), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(N1702), .CP(n42), .CDN(
        n41), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(N1702), .CP(n46), .CDN(
        n11), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(N1702), .CP(n72), .CDN(
        n15), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(N1702), .CP(n58), .CDN(
        n35), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(N1702), .CP(n71), .CDN(n6), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(N1702), .CP(n64), .CDN(n4), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(N1702), .CP(n50), .CDN(
        n36), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(N1702), .CP(n55), .CDN(
        n35), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(N1702), .CP(n54), .CDN(
        n17), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(N1702), .CP(n46), .CDN(
        n13), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(N1702), .CP(n57), .CDN(
        n30), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(N1702), .CP(n48), .CDN(
        n34), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(N1702), .CP(n56), .CDN(
        n33), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(N1702), .CP(n71), .CDN(n31), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(N1702), .CP(n68), .CDN(n9), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(N1702), .CP(n58), .CDN(n3), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(N1702), .CP(n45), .CDN(n16), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(N1702), .CP(n55), .CDN(n9), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(N1702), .CP(n42), .CDN(n23), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(N1702), .CP(n66), .CDN(n4), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(N1702), .CP(n53), .CDN(n21), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(N1702), .CP(n50), .CDN(n6), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(N1702), .CP(n43), .CDN(n3), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N117), .E(N1669), .CP(n46), .CDN(n6), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(N1669), .CP(n70), .CDN(
        n21), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(N1669), .CP(n49), .CDN(n5), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(N1669), .CP(n60), .CDN(
        n36), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(N1669), .CP(n52), .CDN(
        n40), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(N1669), .CP(n61), .CDN(
        n14), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(N1669), .CP(n58), .CDN(
        n37), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(N1669), .CP(n68), .CDN(
        n41), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(N1669), .CP(n73), .CDN(
        n39), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(N1669), .CP(n60), .CDN(
        n38), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(N1669), .CP(n54), .CDN(
        n32), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(N1669), .CP(n73), .CDN(
        n22), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(N1669), .CP(n55), .CDN(n9), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(N1669), .CP(n69), .CDN(
        n23), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(N1669), .CP(n55), .CDN(
        n18), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(N1669), .CP(n64), .CDN(
        n35), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(N1669), .CP(n45), .CDN(
        n41), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(N1669), .CP(n56), .CDN(
        n35), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(N1669), .CP(n69), .CDN(
        n26), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(N1669), .CP(n44), .CDN(
        n14), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(N1669), .CP(n58), .CDN(
        n11), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(N1669), .CP(n67), .CDN(
        n22), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(N1669), .CP(n73), .CDN(n9), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(N1669), .CP(n48), .CDN(n9), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(N1669), .CP(n55), .CDN(n29), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(N1669), .CP(n65), .CDN(n2), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(DataI[6]), .E(N1669), .CP(n68), .CDN(n18), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(N1669), .CP(n44), .CDN(n15), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(N1669), .CP(n42), .CDN(n41), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(N1669), .CP(n64), .CDN(n39), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(N1669), .CP(n53), .CDN(n10), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(N1669), .CP(n50), .CDN(n4), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(N1669), .CP(n43), .CDN(n3), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N117), .E(N1570), .CP(n46), .CDN(n6), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(N1570), .CP(n65), .CDN(
        n27), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(N1570), .CP(n43), .CDN(n2), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(N1570), .CP(n61), .CDN(
        n24), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(N1570), .CP(n60), .CDN(
        n31), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(N1570), .CP(n66), .CDN(
        n36), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(N1570), .CP(n52), .CDN(n5), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(N1570), .CP(n71), .CDN(
        n14), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(N1570), .CP(n43), .CDN(n9), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(N1570), .CP(n52), .CDN(
        n38), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(N1570), .CP(n62), .CDN(n2), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(N1570), .CP(n65), .CDN(n6), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(N1570), .CP(n53), .CDN(n4), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(N1570), .CP(n67), .CDN(n5), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(N1570), .CP(n68), .CDN(n7), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(N1570), .CP(n46), .CDN(
        n25), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(N1570), .CP(n44), .CDN(
        n19), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(DataI[15]), .E(N1570), .CP(n62), .CDN(
        n15), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(DataI[14]), .E(N1570), .CP(n74), .CDN(
        n21), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(DataI[13]), .E(N1570), .CP(n71), .CDN(n4), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(N1570), .CP(n72), .CDN(n8), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(N1570), .CP(n44), .CDN(
        n41), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(N1570), .CP(n55), .CDN(
        n28), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(N1570), .CP(n74), .CDN(n29), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(N1570), .CP(n46), .CDN(n3), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(DataI[7]), .E(N1570), .CP(n59), .CDN(n5), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(DataI[6]), .E(N1570), .CP(n67), .CDN(n17), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(DataI[5]), .E(N1570), .CP(n73), .CDN(n2), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(N1570), .CP(n43), .CDN(n30), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(N1570), .CP(n63), .CDN(n2), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(N1570), .CP(n53), .CDN(n11), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(N1570), .CP(n49), .CDN(n5), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(N1570), .CP(n43), .CDN(n3), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N117), .E(N1537), .CP(n46), .CDN(n5), .Q(
        \Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(N1537), .CP(n65), .CDN(n35), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(N1537), .CP(n62), .CDN(n3), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(N1537), .CP(n47), .CDN(n26), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(N1537), .CP(n45), .CDN(n31), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(N1537), .CP(n74), .CDN(n26), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(N1537), .CP(n52), .CDN(n34), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(N1537), .CP(n50), .CDN(n16), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(N1537), .CP(n45), .CDN(n41), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(N1537), .CP(n44), .CDN(n16), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(N1537), .CP(n42), .CDN(n11), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(N1537), .CP(n55), .CDN(n31), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(N1537), .CP(n47), .CDN(n30), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(N1537), .CP(n57), .CDN(n17), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(N1537), .CP(n44), .CDN(n34), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(N1537), .CP(n61), .CDN(n2), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(N1537), .CP(n48), .CDN(n32), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(DataI[15]), .E(N1537), .CP(n65), .CDN(n33), .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(N1537), .CP(n66), .CDN(n34), .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(N1537), .CP(n71), .CDN(n5), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(N1537), .CP(n64), .CDN(n31), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(N1537), .CP(n62), .CDN(n32), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(N1537), .CP(n63), .CDN(n35), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(N1537), .CP(n59), .CDN(n37), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(N1537), .CP(n60), .CDN(n29), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(DataI[7]), .E(N1537), .CP(n61), .CDN(n18), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(N1537), .CP(n46), .CDN(n6), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(N1537), .CP(n61), .CDN(n41), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(N1537), .CP(n52), .CDN(n19), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(N1537), .CP(n61), .CDN(n32), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(N1537), .CP(n52), .CDN(n12), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(N1537), .CP(n49), .CDN(n18), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(N1537), .CP(n43), .CDN(n3), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N117), .E(N1438), .CP(n46), .CDN(n5), .Q(
        \Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(N1438), .CP(n43), .CDN(n40), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(N1438), .CP(n65), .CDN(n9), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(N1438), .CP(n42), .CDN(n23), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(N1438), .CP(n61), .CDN(n4), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(N1438), .CP(n45), .CDN(n8), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(N1438), .CP(n71), .CDN(n21), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(N1438), .CP(n63), .CDN(n39), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(N1438), .CP(n62), .CDN(n8), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(N1438), .CP(n56), .CDN(n35), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(N1438), .CP(n47), .CDN(n37), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(N1438), .CP(n58), .CDN(n34), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(N1438), .CP(n45), .CDN(n21), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(N1438), .CP(n73), .CDN(n39), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(N1438), .CP(n69), .CDN(n34), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(N1438), .CP(n55), .CDN(n14), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(N1438), .CP(n72), .CDN(n39), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(N1438), .CP(n62), .CDN(n40), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(N1438), .CP(n60), .CDN(n30), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(N1438), .CP(n52), .CDN(n7), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(N1438), .CP(n66), .CDN(
        n174), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(N1438), .CP(n67), .CDN(n32), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(N1438), .CP(n53), .CDN(n31), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(N1438), .CP(n60), .CDN(n33), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(N1438), .CP(n68), .CDN(n32), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(N1438), .CP(n45), .CDN(n35), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(N1438), .CP(n68), .CDN(n25), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(N1438), .CP(n64), .CDN(n27), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(N1438), .CP(n71), .CDN(n22), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(N1438), .CP(n55), .CDN(n40), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(N1438), .CP(n52), .CDN(n40), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(N1438), .CP(n49), .CDN(n6), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(N1438), .CP(n42), .CDN(n2), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N117), .E(N1405), .CP(n45), .CDN(n5), .Q(
        \Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(N1405), .CP(n57), .CDN(n7), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(N1405), .CP(n61), .CDN(n2), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(N1405), .CP(n68), .CDN(n26), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(N1405), .CP(n70), .CDN(n34), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(N1405), .CP(n54), .CDN(n39), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(N1405), .CP(n43), .CDN(n35), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(N1405), .CP(n54), .CDN(n24), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(N1405), .CP(n67), .CDN(n36), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(N1405), .CP(n73), .CDN(n34), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(N1405), .CP(n68), .CDN(n36), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(N1405), .CP(n69), .CDN(n38), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(N1405), .CP(n70), .CDN(n41), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(N1405), .CP(n59), .CDN(n34), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(N1405), .CP(n55), .CDN(n30), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(N1405), .CP(n57), .CDN(
        n174), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(N1405), .CP(n65), .CDN(n37), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(N1405), .CP(n66), .CDN(n22), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(N1405), .CP(n47), .CDN(n22), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(N1405), .CP(n51), .CDN(n28), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(N1405), .CP(n71), .CDN(n21), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(N1405), .CP(n61), .CDN(n34), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(N1405), .CP(n50), .CDN(n17), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(N1405), .CP(n63), .CDN(n36), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(N1405), .CP(n58), .CDN(n36), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(N1405), .CP(n63), .CDN(n31), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(N1405), .CP(n59), .CDN(n4), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(N1405), .CP(n62), .CDN(n19), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(N1405), .CP(n73), .CDN(n26), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(N1405), .CP(n55), .CDN(n39), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(N1405), .CP(n52), .CDN(n15), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(N1405), .CP(n49), .CDN(n33), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(N1405), .CP(n42), .CDN(n2), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N117), .E(N1306), .CP(n45), .CDN(n5), .Q(
        \Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(N1306), .CP(n43), .CDN(n41), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(N1306), .CP(n69), .CDN(n39), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(N1306), .CP(n48), .CDN(n23), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(N1306), .CP(n52), .CDN(n37), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(N1306), .CP(n67), .CDN(n37), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(N1306), .CP(n66), .CDN(n40), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(N1306), .CP(n62), .CDN(n21), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(N1306), .CP(n70), .CDN(n13), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(N1306), .CP(n55), .CDN(n32), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(N1306), .CP(n65), .CDN(n27), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(N1306), .CP(n59), .CDN(n38), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(N1306), .CP(n63), .CDN(n39), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(N1306), .CP(n47), .CDN(n38), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(N1306), .CP(n62), .CDN(n31), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(N1306), .CP(n46), .CDN(n12), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(N1306), .CP(n58), .CDN(n10), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(N1306), .CP(n57), .CDN(n25), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(N1306), .CP(n55), .CDN(n41), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(N1306), .CP(n64), .CDN(n39), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(N1306), .CP(n56), .CDN(n41), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(N1306), .CP(n56), .CDN(n34), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(N1306), .CP(n66), .CDN(n35), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(N1306), .CP(n69), .CDN(n41), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(N1306), .CP(n43), .CDN(n24), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(N1306), .CP(n60), .CDN(n35), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(N1306), .CP(n58), .CDN(n28), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(N1306), .CP(n63), .CDN(n17), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(N1306), .CP(n57), .CDN(n27), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(N1306), .CP(n55), .CDN(n37), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(N1306), .CP(n52), .CDN(n10), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(N1306), .CP(n48), .CDN(n24), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(N1306), .CP(n42), .CDN(n2), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N117), .E(N1273), .CP(n45), .CDN(n5), .Q(
        \Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(N1273), .CP(n60), .CDN(n36), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(N1273), .CP(n65), .CDN(
        n174), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(N1273), .CP(n42), .CDN(n40), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(N1273), .CP(n69), .CDN(n33), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(N1273), .CP(n74), .CDN(n38), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(N1273), .CP(n72), .CDN(n34), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(N1273), .CP(n67), .CDN(n36), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(N1273), .CP(n49), .CDN(n15), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(N1273), .CP(n51), .CDN(n34), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(N1273), .CP(n49), .CDN(n33), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(N1273), .CP(n47), .CDN(n32), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(N1273), .CP(n63), .CDN(n31), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(N1273), .CP(n55), .CDN(n30), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(N1273), .CP(n53), .CDN(n24), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(N1273), .CP(n58), .CDN(n3), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(N1273), .CP(n54), .CDN(
        n174), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(N1273), .CP(n72), .CDN(n38), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(N1273), .CP(n57), .CDN(n25), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(N1273), .CP(n68), .CDN(n36), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(N1273), .CP(n70), .CDN(n41), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(N1273), .CP(n73), .CDN(n31), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(N1273), .CP(n68), .CDN(n32), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(N1273), .CP(n53), .CDN(n16), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(N1273), .CP(n45), .CDN(n40), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(N1273), .CP(n46), .CDN(n32), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(N1273), .CP(n48), .CDN(n6), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(N1273), .CP(n66), .CDN(n18), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(N1273), .CP(n57), .CDN(n24), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(N1273), .CP(n55), .CDN(n36), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(N1273), .CP(n52), .CDN(n9), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(N1273), .CP(n48), .CDN(n28), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(N1273), .CP(n42), .CDN(n2), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(N117), .E(N1999), .CP(n47), .CDN(n7), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(DataI[31]), .E(N1999), .CP(n69), .CDN(
        n11), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(DataI[30]), .E(N1999), .CP(n70), .CDN(
        n28), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(DataI[29]), .E(N1999), .CP(n67), .CDN(
        n28), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(DataI[28]), .E(N1999), .CP(n63), .CDN(
        n22), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(DataI[27]), .E(N1999), .CP(n42), .CDN(
        n25), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(DataI[26]), .E(N1999), .CP(n48), .CDN(
        n29), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(DataI[25]), .E(N1999), .CP(n69), .CDN(
        n14), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(DataI[24]), .E(N1999), .CP(n72), .CDN(
        n17), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(DataI[23]), .E(N1999), .CP(n71), .CDN(
        n29), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(DataI[22]), .E(N1999), .CP(n51), .CDN(
        n31), .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(DataI[21]), .E(N1999), .CP(n65), .CDN(n5), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(DataI[20]), .E(N1999), .CP(n66), .CDN(
        n34), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(DataI[19]), .E(N1999), .CP(n61), .CDN(
        n28), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(DataI[18]), .E(N1999), .CP(n69), .CDN(
        n29), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(DataI[17]), .E(N1999), .CP(n57), .CDN(
        n21), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(DataI[16]), .E(N1999), .CP(n73), .CDN(
        n24), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(DataI[15]), .E(N1999), .CP(n42), .CDN(
        n13), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(DataI[14]), .E(N1999), .CP(n56), .CDN(n3), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(DataI[13]), .E(N1999), .CP(ChipClock), 
        .CDN(n2), .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(DataI[12]), .E(N1999), .CP(n72), .CDN(n7), .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(DataI[11]), .E(N1999), .CP(n67), .CDN(n5), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(DataI[10]), .E(N1999), .CP(n59), .CDN(n4), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(DataI[9]), .E(N1999), .CP(n56), .CDN(n6), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(DataI[8]), .E(N1999), .CP(n57), .CDN(n16), 
        .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(DataI[7]), .E(N1999), .CP(n52), .CDN(n39), 
        .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(DataI[6]), .E(N1999), .CP(n72), .CDN(n13), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(DataI[5]), .E(N1999), .CP(n67), .CDN(n7), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(DataI[4]), .E(N1999), .CP(n48), .CDN(n20), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(DataI[3]), .E(N1999), .CP(n56), .CDN(n37), 
        .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(DataI[2]), .E(N1999), .CP(n54), .CDN(n4), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(DataI[1]), .E(N1999), .CP(n51), .CDN(n41), 
        .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(DataI[0]), .E(N1999), .CP(n44), .CDN(n4), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N117), .E(N1900), .CP(n47), .CDN(n6), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(N1900), .CP(n63), .CDN(
        n39), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(N1900), .CP(n72), .CDN(n4), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(DataI[29]), .E(N1900), .CP(n52), .CDN(n9), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(N1900), .CP(n51), .CDN(
        n10), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(N1900), .CP(n67), .CDN(
        n13), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(N1900), .CP(n72), .CDN(
        n12), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(N1900), .CP(n71), .CDN(
        n14), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(N1900), .CP(n61), .CDN(
        n15), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(N1900), .CP(n60), .CDN(
        n26), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(DataI[22]), .E(N1900), .CP(n59), .CDN(n8), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(N1900), .CP(n73), .CDN(
        n31), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(DataI[20]), .E(N1900), .CP(n68), .CDN(
        n28), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(N1900), .CP(n52), .CDN(
        n29), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(N1900), .CP(n58), .CDN(n2), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(DataI[17]), .E(N1900), .CP(n62), .CDN(
        n27), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(N1900), .CP(n55), .CDN(
        n23), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(DataI[15]), .E(N1900), .CP(n66), .CDN(
        n31), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(N1900), .CP(n61), .CDN(
        n17), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(N1900), .CP(n61), .CDN(n5), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(DataI[12]), .E(N1900), .CP(n49), .CDN(
        n25), .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(N1900), .CP(n45), .CDN(
        n20), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(DataI[10]), .E(N1900), .CP(n46), .CDN(n6), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(DataI[9]), .E(N1900), .CP(n54), .CDN(n36), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(N1900), .CP(n62), .CDN(n2), 
        .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(DataI[7]), .E(N1900), .CP(n51), .CDN(n4), 
        .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(DataI[6]), .E(N1900), .CP(n67), .CDN(n19), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(DataI[5]), .E(N1900), .CP(n57), .CDN(n2), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(DataI[4]), .E(N1900), .CP(n47), .CDN(n22), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(DataI[3]), .E(N1900), .CP(n56), .CDN(n5), 
        .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(DataI[2]), .E(N1900), .CP(n54), .CDN(n19), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(DataI[1]), .E(N1900), .CP(n50), .CDN(n7), 
        .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(DataI[0]), .E(N1900), .CP(n44), .CDN(n4), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(N117), .E(N1867), .CP(n47), .CDN(n6), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(DataI[31]), .E(N1867), .CP(ChipClock), 
        .CDN(n32), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(DataI[30]), .E(N1867), .CP(n68), .CDN(n7), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(N1867), .CP(n73), .CDN(
        n13), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(DataI[28]), .E(N1867), .CP(n52), .CDN(
        n10), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(DataI[27]), .E(N1867), .CP(n73), .CDN(
        n174), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(DataI[26]), .E(N1867), .CP(n62), .CDN(
        n23), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(DataI[25]), .E(N1867), .CP(n44), .CDN(
        n22), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(DataI[24]), .E(N1867), .CP(n71), .CDN(
        n11), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(DataI[23]), .E(N1867), .CP(n55), .CDN(n8), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(DataI[22]), .E(N1867), .CP(n63), .CDN(n8), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(DataI[21]), .E(N1867), .CP(n64), .CDN(
        n19), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(N1867), .CP(n50), .CDN(
        n24), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(DataI[19]), .E(N1867), .CP(n69), .CDN(
        n25), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(DataI[18]), .E(N1867), .CP(n70), .CDN(
        n28), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(N1867), .CP(n65), .CDN(
        n39), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(DataI[16]), .E(N1867), .CP(n51), .CDN(n7), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(N1867), .CP(n59), .CDN(n8), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(DataI[14]), .E(N1867), .CP(n59), .CDN(n8), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(DataI[13]), .E(N1867), .CP(n52), .CDN(
        n38), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(DataI[12]), .E(N1867), .CP(n71), .CDN(n9), .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(DataI[11]), .E(N1867), .CP(n44), .CDN(
        n27), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(N1867), .CP(n61), .CDN(
        n17), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(DataI[9]), .E(N1867), .CP(n49), .CDN(n27), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(DataI[8]), .E(N1867), .CP(n61), .CDN(n24), 
        .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(N1867), .CP(n47), .CDN(n6), 
        .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(DataI[6]), .E(N1867), .CP(n51), .CDN(n21), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(DataI[5]), .E(N1867), .CP(n56), .CDN(n4), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(DataI[4]), .E(N1867), .CP(n51), .CDN(n13), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(N1867), .CP(n56), .CDN(n24), 
        .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(DataI[2]), .E(N1867), .CP(n53), .CDN(n12), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(N1867), .CP(n50), .CDN(n2), 
        .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(DataI[0]), .E(N1867), .CP(n44), .CDN(n3), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N117), .E(N1768), .CP(n47), .CDN(n6), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(DataI[31]), .E(N1768), .CP(n49), .CDN(
        n14), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(DataI[30]), .E(N1768), .CP(n48), .CDN(
        n14), .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(DataI[29]), .E(N1768), .CP(n69), .CDN(
        n14), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(DataI[28]), .E(N1768), .CP(n58), .CDN(
        n14), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(DataI[27]), .E(N1768), .CP(n43), .CDN(
        n14), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(DataI[26]), .E(N1768), .CP(n49), .CDN(
        n14), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(DataI[25]), .E(N1768), .CP(n44), .CDN(
        n13), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(DataI[24]), .E(N1768), .CP(n54), .CDN(
        n13), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(DataI[23]), .E(N1768), .CP(n61), .CDN(
        n13), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(DataI[22]), .E(N1768), .CP(n49), .CDN(
        n13), .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(DataI[21]), .E(N1768), .CP(n60), .CDN(
        n13), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(DataI[20]), .E(N1768), .CP(n61), .CDN(
        n13), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(DataI[19]), .E(N1768), .CP(n56), .CDN(
        n13), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(DataI[18]), .E(N1768), .CP(n58), .CDN(
        n13), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(DataI[17]), .E(N1768), .CP(n54), .CDN(
        n13), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(DataI[16]), .E(N1768), .CP(n43), .CDN(
        n13), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(DataI[15]), .E(N1768), .CP(n51), .CDN(
        n13), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(DataI[14]), .E(N1768), .CP(n45), .CDN(
        n12), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(DataI[13]), .E(N1768), .CP(n71), .CDN(
        n12), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(DataI[12]), .E(N1768), .CP(n59), .CDN(
        n12), .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(DataI[11]), .E(N1768), .CP(n47), .CDN(
        n12), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(DataI[10]), .E(N1768), .CP(n60), .CDN(
        n12), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(DataI[9]), .E(N1768), .CP(n42), .CDN(n12), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(DataI[8]), .E(N1768), .CP(n69), .CDN(n12), 
        .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(DataI[7]), .E(N1768), .CP(n48), .CDN(n15), 
        .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(DataI[6]), .E(N1768), .CP(n56), .CDN(n20), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(DataI[5]), .E(N1768), .CP(n53), .CDN(n5), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(DataI[4]), .E(N1768), .CP(n52), .CDN(n12), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(DataI[3]), .E(N1768), .CP(n59), .CDN(n6), 
        .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(DataI[2]), .E(N1768), .CP(n53), .CDN(n17), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(DataI[1]), .E(N1768), .CP(n50), .CDN(n3), 
        .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(DataI[0]), .E(N1768), .CP(n43), .CDN(n3), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N117), .E(N1735), .CP(n46), .CDN(n6), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(N1735), .CP(n54), .CDN(
        n32), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(N1735), .CP(n53), .CDN(
        n174), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(N1735), .CP(n49), .CDN(n6), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(N1735), .CP(n65), .CDN(
        n22), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(N1735), .CP(n71), .CDN(
        n35), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(N1735), .CP(n64), .CDN(n8), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(N1735), .CP(n62), .CDN(
        n33), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(N1735), .CP(n63), .CDN(
        n29), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(N1735), .CP(n59), .CDN(
        n32), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(N1735), .CP(n60), .CDN(
        n40), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(N1735), .CP(n63), .CDN(
        n37), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(N1735), .CP(n52), .CDN(
        n33), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(N1735), .CP(n57), .CDN(
        n34), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(N1735), .CP(n58), .CDN(
        n12), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(N1735), .CP(n56), .CDN(
        n30), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(N1735), .CP(n66), .CDN(n7), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(N1735), .CP(n74), .CDN(
        n26), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(N1735), .CP(n43), .CDN(
        n11), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(N1735), .CP(n61), .CDN(
        n24), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(N1735), .CP(n42), .CDN(
        n27), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(N1735), .CP(n42), .CDN(
        n36), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(N1735), .CP(n45), .CDN(
        n38), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(N1735), .CP(n72), .CDN(n35), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(N1735), .CP(n74), .CDN(n15), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(N1735), .CP(n72), .CDN(n12), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(N1735), .CP(n68), .CDN(n23), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(N1735), .CP(n54), .CDN(n21), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(N1735), .CP(n50), .CDN(n14), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(N1735), .CP(n60), .CDN(n18), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(N1735), .CP(n53), .CDN(n28), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(N1735), .CP(n50), .CDN(n31), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(N1735), .CP(n43), .CDN(n3), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N117), .E(N1636), .CP(n46), .CDN(n6), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(N1636), .CP(n43), .CDN(
        n36), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(N1636), .CP(n63), .CDN(
        n41), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(N1636), .CP(n51), .CDN(
        n26), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(N1636), .CP(n47), .CDN(
        n19), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(N1636), .CP(n48), .CDN(
        n36), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(N1636), .CP(n46), .CDN(
        n19), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(N1636), .CP(n45), .CDN(
        n40), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(N1636), .CP(n67), .CDN(
        n20), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(N1636), .CP(n74), .CDN(
        n18), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(N1636), .CP(n72), .CDN(
        n40), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(N1636), .CP(n54), .CDN(
        n18), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(N1636), .CP(n45), .CDN(n9), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(N1636), .CP(n60), .CDN(
        n17), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(N1636), .CP(n56), .CDN(n6), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(N1636), .CP(n56), .CDN(
        n29), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(N1636), .CP(n51), .CDN(
        n14), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(DataI[15]), .E(N1636), .CP(n42), .CDN(
        n24), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(DataI[14]), .E(N1636), .CP(n61), .CDN(
        n11), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(N1636), .CP(n65), .CDN(
        n39), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(N1636), .CP(n71), .CDN(
        n33), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(N1636), .CP(n64), .CDN(
        n30), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(N1636), .CP(n62), .CDN(
        n11), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(N1636), .CP(n69), .CDN(n174), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(N1636), .CP(n70), .CDN(n40), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(DataI[7]), .E(N1636), .CP(n62), .CDN(n13), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(DataI[6]), .E(N1636), .CP(n69), .CDN(n8), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(DataI[5]), .E(N1636), .CP(n43), .CDN(n20), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(N1636), .CP(n68), .CDN(n11), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(N1636), .CP(n72), .CDN(n33), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(N1636), .CP(n53), .CDN(n33), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(N1636), .CP(n49), .CDN(n22), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(N1636), .CP(n43), .CDN(n3), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N117), .E(N1603), .CP(n46), .CDN(n6), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(N1603), .CP(ChipClock), 
        .CDN(n15), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(N1603), .CP(ChipClock), 
        .CDN(n14), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(N1603), .CP(n72), .CDN(
        n12), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(N1603), .CP(n67), .CDN(
        n13), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(N1603), .CP(n55), .CDN(
        n10), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(N1603), .CP(n65), .CDN(n9), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(N1603), .CP(n72), .CDN(n3), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(N1603), .CP(n65), .CDN(
        n25), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(N1603), .CP(n57), .CDN(
        n11), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(N1603), .CP(n73), .CDN(
        n21), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(N1603), .CP(n68), .CDN(
        n20), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(N1603), .CP(n69), .CDN(
        n23), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(N1603), .CP(n70), .CDN(
        n22), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(N1603), .CP(n63), .CDN(
        n16), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(N1603), .CP(n69), .CDN(
        n18), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(N1603), .CP(n73), .CDN(
        n17), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(DataI[15]), .E(N1603), .CP(n50), .CDN(
        n19), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(DataI[14]), .E(N1603), .CP(n71), .CDN(
        n20), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(N1603), .CP(n66), .CDN(
        n25), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(N1603), .CP(n57), .CDN(
        n13), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(N1603), .CP(n59), .CDN(
        n25), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(N1603), .CP(n56), .CDN(
        n24), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(N1603), .CP(n58), .CDN(n27), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(N1603), .CP(n53), .CDN(n26), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(DataI[7]), .E(N1603), .CP(n64), .CDN(n10), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(DataI[6]), .E(N1603), .CP(n70), .CDN(n12), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(DataI[5]), .E(N1603), .CP(n44), .CDN(n23), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(N1603), .CP(n54), .CDN(n3), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(N1603), .CP(n46), .CDN(n34), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(N1603), .CP(n53), .CDN(n2), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(N1603), .CP(n49), .CDN(n23), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(N1603), .CP(n43), .CDN(n3), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N117), .E(N1504), .CP(n46), .CDN(n5), .Q(
        \Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(N1504), .CP(n70), .CDN(n18), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(N1504), .CP(n73), .CDN(n11), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(N1504), .CP(n73), .CDN(n25), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(N1504), .CP(n68), .CDN(n20), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(N1504), .CP(n65), .CDN(n23), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(N1504), .CP(n45), .CDN(n22), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(N1504), .CP(n52), .CDN(n18), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(N1504), .CP(n65), .CDN(n15), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(N1504), .CP(n63), .CDN(n14), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(N1504), .CP(n72), .CDN(n12), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(N1504), .CP(n68), .CDN(n13), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(N1504), .CP(n58), .CDN(n10), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(N1504), .CP(n47), .CDN(n38), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(N1504), .CP(n66), .CDN(n29), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(N1504), .CP(n65), .CDN(n23), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(N1504), .CP(n59), .CDN(n5), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(DataI[15]), .E(N1504), .CP(n60), .CDN(n21), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(N1504), .CP(n61), .CDN(n37), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(N1504), .CP(n59), .CDN(n36), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(N1504), .CP(n52), .CDN(n39), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(N1504), .CP(n67), .CDN(n38), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(N1504), .CP(n58), .CDN(n10), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(N1504), .CP(n49), .CDN(n41), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(N1504), .CP(n71), .CDN(n22), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(DataI[7]), .E(N1504), .CP(n71), .CDN(n40), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(N1504), .CP(n60), .CDN(n4), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(N1504), .CP(n58), .CDN(n16), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(N1504), .CP(n69), .CDN(n25), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(N1504), .CP(n67), .CDN(n26), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(N1504), .CP(n52), .CDN(n8), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(N1504), .CP(n49), .CDN(n15), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(N1504), .CP(n43), .CDN(n2), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N117), .E(N1471), .CP(n46), .CDN(n5), .Q(
        \Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(N1471), .CP(n50), .CDN(n36), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(N1471), .CP(n44), .CDN(n30), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(N1471), .CP(n73), .CDN(n11), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(N1471), .CP(n68), .CDN(n9), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(N1471), .CP(n69), .CDN(n15), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(N1471), .CP(n70), .CDN(n32), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(N1471), .CP(n48), .CDN(n28), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(N1471), .CP(n66), .CDN(n33), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(N1471), .CP(n54), .CDN(n12), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(N1471), .CP(n53), .CDN(n37), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(N1471), .CP(n61), .CDN(n38), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(N1471), .CP(n46), .CDN(n39), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(N1471), .CP(n55), .CDN(n39), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(N1471), .CP(n47), .CDN(n41), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(N1471), .CP(n54), .CDN(n34), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(N1471), .CP(n66), .CDN(n27), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(N1471), .CP(n56), .CDN(n33), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(N1471), .CP(n65), .CDN(n34), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(N1471), .CP(n49), .CDN(n30), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(N1471), .CP(n51), .CDN(n14), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(N1471), .CP(n52), .CDN(n31), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(N1471), .CP(n48), .CDN(n3), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(N1471), .CP(n47), .CDN(n29), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(N1471), .CP(n54), .CDN(n22), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(N1471), .CP(n73), .CDN(n29), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(N1471), .CP(n72), .CDN(n31), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(N1471), .CP(n65), .CDN(n32), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(N1471), .CP(n70), .CDN(n16), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(N1471), .CP(n45), .CDN(n19), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(N1471), .CP(n52), .CDN(n11), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(N1471), .CP(n49), .CDN(n11), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(N1471), .CP(n42), .CDN(n2), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N117), .E(N1372), .CP(n45), .CDN(n5), .Q(
        \Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(N1372), .CP(n49), .CDN(n32), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(N1372), .CP(n53), .CDN(n16), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(N1372), .CP(n45), .CDN(n34), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(N1372), .CP(n46), .CDN(n35), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(N1372), .CP(n44), .CDN(n3), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(N1372), .CP(n43), .CDN(n3), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(N1372), .CP(n48), .CDN(n5), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(N1372), .CP(n47), .CDN(n19), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(N1372), .CP(n51), .CDN(n9), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(N1372), .CP(n52), .CDN(n36), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(N1372), .CP(n72), .CDN(n33), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(N1372), .CP(n45), .CDN(n20), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(N1372), .CP(n57), .CDN(n33), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(N1372), .CP(n56), .CDN(n10), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(N1372), .CP(n55), .CDN(n41), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(N1372), .CP(n44), .CDN(n9), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(N1372), .CP(n54), .CDN(n8), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(N1372), .CP(n53), .CDN(n30), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(N1372), .CP(n63), .CDN(n31), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(N1372), .CP(n60), .CDN(n32), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(N1372), .CP(n56), .CDN(n10), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(N1372), .CP(n59), .CDN(n38), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(N1372), .CP(n52), .CDN(n37), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(N1372), .CP(n58), .CDN(n41), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(N1372), .CP(n72), .CDN(n39), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(N1372), .CP(n67), .CDN(n33), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(N1372), .CP(n71), .CDN(n8), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(N1372), .CP(n61), .CDN(n29), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(N1372), .CP(n55), .CDN(n38), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(N1372), .CP(n52), .CDN(n31), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(N1372), .CP(n49), .CDN(n24), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(N1372), .CP(n42), .CDN(n2), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N117), .E(N1339), .CP(n45), .CDN(n5), .Q(
        \Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(N1339), .CP(n50), .CDN(n8), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(N1339), .CP(n49), .CDN(n27), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(N1339), .CP(n68), .CDN(n41), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(N1339), .CP(n67), .CDN(n32), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(N1339), .CP(n69), .CDN(n37), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(N1339), .CP(n44), .CDN(n36), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(N1339), .CP(n59), .CDN(n39), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(N1339), .CP(n59), .CDN(n38), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(N1339), .CP(n52), .CDN(n33), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(N1339), .CP(n43), .CDN(n40), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(N1339), .CP(n47), .CDN(n26), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(N1339), .CP(n67), .CDN(n19), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(N1339), .CP(n64), .CDN(n13), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(N1339), .CP(n43), .CDN(n37), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(N1339), .CP(n70), .CDN(n34), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(N1339), .CP(n49), .CDN(n14), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(N1339), .CP(n70), .CDN(n35), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(N1339), .CP(n50), .CDN(n26), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(N1339), .CP(n49), .CDN(
        n174), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(N1339), .CP(n51), .CDN(n36), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(N1339), .CP(n52), .CDN(n40), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(N1339), .CP(n48), .CDN(n38), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(N1339), .CP(n47), .CDN(n30), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(N1339), .CP(n54), .CDN(n174), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(N1339), .CP(n67), .CDN(n37), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(N1339), .CP(n44), .CDN(n34), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(N1339), .CP(n68), .CDN(n38), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(N1339), .CP(n57), .CDN(n28), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(N1339), .CP(n55), .CDN(n41), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(N1339), .CP(n52), .CDN(n28), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(N1339), .CP(n49), .CDN(n31), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(N1339), .CP(n42), .CDN(n2), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N117), .E(N1240), .CP(n45), .CDN(n5), .Q(
        \Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(N1240), .CP(n67), .CDN(n30), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(N1240), .CP(n45), .CDN(n37), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(N1240), .CP(n57), .CDN(
        n174), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(N1240), .CP(n50), .CDN(n40), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(N1240), .CP(n56), .CDN(n6), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N1240), .CP(n71), .CDN(n2), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(N1240), .CP(n66), .CDN(n37), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(N1240), .CP(n57), .CDN(n25), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(N1240), .CP(n56), .CDN(n39), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(N1240), .CP(n55), .CDN(n35), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(N1240), .CP(n48), .CDN(n6), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(N1240), .CP(n54), .CDN(n32), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(N1240), .CP(n53), .CDN(n32), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(N1240), .CP(n50), .CDN(n31), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(N1240), .CP(n49), .CDN(n30), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(N1240), .CP(n51), .CDN(n15), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(N1240), .CP(n66), .CDN(n33), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(N1240), .CP(n64), .CDN(n31), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(N1240), .CP(n53), .CDN(n40), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(N1240), .CP(n55), .CDN(n38), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(N1240), .CP(n62), .CDN(n28), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(N1240), .CP(n51), .CDN(n5), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(N1240), .CP(n72), .CDN(n20), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(N1240), .CP(n56), .CDN(n37), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(N1240), .CP(n58), .CDN(n36), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(N1240), .CP(n48), .CDN(n30), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(N1240), .CP(n73), .CDN(n7), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(N1240), .CP(n57), .CDN(n3), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(N1240), .CP(n55), .CDN(n7), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(N1240), .CP(n52), .CDN(n29), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(N1240), .CP(n48), .CDN(n23), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(N1240), .CP(n42), .CDN(n2), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(N117), .E(N2263), .CP(n48), .CDN(n7), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(N2263), .CP(n64), .CDN(
        n16), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(N2263), .CP(n70), .CDN(
        n16), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(N2263), .CP(n62), .CDN(
        n16), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(N2263), .CP(n60), .CDN(
        n16), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(N2263), .CP(n71), .CDN(
        n16), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(N2263), .CP(n42), .CDN(
        n16), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(N2263), .CP(n53), .CDN(
        n16), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(N2263), .CP(n50), .CDN(
        n16), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(N2263), .CP(n57), .CDN(
        n15), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(N2263), .CP(n60), .CDN(
        n15), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(N2263), .CP(n70), .CDN(
        n15), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(N2263), .CP(n42), .CDN(
        n15), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(N2263), .CP(n44), .CDN(
        n15), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(N2263), .CP(n61), .CDN(
        n15), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(N2263), .CP(n55), .CDN(
        n15), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(N2263), .CP(n53), .CDN(
        n15), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(N2263), .CP(n73), .CDN(
        n15), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(N2263), .CP(n58), .CDN(
        n15), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(N2263), .CP(n65), .CDN(
        n15), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(N2263), .CP(n60), .CDN(
        n14), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(N2263), .CP(n56), .CDN(
        n14), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(N2263), .CP(ChipClock), 
        .CDN(n14), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(N2263), .CP(n72), .CDN(n14), 
        .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(N2263), .CP(n67), .CDN(n14), 
        .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(N2263), .CP(n73), .CDN(n41), 
        .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(DataI[6]), .E(N2263), .CP(n48), .CDN(n10), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(N2263), .CP(n47), .CDN(n41), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(N2263), .CP(n61), .CDN(n10), 
        .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(N2263), .CP(n57), .CDN(n33), 
        .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(N2263), .CP(n55), .CDN(n13), 
        .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(N2263), .CP(n51), .CDN(n20), 
        .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(N2263), .CP(n45), .CDN(n5), 
        .Q(\Storage[31][0] ) );
  EDFCNQD1 DreadyReg_reg ( .D(Read), .E(ChipEna), .CP(n71), .CDN(n20), .Q(
        DreadyReg) );
  EDFCNQD1 ParityReg_reg ( .D(N116), .E(N2264), .CP(n42), .CDN(n2), .Q(
        ParityErr) );
  EDFCNQD1 \DataOreg_reg[31]  ( .D(N82), .E(N2327), .CP(n53), .CDN(n31), .Q(
        N2330) );
  EDFCNQD1 \DataOreg_reg[30]  ( .D(N83), .E(N2327), .CP(n55), .CDN(n16), .Q(
        N2333) );
  EDFCNQD1 \DataOreg_reg[29]  ( .D(N84), .E(N2327), .CP(n60), .CDN(n15), .Q(
        N2336) );
  EDFCNQD1 \DataOreg_reg[28]  ( .D(N85), .E(N2327), .CP(n43), .CDN(n33), .Q(
        N2339) );
  EDFCNQD1 \DataOreg_reg[27]  ( .D(N86), .E(N2327), .CP(n64), .CDN(n31), .Q(
        N2342) );
  EDFCNQD1 \DataOreg_reg[26]  ( .D(N87), .E(N2327), .CP(n65), .CDN(n31), .Q(
        N2345) );
  EDFCNQD1 \DataOreg_reg[25]  ( .D(N88), .E(N2327), .CP(n59), .CDN(n27), .Q(
        N2348) );
  EDFCNQD1 \DataOreg_reg[24]  ( .D(N89), .E(N2327), .CP(n42), .CDN(n30), .Q(
        N2351) );
  EDFCNQD1 \DataOreg_reg[23]  ( .D(N90), .E(N2327), .CP(n51), .CDN(n9), .Q(
        N2354) );
  EDFCNQD1 \DataOreg_reg[22]  ( .D(N91), .E(N2327), .CP(n58), .CDN(n24), .Q(
        N2357) );
  EDFCNQD1 \DataOreg_reg[21]  ( .D(N92), .E(N2327), .CP(n55), .CDN(n40), .Q(
        N2360) );
  EDFCNQD1 \DataOreg_reg[20]  ( .D(N93), .E(N2327), .CP(n68), .CDN(n13), .Q(
        N2363) );
  EDFCNQD1 \DataOreg_reg[19]  ( .D(N94), .E(N2327), .CP(n46), .CDN(n6), .Q(
        N2366) );
  EDFCNQD1 \DataOreg_reg[18]  ( .D(N95), .E(N2327), .CP(n71), .CDN(n16), .Q(
        N2369) );
  EDFCNQD1 \DataOreg_reg[17]  ( .D(N96), .E(N2327), .CP(n54), .CDN(n18), .Q(
        N2372) );
  EDFCNQD1 \DataOreg_reg[16]  ( .D(N97), .E(N2327), .CP(n53), .CDN(n17), .Q(
        N2375) );
  EDFCNQD1 \DataOreg_reg[15]  ( .D(N98), .E(N2327), .CP(n56), .CDN(n19), .Q(
        N2378) );
  EDFCNQD1 \DataOreg_reg[14]  ( .D(N99), .E(N2327), .CP(n67), .CDN(n21), .Q(
        N2381) );
  EDFCNQD1 \DataOreg_reg[13]  ( .D(N100), .E(N2327), .CP(n43), .CDN(n36), .Q(
        N2384) );
  EDFCNQD1 \DataOreg_reg[12]  ( .D(N101), .E(N2327), .CP(n66), .CDN(n39), .Q(
        N2387) );
  EDFCNQD1 \DataOreg_reg[11]  ( .D(N102), .E(N2327), .CP(n73), .CDN(n41), .Q(
        N2390) );
  EDFCNQD1 \DataOreg_reg[10]  ( .D(N103), .E(N2327), .CP(n70), .CDN(n40), .Q(
        N2393) );
  EDFCNQD1 \DataOreg_reg[9]  ( .D(N104), .E(N2327), .CP(n65), .CDN(n27), .Q(
        N2396) );
  EDFCNQD1 \DataOreg_reg[8]  ( .D(N105), .E(N2327), .CP(n66), .CDN(n21), .Q(
        N2399) );
  EDFCNQD1 \DataOreg_reg[7]  ( .D(N106), .E(N2327), .CP(n47), .CDN(n38), .Q(
        N2402) );
  EDFCNQD1 \DataOreg_reg[6]  ( .D(N107), .E(N2327), .CP(n51), .CDN(n35), .Q(
        N2405) );
  EDFCNQD1 \DataOreg_reg[5]  ( .D(N108), .E(N2327), .CP(n64), .CDN(n26), .Q(
        N2408) );
  EDFCNQD1 \DataOreg_reg[4]  ( .D(N109), .E(N2327), .CP(n57), .CDN(n10), .Q(
        N2411) );
  EDFCNQD1 \DataOreg_reg[3]  ( .D(N110), .E(N2327), .CP(n55), .CDN(n22), .Q(
        N2414) );
  EDFCNQD1 \DataOreg_reg[2]  ( .D(N111), .E(N2327), .CP(n51), .CDN(n4), .Q(
        N2417) );
  EDFCNQD1 \DataOreg_reg[1]  ( .D(N112), .E(N2327), .CP(n48), .CDN(n16), .Q(
        N2420) );
  EDFCNQD1 \DataOreg_reg[0]  ( .D(N113), .E(N2327), .CP(n42), .CDN(n2), .Q(
        N2423) );
  INVD3 U2 ( .I(n1), .ZN(N2327) );
  OA21D1 U3 ( .A1(n568), .A2(n569), .B(n570), .Z(n1) );
  INVD0 U4 ( .I(N75), .ZN(n89) );
  BUFFD0 U5 ( .I(ChipClock), .Z(n74) );
  NR3D2 U6 ( .A1(n568), .A2(Read), .A3(n569), .ZN(N2328) );
  NR2D2P5 U7 ( .A1(n579), .A2(n580), .ZN(N1768) );
  ND3D1 U8 ( .A1(N2328), .A2(n581), .A3(N79), .ZN(n580) );
  NR2D2P5 U9 ( .A1(n572), .A2(n582), .ZN(N1735) );
  ND3D1 U10 ( .A1(N2328), .A2(n583), .A3(N78), .ZN(n582) );
  NR2D2P5 U11 ( .A1(n578), .A2(n580), .ZN(N1801) );
  NR2D2P5 U12 ( .A1(n573), .A2(n582), .ZN(N1702) );
  NR2D2P5 U13 ( .A1(n577), .A2(n580), .ZN(N1834) );
  NR2D2P5 U14 ( .A1(n574), .A2(n582), .ZN(N1669) );
  NR2D2P5 U15 ( .A1(n576), .A2(n580), .ZN(N1867) );
  NR2D2P5 U16 ( .A1(n575), .A2(n582), .ZN(N1636) );
  NR2D2P5 U17 ( .A1(n575), .A2(n580), .ZN(N1900) );
  NR2D2P5 U18 ( .A1(n576), .A2(n582), .ZN(N1603) );
  NR2D2P5 U19 ( .A1(n574), .A2(n580), .ZN(N1933) );
  NR2D2P5 U20 ( .A1(n577), .A2(n582), .ZN(N1570) );
  NR2D2P5 U21 ( .A1(n573), .A2(n580), .ZN(N1966) );
  NR2D2P5 U22 ( .A1(n578), .A2(n582), .ZN(N1537) );
  NR2D2P5 U23 ( .A1(n572), .A2(n580), .ZN(N1999) );
  NR2D2P5 U24 ( .A1(n579), .A2(n582), .ZN(N1504) );
  NR2D2P5 U25 ( .A1(n571), .A2(n579), .ZN(N2032) );
  ND3D1 U26 ( .A1(N78), .A2(N2328), .A3(N79), .ZN(n571) );
  NR2D2P5 U27 ( .A1(n572), .A2(n584), .ZN(N1471) );
  ND3D1 U28 ( .A1(n581), .A2(n583), .A3(N2328), .ZN(n584) );
  NR2D2P5 U29 ( .A1(n571), .A2(n578), .ZN(N2065) );
  NR2D2P5 U30 ( .A1(n573), .A2(n584), .ZN(N1438) );
  NR2D2P5 U31 ( .A1(n571), .A2(n577), .ZN(N2098) );
  NR2D2P5 U32 ( .A1(n574), .A2(n584), .ZN(N1405) );
  NR2D2P5 U33 ( .A1(n571), .A2(n576), .ZN(N2131) );
  NR2D2P5 U34 ( .A1(n575), .A2(n584), .ZN(N1372) );
  NR2D2P5 U35 ( .A1(n571), .A2(n575), .ZN(N2164) );
  NR2D2P5 U36 ( .A1(n576), .A2(n584), .ZN(N1339) );
  NR2D2P5 U37 ( .A1(n571), .A2(n574), .ZN(N2197) );
  NR2D2P5 U38 ( .A1(n577), .A2(n584), .ZN(N1306) );
  NR2D2P5 U39 ( .A1(n571), .A2(n573), .ZN(N2230) );
  NR2D2P5 U40 ( .A1(n578), .A2(n584), .ZN(N1273) );
  NR2D2P5 U41 ( .A1(n571), .A2(n572), .ZN(N2263) );
  NR2D2P5 U42 ( .A1(n579), .A2(n584), .ZN(N1240) );
  INVD0 U43 ( .I(n570), .ZN(N2264) );
  XOR3D1 U44 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n585), .Z(N117) );
  BUFFD1 U45 ( .I(n62), .Z(n52) );
  BUFFD1 U46 ( .I(n63), .Z(n49) );
  BUFFD1 U47 ( .I(n61), .Z(n53) );
  BUFFD1 U48 ( .I(n63), .Z(n50) );
  BUFFD1 U49 ( .I(n64), .Z(n47) );
  BUFFD1 U50 ( .I(n59), .Z(n56) );
  BUFFD1 U51 ( .I(n61), .Z(n54) );
  BUFFD1 U52 ( .I(n62), .Z(n51) );
  BUFFD1 U53 ( .I(n60), .Z(n55) );
  BUFFD1 U54 ( .I(n59), .Z(n57) );
  BUFFD1 U55 ( .I(n64), .Z(n48) );
  BUFFD1 U56 ( .I(n65), .Z(n46) );
  BUFFD1 U57 ( .I(n66), .Z(n43) );
  BUFFD1 U58 ( .I(n66), .Z(n44) );
  BUFFD1 U59 ( .I(n65), .Z(n45) );
  BUFFD1 U60 ( .I(n69), .Z(n63) );
  BUFFD1 U61 ( .I(n70), .Z(n61) );
  BUFFD1 U62 ( .I(n69), .Z(n62) );
  BUFFD1 U63 ( .I(n70), .Z(n60) );
  BUFFD1 U64 ( .I(n70), .Z(n59) );
  BUFFD1 U65 ( .I(n46), .Z(n58) );
  BUFFD1 U66 ( .I(n69), .Z(n64) );
  BUFFD1 U67 ( .I(n33), .Z(n13) );
  BUFFD1 U68 ( .I(n34), .Z(n11) );
  BUFFD1 U69 ( .I(n33), .Z(n12) );
  BUFFD1 U70 ( .I(n34), .Z(n8) );
  BUFFD1 U71 ( .I(n34), .Z(n9) );
  BUFFD1 U72 ( .I(n34), .Z(n10) );
  BUFFD1 U73 ( .I(n34), .Z(n29) );
  BUFFD1 U74 ( .I(n31), .Z(n28) );
  BUFFD1 U75 ( .I(n30), .Z(n26) );
  BUFFD1 U76 ( .I(n30), .Z(n27) );
  BUFFD1 U77 ( .I(n30), .Z(n24) );
  BUFFD1 U78 ( .I(n30), .Z(n25) );
  BUFFD1 U79 ( .I(n31), .Z(n22) );
  BUFFD1 U80 ( .I(n31), .Z(n23) );
  BUFFD1 U81 ( .I(n32), .Z(n19) );
  BUFFD1 U82 ( .I(n31), .Z(n20) );
  BUFFD1 U83 ( .I(n31), .Z(n21) );
  BUFFD1 U84 ( .I(n32), .Z(n17) );
  BUFFD1 U85 ( .I(n32), .Z(n18) );
  BUFFD1 U86 ( .I(n33), .Z(n14) );
  BUFFD1 U87 ( .I(n33), .Z(n15) );
  BUFFD1 U88 ( .I(n32), .Z(n16) );
  INVD1 U89 ( .I(n89), .ZN(n85) );
  INVD1 U90 ( .I(n88), .ZN(n86) );
  INVD1 U91 ( .I(n89), .ZN(n81) );
  INVD1 U92 ( .I(n89), .ZN(n82) );
  INVD1 U93 ( .I(n89), .ZN(n83) );
  INVD1 U94 ( .I(n88), .ZN(n84) );
  INVD1 U95 ( .I(n89), .ZN(n80) );
  INVD1 U96 ( .I(n88), .ZN(n79) );
  INVD1 U97 ( .I(n88), .ZN(n78) );
  INVD1 U98 ( .I(n88), .ZN(n77) );
  INVD1 U99 ( .I(n88), .ZN(n76) );
  INVD1 U100 ( .I(n88), .ZN(n75) );
  INVD1 U101 ( .I(n89), .ZN(n87) );
  INVD1 U102 ( .I(n99), .ZN(n93) );
  INVD1 U103 ( .I(n99), .ZN(n94) );
  INVD1 U104 ( .I(n99), .ZN(n95) );
  INVD1 U105 ( .I(n99), .ZN(n96) );
  INVD1 U106 ( .I(n99), .ZN(n97) );
  INVD1 U107 ( .I(n99), .ZN(n90) );
  INVD1 U108 ( .I(n99), .ZN(n91) );
  INVD1 U109 ( .I(n99), .ZN(n92) );
  INVD1 U110 ( .I(n99), .ZN(n98) );
  BUFFD1 U111 ( .I(n67), .Z(n42) );
  BUFFD1 U112 ( .I(n68), .Z(n67) );
  BUFFD1 U113 ( .I(n68), .Z(n66) );
  BUFFD1 U114 ( .I(n68), .Z(n65) );
  BUFFD1 U115 ( .I(n71), .Z(n70) );
  BUFFD1 U116 ( .I(n71), .Z(n69) );
  BUFFD1 U117 ( .I(n36), .Z(n2) );
  BUFFD1 U118 ( .I(n36), .Z(n3) );
  BUFFD1 U119 ( .I(n35), .Z(n6) );
  BUFFD1 U120 ( .I(n35), .Z(n4) );
  BUFFD1 U121 ( .I(n35), .Z(n5) );
  BUFFD1 U122 ( .I(n35), .Z(n7) );
  BUFFD1 U123 ( .I(n89), .Z(n88) );
  BUFFD1 U124 ( .I(n73), .Z(n71) );
  BUFFD1 U125 ( .I(n72), .Z(n68) );
  BUFFD1 U126 ( .I(n73), .Z(n72) );
  BUFFD1 U127 ( .I(n38), .Z(n34) );
  BUFFD1 U128 ( .I(n28), .Z(n30) );
  BUFFD1 U129 ( .I(n39), .Z(n31) );
  BUFFD1 U130 ( .I(n38), .Z(n33) );
  BUFFD1 U131 ( .I(n39), .Z(n32) );
  INVD1 U132 ( .I(n105), .ZN(n101) );
  INVD1 U133 ( .I(n105), .ZN(n104) );
  INVD1 U134 ( .I(n105), .ZN(n103) );
  INVD1 U135 ( .I(n105), .ZN(n102) );
  BUFFD1 U136 ( .I(n40), .Z(n38) );
  BUFFD1 U137 ( .I(n40), .Z(n39) );
  BUFFD1 U138 ( .I(n74), .Z(n73) );
  BUFFD1 U139 ( .I(n37), .Z(n35) );
  BUFFD1 U140 ( .I(n37), .Z(n36) );
  INVD1 U141 ( .I(n105), .ZN(n100) );
  BUFFD1 U142 ( .I(n174), .Z(n40) );
  BUFFD1 U143 ( .I(n41), .Z(n37) );
  BUFFD1 U144 ( .I(n174), .Z(n41) );
  INVD1 U145 ( .I(N76), .ZN(n99) );
  MUX4ND0 U146 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n78), .S1(n96), .ZN(
        n558) );
  MUX4ND0 U147 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n79), .S1(n95), .ZN(n109) );
  MUX4ND0 U148 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n79), .S1(n98), .ZN(n122) );
  MUX4ND0 U149 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n80), .S1(n98), .ZN(n135) );
  MUX4ND0 U150 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n81), .S1(n98), .ZN(n181) );
  MUX4ND0 U151 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n85), .S1(n98), .ZN(n194) );
  MUX4ND0 U152 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n85), .S1(n98), .ZN(n207) );
  MUX4ND0 U153 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n86), .S1(n98), .ZN(n220) );
  MUX4ND0 U154 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n86), .S1(n98), .ZN(n233) );
  MUX4ND0 U155 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n85), .S1(n98), .ZN(n246) );
  MUX4ND0 U156 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n87), .S1(n98), .ZN(n259) );
  MUX4ND0 U157 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n78), .S1(n98), .ZN(
        n272) );
  MUX4ND0 U158 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n82), .S1(n98), .ZN(
        n285) );
  MUX4ND0 U159 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n80), .S1(n95), .ZN(
        n298) );
  MUX4ND0 U160 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n78), .S1(n98), .ZN(
        n311) );
  MUX4ND0 U161 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n77), .S1(n91), .ZN(
        n324) );
  MUX4ND0 U162 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n76), .S1(n92), .ZN(
        n337) );
  MUX4ND0 U163 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n75), .S1(n90), .ZN(
        n350) );
  MUX4ND0 U164 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n87), .S1(n93), .ZN(
        n363) );
  MUX4ND0 U165 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n75), .S1(n97), .ZN(
        n376) );
  MUX4ND0 U166 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n77), .S1(n96), .ZN(
        n389) );
  MUX4ND0 U167 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n79), .S1(n94), .ZN(
        n402) );
  MUX4ND0 U168 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n80), .S1(n93), .ZN(
        n415) );
  MUX4ND0 U169 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n83), .S1(n95), .ZN(
        n428) );
  MUX4ND0 U170 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n84), .S1(n98), .ZN(
        n441) );
  MUX4ND0 U171 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n80), .S1(N76), .ZN(
        n454) );
  MUX4ND0 U172 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n78), .S1(N76), .ZN(
        n467) );
  MUX4ND0 U173 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n75), .S1(N76), .ZN(
        n480) );
  MUX4ND0 U174 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n76), .S1(N76), .ZN(
        n493) );
  MUX4ND0 U175 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n77), .S1(N76), .ZN(
        n506) );
  MUX4ND0 U176 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n87), .S1(N76), .ZN(
        n519) );
  MUX4ND0 U177 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n82), .S1(N76), .ZN(
        n532) );
  MUX4ND0 U178 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n75), .S1(n95), .ZN(
        n545) );
  INVD1 U179 ( .I(N77), .ZN(n105) );
  MUX4D0 U180 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(N75), .S1(n93), .Z(
        n559) );
  MUX4D0 U181 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n84), .S1(n90), .Z(n110)
         );
  MUX4D0 U182 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n80), .S1(n97), .Z(n123)
         );
  MUX4D0 U183 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n81), .S1(n93), .Z(n136)
         );
  MUX4D0 U184 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n81), .S1(n94), .Z(n182)
         );
  MUX4D0 U185 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n82), .S1(n92), .Z(n195)
         );
  MUX4D0 U186 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n82), .S1(n91), .Z(n208)
         );
  MUX4D0 U187 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n83), .S1(n95), .Z(n221)
         );
  MUX4D0 U188 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n83), .S1(n92), .Z(n234)
         );
  MUX4D0 U189 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n84), .S1(n97), .Z(n247)
         );
  MUX4D0 U190 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n84), .S1(n93), .Z(n260)
         );
  MUX4D0 U191 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n81), .S1(n93), .Z(
        n273) );
  MUX4D0 U192 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n75), .S1(n94), .Z(
        n286) );
  MUX4D0 U193 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n76), .S1(n94), .Z(
        n299) );
  MUX4D0 U194 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n82), .S1(n95), .Z(
        n312) );
  MUX4D0 U195 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n86), .S1(n95), .Z(
        n325) );
  MUX4D0 U196 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n87), .S1(n96), .Z(
        n338) );
  MUX4D0 U197 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n81), .S1(n97), .Z(
        n351) );
  MUX4D0 U198 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n80), .S1(n97), .Z(
        n364) );
  MUX4D0 U199 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n80), .S1(n96), .Z(
        n377) );
  MUX4D0 U200 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n79), .S1(n92), .Z(
        n390) );
  MUX4D0 U201 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n79), .S1(n95), .Z(
        n403) );
  MUX4D0 U202 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n78), .S1(n95), .Z(
        n416) );
  MUX4D0 U203 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n77), .S1(n94), .Z(
        n429) );
  MUX4D0 U204 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n77), .S1(n93), .Z(
        n442) );
  MUX4D0 U205 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n76), .S1(n96), .Z(
        n455) );
  MUX4D0 U206 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n76), .S1(n90), .Z(
        n468) );
  MUX4D0 U207 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n75), .S1(n90), .Z(
        n481) );
  MUX4D0 U208 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n75), .S1(n91), .Z(
        n494) );
  MUX4D0 U209 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n87), .S1(n91), .Z(
        n507) );
  MUX4D0 U210 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n76), .S1(n92), .Z(
        n520) );
  MUX4D0 U211 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n81), .S1(n92), .Z(
        n533) );
  MUX4D0 U212 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n82), .S1(n91), .Z(
        n546) );
  MUX4D0 U213 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(N75), .S1(N76), .Z(
        n561) );
  MUX4D0 U214 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(N75), .S1(n97), .Z(n563)
         );
  MUX4D0 U215 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n79), .S1(n91), .Z(n112)
         );
  MUX4D0 U216 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n78), .S1(n94), .Z(n114)
         );
  MUX4D0 U217 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n82), .S1(n96), .Z(n125)
         );
  MUX4D0 U218 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n81), .S1(n95), .Z(n127)
         );
  MUX4D0 U219 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n81), .S1(n97), .Z(n138)
         );
  MUX4D0 U220 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n81), .S1(n98), .Z(n140)
         );
  MUX4D0 U221 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n81), .S1(n94), .Z(n184)
         );
  MUX4D0 U222 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n81), .S1(n90), .Z(n186)
         );
  MUX4D0 U223 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n82), .S1(n90), .Z(n197)
         );
  MUX4D0 U224 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n82), .S1(n98), .Z(n199)
         );
  MUX4D0 U225 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n82), .S1(n95), .Z(n210)
         );
  MUX4D0 U226 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n83), .S1(n94), .Z(n212)
         );
  MUX4D0 U227 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n83), .S1(n93), .Z(n223)
         );
  MUX4D0 U228 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n83), .S1(n97), .Z(n225)
         );
  MUX4D0 U229 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n83), .S1(n95), .Z(n236)
         );
  MUX4D0 U230 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n84), .S1(n94), .Z(n238)
         );
  MUX4D0 U231 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n84), .S1(n93), .Z(n249)
         );
  MUX4D0 U232 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n84), .S1(n93), .Z(n251)
         );
  MUX4D0 U233 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n80), .S1(n93), .Z(n262)
         );
  MUX4D0 U234 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n77), .S1(n93), .Z(n264)
         );
  MUX4D0 U235 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n76), .S1(n93), .Z(
        n275) );
  MUX4D0 U236 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n75), .S1(n94), .Z(n277)
         );
  MUX4D0 U237 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n77), .S1(n94), .Z(
        n288) );
  MUX4D0 U238 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n83), .S1(n94), .Z(n290)
         );
  MUX4D0 U239 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n81), .S1(n95), .Z(
        n301) );
  MUX4D0 U240 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n80), .S1(n95), .Z(n303)
         );
  MUX4D0 U241 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n85), .S1(n95), .Z(
        n314) );
  MUX4D0 U242 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n86), .S1(n95), .Z(n316)
         );
  MUX4D0 U243 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n87), .S1(n96), .Z(
        n327) );
  MUX4D0 U244 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n82), .S1(n96), .Z(n329)
         );
  MUX4D0 U245 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n79), .S1(n96), .Z(
        n340) );
  MUX4D0 U246 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n84), .S1(n96), .Z(n342)
         );
  MUX4D0 U247 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n83), .S1(n97), .Z(
        n353) );
  MUX4D0 U248 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n80), .S1(n97), .Z(n355)
         );
  MUX4D0 U249 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n80), .S1(n97), .Z(
        n366) );
  MUX4D0 U250 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n80), .S1(n97), .Z(n368)
         );
  MUX4D0 U251 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n79), .S1(n90), .Z(
        n379) );
  MUX4D0 U252 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n79), .S1(n97), .Z(n381)
         );
  MUX4D0 U253 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n79), .S1(n90), .Z(
        n392) );
  MUX4D0 U254 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n79), .S1(n91), .Z(n394)
         );
  MUX4D0 U255 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n78), .S1(n90), .Z(
        n405) );
  MUX4D0 U256 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n78), .S1(n95), .Z(n407)
         );
  MUX4D0 U257 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n78), .S1(n91), .Z(
        n418) );
  MUX4D0 U258 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n78), .S1(n93), .Z(n420)
         );
  MUX4D0 U259 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n77), .S1(n91), .Z(
        n431) );
  MUX4D0 U260 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n77), .S1(n98), .Z(n433)
         );
  MUX4D0 U261 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n77), .S1(n92), .Z(
        n444) );
  MUX4D0 U262 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n77), .S1(n95), .Z(n446)
         );
  MUX4D0 U263 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n76), .S1(n90), .Z(
        n457) );
  MUX4D0 U264 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n76), .S1(n93), .Z(n459)
         );
  MUX4D0 U265 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n76), .S1(n90), .Z(
        n470) );
  MUX4D0 U266 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n75), .S1(n90), .Z(n472)
         );
  MUX4D0 U267 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n75), .S1(n90), .Z(
        n483) );
  MUX4D0 U268 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n75), .S1(n90), .Z(n485)
         );
  MUX4D0 U269 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n75), .S1(n91), .Z(
        n496) );
  MUX4D0 U270 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n85), .S1(n91), .Z(n498)
         );
  MUX4D0 U271 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n86), .S1(n91), .Z(
        n509) );
  MUX4D0 U272 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n78), .S1(n92), .Z(n511)
         );
  MUX4D0 U273 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n83), .S1(n92), .Z(
        n522) );
  MUX4D0 U274 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n84), .S1(n92), .Z(n524)
         );
  MUX4D0 U275 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n80), .S1(n92), .Z(
        n535) );
  MUX4D0 U276 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n79), .S1(n92), .Z(n537)
         );
  MUX4D0 U277 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(N75), .S1(n93), .Z(
        n548) );
  MUX4D0 U278 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(N75), .S1(n98), .Z(n550)
         );
  MUX4D0 U279 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(N75), .S1(n96), .Z(
        n560) );
  MUX4D0 U280 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n83), .S1(n98), .Z(n111)
         );
  MUX4D0 U281 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n84), .S1(n98), .Z(n124)
         );
  MUX4D0 U282 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n81), .S1(n96), .Z(n137)
         );
  MUX4D0 U283 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n81), .S1(n97), .Z(n183)
         );
  MUX4D0 U284 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n82), .S1(n95), .Z(n196)
         );
  MUX4D0 U285 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n82), .S1(n96), .Z(n209)
         );
  MUX4D0 U286 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n83), .S1(n97), .Z(n222)
         );
  MUX4D0 U287 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n83), .S1(n91), .Z(n235)
         );
  MUX4D0 U288 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n84), .S1(n97), .Z(n248)
         );
  MUX4D0 U289 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n76), .S1(n93), .Z(n261)
         );
  MUX4D0 U290 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n87), .S1(n93), .Z(
        n274) );
  MUX4D0 U291 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n87), .S1(n94), .Z(
        n287) );
  MUX4D0 U292 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n86), .S1(n94), .Z(
        n300) );
  MUX4D0 U293 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n79), .S1(n95), .Z(
        n313) );
  MUX4D0 U294 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n81), .S1(n96), .Z(
        n326) );
  MUX4D0 U295 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n77), .S1(n96), .Z(
        n339) );
  MUX4D0 U296 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n81), .S1(n97), .Z(
        n352) );
  MUX4D0 U297 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n80), .S1(n97), .Z(
        n365) );
  MUX4D0 U298 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n80), .S1(n92), .Z(
        n378) );
  MUX4D0 U299 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n79), .S1(n95), .Z(
        n391) );
  MUX4D0 U300 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n78), .S1(n93), .Z(
        n404) );
  MUX4D0 U301 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n78), .S1(n92), .Z(
        n417) );
  MUX4D0 U302 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n77), .S1(n95), .Z(
        n430) );
  MUX4D0 U303 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n77), .S1(n94), .Z(
        n443) );
  MUX4D0 U304 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n76), .S1(n94), .Z(
        n456) );
  MUX4D0 U305 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n76), .S1(n90), .Z(
        n469) );
  MUX4D0 U306 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n75), .S1(n90), .Z(
        n482) );
  MUX4D0 U307 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n75), .S1(n91), .Z(
        n495) );
  MUX4D0 U308 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n79), .S1(n91), .Z(
        n508) );
  MUX4D0 U309 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n80), .S1(n92), .Z(
        n521) );
  MUX4D0 U310 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n78), .S1(n92), .Z(
        n534) );
  MUX4D0 U311 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(N75), .S1(n94), .Z(
        n547) );
  MUX4D0 U312 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(N75), .S1(n96), .Z(
        n562) );
  MUX4D0 U313 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(N75), .S1(n98), .Z(n564)
         );
  MUX4D0 U314 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n78), .S1(n97), .Z(n113)
         );
  MUX4D0 U315 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n81), .S1(n95), .Z(n115)
         );
  MUX4D0 U316 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n84), .S1(n92), .Z(n126)
         );
  MUX4D0 U317 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n82), .S1(N76), .Z(n128)
         );
  MUX4D0 U318 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n81), .S1(n91), .Z(n139)
         );
  MUX4D0 U319 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n81), .S1(n90), .Z(n141)
         );
  MUX4D0 U320 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n81), .S1(n91), .Z(n185)
         );
  MUX4D0 U321 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n82), .S1(n96), .Z(n187)
         );
  MUX4D0 U322 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n82), .S1(n92), .Z(n198)
         );
  MUX4D0 U323 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n82), .S1(n90), .Z(n200)
         );
  MUX4D0 U324 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n82), .S1(n92), .Z(n211)
         );
  MUX4D0 U325 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n83), .S1(n92), .Z(n213)
         );
  MUX4D0 U326 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n83), .S1(n91), .Z(n224)
         );
  MUX4D0 U327 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n83), .S1(n96), .Z(n226)
         );
  MUX4D0 U328 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n84), .S1(n98), .Z(n237)
         );
  MUX4D0 U329 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n84), .S1(n93), .Z(n239)
         );
  MUX4D0 U330 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n84), .S1(n92), .Z(n250)
         );
  MUX4D0 U331 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n84), .S1(n93), .Z(n252)
         );
  MUX4D0 U332 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n86), .S1(n93), .Z(n263)
         );
  MUX4D0 U333 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n85), .S1(n93), .Z(n265)
         );
  MUX4D0 U334 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n87), .S1(n94), .Z(
        n276) );
  MUX4D0 U335 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n84), .S1(n94), .Z(n278)
         );
  MUX4D0 U336 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n85), .S1(n94), .Z(
        n289) );
  MUX4D0 U337 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n77), .S1(n94), .Z(n291)
         );
  MUX4D0 U338 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n78), .S1(n95), .Z(
        n302) );
  MUX4D0 U339 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n79), .S1(n95), .Z(n304)
         );
  MUX4D0 U340 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n83), .S1(n95), .Z(
        n315) );
  MUX4D0 U341 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n84), .S1(n95), .Z(n317)
         );
  MUX4D0 U342 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n84), .S1(n96), .Z(
        n328) );
  MUX4D0 U343 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n82), .S1(n96), .Z(n330)
         );
  MUX4D0 U344 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n83), .S1(n96), .Z(
        n341) );
  MUX4D0 U345 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n84), .S1(n96), .Z(n343)
         );
  MUX4D0 U346 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n80), .S1(n97), .Z(
        n354) );
  MUX4D0 U347 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n80), .S1(n97), .Z(n356)
         );
  MUX4D0 U348 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n80), .S1(n97), .Z(
        n367) );
  MUX4D0 U349 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n80), .S1(n91), .Z(n369)
         );
  MUX4D0 U350 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n79), .S1(n93), .Z(
        n380) );
  MUX4D0 U351 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n79), .S1(n96), .Z(n382)
         );
  MUX4D0 U352 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n79), .S1(n97), .Z(
        n393) );
  MUX4D0 U353 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n79), .S1(n94), .Z(n395)
         );
  MUX4D0 U354 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n78), .S1(n96), .Z(
        n406) );
  MUX4D0 U355 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n78), .S1(n96), .Z(n408)
         );
  MUX4D0 U356 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n78), .S1(n92), .Z(
        n419) );
  MUX4D0 U357 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n78), .S1(n97), .Z(n421)
         );
  MUX4D0 U358 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n77), .S1(n98), .Z(
        n432) );
  MUX4D0 U359 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n77), .S1(n96), .Z(n434)
         );
  MUX4D0 U360 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n77), .S1(n98), .Z(
        n445) );
  MUX4D0 U361 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n76), .S1(n94), .Z(n447)
         );
  MUX4D0 U362 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n76), .S1(n94), .Z(
        n458) );
  MUX4D0 U363 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n76), .S1(n91), .Z(n460)
         );
  MUX4D0 U364 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n76), .S1(n90), .Z(
        n471) );
  MUX4D0 U365 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n75), .S1(n90), .Z(n473)
         );
  MUX4D0 U366 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n75), .S1(n90), .Z(
        n484) );
  MUX4D0 U367 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n75), .S1(n91), .Z(n486)
         );
  MUX4D0 U368 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n75), .S1(n91), .Z(
        n497) );
  MUX4D0 U369 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n76), .S1(n91), .Z(n499)
         );
  MUX4D0 U370 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n77), .S1(n91), .Z(
        n510) );
  MUX4D0 U371 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n83), .S1(n92), .Z(n512)
         );
  MUX4D0 U372 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n77), .S1(n92), .Z(
        n523) );
  MUX4D0 U373 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n76), .S1(n92), .Z(n525)
         );
  MUX4D0 U374 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n75), .S1(n90), .Z(
        n536) );
  MUX4D0 U375 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n76), .S1(n90), .Z(n538)
         );
  MUX4D0 U376 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(N75), .S1(n90), .Z(
        n549) );
  MUX4D0 U377 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n87), .S1(n98), .Z(n551)
         );
  MUX3ND0 U378 ( .I0(n107), .I1(n108), .I2(n109), .S0(n97), .S1(n100), .ZN(
        n106) );
  MUX3ND0 U379 ( .I0(n116), .I1(n117), .I2(n118), .S0(N78), .S1(N79), .ZN(N113) );
  MUX3ND0 U380 ( .I0(n120), .I1(n121), .I2(n122), .S0(n94), .S1(n102), .ZN(
        n119) );
  MUX3ND0 U381 ( .I0(n129), .I1(n130), .I2(n131), .S0(N78), .S1(N79), .ZN(N112) );
  MUX3ND0 U382 ( .I0(n133), .I1(n134), .I2(n135), .S0(n93), .S1(n104), .ZN(
        n132) );
  MUX3ND0 U383 ( .I0(n175), .I1(n176), .I2(n177), .S0(N78), .S1(N79), .ZN(N111) );
  MUX3ND0 U384 ( .I0(n179), .I1(n180), .I2(n181), .S0(n98), .S1(n101), .ZN(
        n178) );
  MUX3ND0 U385 ( .I0(n188), .I1(n189), .I2(n190), .S0(N78), .S1(N79), .ZN(N110) );
  MUX3ND0 U386 ( .I0(n192), .I1(n193), .I2(n194), .S0(n95), .S1(n101), .ZN(
        n191) );
  MUX3ND0 U387 ( .I0(n201), .I1(n202), .I2(n203), .S0(N78), .S1(N79), .ZN(N109) );
  MUX3ND0 U388 ( .I0(n205), .I1(n206), .I2(n207), .S0(n98), .S1(n101), .ZN(
        n204) );
  MUX3ND0 U389 ( .I0(n214), .I1(n215), .I2(n216), .S0(N78), .S1(N79), .ZN(N108) );
  MUX3ND0 U390 ( .I0(n218), .I1(n219), .I2(n220), .S0(n90), .S1(n100), .ZN(
        n217) );
  MUX3ND0 U391 ( .I0(n227), .I1(n228), .I2(n229), .S0(N78), .S1(N79), .ZN(N107) );
  MUX3ND0 U392 ( .I0(n231), .I1(n232), .I2(n233), .S0(n98), .S1(n100), .ZN(
        n230) );
  MUX3ND0 U393 ( .I0(n240), .I1(n241), .I2(n242), .S0(N78), .S1(N79), .ZN(N106) );
  MUX3ND0 U394 ( .I0(n244), .I1(n245), .I2(n246), .S0(n96), .S1(n104), .ZN(
        n243) );
  MUX3ND0 U395 ( .I0(n253), .I1(n254), .I2(n255), .S0(N78), .S1(N79), .ZN(N105) );
  MUX3ND0 U396 ( .I0(n257), .I1(n258), .I2(n259), .S0(n97), .S1(n103), .ZN(
        n256) );
  MUX3ND0 U397 ( .I0(n266), .I1(n267), .I2(n268), .S0(N78), .S1(N79), .ZN(N104) );
  MUX3ND0 U398 ( .I0(n270), .I1(n271), .I2(n272), .S0(n97), .S1(n102), .ZN(
        n269) );
  MUX3ND0 U399 ( .I0(n279), .I1(n280), .I2(n281), .S0(N78), .S1(N79), .ZN(N103) );
  MUX3ND0 U400 ( .I0(n283), .I1(n284), .I2(n285), .S0(n90), .S1(n104), .ZN(
        n282) );
  MUX3ND0 U401 ( .I0(n292), .I1(n293), .I2(n294), .S0(N78), .S1(N79), .ZN(N102) );
  MUX3ND0 U402 ( .I0(n296), .I1(n297), .I2(n298), .S0(n91), .S1(n103), .ZN(
        n295) );
  MUX3ND0 U403 ( .I0(n305), .I1(n306), .I2(n307), .S0(N78), .S1(N79), .ZN(N101) );
  MUX3ND0 U404 ( .I0(n309), .I1(n310), .I2(n311), .S0(N76), .S1(n104), .ZN(
        n308) );
  MUX3ND0 U405 ( .I0(n318), .I1(n319), .I2(n320), .S0(N78), .S1(N79), .ZN(N100) );
  MUX3ND0 U406 ( .I0(n322), .I1(n323), .I2(n324), .S0(n92), .S1(n100), .ZN(
        n321) );
  MUX3ND0 U407 ( .I0(n331), .I1(n332), .I2(n333), .S0(N78), .S1(N79), .ZN(N99)
         );
  MUX3ND0 U408 ( .I0(n335), .I1(n336), .I2(n337), .S0(n96), .S1(n101), .ZN(
        n334) );
  MUX3ND0 U409 ( .I0(n344), .I1(n345), .I2(n346), .S0(N78), .S1(N79), .ZN(N98)
         );
  MUX3ND0 U410 ( .I0(n348), .I1(n349), .I2(n350), .S0(n97), .S1(n104), .ZN(
        n347) );
  MUX3ND0 U411 ( .I0(n357), .I1(n358), .I2(n359), .S0(N78), .S1(N79), .ZN(N97)
         );
  MUX3ND0 U412 ( .I0(n361), .I1(n362), .I2(n363), .S0(n90), .S1(n102), .ZN(
        n360) );
  MUX3ND0 U413 ( .I0(n370), .I1(n371), .I2(n372), .S0(N78), .S1(N79), .ZN(N96)
         );
  MUX3ND0 U414 ( .I0(n374), .I1(n375), .I2(n376), .S0(n94), .S1(n102), .ZN(
        n373) );
  MUX3ND0 U415 ( .I0(n383), .I1(n384), .I2(n385), .S0(N78), .S1(N79), .ZN(N95)
         );
  MUX3ND0 U416 ( .I0(n387), .I1(n388), .I2(n389), .S0(n95), .S1(n104), .ZN(
        n386) );
  MUX3ND0 U417 ( .I0(n396), .I1(n397), .I2(n398), .S0(N78), .S1(N79), .ZN(N94)
         );
  MUX3ND0 U418 ( .I0(n400), .I1(n401), .I2(n402), .S0(n92), .S1(n102), .ZN(
        n399) );
  MUX3ND0 U419 ( .I0(n409), .I1(n410), .I2(n411), .S0(N78), .S1(N79), .ZN(N93)
         );
  MUX3ND0 U420 ( .I0(n413), .I1(n414), .I2(n415), .S0(n94), .S1(n103), .ZN(
        n412) );
  MUX3ND0 U421 ( .I0(n422), .I1(n423), .I2(n424), .S0(N78), .S1(N79), .ZN(N92)
         );
  MUX3ND0 U422 ( .I0(n426), .I1(n427), .I2(n428), .S0(n92), .S1(n103), .ZN(
        n425) );
  MUX3ND0 U423 ( .I0(n435), .I1(n436), .I2(n437), .S0(N78), .S1(N79), .ZN(N91)
         );
  MUX3ND0 U424 ( .I0(n439), .I1(n440), .I2(n441), .S0(n90), .S1(N77), .ZN(n438) );
  MUX3ND0 U425 ( .I0(n448), .I1(n449), .I2(n450), .S0(N78), .S1(N79), .ZN(N90)
         );
  MUX3ND0 U426 ( .I0(n452), .I1(n453), .I2(n454), .S0(n91), .S1(n101), .ZN(
        n451) );
  MUX3ND0 U427 ( .I0(n461), .I1(n462), .I2(n463), .S0(N78), .S1(N79), .ZN(N89)
         );
  MUX3ND0 U428 ( .I0(n465), .I1(n466), .I2(n467), .S0(n98), .S1(N77), .ZN(n464) );
  MUX3ND0 U429 ( .I0(n474), .I1(n475), .I2(n476), .S0(N78), .S1(N79), .ZN(N88)
         );
  MUX3ND0 U430 ( .I0(n478), .I1(n479), .I2(n480), .S0(n93), .S1(N77), .ZN(n477) );
  MUX3ND0 U431 ( .I0(n487), .I1(n488), .I2(n489), .S0(N78), .S1(N79), .ZN(N87)
         );
  MUX3ND0 U432 ( .I0(n491), .I1(n492), .I2(n493), .S0(n91), .S1(N77), .ZN(n490) );
  MUX3ND0 U433 ( .I0(n500), .I1(n501), .I2(n502), .S0(N78), .S1(N79), .ZN(N86)
         );
  MUX3ND0 U434 ( .I0(n504), .I1(n505), .I2(n506), .S0(n94), .S1(N77), .ZN(n503) );
  MUX3ND0 U435 ( .I0(n513), .I1(n514), .I2(n515), .S0(N78), .S1(N79), .ZN(N85)
         );
  MUX3ND0 U436 ( .I0(n517), .I1(n518), .I2(n519), .S0(n96), .S1(N77), .ZN(n516) );
  MUX3ND0 U437 ( .I0(n526), .I1(n527), .I2(n528), .S0(N78), .S1(N79), .ZN(N84)
         );
  MUX3ND0 U438 ( .I0(n530), .I1(n531), .I2(n532), .S0(n93), .S1(N77), .ZN(n529) );
  MUX3ND0 U439 ( .I0(n539), .I1(n540), .I2(n541), .S0(N78), .S1(N79), .ZN(N83)
         );
  MUX3ND0 U440 ( .I0(n543), .I1(n544), .I2(n545), .S0(n93), .S1(n102), .ZN(
        n542) );
  MUX3ND0 U441 ( .I0(n552), .I1(n553), .I2(n554), .S0(N78), .S1(N79), .ZN(N82)
         );
  MUX3ND0 U442 ( .I0(n556), .I1(n557), .I2(n558), .S0(n91), .S1(N77), .ZN(n555) );
  MUX3ND0 U443 ( .I0(n565), .I1(n566), .I2(n567), .S0(N78), .S1(N79), .ZN(N81)
         );
  MUX2ND0 U444 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n85), .ZN(
        n108) );
  MUX2ND0 U445 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n87), .ZN(
        n107) );
  MUX3ND0 U446 ( .I0(n111), .I1(n110), .I2(n106), .S0(n101), .S1(N78), .ZN(
        n118) );
  MUX2ND0 U447 ( .I0(n113), .I1(n112), .S(n104), .ZN(n117) );
  MUX2ND0 U448 ( .I0(n115), .I1(n114), .S(n104), .ZN(n116) );
  MUX2ND0 U449 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n87), .ZN(
        n121) );
  MUX2ND0 U450 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n87), .ZN(
        n120) );
  MUX3ND0 U451 ( .I0(n124), .I1(n123), .I2(n119), .S0(n102), .S1(N78), .ZN(
        n131) );
  MUX2ND0 U452 ( .I0(n126), .I1(n125), .S(n104), .ZN(n130) );
  MUX2ND0 U453 ( .I0(n128), .I1(n127), .S(n104), .ZN(n129) );
  MUX2ND0 U454 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n87), .ZN(
        n134) );
  MUX2ND0 U455 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n87), .ZN(
        n133) );
  MUX3ND0 U456 ( .I0(n137), .I1(n136), .I2(n132), .S0(n101), .S1(N78), .ZN(
        n177) );
  MUX2ND0 U457 ( .I0(n139), .I1(n138), .S(n104), .ZN(n176) );
  MUX2ND0 U458 ( .I0(n141), .I1(n140), .S(n104), .ZN(n175) );
  MUX2ND0 U459 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n87), .ZN(
        n180) );
  MUX2ND0 U460 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n87), .ZN(
        n179) );
  MUX3ND0 U461 ( .I0(n183), .I1(n182), .I2(n178), .S0(n100), .S1(N78), .ZN(
        n190) );
  MUX2ND0 U462 ( .I0(n185), .I1(n184), .S(n104), .ZN(n189) );
  MUX2ND0 U463 ( .I0(n187), .I1(n186), .S(n104), .ZN(n188) );
  MUX2ND0 U464 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n87), .ZN(
        n193) );
  MUX2ND0 U465 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n87), .ZN(
        n192) );
  MUX3ND0 U466 ( .I0(n196), .I1(n195), .I2(n191), .S0(n101), .S1(N78), .ZN(
        n203) );
  MUX2ND0 U467 ( .I0(n198), .I1(n197), .S(n104), .ZN(n202) );
  MUX2ND0 U468 ( .I0(n200), .I1(n199), .S(n104), .ZN(n201) );
  MUX2ND0 U469 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n86), .ZN(
        n206) );
  MUX2ND0 U470 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n87), .ZN(
        n205) );
  MUX3ND0 U471 ( .I0(n209), .I1(n208), .I2(n204), .S0(n103), .S1(N78), .ZN(
        n216) );
  MUX2ND0 U472 ( .I0(n211), .I1(n210), .S(n103), .ZN(n215) );
  MUX2ND0 U473 ( .I0(n213), .I1(n212), .S(n104), .ZN(n214) );
  MUX2ND0 U474 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n86), .ZN(
        n219) );
  MUX2ND0 U475 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n86), .ZN(
        n218) );
  MUX3ND0 U476 ( .I0(n222), .I1(n221), .I2(n217), .S0(n101), .S1(N78), .ZN(
        n229) );
  MUX2ND0 U477 ( .I0(n224), .I1(n223), .S(n103), .ZN(n228) );
  MUX2ND0 U478 ( .I0(n226), .I1(n225), .S(n103), .ZN(n227) );
  MUX2ND0 U479 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n86), .ZN(
        n232) );
  MUX2ND0 U480 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n86), .ZN(
        n231) );
  MUX3ND0 U481 ( .I0(n235), .I1(n234), .I2(n230), .S0(n104), .S1(N78), .ZN(
        n242) );
  MUX2ND0 U482 ( .I0(n237), .I1(n236), .S(n103), .ZN(n241) );
  MUX2ND0 U483 ( .I0(n239), .I1(n238), .S(n103), .ZN(n240) );
  MUX2ND0 U484 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n86), .ZN(
        n245) );
  MUX2ND0 U485 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n86), .ZN(
        n244) );
  MUX3ND0 U486 ( .I0(n248), .I1(n247), .I2(n243), .S0(n101), .S1(N78), .ZN(
        n255) );
  MUX2ND0 U487 ( .I0(n250), .I1(n249), .S(n103), .ZN(n254) );
  MUX2ND0 U488 ( .I0(n252), .I1(n251), .S(n103), .ZN(n253) );
  MUX2ND0 U489 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n86), .ZN(
        n258) );
  MUX2ND0 U490 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n86), .ZN(
        n257) );
  MUX3ND0 U491 ( .I0(n261), .I1(n260), .I2(n256), .S0(n100), .S1(N78), .ZN(
        n268) );
  MUX2ND0 U492 ( .I0(n263), .I1(n262), .S(n103), .ZN(n267) );
  MUX2ND0 U493 ( .I0(n265), .I1(n264), .S(n103), .ZN(n266) );
  MUX2ND0 U494 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n86), .ZN(
        n271) );
  MUX2ND0 U495 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n86), .ZN(
        n270) );
  MUX3ND0 U496 ( .I0(n274), .I1(n273), .I2(n269), .S0(n101), .S1(N78), .ZN(
        n281) );
  MUX2ND0 U497 ( .I0(n276), .I1(n275), .S(n103), .ZN(n280) );
  MUX2ND0 U498 ( .I0(n278), .I1(n277), .S(n103), .ZN(n279) );
  MUX2ND0 U499 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n86), .ZN(
        n284) );
  MUX2ND0 U500 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n86), .ZN(
        n283) );
  MUX3ND0 U501 ( .I0(n287), .I1(n286), .I2(n282), .S0(n100), .S1(N78), .ZN(
        n294) );
  MUX2ND0 U502 ( .I0(n289), .I1(n288), .S(n102), .ZN(n293) );
  MUX2ND0 U503 ( .I0(n291), .I1(n290), .S(n102), .ZN(n292) );
  MUX2ND0 U504 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n86), .ZN(
        n297) );
  MUX2ND0 U505 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n86), .ZN(
        n296) );
  MUX3ND0 U506 ( .I0(n300), .I1(n299), .I2(n295), .S0(n101), .S1(N78), .ZN(
        n307) );
  MUX2ND0 U507 ( .I0(n302), .I1(n301), .S(n104), .ZN(n306) );
  MUX2ND0 U508 ( .I0(n304), .I1(n303), .S(n104), .ZN(n305) );
  MUX2ND0 U509 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n86), .ZN(
        n310) );
  MUX2ND0 U510 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n86), .ZN(
        n309) );
  MUX3ND0 U511 ( .I0(n313), .I1(n312), .I2(n308), .S0(n100), .S1(N78), .ZN(
        n320) );
  MUX2ND0 U512 ( .I0(n315), .I1(n314), .S(n102), .ZN(n319) );
  MUX2ND0 U513 ( .I0(n317), .I1(n316), .S(n104), .ZN(n318) );
  MUX2ND0 U514 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n85), .ZN(
        n323) );
  MUX2ND0 U515 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n85), .ZN(
        n322) );
  MUX3ND0 U516 ( .I0(n326), .I1(n325), .I2(n321), .S0(n100), .S1(N78), .ZN(
        n333) );
  MUX2ND0 U517 ( .I0(n328), .I1(n327), .S(n100), .ZN(n332) );
  MUX2ND0 U518 ( .I0(n330), .I1(n329), .S(n100), .ZN(n331) );
  MUX2ND0 U519 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n85), .ZN(
        n336) );
  MUX2ND0 U520 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n85), .ZN(
        n335) );
  MUX3ND0 U521 ( .I0(n339), .I1(n338), .I2(n334), .S0(n100), .S1(N78), .ZN(
        n346) );
  MUX2ND0 U522 ( .I0(n341), .I1(n340), .S(n101), .ZN(n345) );
  MUX2ND0 U523 ( .I0(n343), .I1(n342), .S(n101), .ZN(n344) );
  MUX2ND0 U524 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n85), .ZN(
        n349) );
  MUX2ND0 U525 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n85), .ZN(
        n348) );
  MUX3ND0 U526 ( .I0(n352), .I1(n351), .I2(n347), .S0(n101), .S1(N78), .ZN(
        n359) );
  MUX2ND0 U527 ( .I0(n354), .I1(n353), .S(n102), .ZN(n358) );
  MUX2ND0 U528 ( .I0(n356), .I1(n355), .S(n104), .ZN(n357) );
  MUX2ND0 U529 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n85), .ZN(
        n362) );
  MUX2ND0 U530 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n85), .ZN(
        n361) );
  MUX3ND0 U531 ( .I0(n365), .I1(n364), .I2(n360), .S0(n101), .S1(N78), .ZN(
        n372) );
  MUX2ND0 U532 ( .I0(n367), .I1(n366), .S(n103), .ZN(n371) );
  MUX2ND0 U533 ( .I0(n369), .I1(n368), .S(n100), .ZN(n370) );
  MUX2ND0 U534 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n85), .ZN(
        n375) );
  MUX2ND0 U535 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n85), .ZN(
        n374) );
  MUX3ND0 U536 ( .I0(n378), .I1(n377), .I2(n373), .S0(n100), .S1(N78), .ZN(
        n385) );
  MUX2ND0 U537 ( .I0(n380), .I1(n379), .S(n103), .ZN(n384) );
  MUX2ND0 U538 ( .I0(n382), .I1(n381), .S(n100), .ZN(n383) );
  MUX2ND0 U539 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n85), .ZN(
        n388) );
  MUX2ND0 U540 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n85), .ZN(
        n387) );
  MUX3ND0 U541 ( .I0(n391), .I1(n390), .I2(n386), .S0(n100), .S1(N78), .ZN(
        n398) );
  MUX2ND0 U542 ( .I0(n393), .I1(n392), .S(n100), .ZN(n397) );
  MUX2ND0 U543 ( .I0(n395), .I1(n394), .S(n100), .ZN(n396) );
  MUX2ND0 U544 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n85), .ZN(
        n401) );
  MUX2ND0 U545 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n85), .ZN(
        n400) );
  MUX3ND0 U546 ( .I0(n404), .I1(n403), .I2(n399), .S0(n101), .S1(N78), .ZN(
        n411) );
  MUX2ND0 U547 ( .I0(n406), .I1(n405), .S(n103), .ZN(n410) );
  MUX2ND0 U548 ( .I0(n408), .I1(n407), .S(n102), .ZN(n409) );
  MUX2ND0 U549 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n82), .ZN(
        n414) );
  MUX2ND0 U550 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n86), .ZN(
        n413) );
  MUX3ND0 U551 ( .I0(n417), .I1(n416), .I2(n412), .S0(n101), .S1(N78), .ZN(
        n424) );
  MUX2ND0 U552 ( .I0(n419), .I1(n418), .S(n104), .ZN(n423) );
  MUX2ND0 U553 ( .I0(n421), .I1(n420), .S(n101), .ZN(n422) );
  MUX2ND0 U554 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n81), .ZN(
        n427) );
  MUX2ND0 U555 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n80), .ZN(
        n426) );
  MUX3ND0 U556 ( .I0(n430), .I1(n429), .I2(n425), .S0(n100), .S1(N78), .ZN(
        n437) );
  MUX2ND0 U557 ( .I0(n432), .I1(n431), .S(n102), .ZN(n436) );
  MUX2ND0 U558 ( .I0(n434), .I1(n433), .S(n103), .ZN(n435) );
  MUX2ND0 U559 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n78), .ZN(
        n440) );
  MUX2ND0 U560 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n85), .ZN(
        n439) );
  MUX3ND0 U561 ( .I0(n443), .I1(n442), .I2(n438), .S0(n100), .S1(N78), .ZN(
        n450) );
  MUX2ND0 U562 ( .I0(n445), .I1(n444), .S(n102), .ZN(n449) );
  MUX2ND0 U563 ( .I0(n447), .I1(n446), .S(n102), .ZN(n448) );
  MUX2ND0 U564 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n75), .ZN(
        n453) );
  MUX2ND0 U565 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n87), .ZN(
        n452) );
  MUX3ND0 U566 ( .I0(n456), .I1(n455), .I2(n451), .S0(n100), .S1(N78), .ZN(
        n463) );
  MUX2ND0 U567 ( .I0(n458), .I1(n457), .S(n102), .ZN(n462) );
  MUX2ND0 U568 ( .I0(n460), .I1(n459), .S(n104), .ZN(n461) );
  MUX2ND0 U569 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n79), .ZN(
        n466) );
  MUX2ND0 U570 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n77), .ZN(
        n465) );
  MUX3ND0 U571 ( .I0(n469), .I1(n468), .I2(n464), .S0(n100), .S1(N78), .ZN(
        n476) );
  MUX2ND0 U572 ( .I0(n471), .I1(n470), .S(n101), .ZN(n475) );
  MUX2ND0 U573 ( .I0(n473), .I1(n472), .S(n102), .ZN(n474) );
  MUX2ND0 U574 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n83), .ZN(
        n479) );
  MUX2ND0 U575 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n76), .ZN(
        n478) );
  MUX3ND0 U576 ( .I0(n482), .I1(n481), .I2(n477), .S0(n101), .S1(N78), .ZN(
        n489) );
  MUX2ND0 U577 ( .I0(n484), .I1(n483), .S(n102), .ZN(n488) );
  MUX2ND0 U578 ( .I0(n486), .I1(n485), .S(n101), .ZN(n487) );
  MUX2ND0 U579 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n82), .ZN(
        n492) );
  MUX2ND0 U580 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n75), .ZN(
        n491) );
  MUX3ND0 U581 ( .I0(n495), .I1(n494), .I2(n490), .S0(n100), .S1(N78), .ZN(
        n502) );
  MUX2ND0 U582 ( .I0(n497), .I1(n496), .S(n103), .ZN(n501) );
  MUX2ND0 U583 ( .I0(n499), .I1(n498), .S(n102), .ZN(n500) );
  MUX2ND0 U584 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n83), .ZN(
        n505) );
  MUX2ND0 U585 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n75), .ZN(
        n504) );
  MUX3ND0 U586 ( .I0(n508), .I1(n507), .I2(n503), .S0(n103), .S1(N78), .ZN(
        n515) );
  MUX2ND0 U587 ( .I0(n510), .I1(n509), .S(n102), .ZN(n514) );
  MUX2ND0 U588 ( .I0(n512), .I1(n511), .S(n100), .ZN(n513) );
  MUX2ND0 U589 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n77), .ZN(
        n518) );
  MUX2ND0 U590 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n78), .ZN(
        n517) );
  MUX3ND0 U591 ( .I0(n521), .I1(n520), .I2(n516), .S0(n103), .S1(N78), .ZN(
        n528) );
  MUX2ND0 U592 ( .I0(n523), .I1(n522), .S(n103), .ZN(n527) );
  MUX2ND0 U593 ( .I0(n525), .I1(n524), .S(n102), .ZN(n526) );
  MUX2ND0 U594 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n82), .ZN(
        n531) );
  MUX2ND0 U595 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n83), .ZN(
        n530) );
  MUX3ND0 U596 ( .I0(n534), .I1(n533), .I2(n529), .S0(n103), .S1(N78), .ZN(
        n541) );
  MUX2ND0 U597 ( .I0(n536), .I1(n535), .S(n102), .ZN(n540) );
  MUX2ND0 U598 ( .I0(n538), .I1(n537), .S(n104), .ZN(n539) );
  MUX2ND0 U599 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n79), .ZN(
        n544) );
  MUX2ND0 U600 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n84), .ZN(
        n543) );
  MUX3ND0 U601 ( .I0(n547), .I1(n546), .I2(n542), .S0(n101), .S1(N78), .ZN(
        n554) );
  MUX2ND0 U602 ( .I0(n549), .I1(n548), .S(n102), .ZN(n553) );
  MUX2ND0 U603 ( .I0(n551), .I1(n550), .S(n102), .ZN(n552) );
  MUX2ND0 U604 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n85), .ZN(
        n557) );
  MUX2ND0 U605 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n85), .ZN(
        n556) );
  MUX3ND0 U606 ( .I0(n560), .I1(n559), .I2(n555), .S0(n101), .S1(N78), .ZN(
        n567) );
  MUX2ND0 U607 ( .I0(n562), .I1(n561), .S(n102), .ZN(n566) );
  MUX2ND0 U608 ( .I0(n564), .I1(n563), .S(N77), .ZN(n565) );
  CKND0 U609 ( .CLK(Reset), .CN(n174) );
  CKND0 U610 ( .CLK(N63), .CN(n173) );
  CKND0 U611 ( .CLK(N62), .CN(n172) );
  CKND0 U612 ( .CLK(N61), .CN(n171) );
  CKND0 U613 ( .CLK(N60), .CN(n170) );
  CKND0 U614 ( .CLK(N59), .CN(n169) );
  CKND0 U615 ( .CLK(N58), .CN(n168) );
  CKND0 U616 ( .CLK(N57), .CN(n167) );
  CKND0 U617 ( .CLK(N56), .CN(n166) );
  CKND0 U618 ( .CLK(N55), .CN(n165) );
  CKND0 U619 ( .CLK(N54), .CN(n164) );
  CKND0 U620 ( .CLK(N53), .CN(n163) );
  CKND0 U621 ( .CLK(N52), .CN(n162) );
  CKND0 U622 ( .CLK(N51), .CN(n161) );
  CKND0 U623 ( .CLK(N50), .CN(n160) );
  CKND0 U624 ( .CLK(N49), .CN(n159) );
  CKND0 U625 ( .CLK(N48), .CN(n158) );
  CKND0 U626 ( .CLK(N47), .CN(n157) );
  CKND0 U627 ( .CLK(N46), .CN(n156) );
  CKND0 U628 ( .CLK(N45), .CN(n155) );
  CKND0 U629 ( .CLK(N44), .CN(n154) );
  CKND0 U630 ( .CLK(N43), .CN(n153) );
  CKND0 U631 ( .CLK(N42), .CN(n152) );
  CKND0 U632 ( .CLK(N41), .CN(n151) );
  CKND0 U633 ( .CLK(N40), .CN(n150) );
  CKND0 U634 ( .CLK(N39), .CN(n149) );
  CKND0 U635 ( .CLK(N38), .CN(n148) );
  CKND0 U636 ( .CLK(N37), .CN(n147) );
  CKND0 U637 ( .CLK(N36), .CN(n146) );
  CKND0 U638 ( .CLK(N35), .CN(n145) );
  CKND0 U639 ( .CLK(N34), .CN(n144) );
  CKND0 U640 ( .CLK(N33), .CN(n143) );
  CKND0 U641 ( .CLK(N32), .CN(n142) );
  CKND2D0 U642 ( .A1(Read), .A2(ChipEna), .ZN(n570) );
  ND3D0 U643 ( .A1(N76), .A2(n87), .A3(N77), .ZN(n572) );
  ND3D0 U644 ( .A1(N76), .A2(n88), .A3(N77), .ZN(n573) );
  ND3D0 U645 ( .A1(n87), .A2(n99), .A3(N77), .ZN(n574) );
  ND3D0 U646 ( .A1(n89), .A2(n99), .A3(N77), .ZN(n575) );
  ND3D0 U647 ( .A1(n87), .A2(n105), .A3(N76), .ZN(n576) );
  ND3D0 U648 ( .A1(n88), .A2(n105), .A3(N76), .ZN(n577) );
  ND3D0 U649 ( .A1(n99), .A2(n105), .A3(n87), .ZN(n578) );
  CKND0 U650 ( .CLK(Write), .CN(n569) );
  CKND0 U651 ( .CLK(N79), .CN(n583) );
  CKND0 U652 ( .CLK(N78), .CN(n581) );
  ND3D0 U653 ( .A1(n99), .A2(n105), .A3(n88), .ZN(n579) );
  XOR3D0 U654 ( .A1(DataI[0]), .A2(n586), .A3(n587), .Z(n585) );
  XOR3D0 U655 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n588), .Z(n587) );
  XOR3D0 U656 ( .A1(n589), .A2(DataI[3]), .A3(n590), .Z(n588) );
  XOR3D0 U657 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n591), .Z(n590) );
  XOR3D0 U658 ( .A1(n592), .A2(DataI[10]), .A3(n593), .Z(n591) );
  XOR3D0 U659 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n594), .Z(n593) );
  XOR3D0 U660 ( .A1(n595), .A2(DataI[17]), .A3(n596), .Z(n594) );
  XNR4D0 U661 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n596) );
  XOR4D0 U662 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n595) );
  XOR4D0 U663 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n592) );
  XOR4D0 U664 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n589) );
  XNR4D0 U665 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n586) );
  XOR4D0 U666 ( .A1(n597), .A2(N110), .A3(n598), .A4(n599), .Z(N116) );
  XNR4D0 U667 ( .A1(N107), .A2(N106), .A3(N109), .A4(N108), .ZN(n599) );
  XNR3D0 U668 ( .A1(N113), .A2(N112), .A3(N111), .ZN(n598) );
  XOR3D0 U669 ( .A1(N105), .A2(N104), .A3(n600), .Z(n597) );
  XOR3D0 U670 ( .A1(N103), .A2(n601), .A3(n602), .Z(n600) );
  XOR3D0 U671 ( .A1(N102), .A2(N101), .A3(n603), .Z(n602) );
  XOR3D0 U672 ( .A1(n604), .A2(N100), .A3(n605), .Z(n603) );
  XOR3D0 U673 ( .A1(N91), .A2(N90), .A3(n606), .Z(n605) );
  XOR3D0 U674 ( .A1(n607), .A2(N89), .A3(n608), .Z(n606) );
  XNR4D0 U675 ( .A1(N82), .A2(N81), .A3(N84), .A4(N83), .ZN(n608) );
  XOR4D0 U676 ( .A1(N86), .A2(N85), .A3(N88), .A4(N87), .Z(n607) );
  XOR4D0 U677 ( .A1(N93), .A2(N92), .A3(N95), .A4(N94), .Z(n604) );
  XNR4D0 U678 ( .A1(N97), .A2(N96), .A3(N99), .A4(N98), .ZN(n601) );
  INR2D0 U679 ( .A1(DreadyReg), .B1(n568), .ZN(Dready) );
  INR2D0 U680 ( .A1(ClockIn), .B1(n568), .ZN(ChipClock) );
  CKND0 U681 ( .CLK(ChipEna), .CN(n568) );
endmodule


module PLLTop ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(Reset) );
  VFO VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(Reset) );
  MultiCounter MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(Reset)
         );
endmodule


module ClockComparator ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   ZeroCounters, N5, N6, \CounterClockN[1] , N7, N8, N9, N19, N20, n2,
         n3, n7, n6, n8, n9, n10;

  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n2), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n2), .QN(n7) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n2), .QN(N7)
         );
  DFSNQD1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n3), .Q(ZeroCounters)
         );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n3), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n3), .Q(
        AdjustFreq[1]) );
  DFCNQD1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n2), .Q(
        \CounterClockN[1] ) );
  CKND0 U3 ( .CLK(Reset), .CN(n3) );
  CKND0 U4 ( .CLK(ZeroCounters), .CN(n2) );
  OAI22D0 U5 ( .A1(n7), .A2(n6), .B1(n8), .B2(N8), .ZN(N20) );
  XNR2D0 U6 ( .A1(N7), .A2(\CounterClockN[1] ), .ZN(N8) );
  IAO21D0 U7 ( .A1(n6), .A2(N5), .B(N9), .ZN(n8) );
  OAI22D0 U8 ( .A1(n6), .A2(n9), .B1(\CounterClockN[1] ), .B2(n10), .ZN(N19)
         );
  NR2D0 U9 ( .A1(N7), .A2(N6), .ZN(n10) );
  CKXOR2D0 U10 ( .A1(n7), .A2(N5), .Z(N6) );
  CKND0 U11 ( .CLK(N9), .CN(n9) );
  NR2D0 U12 ( .A1(N5), .A2(n7), .ZN(N9) );
  INR2D0 U13 ( .A1(\CounterClockN[1] ), .B1(N7), .ZN(n6) );
endmodule


module VFO ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N45, N47, N49, N51, N53, N54, N55, \U3/U3/Z_0 , n23, n24, n25, n26,
         n27, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay83ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay83ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay83ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay83ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay83ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_DW01_incdec_0 r86 ( .A(DivideFactor), .INC_DEC(\U3/U3/Z_0 ), .SUM({N55, 
        N53, N51, N49, N47, N45}) );
  VFO_DW01_inc_0 \ClockOutGen/add_161  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFSNQD1 \DivideFactor_reg[0]  ( .D(n27), .CP(Sample), .SDN(n26), .Q(
        DivideFactor[0]) );
  DFSNQD1 \DivideFactor_reg[4]  ( .D(n24), .CP(Sample), .SDN(n26), .Q(
        DivideFactor[4]) );
  DFSNQD1 \DivideFactor_reg[1]  ( .D(n25), .CP(Sample), .SDN(n26), .Q(
        DivideFactor[1]) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[3]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[0]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n26), 
        .Q(DivideFactor[2]) );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n26), 
        .Q(DivideFactor[5]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[4]) );
  EDFCNQD1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n26), 
        .Q(DivideFactor[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n23), .CP(FastClock), .CDN(n26), .Q(ClockOut)
         );
  OAI31D1 U3 ( .A1(n3), .A2(AdjustFreq[1]), .A3(AdjustFreq[0]), .B(n2), .ZN(
        N54) );
  MUX2D0 U4 ( .I0(DivideFactor[0]), .I1(N45), .S(N54), .Z(n27) );
  CKND0 U5 ( .CLK(Reset), .CN(n26) );
  MUX2D0 U6 ( .I0(DivideFactor[1]), .I1(N47), .S(N54), .Z(n25) );
  MUX2D0 U7 ( .I0(DivideFactor[4]), .I1(N53), .S(N54), .Z(n24) );
  XNR2D0 U8 ( .A1(ClockOut), .A2(n1), .ZN(n23) );
  CKND0 U9 ( .CLK(n2), .CN(\U3/U3/Z_0 ) );
  ND3D0 U10 ( .A1(AdjustFreq[0]), .A2(n3), .A3(AdjustFreq[1]), .ZN(n2) );
  OAI22D0 U11 ( .A1(n4), .A2(n5), .B1(n6), .B2(n7), .ZN(n3) );
  INR3D0 U12 ( .A1(n4), .B1(DivideFactor[5]), .B2(DivideFactor[4]), .ZN(n6) );
  ND4D0 U13 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(n8), .ZN(n4) );
  CKND2D0 U14 ( .A1(n7), .A2(n9), .ZN(n8) );
  CKND0 U15 ( .CLK(AdjustFreq[0]), .CN(n7) );
  AN2D0 U16 ( .A1(N14), .A2(n1), .Z(N21) );
  AN2D0 U17 ( .A1(N13), .A2(n1), .Z(N20) );
  AN2D0 U18 ( .A1(N12), .A2(n1), .Z(N19) );
  AN2D0 U19 ( .A1(N11), .A2(n1), .Z(N18) );
  AN2D0 U20 ( .A1(N10), .A2(n1), .Z(N17) );
  AN2D0 U21 ( .A1(N9), .A2(n1), .Z(N16) );
  OAI21D0 U22 ( .A1(FastDivvy[5]), .A2(n5), .B(n10), .ZN(n1) );
  AO221D0 U23 ( .A1(n9), .A2(FastDivvy[4]), .B1(n5), .B2(FastDivvy[5]), .C(n11), .Z(n10) );
  OA21D0 U24 ( .A1(FastDivvy[4]), .A2(n9), .B(n12), .Z(n11) );
  OAI22D0 U25 ( .A1(DivideFactor[3]), .A2(n13), .B1(n14), .B2(n15), .ZN(n12)
         );
  IOA22D0 U26 ( .B1(n16), .B2(n17), .A1(n13), .A2(DivideFactor[3]), .ZN(n15)
         );
  AOI21D0 U27 ( .A1(n16), .A2(n17), .B(FastDivvy[2]), .ZN(n14) );
  CKND0 U28 ( .CLK(DivideFactor[2]), .CN(n17) );
  OA32D0 U29 ( .A1(n18), .A2(FastDivvy[0]), .A3(n19), .B1(FastDivvy[1]), .B2(
        n20), .Z(n16) );
  CKND0 U30 ( .CLK(DivideFactor[1]), .CN(n20) );
  INR2D0 U31 ( .A1(FastDivvy[1]), .B1(DivideFactor[1]), .ZN(n19) );
  CKND0 U32 ( .CLK(DivideFactor[0]), .CN(n18) );
  CKND0 U33 ( .CLK(FastDivvy[3]), .CN(n13) );
  CKND0 U34 ( .CLK(DivideFactor[4]), .CN(n9) );
  CKND0 U35 ( .CLK(DivideFactor[5]), .CN(n5) );
  CKND0 U36 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U37 ( .A1(WireD[5]), .A2(n26), .ZN(WireD[0]) );
endmodule


module MultiCounter ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  CKND0 U3 ( .CLK(Reset), .CN(n1) );
endmodule


module MultiCounter_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_incdec_0 ( A, INC_DEC, SUM );
  input [5:0] A;
  output [5:0] SUM;
  input INC_DEC;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[1] ,
         \carry[0] ;

  XOR3D1 U1_5 ( .A1(A[5]), .A2(INC_DEC), .A3(\carry[5] ), .Z(SUM[5]) );
  FA1D0 U1_3 ( .A(A[3]), .B(INC_DEC), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  FA1D0 U1_2 ( .A(A[2]), .B(INC_DEC), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  FA1D0 U1_4 ( .A(A[4]), .B(INC_DEC), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  FA1D0 U1_1 ( .A(A[1]), .B(INC_DEC), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  FA1D0 U1_0 ( .A(A[0]), .B(INC_DEC), .CI(\carry[0] ), .CO(\carry[1] ), .S(
        SUM[0]) );
  CKND0 U1 ( .CLK(INC_DEC), .CN(\carry[0] ) );
endmodule


module VFO_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

