/************************************************************************\
|*                                                                      *|
|*    Copyright (c) 2005  Springer. All rights reserved.                *|
|*                                                                      *|
|*  This example code shouyld be used only for illustration purpose     *| 
|*  This material is not to reproduced,  copied,  or used  in any       *|
|*  manner without the authorization of the author's/publishers         *|
|*  written permission                                                  *|
|*                                                                      *|
\************************************************************************/

// Author: Srikanth Vijayaraghavan and Meyyappan Ramanathan


module datapath(

input logic clk,

input logic signed [15:0] d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28, d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61,d62,d63, d64,

input logic dp_enable1, dp_enable2, dp_enable3, dp_enable4, reset,

output logic signed [15:0] do1,do2,do3,do4,do5,do6,do7,do8,do9,do10,do11,do12,do13,do14,do15,do16,do17,do18,do19,do20,do21,do22,do23,do24,do25,do26,do27,do28,do29,do30,do31,do32,do33,do34,do35,do36,do37,do38,do39,do40,do41,do42,do43,do44,do45,do46,do47,do48,do49,do50,do51,do52,do53,do54,do55,do56,do57,do58,do59,do60,do61,do62,do63,do64

);

logic signed [15:0] dw1,dw2,dw3,dw4,dw5,dw6,dw7,dw8,dw9,dw10,dw11,dw12,dw13,dw14,dw15,dw16,dw17,dw18,dw19,dw20,dw21,dw22,dw23,dw24,dw25,dw26,dw27,dw28,dw29,dw30,dw31,dw32,dw33,dw34,dw35,dw36,dw37,dw38,dw39,dw40,dw41,dw42,dw43,dw44,dw45,dw46,dw47,dw48,dw49,dw50,dw51,dw52,dw53,dw54,dw55,dw56,dw57,dw58,dw59,dw60,dw61,dw62,dw63,dw64;

logic signed [15:0] dwl1,dwl2,dwl3,dwl4,dwl5,dwl6,dwl7,dwl8,dwl9,dwl10,dwl11,dwl12,dwl13,dwl14,dwl15,dwl16,dwl17,dwl18,dwl19,dwl20,dwl21,dwl22,dwl23,dwl24,dwl25,dwl26,dwl27,dwl28,dwl29,dwl30,dwl31,dwl32,dwl33,dwl34,dwl35,dwl36,dwl37,dwl38,dwl39,dwl40,dwl41,dwl42,dwl43,dwl44,dwl45,dwl46,dwl47,dwl48,dwl49,dwl50,dwl51,dwl52,dwl53,dwl54,dwl55,dwl56,dwl57,dwl58,dwl59,dwl60,dwl61,dwl62,dwl63,dwl64;

logic signed [15:0] dwlt1, dwlt2, dwlt3, dwlt4, dwlt5, dwlt6, dwlt7, dwlt8, dwlt9, dwlt10, dwlt11, dwlt12, dwlt13, dwlt14, dwlt15, dwlt16, dwlt17, dwlt18, dwlt19, dwlt20, dwlt21, dwlt22, dwlt23, dwlt24, dwlt25, dwlt26, dwlt27, dwlt28, dwlt29, dwlt30, dwlt31, dwlt32, dwlt33, dwlt34, dwlt35, dwlt36, dwlt37, dwlt38, dwlt39, dwlt40, dwlt41, dwlt42, dwlt43, dwlt44, dwlt45, dwlt46, dwlt47, dwlt48, dwlt49, dwlt50, dwlt51, dwlt52, dwlt53, dwlt54, dwlt55, dwlt56, dwlt57, dwlt58, dwlt59, dwlt60, dwlt61, dwlt62, dwlt63, dwlt64;

logic signed [15:0] dwltw1, dwltw2, dwltw3, dwltw4, dwltw5, dwltw6, dwltw7, dwltw8, dwltw9, dwltw10, dwltw11, dwltw12, dwltw13, dwltw14, dwltw15, dwltw16, dwltw17, dwltw18, dwltw19, dwltw20, dwltw21, dwltw22, dwltw23, dwltw24, dwltw25, dwltw26, dwltw27, dwltw28, dwltw29, dwltw30, dwltw31, dwltw32, dwltw33, dwltw34, dwltw35, dwltw36, dwltw37, dwltw38, dwltw39, dwltw40, dwltw41, dwltw42, dwltw43, dwltw44, dwltw45, dwltw46, dwltw47, dwltw48, dwltw49, dwltw50, dwltw51, dwltw52, dwltw53, dwltw54, dwltw55, dwltw56, dwltw57, dwltw58, dwltw59, dwltw60, dwltw61, dwltw62, dwltw63, dwltw64;

logic signed [15:0] dwltwl1, dwltwl2, dwltwl3, dwltwl4, dwltwl5, dwltwl6, dwltwl7, dwltwl8, dwltwl9, dwltwl10, dwltwl11, dwltwl12, dwltwl13, dwltwl14, dwltwl15, dwltwl16, dwltwl17, dwltwl18, dwltwl19, dwltwl20, dwltwl21, dwltwl22, dwltwl23, dwltwl24, dwltwl25, dwltwl26, dwltwl27, dwltwl28, dwltwl29, dwltwl30, dwltwl31, dwltwl32, dwltwl33, dwltwl34, dwltwl35, dwltwl36, dwltwl37, dwltwl38, dwltwl39, dwltwl40, dwltwl41, dwltwl42, dwltwl43, dwltwl44, dwltwl45, dwltwl46, dwltwl47, dwltwl48, dwltwl49, dwltwl50, dwltwl51, dwltwl52, dwltwl53, dwltwl54, dwltwl55, dwltwl56, dwltwl57, dwltwl58, dwltwl59, dwltwl60, dwltwl61, dwltwl62, dwltwl63, dwltwl64;

logic signed [15:0] dwltwlq1, dwltwlq2, dwltwlq3, dwltwlq4, dwltwlq5, dwltwlq6, dwltwlq7, dwltwlq8, dwltwlq9, dwltwlq10, dwltwlq11, dwltwlq12, dwltwlq13, dwltwlq14, dwltwlq15, dwltwlq16, dwltwlq17, dwltwlq18, dwltwlq19, dwltwlq20, dwltwlq21, dwltwlq22, dwltwlq23, dwltwlq24, dwltwlq25, dwltwlq26, dwltwlq27, dwltwlq28, dwltwlq29, dwltwlq30, dwltwlq31, dwltwlq32, dwltwlq33, dwltwlq34, dwltwlq35, dwltwlq36, dwltwlq37, dwltwlq38, dwltwlq39, dwltwlq40, dwltwlq41, dwltwlq42, dwltwlq43, dwltwlq44, dwltwlq45, dwltwlq46, dwltwlq47, dwltwlq48, dwltwlq49, dwltwlq50, dwltwlq51, dwltwlq52, dwltwlq53, dwltwlq54, dwltwlq55, dwltwlq56, dwltwlq57, dwltwlq58, dwltwlq59, dwltwlq60, dwltwlq61, dwltwlq62, dwltwlq63, dwltwlq64;

transform u1 (d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28, d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61,d62,d63,d64,dw1,dw2,dw3,dw4,dw5,dw6,dw7,dw8,dw9,dw10,dw11,dw12,dw13,dw14,dw15,dw16,dw17,dw18,dw19,dw20,dw21,dw22,dw23,dw24,dw25,dw26,dw27,dw28,dw29,dw30,dw31,dw32,dw33,dw34,dw35,dw36,dw37,dw38,dw39,dw40,dw41,dw42,dw43,dw44,dw45,dw46,dw47,dw48,dw49,dw50,dw51,dw52,dw53,dw54,dw55,dw56,dw57,dw58,dw59,dw60,dw61,dw62,dw63,dw64);

pipo u2 (reset, dp_enable1, dw1,dw2,dw3,dw4,dw5,dw6,dw7,dw8,dw9,dw10,dw11,dw12,dw13,dw14,dw15,dw16,dw17,dw18,dw19,dw20,dw21,dw22,dw23,dw24,dw25,dw26,dw27,dw28,dw29,dw30,dw31,dw32,dw33,dw34,dw35,dw36,dw37,dw38,dw39,dw40,dw41,dw42,dw43,dw44,dw45,dw46,dw47,dw48,dw49,dw50,dw51,dw52,dw53,dw54,dw55,dw56,dw57,dw58,dw59,dw60,dw61,dw62,dw63,dw64, dwl1,dwl2,dwl3,dwl4,dwl5,dwl6,dwl7,dwl8,dwl9,dwl10,dwl11,dwl12,dwl13,dwl14,dwl15,dwl16,dwl17,dwl18,dwl19,dwl20,dwl21,dwl22,dwl23,dwl24,dwl25,dwl26,dwl27,dwl28,dwl29,dwl30,dwl31,dwl32,dwl33,dwl34,dwl35,dwl36,dwl37,dwl38,dwl39,dwl40,dwl41,dwl42,dwl43,dwl44,dwl45,dwl46,dwl47,dwl48,dwl49,dwl50,dwl51,dwl52,dwl53,dwl54,dwl55,dwl56,dwl57,dwl58,dwl59,dwl60,dwl61,dwl62,dwl63,dwl64);

transpose u3 (reset, dp_enable2, dwl1,dwl2,dwl3,dwl4,dwl5,dwl6,dwl7,dwl8,dwl9,dwl10,dwl11,dwl12,dwl13,dwl14,dwl15,dwl16,dwl17,dwl18,dwl19,dwl20,dwl21,dwl22,dwl23,dwl24,dwl25,dwl26,dwl27,dwl28,dwl29,dwl30,dwl31,dwl32,dwl33,dwl34,dwl35,dwl36,dwl37,dwl38,dwl39,dwl40,dwl41,dwl42,dwl43,dwl44,dwl45,dwl46,dwl47,dwl48,dwl49,dwl50,dwl51,dwl52,dwl53,dwl54,dwl55,dwl56,dwl57,dwl58,dwl59,dwl60,dwl61,dwl62,dwl63,dwl64,dwlt1, dwlt2, dwlt3, dwlt4, dwlt5, dwlt6, dwlt7, dwlt8, dwlt9, dwlt10, dwlt11, dwlt12, dwlt13, dwlt14, dwlt15, dwlt16, dwlt17, dwlt18, dwlt19, dwlt20, dwlt21, dwlt22, dwlt23, dwlt24, dwlt25, dwlt26, dwlt27, dwlt28, dwlt29, dwlt30, dwlt31, dwlt32, dwlt33, dwlt34, dwlt35, dwlt36, dwlt37, dwlt38, dwlt39, dwlt40, dwlt41, dwlt42, dwlt43, dwlt44, dwlt45, dwlt46, dwlt47, dwlt48, dwlt49, dwlt50, dwlt51, dwlt52, dwlt53, dwlt54, dwlt55,dwlt56, dwlt57, dwlt58, dwlt59, dwlt60, dwlt61, dwlt62, dwlt63, dwlt64);

transform u4 (dwlt1, dwlt2, dwlt3, dwlt4, dwlt5, dwlt6, dwlt7, dwlt8, dwlt9, dwlt10, dwlt11, dwlt12, dwlt13, dwlt14, dwlt15, dwlt16, dwlt17, dwlt18, dwlt19, dwlt20, dwlt21, dwlt22, dwlt23, dwlt24, dwlt25, dwlt26, dwlt27, dwlt28, dwlt29, dwlt30, dwlt31, dwlt32, dwlt33, dwlt34, dwlt35, dwlt36, dwlt37, dwlt38, dwlt39, dwlt40, dwlt41, dwlt42, dwlt43, dwlt44, dwlt45, dwlt46, dwlt47, dwlt48, dwlt49, dwlt50, dwlt51, dwlt52, dwlt53, dwlt54, dwlt55, dwlt56, dwlt57, dwlt58, dwlt59, dwlt60, dwlt61, dwlt62, dwlt63, dwlt64, dwltw1, dwltw2, dwltw3, dwltw4, dwltw5, dwltw6, dwltw7, dwltw8, dwltw9 , dwltw10, dwltw11, dwltw12, dwltw13, dwltw14, dwltw15, dwltw16, dwltw17, dwltw18, dwltw19 , dwltw20, dwltw21, dwltw22, dwltw23, dwltw24, dwltw25, dwltw26, dwltw27, dwltw28, dwltw29 , dwltw30, dwltw31, dwltw32, dwltw33, dwltw34, dwltw35, dwltw36, dwltw37, dwltw38, dwltw39 , dwltw40, dwltw41, dwltw42, dwltw43, dwltw44, dwltw45, dwltw46, dwltw47, dwltw48, dwltw49 , dwltw50, dwltw51, dwltw52, dwltw53, dwltw54, dwltw55, dwltw56, dwltw57, dwltw58, dwltw59 , dwltw60, dwltw61, dwltw62, dwltw63, dwltw64);

pipo u5 (reset, dp_enable3, dwltw1, dwltw2, dwltw3, dwltw4, dwltw5, dwltw6, dwltw7, dwltw8, dwltw9 , dwltw10, dwltw11, dwltw12, dwltw13, dwltw14, dwltw15, dwltw16, dwltw17, dwltw18, dwltw19, dwltw20, dwltw21, dwltw22, dwltw23, dwltw24, dwltw25, dwltw26, dwltw27, dwltw28, dwltw29, dwltw30, dwltw31, dwltw32, dwltw33, dwltw34, dwltw35, dwltw36, dwltw37, dwltw38, dwltw39, dwltw40, dwltw41, dwltw42, dwltw43, dwltw44, dwltw45, dwltw46, dwltw47, dwltw48, dwltw49, dwltw50, dwltw51, dwltw52, dwltw53, dwltw54, dwltw55, dwltw56, dwltw57, dwltw58, dwltw59, dwltw60, dwltw61, dwltw62, dwltw63, dwltw64, dwltwl1, dwltwl2, dwltwl3, dwltwl4, dwltwl5, dwltwl6, dwltwl7, dwltwl8, dwltwl9, dwltwl10, dwltwl11, dwltwl12, dwltwl13, dwltwl14, dwltwl15, dwltwl16, dwltwl17, dwltwl18, dwltwl19, dwltwl20, dwltwl21, dwltwl22, dwltwl23, dwltwl24, dwltwl25, dwltwl26, dwltwl27, dwltwl28, dwltwl29, dwltwl30, dwltwl31, dwltwl32, dwltwl33, dwltwl34, dwltwl35, dwltwl36, dwltwl37, dwltwl38, dwltwl39, dwltwl40, dwltwl41, dwltwl42, dwltwl43, dwltwl44, dwltwl45, dwltwl46, dwltwl47, dwltwl48, dwltwl49, dwltwl50, dwltwl51, dwltwl52, dwltwl53, dwltwl54, dwltwl55, dwltwl56, dwltwl57, dwltwl58, dwltwl59, dwltwl60, dwltwl61, dwltwl62, dwltwl63, dwltwl64 );

quantization u6 (dwltwl1, dwltwl2, dwltwl3, dwltwl4, dwltwl5, dwltwl6, dwltwl7, dwltwl8, dwltwl9, dwltwl10, dwltwl11, dwltwl12, dwltwl13, dwltwl14, dwltwl15, dwltwl16, dwltwl17, dwltwl18, dwltwl19, dwltwl20, dwltwl21, dwltwl22, dwltwl23, dwltwl24, dwltwl25, dwltwl26, dwltwl27, dwltwl28, dwltwl29, dwltwl30, dwltwl31, dwltwl32, dwltwl33, dwltwl34, dwltwl35, dwltwl36, dwltwl37, dwltwl38, dwltwl39, dwltwl40, dwltwl41, dwltwl42, dwltwl43, dwltwl44, dwltwl45, dwltwl46, dwltwl47, dwltwl48, dwltwl49, dwltwl50, dwltwl51, dwltwl52, dwltwl53, dwltwl54, dwltwl55, dwltwl56, dwltwl57, dwltwl58, dwltwl59, dwltwl60, dwltwl61, dwltwl62, dwltwl63, dwltwl64, dwltwlq1, dwltwlq2, dwltwlq3, dwltwlq4, dwltwlq5, dwltwlq6, dwltwlq7, dwltwlq8, dwltwlq9, dwltwlq10, dwltwlq11, dwltwlq12, dwltwlq13, dwltwlq14, dwltwlq15, dwltwlq16, dwltwlq17, dwltwlq18, dwltwlq19, dwltwlq20, dwltwlq21, dwltwlq22, dwltwlq23, dwltwlq24, dwltwlq25, dwltwlq26, dwltwlq27, dwltwlq28, dwltwlq29, dwltwlq30, dwltwlq31, dwltwlq32, dwltwlq33, dwltwlq34, dwltwlq35, dwltwlq36, dwltwlq37, dwltwlq38, dwltwlq39, dwltwlq40, dwltwlq41, dwltwlq42, dwltwlq43, dwltwlq44, dwltwlq45, dwltwlq46, dwltwlq47, dwltwlq48, dwltwlq49, dwltwlq50, dwltwlq51, dwltwlq52, dwltwlq53, dwltwlq54, dwltwlq55, dwltwlq56, dwltwlq57, dwltwlq58, dwltwlq59, dwltwlq60, dwltwlq61, dwltwlq62, dwltwlq63, dwltwlq64);

zigzag u7 (reset, dp_enable4, dwltwlq1, dwltwlq2, dwltwlq3, dwltwlq4, dwltwlq5, dwltwlq6, dwltwlq7, dwltwlq8, dwltwlq9, dwltwlq10, dwltwlq11, dwltwlq12, dwltwlq13, dwltwlq14, dwltwlq15, dwltwlq16, dwltwlq17, dwltwlq18, dwltwlq19, dwltwlq20, dwltwlq21, dwltwlq22, dwltwlq23, dwltwlq24, dwltwlq25, dwltwlq26, dwltwlq27, dwltwlq28, dwltwlq29, dwltwlq30, dwltwlq31, dwltwlq32, dwltwlq33, dwltwlq34, dwltwlq35, dwltwlq36, dwltwlq37, dwltwlq38, dwltwlq39, dwltwlq40, dwltwlq41, dwltwlq42, dwltwlq43, dwltwlq44, dwltwlq45, dwltwlq46, dwltwlq47, dwltwlq48, dwltwlq49, dwltwlq50, dwltwlq51, dwltwlq52, dwltwlq53, dwltwlq54, dwltwlq55, dwltwlq56, dwltwlq57, dwltwlq58, dwltwlq59, dwltwlq60, dwltwlq61, dwltwlq62, dwltwlq63, dwltwlq64, do1,do2,do3,do4,do5,do6,do7,do8,do9,do10,do11,do12,do13,do14,do15,do16,do17,do18,do19,do20,do21,do22,do23,do24,do25,do26,do27,do28,do29,do30,do31,do32,do33,do34,do35,do36,do37,do38,do39,do40,do41,do42,do43,do44,do45,do46,do47,do48,do49,do50,do51,do52,do53,do54,do55,do56,do57,do58,do59,do60,do61,do62,do63,do64); 

endmodule
