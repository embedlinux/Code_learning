library verilog;
use verilog.vl_types.all;
entity dpram_tb is
end dpram_tb;
