
module adder_DW01_add_64_1 ( A, B, CI, SUM, CO );
input  [63:0] A;
input  [63:0] B;
output [63:0] SUM;
input  CI;
output CO;
    wire n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, 
        n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
        n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
        n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
        n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
        n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
        n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
        n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
        n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
        n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
        n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
        n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
        n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
        n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
        n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
        n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
        n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
        n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
        n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
        n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
        n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
        n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
        n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
        n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
        n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
        n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
        n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
        n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
        n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
        n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
        n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
        n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
        n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
        n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
        n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
        n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
        n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
        n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
        n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
        n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
        n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
        n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
        n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
        n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
        n620, n621, n622, n623, n624, n625, n626;
    INV2 U5 ( .O(n343), .I(n188) );
    INV2 U6 ( .O(n219), .I(n218) );
    INV2 U7 ( .O(n375), .I(n171) );
    INV2 U8 ( .O(n209), .I(n208) );
    OR2P U9 ( .O(n49), .I1(n290), .I2(n447) );
    INV2 U10 ( .O(n136), .I(n49) );
    ND4P U11 ( .O(n61), .I1(n336), .I2(n271), .I3(n517), .I4(n518) );
    OAI12 U12 ( .O(n448), .A1(n546), .B1(n366), .B2(n501) );
    NR4P U13 ( .O(n398), .I1(n212), .I2(n50), .I3(n530), .I4(n504) );
    INV1 U14 ( .O(n50), .I(n580) );
    AO12 U15 ( .O(n78), .A1(n502), .B1(n51), .B2(n52) );
    INV2 U16 ( .O(n51), .I(B[38]) );
    INV1 U17 ( .O(n52), .I(A[38]) );
    NR4P U18 ( .O(n400), .I1(n214), .I2(n53), .I3(n544), .I4(n503) );
    INV1 U19 ( .O(n53), .I(n571) );
    OA12 U20 ( .O(n81), .A1(n82), .B1(n54), .B2(n404) );
    INV1 U21 ( .O(n54), .I(n549) );
    OR3 U22 ( .O(n505), .I1(n506), .I2(n507), .I3(n467) );
    AN2 U23 ( .O(n84), .I1(n565), .I2(n554) );
    OR2B1T U24 ( .O(n329), .I1(n558), .B1(n559) );
    INV3 U25 ( .O(n558), .I(n413) );
    OR2B1T U26 ( .O(n330), .I1(n85), .B1(n477) );
    AN2B1P U27 ( .O(n106), .I1(n382), .B1(n325) );
    XOR2 U28 ( .O(SUM[15]), .I1(n107), .I2(n66) );
    AN2B1P U29 ( .O(n202), .I1(n594), .B1(n267) );
    XOR2 U30 ( .O(SUM[49]), .I1(n239), .I2(n482) );
    XNR2 U31 ( .O(SUM[50]), .I1(n196), .I2(n150) );
    AN2B1P U32 ( .O(n197), .I1(n604), .B1(n262) );
    OAI12 U33 ( .O(n112), .A1(n349), .B1(n605), .B2(n607) );
    OAI112 U34 ( .O(n520), .A1(n375), .B1(n395), .C1(n521), .C2(n316) );
    OAI12 U35 ( .O(n137), .A1(n351), .B1(n600), .B2(n602) );
    OA12 U36 ( .O(n449), .A1(n55), .B1(n448), .B2(n136) );
    INV2 U37 ( .O(n55), .I(n450) );
    AO12P U38 ( .O(n479), .A1(n263), .B1(n608), .B2(n56) );
    INV1 U39 ( .O(n56), .I(n138) );
    AO12 U40 ( .O(n478), .A1(n265), .B1(n612), .B2(n57) );
    INV2 U41 ( .O(n57), .I(n139) );
    OAI12T U42 ( .O(n409), .A1(n259), .B1(n599), .B2(n150) );
    MAO222P U43 ( .O(n58), .A1(n618), .B1(B[60]), .C1(A[60]) );
    INV2 U44 ( .O(n619), .I(n58) );
    MOAI1T U45 ( .O(n59), .A1(n289), .A2(n619), .B1(A[61]), .B2(B[61]) );
    INV2 U46 ( .O(n144), .I(n59) );
    OAI112 U47 ( .O(n446), .A1(n294), .B1(n306), .C1(n208), .C2(n118) );
    AO12P U48 ( .O(n145), .A1(n446), .B1(n146), .B2(n69) );
    OA12P U49 ( .O(n60), .A1(n351), .B1(n600), .B2(n602) );
    INV2 U50 ( .O(n603), .I(n60) );
    INV2 U51 ( .O(n600), .I(n409) );
    INV2 U52 ( .O(n351), .I(n185) );
    AO12 U53 ( .O(n551), .A1(n270), .B1(n145), .B2(n393) );
    INV2 U54 ( .O(n393), .I(n533) );
    AN2T U55 ( .O(n290), .I1(n551), .I2(n321) );
    AO12 U56 ( .O(n292), .A1(n270), .B1(n145), .B2(n393) );
    AN3B1T U57 ( .O(n321), .I1(n414), .I2(n317), .B1(n538) );
    INV2 U58 ( .O(n324), .I(n61) );
    ND2F U59 ( .O(n560), .I1(n359), .I2(n329) );
    OAI112T U60 ( .O(n450), .A1(n308), .B1(n312), .C1(n218), .C2(n117) );
    INV2 U61 ( .O(n147), .I(n135) );
    AN2 U62 ( .O(n74), .I1(n535), .I2(n405) );
    AN2 U63 ( .O(n374), .I1(A[13]), .I2(B[13]) );
    AN2 U64 ( .O(n305), .I1(A[29]), .I2(B[29]) );
    AN2 U65 ( .O(n293), .I1(A[28]), .I2(B[28]) );
    AN2 U66 ( .O(n372), .I1(A[38]), .I2(B[38]) );
    AN2 U67 ( .O(n368), .I1(A[26]), .I2(B[26]) );
    AN2 U68 ( .O(n370), .I1(A[22]), .I2(B[22]) );
    AN2 U69 ( .O(n376), .I1(A[42]), .I2(B[42]) );
    AN2 U70 ( .O(n307), .I1(A[44]), .I2(B[44]) );
    AN2 U71 ( .O(n311), .I1(n129), .I2(B[45]) );
    AN2 U72 ( .O(n403), .I1(A[46]), .I2(B[46]) );
    AN2 U73 ( .O(n394), .I1(A[14]), .I2(B[14]) );
    AN2 U74 ( .O(n354), .I1(A[49]), .I2(B[49]) );
    AN2 U75 ( .O(n342), .I1(A[10]), .I2(B[10]) );
    AN2 U76 ( .O(n389), .I1(A[9]), .I2(B[9]) );
    AN2 U77 ( .O(n387), .I1(A[8]), .I2(B[8]) );
    AN2 U78 ( .O(n348), .I1(n128), .I2(B[53]) );
    AN2 U79 ( .O(n344), .I1(A[6]), .I2(B[6]) );
    AN2 U80 ( .O(n356), .I1(n131), .I2(B[57]) );
    AN2 U81 ( .O(n391), .I1(A[4]), .I2(B[4]) );
    AOI12 U82 ( .O(n430), .A1(n433), .B1(n431), .B2(n417) );
    AN2 U83 ( .O(n378), .I1(A[24]), .I2(B[24]) );
    AN2 U84 ( .O(n380), .I1(A[40]), .I2(B[40]) );
    AOI12 U85 ( .O(n420), .A1(n423), .B1(n421), .B2(n418) );
    AN2 U86 ( .O(n352), .I1(n130), .I2(B[55]) );
    OR2P U87 ( .O(n559), .I1(B[3]), .I2(n132) );
    OR2P U88 ( .O(n574), .I1(B[36]), .I2(A[36]) );
    INV2 U89 ( .O(n294), .I(n167) );
    OR2P U90 ( .O(n583), .I1(B[20]), .I2(A[20]) );
    INV2 U91 ( .O(n308), .I(n166) );
    OR2P U92 ( .O(n596), .I1(B[49]), .I2(A[49]) );
    OR2P U93 ( .O(n588), .I1(B[11]), .I2(A[11]) );
    OR2P U94 ( .O(n606), .I1(B[53]), .I2(n128) );
    OR2P U95 ( .O(n614), .I1(B[57]), .I2(n131) );
    AN2 U96 ( .O(n201), .I1(n616), .I2(n269) );
    AN2 U97 ( .O(n195), .I1(n277), .I2(n316) );
    AN2 U98 ( .O(n189), .I1(n534), .I2(n406) );
    AO12 U99 ( .O(n93), .A1(n433), .B1(n456), .B2(n417) );
    AO12 U100 ( .O(n96), .A1(n426), .B1(n452), .B2(n416) );
    AO12 U101 ( .O(n99), .A1(n437), .B1(n457), .B2(n419) );
    AO12 U102 ( .O(n104), .A1(n423), .B1(n451), .B2(n418) );
    AN2 U103 ( .O(n280), .I1(n583), .I2(n302) );
    AN2 U104 ( .O(n194), .I1(n206), .I2(n261) );
    AN2 U105 ( .O(n240), .I1(n548), .I2(n404) );
    AO12 U106 ( .O(n108), .A1(n188), .B1(n465), .B2(n466) );
    AN2 U107 ( .O(n196), .I1(n598), .I2(n259) );
    AN2 U108 ( .O(n283), .I1(n159), .I2(n392) );
    XOR2 U109 ( .O(n114), .I1(A[61]), .I2(B[61]) );
    AN2 U110 ( .O(n198), .I1(n556), .I2(n255) );
    OR2B1 U111 ( .O(n538), .I1(n592), .B1(n402) );
    BUF2 U112 ( .O(n402), .I(n455) );
    OR2 U113 ( .O(n549), .I1(B[47]), .I2(A[47]) );
    OR2B1 U114 ( .O(n468), .I1(n392), .B1(n160) );
    AN2T U115 ( .O(n62), .I1(n588), .I2(n466) );
    INV3 U116 ( .O(n469), .I(n62) );
    OR2 U117 ( .O(n519), .I1(B[12]), .I2(A[12]) );
    OR2 U118 ( .O(n578), .I1(B[27]), .I2(A[27]) );
    INV2 U119 ( .O(n503), .I(n207) );
    BUF2 U120 ( .O(n207), .I(n569) );
    OR2 U121 ( .O(n569), .I1(B[43]), .I2(A[43]) );
    OR2 U122 ( .O(n516), .I1(B[9]), .I2(A[9]) );
    AN2T U123 ( .O(n63), .I1(n553), .I2(n554) );
    INV3 U124 ( .O(n467), .I(n63) );
    OR2 U125 ( .O(n561), .I1(B[4]), .I2(A[4]) );
    OR2P U126 ( .O(n64), .I1(B[59]), .I2(n133) );
    INV3 U127 ( .O(n85), .I(n64) );
    BUF2 U128 ( .O(n286), .I(n305) );
    AN2 U129 ( .O(n281), .I1(n574), .I2(n300) );
    INV2 U130 ( .O(n529), .I(n583) );
    BUF2 U131 ( .O(n287), .I(n311) );
    OA12P U132 ( .O(n65), .A1(n332), .B1(n285), .B2(n525) );
    INV1 U133 ( .O(n494), .I(n65) );
    INV3 U134 ( .O(n404), .I(n176) );
    BUF2 U135 ( .O(n176), .I(n403) );
    OR2 U136 ( .O(n66), .I1(n178), .I2(n464) );
    INV2 U137 ( .O(n395), .I(n178) );
    AN2 U138 ( .O(n234), .I1(n587), .I2(n395) );
    AN2 U139 ( .O(n227), .I1(n158), .I2(n388) );
    BUF2 U140 ( .O(n158), .I(n562) );
    OR2B1 U141 ( .O(n111), .I1(n84), .B1(n345) );
    INV2 U142 ( .O(n507), .I(n384) );
    BUF2 U143 ( .O(n384), .I(n160) );
    AO12 U144 ( .O(n113), .A1(n184), .B1(n479), .B2(n610) );
    INV2 U145 ( .O(n353), .I(n184) );
    INV2 U146 ( .O(n506), .I(n159) );
    BUF2 U147 ( .O(n159), .I(n561) );
    AN2P U148 ( .O(n67), .I1(n339), .I2(n555) );
    INV1 U149 ( .O(n115), .I(n67) );
    INV2 U150 ( .O(n458), .I(n555) );
    OR2 U151 ( .O(n444), .I1(n497), .I2(n495) );
    BUF2 U152 ( .O(n206), .I(n584) );
    OAI12P U153 ( .O(n495), .A1(n261), .B1(n496), .B2(n438) );
    INV1 U154 ( .O(n526), .I(n497) );
    AN2 U155 ( .O(n532), .I1(n209), .I2(n398) );
    INV2 U156 ( .O(n399), .I(n398) );
    INV3 U157 ( .O(n528), .I(n217) );
    INV3 U158 ( .O(n217), .I(n216) );
    INV2 U159 ( .O(n527), .I(n436) );
    AN2P U160 ( .O(n68), .I1(n277), .I2(n415) );
    INV1 U161 ( .O(n442), .I(n68) );
    OR2P U162 ( .O(n415), .I1(B[13]), .I2(A[13]) );
    BUF2 U163 ( .O(n277), .I(n519) );
    OR2B1 U164 ( .O(n470), .I1(n388), .B1(n385) );
    BUF2 U165 ( .O(n385), .I(n516) );
    INV2 U166 ( .O(n69), .I(n445) );
    ND2P U167 ( .O(n146), .I1(n552), .I2(n147) );
    INV2 U168 ( .O(n504), .I(n203) );
    BUF2 U169 ( .O(n203), .I(n578) );
    INV3 U170 ( .O(n306), .I(n286) );
    OR2P U171 ( .O(n317), .I1(B[35]), .I2(A[35]) );
    OR2P U172 ( .O(n539), .I1(B[32]), .I2(A[32]) );
    INV2 U173 ( .O(n592), .I(n539) );
    AO12 U174 ( .O(n428), .A1(n70), .B1(n455), .B2(n333) );
    INV1 U175 ( .O(n70), .I(n323) );
    INV2 U176 ( .O(n334), .I(n333) );
    INV2 U177 ( .O(n530), .I(n432) );
    INV3 U178 ( .O(n531), .I(n213) );
    INV3 U179 ( .O(n213), .I(n212) );
    INV2 U180 ( .O(n379), .I(n165) );
    BUF2 U181 ( .O(n165), .I(n378) );
    INV3 U182 ( .O(n542), .I(n211) );
    INV3 U183 ( .O(n211), .I(n210) );
    INV3 U184 ( .O(n221), .I(n220) );
    AN2 U185 ( .O(n522), .I1(n584), .I2(n319) );
    INV3 U186 ( .O(n319), .I(n318) );
    INV2 U187 ( .O(n496), .I(n206) );
    INV2 U188 ( .O(n544), .I(n422) );
    INV3 U189 ( .O(n545), .I(n215) );
    INV3 U190 ( .O(n215), .I(n214) );
    INV2 U191 ( .O(n381), .I(n164) );
    BUF2 U192 ( .O(n164), .I(n380) );
    AN2 U193 ( .O(n546), .I1(n219), .I2(n400) );
    INV2 U194 ( .O(n401), .I(n400) );
    BUF2 U195 ( .O(n166), .I(n307) );
    INV3 U196 ( .O(n312), .I(n287) );
    INV2 U197 ( .O(n498), .I(n204) );
    BUF2 U198 ( .O(n204), .I(n581) );
    OR2 U199 ( .O(n581), .I1(B[23]), .I2(A[23]) );
    OR2P U200 ( .O(n71), .I1(n73), .I2(n72) );
    INV2 U201 ( .O(n367), .I(n71) );
    OR2 U202 ( .O(n72), .I1(n527), .I2(n498) );
    OR2 U203 ( .O(n73), .I1(n528), .I2(n529) );
    AN2 U204 ( .O(n127), .I1(n586), .I2(n587) );
    OR2B1 U205 ( .O(n517), .I1(n343), .B1(n512) );
    OR2 U206 ( .O(n518), .I1(n390), .I2(n469) );
    OR2 U207 ( .O(n271), .I1(n469), .I2(n470) );
    INV2 U208 ( .O(n512), .I(n469) );
    AN2P U209 ( .O(n513), .I1(n386), .I2(n562) );
    INV2 U210 ( .O(n515), .I(n158) );
    INV2 U211 ( .O(n514), .I(n386) );
    BUF3 U212 ( .O(n386), .I(n385) );
    INV2 U213 ( .O(n406), .I(n405) );
    AN2 U214 ( .O(n75), .I1(n414), .I2(n76) );
    INV2 U215 ( .O(n76), .I(n453) );
    INV2 U216 ( .O(n543), .I(n574) );
    OR2P U217 ( .O(n417), .I1(B[26]), .I2(A[26]) );
    OR2P U218 ( .O(n416), .I1(B[38]), .I2(A[38]) );
    INV2 U219 ( .O(n502), .I(n205) );
    BUF2 U220 ( .O(n205), .I(n572) );
    OR2 U221 ( .O(n572), .I1(B[39]), .I2(A[39]) );
    INV3 U222 ( .O(n373), .I(n174) );
    BUF2 U223 ( .O(n174), .I(n372) );
    OR2P U224 ( .O(n77), .I1(n79), .I2(n78) );
    INV2 U225 ( .O(n366), .I(n77) );
    OR2 U226 ( .O(n79), .I1(n542), .I2(n543) );
    OR2P U227 ( .O(n419), .I1(B[22]), .I2(A[22]) );
    OR2P U228 ( .O(n418), .I1(B[42]), .I2(A[42]) );
    INV3 U229 ( .O(n377), .I(n175) );
    BUF2 U230 ( .O(n175), .I(n376) );
    AN2 U231 ( .O(n459), .I1(n319), .I2(n626) );
    OAI12P U232 ( .O(n626), .A1(n298), .B1(n274), .B2(n65) );
    AN2 U233 ( .O(n464), .I1(n587), .I2(n80) );
    INV2 U234 ( .O(n80), .I(n461) );
    INV1 U235 ( .O(n82), .I(n325) );
    OR2P U236 ( .O(n382), .I1(B[47]), .I2(A[47]) );
    INV2 U237 ( .O(n602), .I(n601) );
    ND4P U238 ( .O(n83), .I1(n510), .I2(n511), .I3(n338), .I4(n272) );
    INV2 U239 ( .O(n509), .I(n83) );
    OR2 U240 ( .O(n510), .I1(n345), .I2(n363) );
    OR2 U241 ( .O(n511), .I1(n408), .I2(n363) );
    INV3 U242 ( .O(n345), .I(n187) );
    BUF2 U243 ( .O(n187), .I(n344) );
    OR2 U244 ( .O(n272), .I1(n467), .I2(n468) );
    BUF2 U245 ( .O(n363), .I(n467) );
    OAI12P U246 ( .O(n565), .A1(n408), .B1(n507), .B2(n564) );
    INV2 U247 ( .O(n611), .I(n610) );
    XNR2 U248 ( .O(SUM[24]), .I1(n86), .I2(n624) );
    AN2 U249 ( .O(n86), .I1(n327), .I2(n379) );
    XNR2 U250 ( .O(SUM[16]), .I1(n87), .I2(n285) );
    AN2 U251 ( .O(n87), .I1(n221), .I2(n332) );
    INV2 U252 ( .O(n341), .I(n340) );
    XOR2 U253 ( .O(SUM[55]), .I1(n237), .I2(n411) );
    AN2 U254 ( .O(n237), .I1(n610), .I2(n353) );
    XOR2 U255 ( .O(SUM[13]), .I1(n233), .I2(n462) );
    AN2 U256 ( .O(n233), .I1(n415), .I2(n375) );
    XNR2 U257 ( .O(SUM[58]), .I1(n201), .I2(n152) );
    XNR2 U258 ( .O(SUM[12]), .I1(n195), .I2(n148) );
    OR2 U259 ( .O(n88), .I1(n85), .I2(n180) );
    INV3 U260 ( .O(n361), .I(n180) );
    XOR2 U261 ( .O(SUM[32]), .I1(n282), .I2(n320) );
    INV1 U262 ( .O(n488), .I(n320) );
    AN2 U263 ( .O(n282), .I1(n539), .I2(n334) );
    XOR2 U264 ( .O(SUM[33]), .I1(n230), .I2(n454) );
    AN2 U265 ( .O(n230), .I1(n402), .I2(n323) );
    XOR2 U266 ( .O(SUM[31]), .I1(n232), .I2(n489) );
    AN2 U267 ( .O(n232), .I1(n535), .I2(n347) );
    XNR2 U268 ( .O(SUM[34]), .I1(n89), .I2(n453) );
    AN2 U269 ( .O(n89), .I1(n414), .I2(n365) );
    BUF2 U270 ( .O(n170), .I(n364) );
    XNR2 U271 ( .O(SUM[30]), .I1(n189), .I2(n123) );
    XOR2 U272 ( .O(SUM[35]), .I1(n242), .I2(n90) );
    OR2 U273 ( .O(n90), .I1(n75), .I2(n170) );
    AN2 U274 ( .O(n242), .I1(n317), .I2(n154) );
    XOR2 U275 ( .O(SUM[29]), .I1(n223), .I2(n625) );
    BUF2 U276 ( .O(n167), .I(n293) );
    AN2 U277 ( .O(n223), .I1(n536), .I2(n306) );
    XNR2 U278 ( .O(SUM[36]), .I1(n281), .I2(n487) );
    XNR2 U279 ( .O(SUM[28]), .I1(n91), .I2(n122) );
    AN2 U280 ( .O(n91), .I1(n209), .I2(n294) );
    XNR2 U281 ( .O(SUM[37]), .I1(n92), .I2(n121) );
    AN2 U282 ( .O(n92), .I1(n211), .I2(n314) );
    XOR2 U283 ( .O(SUM[27]), .I1(n190), .I2(n93) );
    INV3 U284 ( .O(n369), .I(n172) );
    BUF2 U285 ( .O(n172), .I(n368) );
    AN2 U286 ( .O(n190), .I1(n203), .I2(n251) );
    XOR2 U287 ( .O(SUM[38]), .I1(n94), .I2(n452) );
    AN2 U288 ( .O(n94), .I1(n416), .I2(n373) );
    OAI12P U289 ( .O(n452), .A1(n314), .B1(n542), .B2(n121) );
    XOR2 U290 ( .O(SUM[26]), .I1(n95), .I2(n456) );
    AN2 U291 ( .O(n95), .I1(n417), .I2(n369) );
    OAI12P U292 ( .O(n456), .A1(n296), .B1(n531), .B2(n125) );
    XOR2 U293 ( .O(SUM[39]), .I1(n191), .I2(n96) );
    AN2 U294 ( .O(n191), .I1(n205), .I2(n253) );
    XNR2 U295 ( .O(SUM[25]), .I1(n97), .I2(n125) );
    AN2 U296 ( .O(n97), .I1(n213), .I2(n296) );
    XNR2 U297 ( .O(SUM[40]), .I1(n98), .I2(n621) );
    AN2 U298 ( .O(n98), .I1(n326), .I2(n381) );
    XOR2 U299 ( .O(SUM[23]), .I1(n192), .I2(n99) );
    INV3 U300 ( .O(n371), .I(n173) );
    BUF2 U301 ( .O(n173), .I(n370) );
    AN2 U302 ( .O(n192), .I1(n204), .I2(n257) );
    XNR2 U303 ( .O(SUM[41]), .I1(n100), .I2(n126) );
    AN2 U304 ( .O(n100), .I1(n215), .I2(n304) );
    XOR2 U305 ( .O(SUM[22]), .I1(n101), .I2(n457) );
    AN2 U306 ( .O(n101), .I1(n419), .I2(n371) );
    OAI12P U307 ( .O(n457), .A1(n310), .B1(n528), .B2(n124) );
    XOR2 U308 ( .O(SUM[42]), .I1(n102), .I2(n451) );
    AN2 U309 ( .O(n102), .I1(n418), .I2(n377) );
    OAI12P U310 ( .O(n451), .A1(n304), .B1(n545), .B2(n126) );
    XNR2 U311 ( .O(SUM[21]), .I1(n103), .I2(n124) );
    AN2 U312 ( .O(n103), .I1(n217), .I2(n310) );
    XOR2 U313 ( .O(SUM[43]), .I1(n193), .I2(n104) );
    AN2 U314 ( .O(n193), .I1(n207), .I2(n249) );
    XNR2 U315 ( .O(SUM[20]), .I1(n280), .I2(n492) );
    XNR2 U316 ( .O(SUM[44]), .I1(n105), .I2(n119) );
    AN2 U317 ( .O(n105), .I1(n219), .I2(n308) );
    XNR2 U318 ( .O(SUM[19]), .I1(n194), .I2(n460) );
    XOR2 U319 ( .O(SUM[45]), .I1(n222), .I2(n622) );
    AN2 U320 ( .O(n222), .I1(n550), .I2(n312) );
    XOR2 U321 ( .O(SUM[18]), .I1(n231), .I2(n626) );
    INV3 U322 ( .O(n274), .I(n273) );
    AN2 U323 ( .O(n231), .I1(n319), .I2(n397) );
    XNR2 U324 ( .O(SUM[46]), .I1(n240), .I2(n120) );
    INV3 U325 ( .O(n525), .I(n221) );
    XOR2 U326 ( .O(SUM[47]), .I1(n106), .I2(n483) );
    AN2 U327 ( .O(n107), .I1(n586), .I2(n341) );
    XOR2 U328 ( .O(SUM[48]), .I1(n202), .I2(n593) );
    XNR2 U329 ( .O(SUM[14]), .I1(n234), .I2(n461) );
    BUF2 U330 ( .O(n178), .I(n394) );
    AN2 U331 ( .O(n239), .I1(n596), .I2(n355) );
    XOR2 U332 ( .O(SUM[11]), .I1(n228), .I2(n108) );
    AN2 U333 ( .O(n228), .I1(n588), .I2(n336) );
    XOR2 U334 ( .O(SUM[10]), .I1(n225), .I2(n465) );
    OAI12P U335 ( .O(n465), .A1(n390), .B1(n563), .B2(n514) );
    AN2 U336 ( .O(n225), .I1(n466), .I2(n343) );
    OR2 U337 ( .O(n109), .I1(n110), .I2(n185) );
    INV1 U338 ( .O(n110), .I(n601) );
    XOR2 U339 ( .O(SUM[9]), .I1(n235), .I2(n471) );
    AN2 U340 ( .O(n235), .I1(n386), .I2(n390) );
    XOR2 U341 ( .O(SUM[52]), .I1(n197), .I2(n137) );
    XNR2 U342 ( .O(SUM[8]), .I1(n227), .I2(n247) );
    XOR2 U343 ( .O(SUM[53]), .I1(n236), .I2(n480) );
    AN2 U344 ( .O(n236), .I1(n606), .I2(n349) );
    XOR2 U345 ( .O(SUM[7]), .I1(n229), .I2(n111) );
    AN2 U346 ( .O(n229), .I1(n553), .I2(n338) );
    XOR2 U347 ( .O(SUM[54]), .I1(n200), .I2(n112) );
    AN2 U348 ( .O(n200), .I1(n608), .I2(n264) );
    XOR2 U349 ( .O(SUM[6]), .I1(n226), .I2(n565) );
    AN2 U350 ( .O(n226), .I1(n554), .I2(n345) );
    XOR2 U351 ( .O(SUM[56]), .I1(n199), .I2(n113) );
    AN2 U352 ( .O(n199), .I1(n612), .I2(n266) );
    XOR2 U353 ( .O(SUM[5]), .I1(n241), .I2(n412) );
    AN2 U354 ( .O(n241), .I1(n384), .I2(n408) );
    XOR2 U355 ( .O(SUM[57]), .I1(n238), .I2(n140) );
    AN2 U356 ( .O(n238), .I1(n614), .I2(n357) );
    XNR2 U357 ( .O(SUM[4]), .I1(n283), .I2(n481) );
    XNR2 U358 ( .O(SUM[60]), .I1(n475), .I2(n618) );
    XNR2 U359 ( .O(SUM[61]), .I1(n114), .I2(n149) );
    XNR2 U360 ( .O(SUM[2]), .I1(n198), .I2(n116) );
    XOR2 U361 ( .O(SUM[1]), .I1(n362), .I2(n115) );
    AN2 U362 ( .O(SUM[0]), .I1(n362), .I2(n284) );
    OR2 U363 ( .O(n284), .I1(B[0]), .I2(A[0]) );
    BUF2 U364 ( .O(n171), .I(n374) );
    INV3 U365 ( .O(n388), .I(n179) );
    BUF2 U366 ( .O(n179), .I(n387) );
    OAI12P U367 ( .O(n445), .A1(n532), .B1(n367), .B2(n497) );
    NR2T U368 ( .O(n523), .I1(n274), .I2(n525) );
    OAI12 U369 ( .O(n439), .A1(n298), .B1(n524), .B2(n332) );
    INV3 U370 ( .O(n392), .I(n177) );
    BUF2 U371 ( .O(n177), .I(n391) );
    AOI12 U372 ( .O(n434), .A1(n437), .B1(n435), .B2(n419) );
    INV2 U373 ( .O(n521), .I(n463) );
    INV3 U374 ( .O(n390), .I(n163) );
    BUF2 U375 ( .O(n163), .I(n389) );
    AOI12 U376 ( .O(n427), .A1(n364), .B1(n428), .B2(n429) );
    AOI12 U377 ( .O(n424), .A1(n426), .B1(n425), .B2(n416) );
    AOI12 U378 ( .O(n438), .A1(n396), .B1(n439), .B2(n319) );
    INV2 U379 ( .O(n607), .I(n606) );
    BUF3 U380 ( .O(n157), .I(n155) );
    INV2 U381 ( .O(n615), .I(n614) );
    OAI12 U382 ( .O(n489), .A1(n406), .B1(n575), .B2(n123) );
    OAI12 U383 ( .O(n483), .A1(n404), .B1(n566), .B2(n120) );
    BUF2 U384 ( .O(n188), .I(n342) );
    INV2 U385 ( .O(n597), .I(n596) );
    INV2 U386 ( .O(n355), .I(n183) );
    BUF2 U387 ( .O(n183), .I(n354) );
    INV3 U388 ( .O(n349), .I(n186) );
    BUF2 U389 ( .O(n186), .I(n348) );
    INV2 U390 ( .O(n564), .I(n412) );
    BUF2 U391 ( .O(n412), .I(n476) );
    BUF2 U392 ( .O(n184), .I(n352) );
    INV2 U393 ( .O(n357), .I(n182) );
    BUF2 U394 ( .O(n182), .I(n356) );
    BUF3 U395 ( .O(n155), .I(B[1]) );
    OA12P U396 ( .O(n116), .A1(n339), .B1(n328), .B2(n458) );
    OA12P U397 ( .O(n117), .A1(n249), .B1(n503), .B2(n420) );
    OA12P U398 ( .O(n118), .A1(n251), .B1(n504), .B2(n430) );
    OA12P U399 ( .O(n119), .A1(n117), .B1(n621), .B2(n401) );
    OA12P U400 ( .O(n120), .A1(n312), .B1(n567), .B2(n484) );
    OA12P U401 ( .O(n121), .A1(n300), .B1(n543), .B2(n487) );
    OA12P U402 ( .O(n122), .A1(n118), .B1(n624), .B2(n399) );
    OA12P U403 ( .O(n123), .A1(n306), .B1(n576), .B2(n490) );
    OA12P U404 ( .O(n124), .A1(n302), .B1(n529), .B2(n492) );
    AOI12P U405 ( .O(n125), .A1(n165), .B1(n491), .B2(n327) );
    AOI12P U406 ( .O(n126), .A1(n164), .B1(n485), .B2(n326) );
    AN2T U407 ( .O(n325), .I1(A[47]), .I2(B[47]) );
    INV2 U408 ( .O(n323), .I(n322) );
    INV2 U409 ( .O(n365), .I(n170) );
    AN2T U410 ( .O(n364), .I1(A[34]), .I2(B[34]) );
    ND2T U411 ( .O(n328), .I1(B[0]), .I2(A[0]) );
    AN2T U412 ( .O(n254), .I1(A[2]), .I2(B[2]) );
    AN2T U413 ( .O(n263), .I1(A[54]), .I2(B[54]) );
    AN2T U414 ( .O(n258), .I1(A[50]), .I2(B[50]) );
    AN2T U415 ( .O(n265), .I1(A[56]), .I2(B[56]) );
    AN2T U416 ( .O(n268), .I1(A[58]), .I2(B[58]) );
    AN2T U417 ( .O(n248), .I1(A[43]), .I2(B[43]) );
    AN2T U418 ( .O(n250), .I1(A[27]), .I2(B[27]) );
    AN2T U419 ( .O(n252), .I1(A[39]), .I2(B[39]) );
    AN2T U420 ( .O(n260), .I1(A[19]), .I2(B[19]) );
    AN2T U421 ( .O(n256), .I1(A[23]), .I2(B[23]) );
    AO12T U422 ( .O(n480), .A1(n262), .B1(n603), .B2(n604) );
    AN2T U423 ( .O(n262), .I1(A[52]), .I2(B[52]) );
    AN2T U424 ( .O(n267), .I1(A[48]), .I2(B[48]) );
    AO12T U425 ( .O(n482), .A1(n267), .B1(n593), .B2(n594) );
    BUF2 U426 ( .O(n128), .I(A[53]) );
    BUF2 U427 ( .O(n129), .I(A[45]) );
    BUF2 U428 ( .O(n130), .I(A[55]) );
    BUF2 U429 ( .O(n131), .I(A[57]) );
    BUF2 U430 ( .O(n132), .I(A[3]) );
    BUF2 U431 ( .O(n133), .I(A[59]) );
    BUF2 U432 ( .O(n134), .I(A[1]) );
    BUF2 U433 ( .O(n135), .I(n444) );
    OA12P U434 ( .O(n138), .A1(n349), .B1(n605), .B2(n607) );
    OA12P U435 ( .O(n139), .A1(n353), .B1(n609), .B2(n611) );
    BUF4 U436 ( .O(n413), .I(n486) );
    ND2T U437 ( .O(n618), .I1(n330), .I2(n361) );
    INV2 U438 ( .O(n605), .I(n480) );
    INV2 U439 ( .O(n595), .I(n482) );
    INV2 U440 ( .O(n609), .I(n411) );
    BUF2 U441 ( .O(n411), .I(n479) );
    DELA U442 ( .O(n140), .I(n410) );
    INV2 U443 ( .O(n613), .I(n410) );
    BUF2 U444 ( .O(n410), .I(n478) );
    DELA U445 ( .O(n141), .I(n291) );
    OAI12 U446 ( .O(n590), .A1(n127), .B1(n441), .B2(n520) );
    DELA U447 ( .O(n142), .I(n383) );
    OA12P U448 ( .O(n151), .A1(n324), .B1(n383), .B2(n246) );
    BUF2 U449 ( .O(n247), .I(n142) );
    OA12P U450 ( .O(n383), .A1(n509), .B1(n505), .B2(n481) );
    DELA U451 ( .O(n143), .I(n552) );
    INV2 U452 ( .O(n289), .I(n288) );
    INV1 U453 ( .O(n443), .I(n143) );
    MOAI1T U454 ( .O(n473), .A1(n279), .A2(n144), .B1(A[62]), .B2(B[62]) );
    OAI12P U455 ( .O(n593), .A1(n81), .B1(n449), .B2(n547) );
    OA12T U456 ( .O(n148), .A1(n324), .B1(n247), .B2(n246) );
    BUF1 U457 ( .O(n149), .I(n619) );
    OA12P U458 ( .O(n150), .A1(n355), .B1(n595), .B2(n597) );
    OA12P U459 ( .O(n152), .A1(n357), .B1(n613), .B2(n615) );
    OAI12P U460 ( .O(n486), .A1(n255), .B1(n116), .B2(n557) );
    OAI12P U461 ( .O(n462), .A1(n316), .B1(n148), .B2(n589) );
    OR2P U462 ( .O(n556), .I1(B[2]), .I2(A[2]) );
    OR2P U463 ( .O(n616), .I1(B[58]), .I2(A[58]) );
    OR2P U464 ( .O(n604), .I1(B[52]), .I2(A[52]) );
    OR2P U465 ( .O(n598), .I1(B[50]), .I2(A[50]) );
    OR2P U466 ( .O(n608), .I1(B[54]), .I2(A[54]) );
    OR2P U467 ( .O(n594), .I1(B[48]), .I2(A[48]) );
    OR2P U468 ( .O(n612), .I1(B[56]), .I2(A[56]) );
    OR2P U469 ( .O(n553), .I1(B[7]), .I2(A[7]) );
    AN2T U470 ( .O(n153), .I1(A[35]), .I2(B[35]) );
    INV2 U471 ( .O(n154), .I(n153) );
    BUF2 U472 ( .O(n156), .I(n134) );
    XNR2 U473 ( .O(n475), .I1(A[60]), .I2(B[60]) );
    XNR2 U474 ( .O(n474), .I1(A[62]), .I2(B[62]) );
    OR2 U475 ( .O(n429), .I1(B[34]), .I2(A[34]) );
    OR2P U476 ( .O(n432), .I1(B[26]), .I2(A[26]) );
    OR2P U477 ( .O(n422), .I1(B[42]), .I2(A[42]) );
    OR2P U478 ( .O(n463), .I1(B[13]), .I2(A[13]) );
    OR2P U479 ( .O(n436), .I1(B[22]), .I2(A[22]) );
    OR2P U480 ( .O(n537), .I1(B[35]), .I2(A[35]) );
    INV2 U481 ( .O(n540), .I(n499) );
    OR2P U482 ( .O(n587), .I1(B[14]), .I2(A[14]) );
    OR2P U483 ( .O(n562), .I1(B[8]), .I2(A[8]) );
    INV3 U484 ( .O(n316), .I(n315) );
    AN2T U485 ( .O(n315), .I1(A[12]), .I2(B[12]) );
    BUF2 U486 ( .O(n160), .I(n508) );
    OR2 U487 ( .O(n508), .I1(B[5]), .I2(A[5]) );
    BUF2 U488 ( .O(n161), .I(n335) );
    AN2 U489 ( .O(n335), .I1(A[11]), .I2(B[11]) );
    BUF2 U490 ( .O(n162), .I(n337) );
    AN2 U491 ( .O(n337), .I1(A[7]), .I2(B[7]) );
    ND2P U492 ( .O(n447), .I1(n540), .I2(n541) );
    INV2 U493 ( .O(n397), .I(n396) );
    INV1 U494 ( .O(n347), .I(n346) );
    AN2T U495 ( .O(n168), .I1(n522), .I2(n523) );
    INV2 U496 ( .O(n169), .I(n168) );
    BUF3 U497 ( .O(n180), .I(n360) );
    AN2P U498 ( .O(n360), .I1(n133), .I2(B[59]) );
    BUF3 U499 ( .O(n181), .I(n358) );
    AN2P U500 ( .O(n358), .I1(n132), .I2(B[3]) );
    BUF3 U501 ( .O(n185), .I(n350) );
    AN2P U502 ( .O(n350), .I1(A[51]), .I2(B[51]) );
    OR2P U503 ( .O(n584), .I1(B[19]), .I2(A[19]) );
    INV3 U504 ( .O(n208), .I(n577) );
    OR2P U505 ( .O(n577), .I1(B[28]), .I2(A[28]) );
    INV3 U506 ( .O(n210), .I(n573) );
    OR2P U507 ( .O(n573), .I1(B[37]), .I2(A[37]) );
    INV3 U508 ( .O(n212), .I(n579) );
    OR2P U509 ( .O(n579), .I1(B[25]), .I2(A[25]) );
    INV3 U510 ( .O(n214), .I(n570) );
    OR2P U511 ( .O(n570), .I1(B[41]), .I2(A[41]) );
    INV3 U512 ( .O(n216), .I(n582) );
    OR2P U513 ( .O(n582), .I1(B[21]), .I2(A[21]) );
    INV3 U514 ( .O(n218), .I(n568) );
    OR2P U515 ( .O(n568), .I1(B[44]), .I2(A[44]) );
    INV3 U516 ( .O(n220), .I(n591) );
    OR2P U517 ( .O(n591), .I1(A[16]), .I2(B[16]) );
    BUF1 U518 ( .O(n224), .I(n493) );
    BUF2 U519 ( .O(n327), .I(n580) );
    BUF2 U520 ( .O(n326), .I(n571) );
    AN2P U521 ( .O(n243), .I1(n559), .I2(n359) );
    INV1 U522 ( .O(n244), .I(n243) );
    OR2P U523 ( .O(n623), .I1(n443), .I2(n495) );
    AN2T U524 ( .O(n245), .I1(n512), .I2(n513) );
    INV2 U525 ( .O(n246), .I(n245) );
    INV2 U526 ( .O(n249), .I(n248) );
    INV2 U527 ( .O(n251), .I(n250) );
    INV2 U528 ( .O(n253), .I(n252) );
    INV2 U529 ( .O(n255), .I(n254) );
    INV2 U530 ( .O(n257), .I(n256) );
    INV2 U531 ( .O(n259), .I(n258) );
    INV2 U532 ( .O(n261), .I(n260) );
    INV2 U533 ( .O(n264), .I(n263) );
    INV2 U534 ( .O(n266), .I(n265) );
    INV2 U535 ( .O(n269), .I(n268) );
    BUF2 U536 ( .O(n320), .I(n292) );
    OR2P U537 ( .O(n270), .I1(n346), .I2(n74) );
    AN2T U538 ( .O(n331), .I1(A[16]), .I2(B[16]) );
    AN2T U539 ( .O(n333), .I1(A[32]), .I2(B[32]) );
    ND2T U540 ( .O(n339), .I1(n156), .I2(n157) );
    OAI12 U541 ( .O(n431), .A1(n296), .B1(n531), .B2(n379) );
    OAI12 U542 ( .O(n435), .A1(n310), .B1(n528), .B2(n302) );
    OAI12 U543 ( .O(n425), .A1(n314), .B1(n542), .B2(n300) );
    INV3 U544 ( .O(n273), .I(n524) );
    INV3 U545 ( .O(n524), .I(n585) );
    OAI12 U546 ( .O(n421), .A1(n304), .B1(n545), .B2(n381) );
    DELA U547 ( .O(n275), .I(n290) );
    BUF2 U548 ( .O(n276), .I(n442) );
    INV1 U549 ( .O(n589), .I(n277) );
    OR2P U550 ( .O(n278), .I1(B[62]), .I2(A[62]) );
    INV2 U551 ( .O(n279), .I(n278) );
    OR2P U552 ( .O(n586), .I1(B[15]), .I2(A[15]) );
    BUF2 U553 ( .O(n285), .I(n141) );
    OR2P U554 ( .O(n288), .I1(B[61]), .I2(A[61]) );
    AN2T U555 ( .O(n291), .I1(n590), .I2(n341) );
    AN2T U556 ( .O(n295), .I1(B[25]), .I2(A[25]) );
    INV3 U557 ( .O(n296), .I(n295) );
    AN2T U558 ( .O(n297), .I1(A[17]), .I2(B[17]) );
    INV3 U559 ( .O(n298), .I(n297) );
    AN2T U560 ( .O(n299), .I1(A[36]), .I2(B[36]) );
    INV3 U561 ( .O(n300), .I(n299) );
    AN2T U562 ( .O(n301), .I1(A[20]), .I2(B[20]) );
    INV3 U563 ( .O(n302), .I(n301) );
    AN2T U564 ( .O(n303), .I1(B[41]), .I2(A[41]) );
    INV3 U565 ( .O(n304), .I(n303) );
    AN2T U566 ( .O(n309), .I1(A[21]), .I2(B[21]) );
    INV3 U567 ( .O(n310), .I(n309) );
    AN2T U568 ( .O(n313), .I1(A[37]), .I2(B[37]) );
    INV3 U569 ( .O(n314), .I(n313) );
    INV3 U570 ( .O(n318), .I(n440) );
    OR2P U571 ( .O(n440), .I1(B[18]), .I2(A[18]) );
    OR2P U572 ( .O(n535), .I1(B[31]), .I2(A[31]) );
    AN2T U573 ( .O(n322), .I1(A[33]), .I2(B[33]) );
    INV2 U574 ( .O(n576), .I(n536) );
    OR2P U575 ( .O(n571), .I1(B[40]), .I2(A[40]) );
    OR2P U576 ( .O(n580), .I1(B[24]), .I2(A[24]) );
    INV3 U577 ( .O(n332), .I(n331) );
    INV3 U578 ( .O(n408), .I(n407) );
    INV2 U579 ( .O(n336), .I(n161) );
    INV2 U580 ( .O(n338), .I(n162) );
    AN2T U581 ( .O(n340), .I1(A[15]), .I2(B[15]) );
    XNR2 U582 ( .O(n472), .I1(A[63]), .I2(B[63]) );
    AN2T U583 ( .O(n346), .I1(A[31]), .I2(B[31]) );
    INV4 U584 ( .O(n359), .I(n181) );
    BUF2 U585 ( .O(n362), .I(n328) );
    INV2 U586 ( .O(n433), .I(n369) );
    INV2 U587 ( .O(n437), .I(n371) );
    INV2 U588 ( .O(n426), .I(n373) );
    INV2 U589 ( .O(n423), .I(n377) );
    OR2P U590 ( .O(n620), .I1(n275), .I2(n499) );
    INV2 U591 ( .O(n567), .I(n550) );
    ND3T U592 ( .O(n547), .I1(n548), .I2(n382), .I3(n550) );
    INV3 U593 ( .O(n481), .I(n560) );
    INV3 U594 ( .O(n487), .I(n620) );
    INV3 U595 ( .O(n492), .I(n623) );
    AN2B1P U596 ( .O(n460), .I1(n397), .B1(n459) );
    XNR2 U597 ( .O(SUM[63]), .I1(n472), .I2(n473) );
    XOR2 U598 ( .O(SUM[62]), .I1(n474), .I2(n144) );
    OR2P U599 ( .O(n414), .I1(B[34]), .I2(A[34]) );
    ND3T U600 ( .O(n533), .I1(n534), .I2(n535), .I3(n536) );
    AN2T U601 ( .O(n396), .I1(A[18]), .I2(B[18]) );
    OR2P U602 ( .O(n455), .I1(B[33]), .I2(A[33]) );
    INV3 U603 ( .O(n541), .I(n501) );
    OAI12T U604 ( .O(n501), .A1(n253), .B1(n502), .B2(n424) );
    OAI12T U605 ( .O(n497), .A1(n257), .B1(n498), .B2(n434) );
    AN2T U606 ( .O(n405), .I1(A[30]), .I2(B[30]) );
    OAI12T U607 ( .O(n622), .A1(n308), .B1(n218), .B2(n119) );
    AN2T U608 ( .O(n407), .I1(A[5]), .I2(B[5]) );
    OAI12T U609 ( .O(n625), .A1(n294), .B1(n208), .B2(n122) );
    OAI12T U610 ( .O(n499), .A1(n154), .B1(n500), .B2(n427) );
    XNR2 U611 ( .O(SUM[17]), .I1(n224), .I2(n494) );
    XNR2 U612 ( .O(SUM[51]), .I1(n109), .I2(n409) );
    XNR2 U613 ( .O(SUM[59]), .I1(n88), .I2(n477) );
    OAI12P U614 ( .O(n477), .A1(n269), .B1(n152), .B2(n617) );
    OAI12P U615 ( .O(n476), .A1(n392), .B1(n481), .B2(n506) );
    XNR2 U616 ( .O(SUM[3]), .I1(n244), .I2(n413) );
    OAI12T U617 ( .O(n471), .A1(n388), .B1(n247), .B2(n515) );
    AOI12T U618 ( .O(n453), .A1(n322), .B1(n454), .B2(n402) );
    OAI12P U619 ( .O(n454), .A1(n334), .B1(n488), .B2(n592) );
    AOI12T U620 ( .O(n461), .A1(n171), .B1(n462), .B2(n415) );
    OAI12T U621 ( .O(n485), .A1(n541), .B1(n487), .B2(n77) );
    OAI12T U622 ( .O(n491), .A1(n526), .B1(n492), .B2(n71) );
    NR2T U623 ( .O(n441), .I1(n276), .I2(n151) );
    OR2T U624 ( .O(n552), .I1(n169), .I2(n291) );
    OR2T U625 ( .O(n554), .I1(B[6]), .I2(A[6]) );
    OR2T U626 ( .O(n555), .I1(n155), .I2(n134) );
    INV2 U627 ( .O(n557), .I(n556) );
    INV2 U628 ( .O(n563), .I(n471) );
    OR2T U629 ( .O(n548), .I1(B[46]), .I2(A[46]) );
    INV2 U630 ( .O(n566), .I(n548) );
    OR2T U631 ( .O(n550), .I1(B[45]), .I2(n129) );
    INV2 U632 ( .O(n500), .I(n537) );
    OR2T U633 ( .O(n534), .I1(B[30]), .I2(A[30]) );
    INV2 U634 ( .O(n575), .I(n534) );
    OR2T U635 ( .O(n536), .I1(B[29]), .I2(A[29]) );
    OR2T U636 ( .O(n585), .I1(B[17]), .I2(A[17]) );
    OR2T U637 ( .O(n466), .I1(B[10]), .I2(A[10]) );
    INV2 U638 ( .O(n599), .I(n598) );
    OR2T U639 ( .O(n601), .I1(B[51]), .I2(A[51]) );
    OR2T U640 ( .O(n610), .I1(B[55]), .I2(n130) );
    INV2 U641 ( .O(n617), .I(n616) );
    INV2 U642 ( .O(n621), .I(n485) );
    INV2 U643 ( .O(n484), .I(n622) );
    INV2 U644 ( .O(n624), .I(n491) );
    INV2 U645 ( .O(n490), .I(n625) );
    ND2 U646 ( .O(n493), .I1(n585), .I2(n298) );
endmodule


module adder ( clk, rst_n, a, b, s );
input  [63:0] a;
input  [63:0] b;
output [63:0] s;
input  clk, rst_n;
    wire n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
        n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
        n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
        n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
        n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
        n919, n920, n921, n922, \cnt[2] , \cnt[1] , \am[63] , \am[62] , 
        \am[61] , \am[60] , \am[59] , \am[58] , \am[57] , \am[56] , \am[55] , 
        \am[54] , \am[53] , \am[52] , \am[51] , \am[50] , \am[49] , \am[48] , 
        \am[47] , \am[46] , \am[45] , \am[44] , \am[43] , \am[42] , \am[41] , 
        \am[40] , \am[39] , \am[38] , \am[37] , \am[36] , \am[35] , \am[34] , 
        \am[33] , \am[32] , \am[31] , \am[30] , \am[29] , \am[28] , \am[27] , 
        \am[26] , \am[25] , \am[24] , \am[23] , \am[22] , \am[21] , \am[20] , 
        \am[19] , \am[18] , \am[17] , \am[16] , \am[15] , \am[14] , \am[13] , 
        \am[12] , \am[11] , \am[10] , \am[9] , \am[8] , \am[7] , \am[6] , 
        \am[5] , \am[4] , \am[3] , \am[2] , \am[1] , \am[0] , \bm[63] , 
        \bm[62] , \bm[61] , \bm[60] , \bm[59] , \bm[58] , \bm[57] , \bm[56] , 
        \bm[55] , \bm[54] , \bm[53] , \bm[52] , \bm[51] , \bm[50] , \bm[49] , 
        \bm[48] , \bm[47] , \bm[46] , \bm[45] , \bm[44] , \bm[43] , \bm[42] , 
        \bm[41] , \bm[40] , \bm[39] , \bm[38] , \bm[37] , \bm[36] , \bm[35] , 
        \bm[34] , \bm[33] , \bm[32] , \bm[31] , \bm[30] , \bm[29] , \bm[28] , 
        \bm[27] , \bm[26] , \bm[25] , \bm[24] , \bm[23] , \bm[22] , \bm[21] , 
        \bm[20] , \bm[19] , \bm[18] , \bm[17] , \bm[16] , \bm[15] , \bm[14] , 
        \bm[13] , \bm[12] , \bm[11] , \bm[10] , \bm[9] , \bm[8] , \bm[7] , 
        \bm[6] , \bm[5] , \bm[4] , \bm[3] , \bm[2] , \bm[1] , \bm[0] , N6, N7, 
        N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, 
        N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, 
        N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, 
        N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, 
        N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, 
        N746, N747, N748, N749, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
        n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
        n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
        n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
        n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
        n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
        n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
        n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
        n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
        n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
        n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
        n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
        n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
        n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
        n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
        n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
        n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
        n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
        n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
        n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
        n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
        n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
        n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
        n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
        n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
        n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
        n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
        n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
        n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
        n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
        n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
        n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
        n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
        n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
        n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
        n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
        n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
        n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
        n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
        n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
        n521, n522, n523, n524, n525, n526, n591, n592, n593, n594, n595, n596, 
        n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
        n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
        n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
        n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
        n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
        n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
        n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
        n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
        n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
        n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
        n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
        n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
        n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
        n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
        n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
        n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
        n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
        n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
        n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
        n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
        n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
        n849, n850, n851, n852, n853, n854, n855, n856, n858, n859;
    BUF2 U3 ( .O(n507), .I(\am[47] ) );
    BUF2 U5 ( .O(n526), .I(n517) );
    ND2P U6 ( .O(n859), .I1(n516), .I2(n526) );
    DFFRBN \bm_reg[20]  ( .Q(\bm[20] ), .QB(n398), .D(n838), .CK(clk), .RB(
        n711) );
    DFFRBN \am_reg[42]  ( .Q(\am[42] ), .QB(n9), .D(n7), .CK(clk), .RB(n701)
         );
    DFFRBP \am_reg[4]  ( .Q(\am[4] ), .D(n154), .CK(clk), .RB(n703) );
    DFFRBP \am_reg[9]  ( .Q(\am[9] ), .D(n169), .CK(clk), .RB(n676) );
    BUF3 U7 ( .O(n514), .I(\bm[47] ) );
    BUF3 U8 ( .O(n449), .I(\bm[35] ) );
    BUF3 U9 ( .O(n491), .I(\am[0] ) );
    BUF3 U10 ( .O(n497), .I(\am[26] ) );
    BUF3 U11 ( .O(n498), .I(\am[22] ) );
    BUF2 U12 ( .O(n499), .I(\am[38] ) );
    BUF3 U13 ( .O(n500), .I(\am[13] ) );
    BUF2 U14 ( .O(n501), .I(\am[42] ) );
    BUF2 U15 ( .O(n799), .I(n808) );
    DELA U16 ( .O(n378), .I(n405) );
    BUF3 U17 ( .O(n682), .I(n769) );
    BUF3 U18 ( .O(n704), .I(n741) );
    BUF3 U19 ( .O(n705), .I(n805) );
    BUF3 U20 ( .O(n716), .I(n753) );
    BUF3 U21 ( .O(n714), .I(n754) );
    BUF3 U22 ( .O(n673), .I(n774) );
    BUF3 U23 ( .O(n715), .I(n754) );
    BUF2 U24 ( .O(n754), .I(n800) );
    BUF3 U25 ( .O(n708), .I(n757) );
    BUF3 U26 ( .O(n720), .I(n751) );
    BUF3 U27 ( .O(n721), .I(n751) );
    BUF2 U28 ( .O(n751), .I(n801) );
    BUF3 U29 ( .O(n670), .I(n775) );
    BUF3 U30 ( .O(n685), .I(n768) );
    BUF3 U31 ( .O(n677), .I(n772) );
    BUF3 U32 ( .O(n695), .I(n763) );
    BUF3 U33 ( .O(n763), .I(n797) );
    BUF3 U34 ( .O(n684), .I(n768) );
    BUF2 U35 ( .O(n768), .I(n795) );
    BUF3 U36 ( .O(n661), .I(n780) );
    BUF3 U37 ( .O(n722), .I(n750) );
    BUF3 U38 ( .O(n669), .I(n776) );
    BUF3 U39 ( .O(n681), .I(n770) );
    BUF3 U40 ( .O(n712), .I(n755) );
    BUF3 U41 ( .O(n709), .I(n757) );
    BUF2 U42 ( .O(n757), .I(n799) );
    BUF3 U43 ( .O(n699), .I(n761) );
    BUF3 U44 ( .O(n665), .I(n778) );
    BUF3 U45 ( .O(n711), .I(n756) );
    BUF3 U46 ( .O(n730), .I(n746) );
    BUF3 U47 ( .O(n653), .I(n784) );
    BUF3 U48 ( .O(n654), .I(n783) );
    BUF3 U49 ( .O(n731), .I(n746) );
    BUF2 U50 ( .O(n746), .I(n803) );
    BUF3 U51 ( .O(n652), .I(n784) );
    BUF2 U52 ( .O(n784), .I(n790) );
    BUF3 U53 ( .O(n728), .I(n747) );
    BUF3 U54 ( .O(n732), .I(n745) );
    BUF3 U55 ( .O(n656), .I(n782) );
    BUF3 U56 ( .O(n727), .I(n748) );
    BUF3 U57 ( .O(n733), .I(n745) );
    BUF2 U58 ( .O(n745), .I(n803) );
    BUF3 U59 ( .O(n803), .I(n806) );
    BUF3 U60 ( .O(n650), .I(n785) );
    BUF3 U61 ( .O(n726), .I(n748) );
    BUF2 U62 ( .O(n748), .I(n802) );
    BUF3 U63 ( .O(n655), .I(n783) );
    BUF2 U64 ( .O(n783), .I(n790) );
    BUF3 U65 ( .O(n790), .I(n812) );
    BUF3 U66 ( .O(n725), .I(n749) );
    BUF3 U67 ( .O(n734), .I(n744) );
    BUF3 U68 ( .O(n658), .I(n781) );
    BUF3 U69 ( .O(n649), .I(n786) );
    BUF3 U70 ( .O(n659), .I(n781) );
    BUF2 U71 ( .O(n781), .I(n791) );
    BUF3 U72 ( .O(n667), .I(n777) );
    BUF3 U73 ( .O(n648), .I(n786) );
    BUF2 U74 ( .O(n786), .I(n789) );
    BUF3 U75 ( .O(n736), .I(n743) );
    BUF3 U76 ( .O(n739), .I(n742) );
    BUF3 U77 ( .O(n647), .I(n787) );
    BUF3 U78 ( .O(n646), .I(n787) );
    BUF2 U79 ( .O(n787), .I(n789) );
    BUF3 U80 ( .O(n789), .I(n809) );
    BUF3 U81 ( .O(n737), .I(n743) );
    BUF2 U82 ( .O(n743), .I(n804) );
    BUF3 U83 ( .O(n735), .I(n744) );
    BUF2 U84 ( .O(n744), .I(n804) );
    BUF3 U85 ( .O(n804), .I(n805) );
    BUF3 U86 ( .O(n651), .I(n785) );
    BUF2 U87 ( .O(n785), .I(n790) );
    BUF3 U88 ( .O(n645), .I(n788) );
    BUF3 U89 ( .O(n729), .I(n747) );
    BUF2 U90 ( .O(n747), .I(n803) );
    BUF3 U91 ( .O(n738), .I(n742) );
    BUF2 U92 ( .O(n742), .I(n804) );
    BUF3 U93 ( .O(n657), .I(n782) );
    BUF2 U94 ( .O(n782), .I(n791) );
    BUF3 U95 ( .O(n791), .I(n812) );
    BUF3 U96 ( .O(n724), .I(n749) );
    BUF2 U97 ( .O(n749), .I(n802) );
    BUF3 U98 ( .O(n802), .I(n806) );
    BUF3 U99 ( .O(n686), .I(n767) );
    BUF3 U100 ( .O(n740), .I(n741) );
    BUF3 U101 ( .O(n680), .I(n770) );
    BUF2 U102 ( .O(n770), .I(n795) );
    BUF3 U103 ( .O(n795), .I(n810) );
    BUF3 U104 ( .O(n702), .I(n759) );
    BUF3 U105 ( .O(n679), .I(n771) );
    BUF3 U106 ( .O(n703), .I(n759) );
    BUF2 U107 ( .O(n759), .I(n798) );
    BUF3 U108 ( .O(n707), .I(n758) );
    BUF3 U109 ( .O(n692), .I(n764) );
    BUF3 U110 ( .O(n700), .I(n760) );
    BUF3 U111 ( .O(n694), .I(n763) );
    BUF3 U112 ( .O(n666), .I(n777) );
    BUF2 U113 ( .O(n777), .I(n792) );
    BUF3 U114 ( .O(n672), .I(n774) );
    BUF2 U115 ( .O(n774), .I(n793) );
    BUF3 U116 ( .O(n710), .I(n756) );
    BUF2 U117 ( .O(n756), .I(n800) );
    BUF3 U118 ( .O(n800), .I(n807) );
    BUF3 U119 ( .O(n664), .I(n778) );
    BUF2 U120 ( .O(n778), .I(n792) );
    BUF3 U121 ( .O(n792), .I(n811) );
    BUF3 U122 ( .O(n663), .I(n779) );
    BUF3 U123 ( .O(n718), .I(n752) );
    BUF3 U124 ( .O(n662), .I(n779) );
    BUF2 U125 ( .O(n779), .I(n792) );
    BUF3 U126 ( .O(n690), .I(n765) );
    BUF3 U127 ( .O(n693), .I(n764) );
    BUF2 U128 ( .O(n764), .I(n797) );
    BUF3 U129 ( .O(n797), .I(n809) );
    BUF3 U130 ( .O(n689), .I(n766) );
    BUF3 U131 ( .O(n698), .I(n761) );
    BUF2 U132 ( .O(n761), .I(n798) );
    BUF3 U133 ( .O(n798), .I(n808) );
    BUF3 U134 ( .O(n696), .I(n762) );
    BUF3 U135 ( .O(n678), .I(n771) );
    BUF2 U136 ( .O(n771), .I(n794) );
    BUF3 U137 ( .O(n676), .I(n772) );
    BUF2 U138 ( .O(n772), .I(n794) );
    BUF3 U139 ( .O(n794), .I(n810) );
    BUF3 U140 ( .O(n706), .I(n758) );
    BUF2 U141 ( .O(n758), .I(n799) );
    DFFRBP \am_reg[62]  ( .Q(\am[62] ), .D(n348), .CK(clk), .RB(n706) );
    BUF3 U142 ( .O(n723), .I(n750) );
    BUF2 U143 ( .O(n750), .I(n802) );
    BUF2 U144 ( .O(n806), .I(n815) );
    BUF3 U145 ( .O(n660), .I(n780) );
    BUF2 U146 ( .O(n780), .I(n791) );
    BUF2 U147 ( .O(n812), .I(n813) );
    BUF3 U148 ( .O(n719), .I(n752) );
    BUF2 U149 ( .O(n752), .I(n801) );
    BUF3 U150 ( .O(n801), .I(n807) );
    BUF3 U151 ( .O(n688), .I(n766) );
    BUF2 U152 ( .O(n766), .I(n796) );
    BUF3 U153 ( .O(n674), .I(n773) );
    BUF3 U154 ( .O(n691), .I(n765) );
    BUF2 U155 ( .O(n765), .I(n796) );
    BUF3 U156 ( .O(n796), .I(n809) );
    BUF3 U157 ( .O(n675), .I(n773) );
    BUF2 U158 ( .O(n773), .I(n794) );
    BUF2 U159 ( .O(n760), .I(n798) );
    BUF2 U160 ( .O(n808), .I(n814) );
    BUF3 U161 ( .O(n814), .I(n816) );
    BUF3 U162 ( .O(n717), .I(n753) );
    BUF2 U163 ( .O(n753), .I(n801) );
    BUF3 U164 ( .O(n697), .I(n762) );
    BUF2 U165 ( .O(n762), .I(n797) );
    BUF3 U166 ( .O(n713), .I(n755) );
    BUF2 U167 ( .O(n755), .I(n800) );
    BUF2 U168 ( .O(n807), .I(n815) );
    BUF3 U169 ( .O(n815), .I(n816) );
    BUF3 U170 ( .O(n687), .I(n767) );
    BUF2 U171 ( .O(n767), .I(n796) );
    BUF3 U172 ( .O(n671), .I(n775) );
    BUF2 U173 ( .O(n775), .I(n793) );
    BUF3 U174 ( .O(n793), .I(n811) );
    BUF3 U175 ( .O(n683), .I(n769) );
    BUF2 U176 ( .O(n769), .I(n795) );
    BUF2 U177 ( .O(n810), .I(n814) );
    BUF3 U178 ( .O(n668), .I(n776) );
    BUF2 U179 ( .O(n776), .I(n793) );
    BUF2 U180 ( .O(n811), .I(n813) );
    XOR2P U181 ( .O(N6), .I1(n516), .I2(n517) );
    BUF3 U182 ( .O(n644), .I(n788) );
    BUF2 U183 ( .O(n788), .I(n789) );
    BUF2 U184 ( .O(n816), .I(rst_n) );
    BUF2 U185 ( .O(n474), .I(\bm[30] ) );
    BUF2 U186 ( .O(n475), .I(\bm[32] ) );
    BUF2 U187 ( .O(n476), .I(\bm[20] ) );
    BUF2 U188 ( .O(n477), .I(\bm[36] ) );
    BUF2 U189 ( .O(n478), .I(\bm[17] ) );
    BUF3 U190 ( .O(n512), .I(\am[35] ) );
    BUF2 U191 ( .O(n805), .I(n815) );
    BUF2 U192 ( .O(n813), .I(rst_n) );
    BUF4 U193 ( .O(n809), .I(n814) );
    BUF2 U194 ( .O(n741), .I(n701) );
    BUF4 U195 ( .O(n448), .I(\bm[0] ) );
    MXL2P U196 ( .OB(n7), .S(n600), .A(n9), .B(n8) );
    INV2 U197 ( .O(n8), .I(a[42]) );
    MXL2P U198 ( .OB(n10), .S(n600), .A(n12), .B(n11) );
    INV2 U199 ( .O(n11), .I(a[43]) );
    DFFRBP \am_reg[43]  ( .Q(\am[43] ), .QB(n12), .D(n10), .CK(clk), .RB(n682)
         );
    MXL2P U200 ( .OB(n13), .S(n623), .A(n419), .B(N749) );
    INV2 U201 ( .O(n14), .I(n13) );
    MXL2P U202 ( .OB(n15), .S(n626), .A(n905), .B(N703) );
    INV2 U203 ( .O(n16), .I(n15) );
    MXL2P U204 ( .OB(n17), .S(n628), .A(n861), .B(N747) );
    INV2 U205 ( .O(n18), .I(n17) );
    MXL2P U206 ( .OB(n19), .S(n620), .A(n898), .B(N710) );
    INV2 U207 ( .O(n20), .I(n19) );
    MXL2P U208 ( .OB(n21), .S(n599), .A(n882), .B(N726) );
    INV2 U209 ( .O(n22), .I(n21) );
    MXL2P U210 ( .OB(n23), .S(n616), .A(n875), .B(N733) );
    INV2 U211 ( .O(n24), .I(n23) );
    MXL2P U212 ( .OB(n25), .S(n623), .A(n873), .B(N735) );
    INV2 U213 ( .O(n26), .I(n25) );
    MXL2P U214 ( .OB(n27), .S(n831), .A(n889), .B(N719) );
    INV2 U215 ( .O(n28), .I(n27) );
    MXL2P U216 ( .OB(n29), .S(n620), .A(n871), .B(N737) );
    INV2 U217 ( .O(n30), .I(n29) );
    MXL2P U218 ( .OB(n31), .S(n628), .A(n891), .B(N717) );
    INV2 U219 ( .O(n32), .I(n31) );
    MXL2P U220 ( .OB(n33), .S(n620), .A(n869), .B(N739) );
    INV2 U221 ( .O(n34), .I(n33) );
    MXL2P U222 ( .OB(n35), .S(n627), .A(n909), .B(N699) );
    INV2 U223 ( .O(n36), .I(n35) );
    MXL2P U224 ( .OB(n37), .S(n828), .A(n867), .B(N741) );
    INV2 U225 ( .O(n38), .I(n37) );
    MXL2P U226 ( .OB(n39), .S(n829), .A(n913), .B(N695) );
    INV2 U227 ( .O(n40), .I(n39) );
    MXL2P U228 ( .OB(n41), .S(n395), .A(n865), .B(N743) );
    INV2 U229 ( .O(n42), .I(n41) );
    MXL2P U230 ( .OB(n43), .S(n828), .A(n917), .B(N691) );
    INV2 U231 ( .O(n44), .I(n43) );
    MXL2P U232 ( .OB(n45), .S(n616), .A(n863), .B(N745) );
    INV2 U233 ( .O(n46), .I(n45) );
    MXL2P U234 ( .OB(n47), .S(n625), .A(n919), .B(N689) );
    INV2 U235 ( .O(n48), .I(n47) );
    MXL2P U236 ( .OB(n49), .S(n626), .A(n862), .B(N746) );
    INV2 U237 ( .O(n50), .I(n49) );
    MXL2P U238 ( .OB(n51), .S(n623), .A(n860), .B(N748) );
    INV2 U239 ( .O(n52), .I(n51) );
    MXL2P U240 ( .OB(n53), .S(n819), .A(n921), .B(N687) );
    INV2 U241 ( .O(n54), .I(n53) );
    MXL2P U242 ( .OB(n55), .S(n643), .A(n897), .B(N711) );
    INV2 U243 ( .O(n56), .I(n55) );
    MXL2P U244 ( .OB(n57), .S(n643), .A(n894), .B(N714) );
    INV2 U245 ( .O(n58), .I(n57) );
    MXL2P U246 ( .OB(n59), .S(n617), .A(n901), .B(N707) );
    INV2 U247 ( .O(n60), .I(n59) );
    MXL2P U248 ( .OB(n61), .S(n624), .A(n885), .B(N723) );
    INV2 U249 ( .O(n62), .I(n61) );
    MXL2P U250 ( .OB(n63), .S(n617), .A(n906), .B(N702) );
    INV2 U251 ( .O(n64), .I(n63) );
    MXL2P U252 ( .OB(n65), .S(n621), .A(n881), .B(N727) );
    INV2 U253 ( .O(n66), .I(n65) );
    MXL2P U254 ( .OB(n67), .S(n626), .A(n907), .B(N701) );
    INV2 U255 ( .O(n68), .I(n67) );
    MXL2P U256 ( .OB(n69), .S(n618), .A(n878), .B(N730) );
    INV2 U257 ( .O(n70), .I(n69) );
    MXL2P U258 ( .OB(n71), .S(n623), .A(n888), .B(N720) );
    INV2 U259 ( .O(n72), .I(n71) );
    MXL2P U260 ( .OB(n73), .S(n829), .A(n884), .B(N724) );
    INV2 U261 ( .O(n74), .I(n73) );
    MXL2P U262 ( .OB(n75), .S(n828), .A(n896), .B(N712) );
    INV2 U263 ( .O(n76), .I(n75) );
    MXL2P U264 ( .OB(n77), .S(n627), .A(n880), .B(N728) );
    INV2 U265 ( .O(n78), .I(n77) );
    MXL2P U266 ( .OB(n79), .S(n386), .A(n900), .B(N708) );
    INV2 U267 ( .O(n80), .I(n79) );
    MXL2P U268 ( .OB(n81), .S(n624), .A(n895), .B(N713) );
    INV2 U269 ( .O(n82), .I(n81) );
    MXL2P U270 ( .OB(n83), .S(n628), .A(n899), .B(N709) );
    INV2 U271 ( .O(n84), .I(n83) );
    MXL2P U272 ( .OB(n85), .S(n496), .A(n893), .B(N715) );
    INV2 U273 ( .O(n86), .I(n85) );
    MXL2P U274 ( .OB(n87), .S(n617), .A(n902), .B(N706) );
    INV2 U275 ( .O(n88), .I(n87) );
    MXL2P U276 ( .OB(n89), .S(n616), .A(n892), .B(N716) );
    INV2 U277 ( .O(n90), .I(n89) );
    MXL2P U278 ( .OB(n91), .S(n831), .A(n903), .B(N705) );
    INV2 U279 ( .O(n92), .I(n91) );
    MXL2P U280 ( .OB(n93), .S(n618), .A(n890), .B(N718) );
    INV2 U281 ( .O(n94), .I(n93) );
    MXL2P U282 ( .OB(n95), .S(n627), .A(n904), .B(N704) );
    INV2 U283 ( .O(n96), .I(n95) );
    MXL2P U284 ( .OB(n97), .S(n606), .A(n887), .B(N721) );
    INV2 U285 ( .O(n98), .I(n97) );
    MXL2P U286 ( .OB(n99), .S(n606), .A(n908), .B(N700) );
    INV2 U287 ( .O(n100), .I(n99) );
    MXL2P U288 ( .OB(n101), .S(n395), .A(n886), .B(N722) );
    INV2 U289 ( .O(n102), .I(n101) );
    MXL2P U290 ( .OB(n103), .S(n828), .A(n910), .B(N698) );
    INV2 U291 ( .O(n104), .I(n103) );
    MXL2P U292 ( .OB(n105), .S(n614), .A(n883), .B(N725) );
    INV2 U293 ( .O(n106), .I(n105) );
    MXL2P U294 ( .OB(n107), .S(n614), .A(n911), .B(N697) );
    INV2 U295 ( .O(n108), .I(n107) );
    MXL2P U296 ( .OB(n109), .S(n621), .A(n879), .B(N729) );
    INV2 U297 ( .O(n110), .I(n109) );
    MXL2P U298 ( .OB(n111), .S(n625), .A(n912), .B(N696) );
    INV2 U299 ( .O(n112), .I(n111) );
    MXL2P U300 ( .OB(n113), .S(n624), .A(n877), .B(N731) );
    INV2 U301 ( .O(n114), .I(n113) );
    MXL2P U302 ( .OB(n115), .S(n606), .A(n914), .B(N694) );
    INV2 U303 ( .O(n116), .I(n115) );
    MXL2P U304 ( .OB(n117), .S(n624), .A(n876), .B(N732) );
    INV2 U305 ( .O(n118), .I(n117) );
    MXL2P U306 ( .OB(n119), .S(n626), .A(n915), .B(N693) );
    INV2 U307 ( .O(n120), .I(n119) );
    MXL2P U308 ( .OB(n121), .S(n627), .A(n872), .B(N736) );
    INV2 U309 ( .O(n122), .I(n121) );
    MXL2P U310 ( .OB(n123), .S(n827), .A(n916), .B(N692) );
    INV2 U311 ( .O(n124), .I(n123) );
    MXL2P U312 ( .OB(n125), .S(n395), .A(n868), .B(N740) );
    INV2 U313 ( .O(n126), .I(n125) );
    MXL2P U314 ( .OB(n127), .S(n600), .A(n918), .B(N690) );
    INV2 U315 ( .O(n128), .I(n127) );
    MXL2P U316 ( .OB(n129), .S(n614), .A(n866), .B(N742) );
    INV2 U317 ( .O(n130), .I(n129) );
    MXL2P U318 ( .OB(n131), .S(n625), .A(n920), .B(N688) );
    INV2 U319 ( .O(n132), .I(n131) );
    MXL2P U320 ( .OB(n133), .S(n628), .A(n864), .B(N744) );
    INV2 U321 ( .O(n134), .I(n133) );
    MXL2P U322 ( .OB(n135), .S(n621), .A(n874), .B(N734) );
    INV2 U323 ( .O(n136), .I(n135) );
    MXL2P U324 ( .OB(n137), .S(n625), .A(n870), .B(N738) );
    INV2 U325 ( .O(n138), .I(n137) );
    MXL2P U326 ( .OB(n139), .S(n819), .A(n922), .B(N686) );
    INV2 U327 ( .O(n140), .I(n139) );
    MXL2P U328 ( .OB(n141), .S(n829), .A(\am[1] ), .B(a[1]) );
    INV2 U329 ( .O(n142), .I(n141) );
    MXL2P U330 ( .OB(n143), .S(n609), .A(\am[0] ), .B(a[0]) );
    INV2 U331 ( .O(n144), .I(n143) );
    MXL2P U332 ( .OB(n145), .S(n413), .A(\am[2] ), .B(a[2]) );
    INV2 U333 ( .O(n146), .I(n145) );
    MXL2P U334 ( .OB(n147), .S(n819), .A(\bm[63] ), .B(b[63]) );
    INV2 U335 ( .O(n148), .I(n147) );
    MXL2P U336 ( .OB(n149), .S(n594), .A(\am[3] ), .B(a[3]) );
    INV2 U337 ( .O(n150), .I(n149) );
    MXL2P U338 ( .OB(n151), .S(n608), .A(\bm[62] ), .B(b[62]) );
    INV2 U339 ( .O(n152), .I(n151) );
    MXL2P U340 ( .OB(n153), .S(n608), .A(\am[4] ), .B(a[4]) );
    INV2 U341 ( .O(n154), .I(n153) );
    MXL2P U342 ( .OB(n155), .S(n610), .A(\bm[61] ), .B(b[61]) );
    INV2 U343 ( .O(n156), .I(n155) );
    MXL2P U344 ( .OB(n157), .S(n826), .A(\am[5] ), .B(a[5]) );
    INV2 U345 ( .O(n158), .I(n157) );
    MXL2P U346 ( .OB(n159), .S(n619), .A(\bm[60] ), .B(b[60]) );
    INV2 U347 ( .O(n160), .I(n159) );
    BUF2 U348 ( .O(n161), .I(n847) );
    MXL2P U349 ( .OB(n162), .S(n593), .A(\bm[59] ), .B(b[59]) );
    INV2 U350 ( .O(n163), .I(n162) );
    MXL2P U351 ( .OB(n164), .S(n612), .A(\am[8] ), .B(a[8]) );
    INV2 U352 ( .O(n165), .I(n164) );
    MXL2P U353 ( .OB(n166), .S(n604), .A(\bm[58] ), .B(b[58]) );
    INV2 U354 ( .O(n167), .I(n166) );
    MXL2P U355 ( .OB(n168), .S(n619), .A(\am[9] ), .B(a[9]) );
    INV2 U356 ( .O(n169), .I(n168) );
    BUF1 U357 ( .O(n170), .I(n846) );
    MUX2 U358 ( .O(n846), .S(n823), .A(\bm[57] ), .B(b[57]) );
    MXL2P U359 ( .OB(n171), .S(n826), .A(\am[10] ), .B(a[10]) );
    INV2 U360 ( .O(n172), .I(n171) );
    MXL2P U361 ( .OB(n173), .S(n610), .A(\bm[55] ), .B(b[55]) );
    INV2 U362 ( .O(n174), .I(n173) );
    BUF2 U363 ( .O(n175), .I(n849) );
    MXL2P U364 ( .OB(n176), .S(n821), .A(\bm[54] ), .B(b[54]) );
    INV2 U365 ( .O(n177), .I(n176) );
    MXL2P U366 ( .OB(n178), .S(n827), .A(\am[12] ), .B(a[12]) );
    INV2 U367 ( .O(n179), .I(n178) );
    MXL2P U368 ( .OB(n180), .S(n638), .A(\bm[53] ), .B(b[53]) );
    INV2 U369 ( .O(n181), .I(n180) );
    MXL2P U370 ( .OB(n182), .S(n593), .A(n500), .B(a[13]) );
    INV2 U371 ( .O(n183), .I(n182) );
    MXL2P U372 ( .OB(n184), .S(n603), .A(\bm[52] ), .B(b[52]) );
    INV2 U373 ( .O(n185), .I(n184) );
    MXL2P U374 ( .OB(n186), .S(n609), .A(\am[14] ), .B(a[14]) );
    INV2 U375 ( .O(n187), .I(n186) );
    MXL2P U376 ( .OB(n188), .S(n358), .A(\bm[51] ), .B(b[51]) );
    INV2 U377 ( .O(n189), .I(n188) );
    MXL2P U378 ( .OB(n190), .S(n640), .A(\am[15] ), .B(a[15]) );
    INV2 U379 ( .O(n191), .I(n190) );
    MXL2P U380 ( .OB(n192), .S(n835), .A(\bm[50] ), .B(b[50]) );
    INV2 U381 ( .O(n193), .I(n192) );
    MXL2P U382 ( .OB(n194), .S(n640), .A(\am[16] ), .B(a[16]) );
    INV2 U383 ( .O(n195), .I(n194) );
    MXL2P U384 ( .OB(n196), .S(n594), .A(\bm[49] ), .B(b[49]) );
    INV2 U385 ( .O(n197), .I(n196) );
    MXL2P U386 ( .OB(n198), .S(n610), .A(n459), .B(a[17]) );
    INV2 U387 ( .O(n199), .I(n198) );
    MXL2P U388 ( .OB(n200), .S(n615), .A(\bm[48] ), .B(b[48]) );
    INV2 U389 ( .O(n201), .I(n200) );
    MXL2P U390 ( .OB(n202), .S(n622), .A(\am[18] ), .B(a[18]) );
    INV2 U391 ( .O(n203), .I(n202) );
    MXL2P U392 ( .OB(n204), .S(n383), .A(\bm[47] ), .B(b[47]) );
    INV2 U393 ( .O(n205), .I(n204) );
    MXL2P U394 ( .OB(n206), .S(n593), .A(\am[19] ), .B(a[19]) );
    INV2 U395 ( .O(n207), .I(n206) );
    MXL2P U396 ( .OB(n208), .S(n827), .A(\bm[46] ), .B(b[46]) );
    INV2 U397 ( .O(n209), .I(n208) );
    MXL2P U398 ( .OB(n210), .S(n639), .A(n455), .B(a[20]) );
    INV2 U399 ( .O(n211), .I(n210) );
    MXL2P U400 ( .OB(n212), .S(n643), .A(\bm[44] ), .B(b[44]) );
    INV2 U401 ( .O(n213), .I(n212) );
    MXL2P U402 ( .OB(n214), .S(n643), .A(\am[21] ), .B(a[21]) );
    INV2 U403 ( .O(n215), .I(n214) );
    MXL2P U404 ( .OB(n216), .S(n642), .A(\bm[43] ), .B(b[43]) );
    INV2 U405 ( .O(n217), .I(n216) );
    MXL2P U406 ( .OB(n218), .S(n608), .A(n498), .B(a[22]) );
    INV2 U407 ( .O(n219), .I(n218) );
    MXL2P U408 ( .OB(n220), .S(n619), .A(n510), .B(b[42]) );
    INV2 U409 ( .O(n221), .I(n220) );
    MXL2P U410 ( .OB(n222), .S(n622), .A(\am[23] ), .B(a[23]) );
    INV2 U411 ( .O(n223), .I(n222) );
    MXL2P U412 ( .OB(n224), .S(n822), .A(\bm[41] ), .B(b[41]) );
    INV2 U413 ( .O(n225), .I(n224) );
    MXL2P U414 ( .OB(n226), .S(n822), .A(\am[24] ), .B(a[24]) );
    INV2 U415 ( .O(n227), .I(n226) );
    MXL2P U416 ( .OB(n228), .S(n618), .A(n513), .B(b[38]) );
    INV2 U417 ( .O(n229), .I(n228) );
    MXL2P U418 ( .OB(n230), .S(n619), .A(\am[25] ), .B(a[25]) );
    INV2 U419 ( .O(n231), .I(n230) );
    MXL2P U420 ( .OB(n232), .S(n599), .A(n437), .B(b[37]) );
    INV2 U421 ( .O(n233), .I(n232) );
    MXL2P U422 ( .OB(n234), .S(n383), .A(n497), .B(a[26]) );
    INV2 U423 ( .O(n235), .I(n234) );
    MXL2P U424 ( .OB(n236), .S(n620), .A(\bm[36] ), .B(b[36]) );
    INV2 U425 ( .O(n237), .I(n236) );
    MXL2P U426 ( .OB(n238), .S(n618), .A(\am[27] ), .B(a[27]) );
    INV2 U427 ( .O(n239), .I(n238) );
    MXL2P U428 ( .OB(n240), .S(n641), .A(\bm[35] ), .B(b[35]) );
    INV2 U429 ( .O(n241), .I(n240) );
    MXL2P U430 ( .OB(n242), .S(n612), .A(\am[28] ), .B(a[28]) );
    INV2 U431 ( .O(n243), .I(n242) );
    MXL2P U432 ( .OB(n244), .S(n603), .A(\bm[34] ), .B(b[34]) );
    INV2 U433 ( .O(n245), .I(n244) );
    MXL2P U434 ( .OB(n246), .S(n377), .A(n592), .B(a[30]) );
    INV2 U435 ( .O(n247), .I(n246) );
    MXL2P U436 ( .OB(n248), .S(n594), .A(n439), .B(b[33]) );
    INV2 U437 ( .O(n249), .I(n248) );
    MXL2P U438 ( .OB(n250), .S(n594), .A(\am[31] ), .B(a[31]) );
    INV2 U439 ( .O(n251), .I(n250) );
    MXL2P U440 ( .OB(n252), .S(n406), .A(\bm[32] ), .B(b[32]) );
    INV2 U441 ( .O(n253), .I(n252) );
    BUF2 U442 ( .O(n254), .I(n851) );
    MXL2P U443 ( .OB(n255), .S(n613), .A(n441), .B(b[31]) );
    INV2 U444 ( .O(n256), .I(n255) );
    MXL2P U445 ( .OB(n257), .S(n394), .A(\am[34] ), .B(a[34]) );
    INV2 U446 ( .O(n258), .I(n257) );
    MXL2P U447 ( .OB(n259), .S(n603), .A(\bm[30] ), .B(b[30]) );
    INV2 U448 ( .O(n260), .I(n259) );
    MXL2P U449 ( .OB(n261), .S(n642), .A(\am[35] ), .B(a[35]) );
    INV2 U450 ( .O(n262), .I(n261) );
    MXL2P U451 ( .OB(n263), .S(n599), .A(\bm[28] ), .B(b[28]) );
    INV2 U452 ( .O(n264), .I(n263) );
    MXL2P U453 ( .OB(n265), .S(n641), .A(n461), .B(a[36]) );
    INV2 U454 ( .O(n266), .I(n265) );
    MXL2P U455 ( .OB(n267), .S(n394), .A(\bm[27] ), .B(b[27]) );
    INV2 U456 ( .O(n268), .I(n267) );
    MXL2P U457 ( .OB(n269), .S(n425), .A(\am[38] ), .B(a[38]) );
    INV2 U458 ( .O(n270), .I(n269) );
    MXL2P U459 ( .OB(n271), .S(n610), .A(n509), .B(b[26]) );
    INV2 U460 ( .O(n272), .I(n271) );
    MXL2P U461 ( .OB(n273), .S(n603), .A(\am[39] ), .B(a[39]) );
    INV2 U462 ( .O(n274), .I(n273) );
    MXL2P U463 ( .OB(n275), .S(n508), .A(\bm[25] ), .B(b[25]) );
    INV2 U464 ( .O(n276), .I(n275) );
    MXL2P U465 ( .OB(n277), .S(n826), .A(\am[41] ), .B(a[41]) );
    INV2 U466 ( .O(n278), .I(n277) );
    BUF1 U467 ( .O(n279), .I(n839) );
    MUX2 U468 ( .O(n839), .S(n824), .A(\bm[23] ), .B(b[23]) );
    MXL2P U469 ( .OB(n280), .S(n827), .A(n515), .B(b[22]) );
    INV2 U470 ( .O(n281), .I(n280) );
    MXL2P U471 ( .OB(n282), .S(n641), .A(n447), .B(b[21]) );
    INV2 U472 ( .O(n283), .I(n282) );
    MXL2P U473 ( .OB(n284), .S(n607), .A(\am[45] ), .B(a[45]) );
    INV2 U474 ( .O(n285), .I(n284) );
    MXL2P U475 ( .OB(n286), .S(n604), .A(\bm[19] ), .B(b[19]) );
    INV2 U476 ( .O(n287), .I(n286) );
    MXL2P U477 ( .OB(n288), .S(n641), .A(n428), .B(a[46]) );
    INV2 U478 ( .O(n289), .I(n288) );
    MXL2P U479 ( .OB(n290), .S(n386), .A(n443), .B(b[18]) );
    INV2 U480 ( .O(n291), .I(n290) );
    MXL2P U481 ( .OB(n292), .S(n615), .A(\am[47] ), .B(a[47]) );
    INV2 U482 ( .O(n293), .I(n292) );
    MXL2P U483 ( .OB(n294), .S(n604), .A(\bm[17] ), .B(b[17]) );
    INV2 U484 ( .O(n295), .I(n294) );
    BUF1 U485 ( .O(n296), .I(n855) );
    MUX2 U486 ( .O(n855), .S(n821), .A(\am[48] ), .B(a[48]) );
    MXL2P U487 ( .OB(n297), .S(n609), .A(\bm[16] ), .B(b[16]) );
    INV2 U488 ( .O(n298), .I(n297) );
    MXL2P U489 ( .OB(n299), .S(n599), .A(n430), .B(a[49]) );
    INV2 U490 ( .O(n300), .I(n299) );
    MXL2P U491 ( .OB(n301), .S(n593), .A(n445), .B(b[15]) );
    INV2 U492 ( .O(n302), .I(n301) );
    MXL2P U493 ( .OB(n303), .S(n612), .A(n432), .B(a[51]) );
    INV2 U494 ( .O(n304), .I(n303) );
    MXL2P U495 ( .OB(n305), .S(n413), .A(\bm[14] ), .B(b[14]) );
    INV2 U496 ( .O(n306), .I(n305) );
    MXL2P U497 ( .OB(n307), .S(n608), .A(\am[52] ), .B(a[52]) );
    INV2 U498 ( .O(n308), .I(n307) );
    MXL2P U499 ( .OB(n309), .S(n642), .A(n511), .B(b[13]) );
    INV2 U500 ( .O(n310), .I(n309) );
    MXL2P U501 ( .OB(n311), .S(n824), .A(\am[53] ), .B(a[53]) );
    INV2 U502 ( .O(n312), .I(n311) );
    MXL2P U503 ( .OB(n313), .S(n508), .A(\bm[12] ), .B(b[12]) );
    INV2 U504 ( .O(n314), .I(n313) );
    MXL2P U505 ( .OB(n315), .S(n604), .A(\am[54] ), .B(a[54]) );
    INV2 U506 ( .O(n316), .I(n315) );
    MXL2P U507 ( .OB(n317), .S(n518), .A(n453), .B(b[11]) );
    INV2 U508 ( .O(n318), .I(n317) );
    MXL2P U509 ( .OB(n319), .S(n829), .A(\am[55] ), .B(a[55]) );
    INV2 U510 ( .O(n320), .I(n319) );
    MXL2P U511 ( .OB(n321), .S(n825), .A(\bm[10] ), .B(b[10]) );
    INV2 U512 ( .O(n322), .I(n321) );
    MXL2P U513 ( .OB(n323), .S(n831), .A(\am[56] ), .B(a[56]) );
    INV2 U514 ( .O(n324), .I(n323) );
    MXL2P U515 ( .OB(n325), .S(n496), .A(\bm[9] ), .B(b[9]) );
    INV2 U516 ( .O(n326), .I(n325) );
    MXL2P U517 ( .OB(n327), .S(n819), .A(\am[57] ), .B(a[57]) );
    INV2 U518 ( .O(n328), .I(n327) );
    MXL2P U519 ( .OB(n329), .S(n831), .A(\bm[8] ), .B(b[8]) );
    INV2 U520 ( .O(n330), .I(n329) );
    MXL2P U521 ( .OB(n331), .S(n826), .A(\am[58] ), .B(a[58]) );
    INV2 U522 ( .O(n332), .I(n331) );
    MXL2P U523 ( .OB(n333), .S(n612), .A(\bm[7] ), .B(b[7]) );
    INV2 U524 ( .O(n334), .I(n333) );
    MXL2P U525 ( .OB(n335), .S(n362), .A(\am[59] ), .B(a[59]) );
    INV2 U526 ( .O(n336), .I(n335) );
    MXL2P U527 ( .OB(n337), .S(n377), .A(\bm[6] ), .B(b[6]) );
    INV2 U528 ( .O(n338), .I(n337) );
    MXL2P U529 ( .OB(n339), .S(n615), .A(\am[60] ), .B(a[60]) );
    INV2 U530 ( .O(n340), .I(n339) );
    MXL2P U531 ( .OB(n341), .S(n622), .A(\bm[4] ), .B(b[4]) );
    INV2 U532 ( .O(n342), .I(n341) );
    MXL2P U533 ( .OB(n343), .S(n607), .A(\am[61] ), .B(a[61]) );
    INV2 U534 ( .O(n344), .I(n343) );
    MXL2P U535 ( .OB(n345), .S(n825), .A(\bm[3] ), .B(b[3]) );
    INV2 U536 ( .O(n346), .I(n345) );
    MXL2P U537 ( .OB(n347), .S(n825), .A(n494), .B(a[62]) );
    INV2 U538 ( .O(n348), .I(n347) );
    MXL2P U539 ( .OB(n349), .S(n621), .A(\bm[2] ), .B(b[2]) );
    INV2 U540 ( .O(n350), .I(n349) );
    MXL2P U541 ( .OB(n351), .S(n638), .A(\am[63] ), .B(a[63]) );
    INV2 U542 ( .O(n352), .I(n351) );
    MXL2P U543 ( .OB(n353), .S(n358), .A(n448), .B(b[0]) );
    INV2 U544 ( .O(n354), .I(n353) );
    MXL2P U545 ( .OB(n355), .S(n518), .A(\am[44] ), .B(a[44]) );
    INV2 U546 ( .O(n356), .I(n355) );
    INV3 U547 ( .O(n426), .I(n425) );
    DFFRBP \am_reg[53]  ( .Q(\am[53] ), .D(n312), .CK(clk), .RB(n704) );
    DFFRBP \am_reg[45]  ( .Q(\am[45] ), .D(n285), .CK(clk), .RB(n682) );
    DFFRBP \am_reg[55]  ( .Q(\am[55] ), .D(n320), .CK(clk), .RB(n704) );
    DFFRBP \am_reg[57]  ( .Q(\am[57] ), .D(n328), .CK(clk), .RB(n705) );
    DFFRBP \am_reg[3]  ( .Q(\am[3] ), .D(n150), .CK(clk), .RB(n683) );
    DFFRBP \am_reg[59]  ( .Q(\am[59] ), .D(n336), .CK(clk), .RB(n705) );
    DFFRBP \am_reg[1]  ( .Q(\am[1] ), .D(n142), .CK(clk), .RB(n689) );
    INV3 U548 ( .O(n834), .I(n490) );
    INV4 U549 ( .O(n391), .I(n406) );
    INV4 U550 ( .O(n357), .I(n824) );
    INV2 U551 ( .O(n358), .I(n633) );
    MXL2P U552 ( .OB(n840), .S(n639), .A(n360), .B(n359) );
    INV2 U553 ( .O(n359), .I(b[24]) );
    DFFRBP \bm_reg[24]  ( .Q(\bm[24] ), .QB(n360), .D(n840), .CK(clk), .RB(
        n712) );
    ND3T U554 ( .O(n818), .I1(n361), .I2(n516), .I3(\cnt[2] ) );
    INV2 U555 ( .O(n361), .I(n405) );
    DFFRBN \bm_reg[29]  ( .Q(\bm[29] ), .QB(n365), .D(n841), .CK(clk), .RB(
        n670) );
    INV1 U556 ( .O(n362), .I(n525) );
    INV2 U557 ( .O(n363), .I(n422) );
    BUF4 U558 ( .O(n422), .I(n371) );
    MXL2P U559 ( .OB(n841), .S(n820), .A(n365), .B(n364) );
    INV2 U560 ( .O(n364), .I(b[29]) );
    INV4 U561 ( .O(n394), .I(n387) );
    INV2 U562 ( .O(n366), .I(n370) );
    INV4 U563 ( .O(n370), .I(n421) );
    MXL2P U564 ( .OB(n852), .S(n825), .A(n368), .B(n367) );
    INV2 U565 ( .O(n367), .I(a[33]) );
    DFFRBP \am_reg[33]  ( .Q(\am[33] ), .QB(n368), .D(n852), .CK(clk), .RB(
        n698) );
    INV3 U566 ( .O(n369), .I(n613) );
    INV4 U567 ( .O(n613), .I(n633) );
    BUF4 U568 ( .O(n421), .I(n601) );
    BUF4 U569 ( .O(n371), .I(n601) );
    INV4 U570 ( .O(n833), .I(n835) );
    INV3 U571 ( .O(n372), .I(n820) );
    INV3 U572 ( .O(n377), .I(n376) );
    MXL2P U573 ( .OB(n836), .S(n613), .A(n418), .B(n373) );
    INV2 U574 ( .O(n373), .I(b[1]) );
    MXL2P U575 ( .OB(n842), .S(n376), .A(n374), .B(n375) );
    INV2 U576 ( .O(n374), .I(b[39]) );
    BUF4 U577 ( .O(n376), .I(n407) );
    DFFRBP \bm_reg[39]  ( .Q(\bm[39] ), .QB(n375), .D(n842), .CK(clk), .RB(
        n716) );
    MXL2P U578 ( .OB(n843), .S(n376), .A(n379), .B(n380) );
    BUF2 U579 ( .O(n410), .I(n820) );
    INV4 U580 ( .O(n407), .I(n403) );
    BUF4 U581 ( .O(n403), .I(n601) );
    INV4 U582 ( .O(n387), .I(n390) );
    BUF4 U583 ( .O(n390), .I(n366) );
    INV2 U584 ( .O(n379), .I(b[40]) );
    DFFRBP \bm_reg[40]  ( .Q(\bm[40] ), .QB(n380), .D(n843), .CK(clk), .RB(
        n716) );
    MXL2P U585 ( .OB(n848), .S(n622), .A(n382), .B(n381) );
    INV2 U586 ( .O(n381), .I(a[7]) );
    DFFRBP \am_reg[7]  ( .Q(\am[7] ), .QB(n382), .D(n848), .CK(clk), .RB(n676)
         );
    INV2 U587 ( .O(n383), .I(n396) );
    BUF4 U588 ( .O(n413), .I(n642) );
    MXL2P U589 ( .OB(n845), .S(n404), .A(n385), .B(n384) );
    INV2 U590 ( .O(n384), .I(b[56]) );
    DFFRBP \bm_reg[56]  ( .Q(\bm[56] ), .QB(n385), .D(n845), .CK(clk), .RB(
        n663) );
    INV2 U591 ( .O(n386), .I(n387) );
    MXL2P U592 ( .OB(n853), .S(n390), .A(n389), .B(n388) );
    INV2 U593 ( .O(n388), .I(a[37]) );
    DFFRBP \am_reg[37]  ( .Q(\am[37] ), .QB(n389), .D(n853), .CK(clk), .RB(
        n699) );
    BUF4 U594 ( .O(n404), .I(n421) );
    BUF4 U595 ( .O(n518), .I(n496) );
    INV4 U596 ( .O(n496), .I(n409) );
    MXL2P U597 ( .OB(n837), .S(n609), .A(n393), .B(n392) );
    INV2 U598 ( .O(n392), .I(b[5]) );
    DFFRBP \bm_reg[5]  ( .Q(\bm[5] ), .QB(n393), .D(n837), .CK(clk), .RB(n662)
         );
    BUF4 U599 ( .O(n634), .I(n834) );
    BUF3 U600 ( .O(n395), .I(n600) );
    BUF3 U601 ( .O(n409), .I(n363) );
    BUF3 U602 ( .O(n396), .I(n834) );
    MXL2P U603 ( .OB(n838), .S(n496), .A(n398), .B(n397) );
    INV2 U604 ( .O(n397), .I(b[20]) );
    MXL2P U605 ( .OB(n850), .S(n617), .A(n433), .B(n399) );
    INV2 U606 ( .O(n399), .I(a[29]) );
    MXL2P U607 ( .OB(n844), .S(n616), .A(n401), .B(n400) );
    INV2 U608 ( .O(n400), .I(b[45]) );
    INV2 U609 ( .O(n402), .I(n490) );
    JKFRBN \cnt_reg[0]  ( .QB(n858), .J(1'b1), .K(1'b1), .CK(clk), .RB(n763)
         );
    BUF2 U610 ( .O(n405), .I(n451) );
    BUF1 U611 ( .O(n451), .I(n858) );
    BUF3 U612 ( .O(n629), .I(n818) );
    BUF4 U613 ( .O(n406), .I(n403) );
    INV4 U614 ( .O(n408), .I(n631) );
    BUF3 U615 ( .O(n522), .I(n635) );
    INV4 U616 ( .O(n525), .I(n404) );
    MXL2P U617 ( .OB(n854), .S(n377), .A(n412), .B(n411) );
    INV2 U618 ( .O(n411), .I(a[40]) );
    DFFRBP \am_reg[40]  ( .Q(\am[40] ), .QB(n412), .D(n854), .CK(clk), .RB(
        n700) );
    INV4 U619 ( .O(n631), .I(n371) );
    BUF2 U620 ( .O(n414), .I(n523) );
    MXL2P U621 ( .OB(n856), .S(n606), .A(n416), .B(n415) );
    INV2 U622 ( .O(n415), .I(a[50]) );
    DFFRBP \am_reg[50]  ( .Q(\am[50] ), .QB(n416), .D(n856), .CK(clk), .RB(
        n680) );
    BUF3 U623 ( .O(n417), .I(n631) );
    BUF4 U624 ( .O(n490), .I(n523) );
    DFFRBP \bm_reg[1]  ( .Q(\bm[1] ), .QB(n418), .D(n836), .CK(clk), .RB(n673)
         );
    BUF3 U625 ( .O(n504), .I(\bm[60] ) );
    QDFFRBP \s_reg[63]  ( .Q(n419), .D(n14), .CK(clk), .RB(n646) );
    MUX2P U626 ( .O(n849), .S(n823), .A(\am[11] ), .B(a[11]) );
    BUF4 U627 ( .O(n502), .I(\bm[61] ) );
    BUF4 U628 ( .O(n633), .I(n611) );
    INV1 U629 ( .O(n420), .I(n378) );
    BUF3 U630 ( .O(n423), .I(n391) );
    INV3 U631 ( .O(n424), .I(n639) );
    INV4 U632 ( .O(n639), .I(n357) );
    INV3 U633 ( .O(n425), .I(n833) );
    INV1 U634 ( .O(n428), .I(n427) );
    DFFRBP \am_reg[46]  ( .Q(\am[46] ), .QB(n427), .D(n289), .CK(clk), .RB(
        n702) );
    INV1 U635 ( .O(n430), .I(n429) );
    DFFRBP \am_reg[49]  ( .Q(\am[49] ), .QB(n429), .D(n300), .CK(clk), .RB(
        n681) );
    INV1 U636 ( .O(n432), .I(n431) );
    DFFRBP \am_reg[51]  ( .Q(\am[51] ), .QB(n431), .D(n304), .CK(clk), .RB(
        n703) );
    DFFRBP \am_reg[29]  ( .Q(\am[29] ), .QB(n433), .D(n850), .CK(clk), .RB(
        n686) );
    INV1 U637 ( .O(n435), .I(n434) );
    DFFRBP \am_reg[6]  ( .Q(\am[6] ), .QB(n434), .D(n161), .CK(clk), .RB(n707)
         );
    INV1 U638 ( .O(n437), .I(n436) );
    DFFRBP \bm_reg[37]  ( .Q(\bm[37] ), .QB(n436), .D(n233), .CK(clk), .RB(
        n715) );
    INV1 U639 ( .O(n439), .I(n438) );
    DFFRBP \bm_reg[33]  ( .Q(\bm[33] ), .QB(n438), .D(n249), .CK(clk), .RB(
        n714) );
    INV1 U640 ( .O(n441), .I(n440) );
    DFFRBP \bm_reg[31]  ( .Q(\bm[31] ), .QB(n440), .D(n256), .CK(clk), .RB(
        n714) );
    INV1 U641 ( .O(n443), .I(n442) );
    DFFRBP \bm_reg[18]  ( .Q(\bm[18] ), .QB(n442), .D(n291), .CK(clk), .RB(
        n673) );
    INV1 U642 ( .O(n445), .I(n444) );
    DFFRBP \bm_reg[15]  ( .Q(\bm[15] ), .QB(n444), .D(n302), .CK(clk), .RB(
        n709) );
    INV1 U643 ( .O(n447), .I(n446) );
    DFFRBP \bm_reg[21]  ( .Q(\bm[21] ), .QB(n446), .D(n283), .CK(clk), .RB(
        n672) );
    DFFRBP \bm_reg[0]  ( .Q(\bm[0] ), .D(n354), .CK(clk), .RB(n708) );
    DFFRBP \bm_reg[35]  ( .Q(\bm[35] ), .D(n241), .CK(clk), .RB(n715) );
    INV2 U644 ( .O(n450), .I(n521) );
    BUF4 U645 ( .O(n521), .I(n832) );
    DFFRBP \am_reg[63]  ( .Q(\am[63] ), .D(n352), .CK(clk), .RB(n677) );
    BUF2 U646 ( .O(n517), .I(n420) );
    INV1 U647 ( .O(n453), .I(n452) );
    DFFRBP \bm_reg[11]  ( .Q(\bm[11] ), .QB(n452), .D(n318), .CK(clk), .RB(
        n708) );
    INV1 U648 ( .O(n455), .I(n454) );
    DFFRBP \am_reg[20]  ( .Q(\am[20] ), .QB(n454), .D(n211), .CK(clk), .RB(
        n695) );
    INV1 U649 ( .O(n457), .I(n456) );
    DFFRBP \am_reg[32]  ( .Q(\am[32] ), .QB(n456), .D(n254), .CK(clk), .RB(
        n685) );
    INV1 U650 ( .O(n459), .I(n458) );
    DFFRBP \am_reg[17]  ( .Q(\am[17] ), .QB(n458), .D(n199), .CK(clk), .RB(
        n694) );
    INV1 U651 ( .O(n461), .I(n460) );
    DFFRBP \am_reg[36]  ( .Q(\am[36] ), .QB(n460), .D(n266), .CK(clk), .RB(
        n684) );
    INV2 U652 ( .O(n822), .I(n605) );
    BUF2 U653 ( .O(n462), .I(\bm[29] ) );
    BUF2 U654 ( .O(n463), .I(\bm[10] ) );
    DFFRBP \bm_reg[10]  ( .Q(\bm[10] ), .D(n322), .CK(clk), .RB(n675) );
    BUF2 U655 ( .O(n464), .I(\bm[53] ) );
    DFFRBP \bm_reg[53]  ( .Q(\bm[53] ), .D(n181), .CK(clk), .RB(n720) );
    BUF2 U656 ( .O(n465), .I(\bm[3] ) );
    DFFRBP \bm_reg[3]  ( .Q(\bm[3] ), .D(n346), .CK(clk), .RB(n691) );
    BUF2 U657 ( .O(n466), .I(\bm[57] ) );
    DFFRBP \bm_reg[57]  ( .Q(\bm[57] ), .D(n170), .CK(clk), .RB(n721) );
    BUF2 U658 ( .O(n467), .I(\bm[49] ) );
    DFFRBP \bm_reg[49]  ( .Q(\bm[49] ), .D(n197), .CK(clk), .RB(n665) );
    BUF2 U659 ( .O(n468), .I(\bm[46] ) );
    DFFRBP \bm_reg[46]  ( .Q(\bm[46] ), .D(n209), .CK(clk), .RB(n718) );
    BUF2 U660 ( .O(n469), .I(\bm[51] ) );
    DFFRBP \bm_reg[51]  ( .Q(\bm[51] ), .D(n189), .CK(clk), .RB(n719) );
    DFFRBP \bm_reg[45]  ( .Q(\bm[45] ), .QB(n401), .D(n844), .CK(clk), .RB(
        n666) );
    BUF2 U661 ( .O(n470), .I(\bm[55] ) );
    DFFRBP \bm_reg[55]  ( .Q(\bm[55] ), .D(n174), .CK(clk), .RB(n720) );
    BUF2 U662 ( .O(n471), .I(\bm[6] ) );
    DFFRBP \bm_reg[6]  ( .Q(\bm[6] ), .D(n338), .CK(clk), .RB(n723) );
    BUF2 U663 ( .O(n472), .I(\bm[59] ) );
    DFFRBP \bm_reg[59]  ( .Q(\bm[59] ), .D(n163), .CK(clk), .RB(n721) );
    BUF2 U664 ( .O(n473), .I(n372) );
    BUF3 U665 ( .O(n479), .I(n630) );
    BUF3 U666 ( .O(n503), .I(n833) );
    DFFRBP \bm_reg[30]  ( .Q(\bm[30] ), .D(n260), .CK(clk), .RB(n670) );
    DFFRBP \bm_reg[32]  ( .Q(\bm[32] ), .D(n253), .CK(clk), .RB(n669) );
    DFFRBP \bm_reg[36]  ( .Q(\bm[36] ), .D(n237), .CK(clk), .RB(n668) );
    DFFRBP \bm_reg[17]  ( .Q(\bm[17] ), .D(n295), .CK(clk), .RB(n710) );
    BUF3 U667 ( .O(n480), .I(n833) );
    INV3 U668 ( .O(n481), .I(n518) );
    INV3 U669 ( .O(n597), .I(n394) );
    BUF4 U670 ( .O(n635), .I(n636) );
    INV3 U671 ( .O(n602), .I(n830) );
    INV3 U672 ( .O(n482), .I(n830) );
    INV4 U673 ( .O(n830), .I(n635) );
    BUF3 U674 ( .O(n483), .I(n372) );
    BUF3 U675 ( .O(n484), .I(n832) );
    BUF3 U676 ( .O(n485), .I(n632) );
    BUF3 U677 ( .O(n486), .I(n632) );
    BUF2 U678 ( .O(n632), .I(n832) );
    BUF3 U679 ( .O(n487), .I(n396) );
    BUF3 U680 ( .O(n488), .I(n634) );
    BUF2 U681 ( .O(n489), .I(\am[34] ) );
    DFFRBP \am_reg[34]  ( .Q(\am[34] ), .D(n258), .CK(clk), .RB(n685) );
    DFFRBP \am_reg[0]  ( .Q(\am[0] ), .D(n144), .CK(clk), .RB(n740) );
    BUF3 U682 ( .O(n492), .I(\am[61] ) );
    DFFRBP \am_reg[61]  ( .Q(\am[61] ), .D(n344), .CK(clk), .RB(n677) );
    INV3 U683 ( .O(n493), .I(\am[62] ) );
    INV4 U684 ( .O(n494), .I(n493) );
    BUF3 U685 ( .O(n495), .I(\am[60] ) );
    DFFRBP \am_reg[60]  ( .Q(\am[60] ), .D(n340), .CK(clk), .RB(n706) );
    DFFRBP \bm_reg[63]  ( .Q(\bm[63] ), .D(n148), .CK(clk), .RB(n661) );
    DFFRBP \am_reg[26]  ( .Q(\am[26] ), .D(n235), .CK(clk), .RB(n696) );
    DFFRBP \am_reg[22]  ( .Q(\am[22] ), .D(n219), .CK(clk), .RB(n695) );
    DFFRBP \am_reg[38]  ( .Q(\am[38] ), .D(n270), .CK(clk), .RB(n684) );
    DFFRBP \am_reg[13]  ( .Q(\am[13] ), .D(n183), .CK(clk), .RB(n693) );
    DFFRBP \bm_reg[61]  ( .Q(\bm[61] ), .D(n156), .CK(clk), .RB(n661) );
    DFFRBP \bm_reg[60]  ( .Q(\bm[60] ), .D(n160), .CK(clk), .RB(n722) );
    BUF3 U686 ( .O(n505), .I(\bm[62] ) );
    DFFRBP \bm_reg[62]  ( .Q(\bm[62] ), .D(n152), .CK(clk), .RB(n722) );
    BUF3 U687 ( .O(n506), .I(\bm[34] ) );
    DFFRBP \bm_reg[34]  ( .Q(\bm[34] ), .D(n245), .CK(clk), .RB(n669) );
    DFFRBP \am_reg[47]  ( .Q(\am[47] ), .D(n293), .CK(clk), .RB(n681) );
    XNR2P U688 ( .O(N7), .I1(\cnt[2] ), .I2(n859) );
    INV2 U689 ( .O(n508), .I(n520) );
    BUF4 U690 ( .O(n520), .I(n832) );
    BUF4 U691 ( .O(n509), .I(\bm[26] ) );
    DFFRBP \bm_reg[26]  ( .Q(\bm[26] ), .D(n272), .CK(clk), .RB(n712) );
    BUF4 U692 ( .O(n510), .I(\bm[42] ) );
    DFFRBP \bm_reg[42]  ( .Q(\bm[42] ), .D(n221), .CK(clk), .RB(n717) );
    BUF4 U693 ( .O(n511), .I(\bm[13] ) );
    DFFRBP \bm_reg[13]  ( .Q(\bm[13] ), .D(n310), .CK(clk), .RB(n709) );
    DFFRBP \am_reg[35]  ( .Q(\am[35] ), .D(n262), .CK(clk), .RB(n699) );
    BUF4 U694 ( .O(n513), .I(\bm[38] ) );
    DFFRBP \bm_reg[38]  ( .Q(\bm[38] ), .D(n229), .CK(clk), .RB(n692) );
    DFFRBP \bm_reg[47]  ( .Q(\bm[47] ), .D(n205), .CK(clk), .RB(n665) );
    BUF4 U695 ( .O(n515), .I(\bm[22] ) );
    DFFRBP \bm_reg[22]  ( .Q(\bm[22] ), .D(n281), .CK(clk), .RB(n711) );
    BUF4 U696 ( .O(n516), .I(\cnt[1] ) );
    INV4 U697 ( .O(n817), .I(n391) );
    INV3 U698 ( .O(n519), .I(n414) );
    INV3 U699 ( .O(n640), .I(n369) );
    INV4 U700 ( .O(n523), .I(n407) );
    INV3 U701 ( .O(n524), .I(n413) );
    BUF3 U702 ( .O(s[24]), .I(n898) );
    DFFRBP \s_reg[24]  ( .Q(n898), .D(n20), .CK(clk), .RB(n728) );
    BUF3 U703 ( .O(s[16]), .I(n906) );
    DFFRBP \s_reg[16]  ( .Q(n906), .D(n64), .CK(clk), .RB(n658) );
    BUF3 U704 ( .O(s[55]), .I(n867) );
    DFFRBP \s_reg[55]  ( .Q(n867), .D(n38), .CK(clk), .RB(n736) );
    BUF3 U705 ( .O(s[13]), .I(n909) );
    DFFRBP \s_reg[13]  ( .Q(n909), .D(n36), .CK(clk), .RB(n725) );
    BUF3 U706 ( .O(s[58]), .I(n864) );
    DFFRBP \s_reg[58]  ( .Q(n864), .D(n134), .CK(clk), .RB(n649) );
    BUF3 U707 ( .O(s[12]), .I(n910) );
    DFFRBP \s_reg[12]  ( .Q(n910), .D(n104), .CK(clk), .RB(n659) );
    BUF3 U708 ( .O(s[59]), .I(n863) );
    DFFRBP \s_reg[59]  ( .Q(n863), .D(n46), .CK(clk), .RB(n737) );
    BUF3 U709 ( .O(s[32]), .I(n890) );
    DFFRBP \s_reg[32]  ( .Q(n890), .D(n94), .CK(clk), .RB(n653) );
    BUF3 U710 ( .O(s[33]), .I(n889) );
    DFFRBP \s_reg[33]  ( .Q(n889), .D(n28), .CK(clk), .RB(n730) );
    BUF3 U711 ( .O(s[31]), .I(n891) );
    DFFRBP \s_reg[31]  ( .Q(n891), .D(n32), .CK(clk), .RB(n730) );
    BUF3 U712 ( .O(s[34]), .I(n888) );
    DFFRBP \s_reg[34]  ( .Q(n888), .D(n72), .CK(clk), .RB(n653) );
    BUF3 U713 ( .O(s[30]), .I(n892) );
    DFFRBP \s_reg[30]  ( .Q(n892), .D(n90), .CK(clk), .RB(n654) );
    BUF3 U714 ( .O(s[35]), .I(n887) );
    DFFRBP \s_reg[35]  ( .Q(n887), .D(n98), .CK(clk), .RB(n731) );
    BUF3 U715 ( .O(s[29]), .I(n893) );
    DFFRBP \s_reg[29]  ( .Q(n893), .D(n86), .CK(clk), .RB(n654) );
    BUF3 U716 ( .O(s[36]), .I(n886) );
    DFFRBP \s_reg[36]  ( .Q(n886), .D(n102), .CK(clk), .RB(n652) );
    BUF3 U717 ( .O(s[28]), .I(n894) );
    DFFRBP \s_reg[28]  ( .Q(n894), .D(n58), .CK(clk), .RB(n729) );
    BUF3 U718 ( .O(s[37]), .I(n885) );
    DFFRBP \s_reg[37]  ( .Q(n885), .D(n62), .CK(clk), .RB(n731) );
    BUF3 U719 ( .O(s[27]), .I(n895) );
    DFFRBP \s_reg[27]  ( .Q(n895), .D(n82), .CK(clk), .RB(n655) );
    BUF3 U720 ( .O(s[38]), .I(n884) );
    DFFRBP \s_reg[38]  ( .Q(n884), .D(n74), .CK(clk), .RB(n652) );
    BUF3 U721 ( .O(s[26]), .I(n896) );
    DFFRBP \s_reg[26]  ( .Q(n896), .D(n76), .CK(clk), .RB(n728) );
    BUF3 U722 ( .O(s[39]), .I(n883) );
    DFFRBP \s_reg[39]  ( .Q(n883), .D(n106), .CK(clk), .RB(n732) );
    BUF3 U723 ( .O(s[25]), .I(n897) );
    DFFRBP \s_reg[25]  ( .Q(n897), .D(n56), .CK(clk), .RB(n667) );
    BUF3 U724 ( .O(s[40]), .I(n882) );
    DFFRBP \s_reg[40]  ( .Q(n882), .D(n22), .CK(clk), .RB(n732) );
    BUF3 U725 ( .O(s[23]), .I(n899) );
    DFFRBP \s_reg[23]  ( .Q(n899), .D(n84), .CK(clk), .RB(n656) );
    BUF3 U726 ( .O(s[41]), .I(n881) );
    DFFRBP \s_reg[41]  ( .Q(n881), .D(n66), .CK(clk), .RB(n651) );
    BUF3 U727 ( .O(s[22]), .I(n900) );
    DFFRBP \s_reg[22]  ( .Q(n900), .D(n80), .CK(clk), .RB(n727) );
    BUF3 U728 ( .O(s[42]), .I(n880) );
    DFFRBP \s_reg[42]  ( .Q(n880), .D(n78), .CK(clk), .RB(n733) );
    BUF3 U729 ( .O(s[21]), .I(n901) );
    DFFRBP \s_reg[21]  ( .Q(n901), .D(n60), .CK(clk), .RB(n656) );
    BUF3 U730 ( .O(s[43]), .I(n879) );
    DFFRBP \s_reg[43]  ( .Q(n879), .D(n110), .CK(clk), .RB(n650) );
    BUF3 U731 ( .O(s[20]), .I(n902) );
    DFFRBP \s_reg[20]  ( .Q(n902), .D(n88), .CK(clk), .RB(n727) );
    BUF3 U732 ( .O(s[44]), .I(n878) );
    DFFRBP \s_reg[44]  ( .Q(n878), .D(n70), .CK(clk), .RB(n733) );
    BUF3 U733 ( .O(s[19]), .I(n903) );
    DFFRBP \s_reg[19]  ( .Q(n903), .D(n92), .CK(clk), .RB(n726) );
    BUF3 U734 ( .O(s[45]), .I(n877) );
    DFFRBP \s_reg[45]  ( .Q(n877), .D(n114), .CK(clk), .RB(n650) );
    BUF3 U735 ( .O(s[18]), .I(n904) );
    DFFRBP \s_reg[18]  ( .Q(n904), .D(n96), .CK(clk), .RB(n657) );
    BUF3 U736 ( .O(s[46]), .I(n876) );
    DFFRBP \s_reg[46]  ( .Q(n876), .D(n118), .CK(clk), .RB(n734) );
    BUF3 U737 ( .O(s[17]), .I(n905) );
    DFFRBP \s_reg[17]  ( .Q(n905), .D(n16), .CK(clk), .RB(n726) );
    BUF3 U738 ( .O(s[47]), .I(n875) );
    DFFRBP \s_reg[47]  ( .Q(n875), .D(n24), .CK(clk), .RB(n655) );
    BUF3 U739 ( .O(s[15]), .I(n907) );
    DFFRBP \s_reg[15]  ( .Q(n907), .D(n68), .CK(clk), .RB(n725) );
    BUF3 U740 ( .O(s[48]), .I(n874) );
    DFFRBP \s_reg[48]  ( .Q(n874), .D(n136), .CK(clk), .RB(n734) );
    BUF3 U741 ( .O(s[14]), .I(n908) );
    DFFRBP \s_reg[14]  ( .Q(n908), .D(n100), .CK(clk), .RB(n658) );
    BUF3 U742 ( .O(s[49]), .I(n873) );
    DFFRBP \s_reg[49]  ( .Q(n873), .D(n26), .CK(clk), .RB(n649) );
    BUF3 U743 ( .O(s[11]), .I(n911) );
    DFFRBP \s_reg[11]  ( .Q(n911), .D(n108), .CK(clk), .RB(n724) );
    BUF3 U744 ( .O(s[50]), .I(n872) );
    DFFRBP \s_reg[50]  ( .Q(n872), .D(n122), .CK(clk), .RB(n648) );
    BUF3 U745 ( .O(s[10]), .I(n912) );
    DFFRBP \s_reg[10]  ( .Q(n912), .D(n112), .CK(clk), .RB(n659) );
    BUF3 U746 ( .O(s[51]), .I(n871) );
    DFFRBP \s_reg[51]  ( .Q(n871), .D(n30), .CK(clk), .RB(n735) );
    BUF3 U747 ( .O(s[9]), .I(n913) );
    DFFRBP \s_reg[9]  ( .Q(n913), .D(n40), .CK(clk), .RB(n667) );
    BUF3 U748 ( .O(s[52]), .I(n870) );
    DFFRBP \s_reg[52]  ( .Q(n870), .D(n138), .CK(clk), .RB(n648) );
    BUF3 U749 ( .O(s[8]), .I(n914) );
    DFFRBP \s_reg[8]  ( .Q(n914), .D(n116), .CK(clk), .RB(n739) );
    BUF3 U750 ( .O(s[53]), .I(n869) );
    DFFRBP \s_reg[53]  ( .Q(n869), .D(n34), .CK(clk), .RB(n736) );
    BUF3 U751 ( .O(s[7]), .I(n915) );
    DFFRBP \s_reg[7]  ( .Q(n915), .D(n120), .CK(clk), .RB(n645) );
    BUF3 U752 ( .O(s[54]), .I(n868) );
    DFFRBP \s_reg[54]  ( .Q(n868), .D(n126), .CK(clk), .RB(n647) );
    BUF3 U753 ( .O(s[6]), .I(n916) );
    DFFRBP \s_reg[6]  ( .Q(n916), .D(n124), .CK(clk), .RB(n739) );
    BUF3 U754 ( .O(s[56]), .I(n866) );
    DFFRBP \s_reg[56]  ( .Q(n866), .D(n130), .CK(clk), .RB(n647) );
    BUF3 U755 ( .O(s[5]), .I(n917) );
    DFFRBP \s_reg[5]  ( .Q(n917), .D(n44), .CK(clk), .RB(n646) );
    BUF3 U756 ( .O(s[57]), .I(n865) );
    DFFRBP \s_reg[57]  ( .Q(n865), .D(n42), .CK(clk), .RB(n737) );
    BUF3 U757 ( .O(s[4]), .I(n918) );
    DFFRBP \s_reg[4]  ( .Q(n918), .D(n128), .CK(clk), .RB(n735) );
    BUF3 U758 ( .O(s[60]), .I(n862) );
    DFFRBP \s_reg[60]  ( .Q(n862), .D(n50), .CK(clk), .RB(n738) );
    BUF3 U759 ( .O(s[3]), .I(n919) );
    DFFRBP \s_reg[3]  ( .Q(n919), .D(n48), .CK(clk), .RB(n651) );
    BUF3 U760 ( .O(s[61]), .I(n861) );
    DFFRBP \s_reg[61]  ( .Q(n861), .D(n18), .CK(clk), .RB(n645) );
    BUF3 U761 ( .O(s[2]), .I(n920) );
    DFFRBP \s_reg[2]  ( .Q(n920), .D(n132), .CK(clk), .RB(n729) );
    BUF3 U762 ( .O(s[62]), .I(n860) );
    DFFRBP \s_reg[62]  ( .Q(n860), .D(n52), .CK(clk), .RB(n738) );
    BUF3 U763 ( .O(s[1]), .I(n921) );
    DFFRBP \s_reg[1]  ( .Q(n921), .D(n54), .CK(clk), .RB(n657) );
    BUF3 U764 ( .O(s[63]), .I(n419) );
    BUF3 U765 ( .O(s[0]), .I(n922) );
    DFFRBP \s_reg[0]  ( .Q(n922), .D(n140), .CK(clk), .RB(n724) );
    INV1 U766 ( .O(n592), .I(n591) );
    DFFRBP \am_reg[30]  ( .Q(\am[30] ), .QB(n591), .D(n247), .CK(clk), .RB(
        n686) );
    INV4 U767 ( .O(n593), .I(n479) );
    INV4 U768 ( .O(n630), .I(n422) );
    INV4 U769 ( .O(n594), .I(n482) );
    INV4 U770 ( .O(n595), .I(n605) );
    INV3 U771 ( .O(n596), .I(n595) );
    INV3 U772 ( .O(n598), .I(n595) );
    INV4 U773 ( .O(n600), .I(n481) );
    INV4 U774 ( .O(n599), .I(n596) );
    INV4 U775 ( .O(n601), .I(n629) );
    INV4 U776 ( .O(n603), .I(n503) );
    INV4 U777 ( .O(n604), .I(n602) );
    BUF4 U778 ( .O(n605), .I(n402) );
    INV4 U779 ( .O(n607), .I(n486) );
    INV4 U780 ( .O(n606), .I(n484) );
    INV4 U781 ( .O(n608), .I(n424) );
    INV4 U782 ( .O(n609), .I(n423) );
    INV4 U783 ( .O(n610), .I(n480) );
    INV4 U784 ( .O(n611), .I(n823) );
    INV4 U785 ( .O(n612), .I(n611) );
    INV3 U786 ( .O(n615), .I(n426) );
    INV3 U787 ( .O(n614), .I(n473) );
    MUX2P U788 ( .O(n851), .S(n637), .A(n457), .B(a[32]) );
    BUF4 U789 ( .O(n616), .I(n607) );
    BUF4 U790 ( .O(n617), .I(n607) );
    BUF4 U791 ( .O(n618), .I(n450) );
    BUF4 U792 ( .O(n619), .I(n640) );
    BUF4 U793 ( .O(n620), .I(n638) );
    BUF4 U794 ( .O(n621), .I(n638) );
    BUF4 U795 ( .O(n622), .I(n523) );
    BUF4 U796 ( .O(n623), .I(n637) );
    BUF4 U797 ( .O(n624), .I(n637) );
    BUF4 U798 ( .O(n625), .I(n821) );
    BUF4 U799 ( .O(n626), .I(n821) );
    BUF4 U800 ( .O(n627), .I(n410) );
    BUF4 U801 ( .O(n628), .I(n410) );
    MUX2P U802 ( .O(n847), .S(n637), .A(n435), .B(a[6]) );
    INV4 U803 ( .O(n636), .I(n817) );
    INV4 U804 ( .O(n835), .I(n417) );
    INV4 U805 ( .O(n638), .I(n519) );
    INV4 U806 ( .O(n637), .I(n521) );
    INV4 U807 ( .O(n832), .I(n408) );
    INV4 U808 ( .O(n641), .I(n524) );
    INV4 U809 ( .O(n642), .I(n525) );
    INV4 U810 ( .O(n643), .I(n488) );
    DFFRBT \am_reg[58]  ( .Q(\am[58] ), .D(n332), .CK(clk), .RB(n678) );
    DFFRBT \am_reg[11]  ( .Q(\am[11] ), .D(n175), .CK(clk), .RB(n740) );
    DFFRBT \am_reg[56]  ( .Q(\am[56] ), .D(n324), .CK(clk), .RB(n679) );
    DFFRBT \am_reg[52]  ( .Q(\am[52] ), .D(n308), .CK(clk), .RB(n680) );
    DFFRBT \am_reg[48]  ( .Q(\am[48] ), .D(n296), .CK(clk), .RB(n702) );
    DFFRBT \am_reg[54]  ( .Q(\am[54] ), .D(n316), .CK(clk), .RB(n679) );
    DFFRBT \am_reg[2]  ( .Q(\am[2] ), .D(n146), .CK(clk), .RB(n697) );
    DFFRBT \am_reg[14]  ( .Q(\am[14] ), .D(n187), .CK(clk), .RB(n690) );
    DFFRBT \am_reg[8]  ( .Q(\am[8] ), .D(n165), .CK(clk), .RB(n707) );
    DFFRBT \am_reg[10]  ( .Q(\am[10] ), .D(n172), .CK(clk), .RB(n692) );
    DFFRBT \am_reg[27]  ( .Q(\am[27] ), .D(n239), .CK(clk), .RB(n687) );
    DFFRBT \am_reg[23]  ( .Q(\am[23] ), .D(n223), .CK(clk), .RB(n688) );
    DFFRBT \am_reg[39]  ( .Q(\am[39] ), .D(n274), .CK(clk), .RB(n700) );
    DFFRBT \am_reg[19]  ( .Q(\am[19] ), .D(n207), .CK(clk), .RB(n694) );
    DFFRBT \bm_reg[43]  ( .Q(\bm[43] ), .D(n217), .CK(clk), .RB(n666) );
    DFFRBT \bm_reg[27]  ( .Q(\bm[27] ), .D(n268), .CK(clk), .RB(n671) );
    DFFRBT \bm_reg[2]  ( .Q(\bm[2] ), .D(n350), .CK(clk), .RB(n713) );
    DFFRBT \bm_reg[23]  ( .Q(\bm[23] ), .D(n279), .CK(clk), .RB(n672) );
    DFFRBT \bm_reg[50]  ( .Q(\bm[50] ), .D(n193), .CK(clk), .RB(n664) );
    DFFRBT \bm_reg[19]  ( .Q(\bm[19] ), .D(n287), .CK(clk), .RB(n710) );
    DFFRBT \bm_reg[52]  ( .Q(\bm[52] ), .D(n185), .CK(clk), .RB(n664) );
    DFFRBT \bm_reg[54]  ( .Q(\bm[54] ), .D(n177), .CK(clk), .RB(n663) );
    DFFRBT \bm_reg[48]  ( .Q(\bm[48] ), .D(n201), .CK(clk), .RB(n718) );
    DFFRBT \bm_reg[58]  ( .Q(\bm[58] ), .D(n167), .CK(clk), .RB(n662) );
    DFFRBT \am_reg[16]  ( .Q(\am[16] ), .D(n195), .CK(clk), .RB(n690) );
    DFFRBT \am_reg[15]  ( .Q(\am[15] ), .D(n191), .CK(clk), .RB(n693) );
    DFFRBT \am_reg[18]  ( .Q(\am[18] ), .D(n203), .CK(clk), .RB(n689) );
    DFFRBT \am_reg[31]  ( .Q(\am[31] ), .D(n251), .CK(clk), .RB(n698) );
    DFFRBT \am_reg[24]  ( .Q(\am[24] ), .D(n227), .CK(clk), .RB(n696) );
    DFFRBT \bm_reg[16]  ( .Q(\bm[16] ), .D(n298), .CK(clk), .RB(n674) );
    DFFRBT \bm_reg[7]  ( .Q(\bm[7] ), .D(n334), .CK(clk), .RB(n660) );
    DFFRBT \am_reg[5]  ( .Q(\am[5] ), .D(n158), .CK(clk), .RB(n678) );
    DFFRBT \bm_reg[8]  ( .Q(\bm[8] ), .D(n330), .CK(clk), .RB(n723) );
    DFFRBT \bm_reg[9]  ( .Q(\bm[9] ), .D(n326), .CK(clk), .RB(n660) );
    DFFRBT \bm_reg[4]  ( .Q(\bm[4] ), .D(n342), .CK(clk), .RB(n719) );
    DFFRBT \am_reg[21]  ( .Q(\am[21] ), .D(n215), .CK(clk), .RB(n688) );
    DFFRBT \bm_reg[14]  ( .Q(\bm[14] ), .D(n306), .CK(clk), .RB(n674) );
    DFFRBT \bm_reg[12]  ( .Q(\bm[12] ), .D(n314), .CK(clk), .RB(n675) );
    DFFRBT \am_reg[12]  ( .Q(\am[12] ), .D(n179), .CK(clk), .RB(n691) );
    DFFRBT \bm_reg[44]  ( .Q(\bm[44] ), .D(n213), .CK(clk), .RB(n717) );
    DFFRBT \am_reg[44]  ( .Q(\am[44] ), .D(n356), .CK(clk), .RB(n701) );
    DFFRBT \bm_reg[28]  ( .Q(\bm[28] ), .D(n264), .CK(clk), .RB(n713) );
    DFFRBT \am_reg[28]  ( .Q(\am[28] ), .D(n243), .CK(clk), .RB(n697) );
    DFFRBT \bm_reg[25]  ( .Q(\bm[25] ), .D(n276), .CK(clk), .RB(n671) );
    DFFRBT \am_reg[25]  ( .Q(\am[25] ), .D(n231), .CK(clk), .RB(n687) );
    DFFRBT \bm_reg[41]  ( .Q(\bm[41] ), .D(n225), .CK(clk), .RB(n668) );
    DFFRBT \am_reg[41]  ( .Q(\am[41] ), .D(n278), .CK(clk), .RB(n683) );
    BUF4 U811 ( .O(n701), .I(n760) );
    adder_DW01_add_64_1 add_52 ( .A({\am[63] , n494, n492, n495, \am[59] , 
        \am[58] , \am[57] , \am[56] , \am[55] , \am[54] , \am[53] , \am[52] , 
        \am[51] , \am[50] , \am[49] , \am[48] , n507, \am[46] , \am[45] , 
        \am[44] , \am[43] , n501, \am[41] , \am[40] , \am[39] , n499, \am[37] , 
        \am[36] , n512, n489, \am[33] , \am[32] , \am[31] , \am[30] , \am[29] , 
        \am[28] , \am[27] , n497, \am[25] , \am[24] , \am[23] , n498, \am[21] , 
        \am[20] , \am[19] , \am[18] , \am[17] , \am[16] , \am[15] , \am[14] , 
        n500, \am[12] , \am[11] , \am[10] , \am[9] , \am[8] , \am[7] , \am[6] , 
        \am[5] , \am[4] , \am[3] , \am[2] , \am[1] , n491}), .B({\bm[63] , 
        n505, n502, n504, n472, \bm[58] , n466, \bm[56] , n470, \bm[54] , n464, 
        \bm[52] , n469, \bm[50] , n467, \bm[48] , n514, n468, \bm[45] , 
        \bm[44] , \bm[43] , n510, \bm[41] , \bm[40] , \bm[39] , n513, \bm[37] , 
        n477, n449, n506, \bm[33] , n475, \bm[31] , n474, n462, \bm[28] , 
        \bm[27] , n509, \bm[25] , \bm[24] , \bm[23] , n515, \bm[21] , n476, 
        \bm[19] , \bm[18] , n478, \bm[16] , \bm[15] , \bm[14] , n511, \bm[12] , 
        \bm[11] , n463, \bm[9] , \bm[8] , \bm[7] , n471, \bm[5] , \bm[4] , 
        n465, \bm[2] , \bm[1] , n448}), .CI(1'b0), .SUM({N749, N748, N747, 
        N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, 
        N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, 
        N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, 
        N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, 
        N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, 
        N686}) );
    INV4 U812 ( .O(n819), .I(n634) );
    INV4 U813 ( .O(n820), .I(n522) );
    INV4 U814 ( .O(n821), .I(n520) );
    INV4 U815 ( .O(n823), .I(n370) );
    INV4 U816 ( .O(n824), .I(n636) );
    INV4 U817 ( .O(n825), .I(n597) );
    INV4 U818 ( .O(n826), .I(n630) );
    INV4 U819 ( .O(n827), .I(n598) );
    INV4 U820 ( .O(n828), .I(n483) );
    INV4 U821 ( .O(n829), .I(n485) );
    INV4 U822 ( .O(n831), .I(n487) );
    QDFFRBP \cnt_reg[1]  ( .Q(\cnt[1] ), .D(N6), .CK(clk), .RB(n644) );
    QDFFRBP \cnt_reg[2]  ( .Q(\cnt[2] ), .D(N7), .CK(clk), .RB(n644) );
endmodule

