// For SDF Simulation:
`timescale 1ns/10ps

module FIFOTop ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, ClkW, Reseter
 );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

// For SDF Simulation:
initial $sdf_annotate("FIFOTopNetlist.sdf");

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), .WriteReq(WriteIn), 
        .ClkR(ClkR), .ClkW(ClkW), .Reset(n1) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({n34, n33, n32, n31, 
        n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, n18, n17, 
        n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3}), 
        .AddrR(SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n2), .Write(SM_MemWriteCmd), .Reset(n1) );
  CKBXD0 U2 ( .I(Reseter), .Z(n1) );
  BUFFD1 U3 ( .I(Din[28]), .Z(n31) );
  BUFFD1 U4 ( .I(Din[30]), .Z(n33) );
  BUFFD1 U5 ( .I(Din[31]), .Z(n34) );
  BUFFD1 U6 ( .I(Din[0]), .Z(n3) );
  BUFFD1 U7 ( .I(Din[1]), .Z(n4) );
  BUFFD1 U8 ( .I(Din[2]), .Z(n5) );
  BUFFD1 U9 ( .I(Din[3]), .Z(n6) );
  BUFFD1 U10 ( .I(Din[4]), .Z(n7) );
  BUFFD1 U11 ( .I(Din[5]), .Z(n8) );
  BUFFD1 U12 ( .I(Din[6]), .Z(n9) );
  BUFFD1 U13 ( .I(Din[7]), .Z(n10) );
  BUFFD1 U14 ( .I(Din[8]), .Z(n11) );
  BUFFD1 U15 ( .I(Din[9]), .Z(n12) );
  BUFFD1 U16 ( .I(Din[10]), .Z(n13) );
  BUFFD1 U17 ( .I(Din[11]), .Z(n14) );
  BUFFD1 U18 ( .I(Din[12]), .Z(n15) );
  BUFFD1 U19 ( .I(Din[13]), .Z(n16) );
  BUFFD1 U20 ( .I(Din[14]), .Z(n17) );
  BUFFD1 U21 ( .I(Din[15]), .Z(n18) );
  BUFFD1 U22 ( .I(Din[16]), .Z(n19) );
  BUFFD1 U23 ( .I(Din[17]), .Z(n20) );
  BUFFD1 U24 ( .I(Din[18]), .Z(n21) );
  BUFFD1 U25 ( .I(Din[19]), .Z(n22) );
  BUFFD1 U26 ( .I(Din[20]), .Z(n23) );
  BUFFD1 U27 ( .I(Din[21]), .Z(n24) );
  BUFFD1 U28 ( .I(Din[22]), .Z(n25) );
  BUFFD1 U29 ( .I(Din[23]), .Z(n26) );
  BUFFD1 U30 ( .I(Din[24]), .Z(n27) );
  BUFFD1 U31 ( .I(Din[25]), .Z(n28) );
  BUFFD1 U32 ( .I(Din[26]), .Z(n29) );
  BUFFD1 U33 ( .I(Din[27]), .Z(n30) );
  BUFFD1 U34 ( .I(Din[29]), .Z(n32) );
  BUFFD1 U35 ( .I(SM_MemReadCmd), .Z(n2) );
  TIEH U36 ( .Z(\*Logic1* ) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n156, StateClockRaw, StateClock, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N169, N171, N172, N173, N321, N323, N324, N325, n73, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n107, \add_389/carry[2] , \add_389/carry[3] , \add_389/carry[4] ,
         \add_308/carry[2] , \add_308/carry[3] , \add_308/carry[4] , n1, n2,
         n18, n19, n21, n22, n24, n26, n28, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n74, n86, n88, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  assign WriteAddr[0] = N321;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n93), .CPN(StateClock), .Q(FullFIFO), .QN(n76) );
  DFND1 EmptyFIFOr_reg ( .D(n1), .CPN(StateClock), .Q(EmptyFIFO) );
  FIFOStateM_AWid5_DW01_inc_0 r151 ( .A({WriteAddr[4:1], N321}), .SUM({N70, 
        N69, N68, N67, N66}) );
  FIFOStateM_AWid5_DW01_inc_1 r150 ( .A(ReadAddr), .SUM({N47, N46, N45, N44, 
        N43}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n107), .CPN(StateClock), .CDN(n18), .QN(n89)
         );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n104), .CPN(StateClock), .CDN(n18), .QN(n87) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n97), .CPN(StateClock), .CDN(n18), .QN(n80)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n94), .CPN(StateClock), .CDN(n19), .QN(n77)
         );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n92), .CPN(StateClock), .CDN(n19), .QN(n75)
         );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n90), .CPN(StateClock), .CDN(n19), .QN(n73)
         );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n99), .CPN(StateClock), .CDN(n18), .QN(n82)
         );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n98), .CPN(StateClock), .CDN(n18), .QN(n81)
         );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n96), .CPN(StateClock), .CDN(n18), .QN(n79)
         );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n95), .CPN(StateClock), .CDN(n19), .QN(n78)
         );
  DFNCND1 \NextState_reg[1]  ( .D(n102), .CPN(StateClock), .CDN(n18), .Q(
        NextState[1]), .QN(n85) );
  DFNCND1 \NextState_reg[2]  ( .D(n101), .CPN(StateClock), .CDN(n18), .Q(
        NextState[2]), .QN(n84) );
  DFNCND1 \NextState_reg[0]  ( .D(n100), .CPN(StateClock), .CDN(n18), .Q(
        NextState[0]), .QN(n83) );
  DFNCND1 ReadCmdr_reg ( .D(n105), .CPN(StateClock), .CDN(n18), .Q(ReadCmd) );
  DFNCND1 WriteCmdr_reg ( .D(n103), .CPN(StateClock), .CDN(n18), .Q(WriteCmd)
         );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n19), 
        .Q(CurState[1]) );
  EDFCNQD1 \ReadAr_reg[3]  ( .D(N51), .E(N52), .CP(StateClock), .CDN(n19), .Q(
        n156) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n19), 
        .Q(CurState[0]) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n19), 
        .Q(CurState[2]) );
  EDFCNQD1 \ReadAr_reg[0]  ( .D(N48), .E(N52), .CP(StateClock), .CDN(n19), .Q(
        N169) );
  EDFCNQD1 \ReadAr_reg[1]  ( .D(N49), .E(N52), .CP(StateClock), .CDN(n19), .Q(
        \add_308/carry[2] ) );
  EDFCND1 \ReadAr_reg[4]  ( .D(N53), .E(N52), .CP(StateClock), .CDN(n18), .QN(
        n30) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N50), .E(N52), .CP(StateClock), .CDN(n19), .QN(
        n26) );
  EDFCND1 \WriteAr_reg[4]  ( .D(N75), .E(N76), .CP(StateClock), .CDN(n19), .Q(
        WriteAddr[4]), .QN(n31) );
  EDFCND1 \WriteAr_reg[3]  ( .D(N74), .E(N76), .CP(StateClock), .CDN(n19), .Q(
        WriteAddr[3]), .QN(n34) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N73), .E(N76), .CP(StateClock), .CDN(n18), .Q(
        WriteAddr[2]), .QN(n33) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N72), .E(N76), .CP(StateClock), .CDN(n19), .Q(
        \add_389/carry[2] ), .QN(n2) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N71), .E(N76), .CP(StateClock), .CDN(n18), .Q(
        N321), .QN(n54) );
  BUFFD0 U3 ( .I(n91), .Z(n1) );
  INVD1 U4 ( .I(Reset), .ZN(n19) );
  CKBD0 U5 ( .CLK(\add_389/carry[2] ), .C(WriteAddr[1]) );
  INVD1 U6 ( .I(N43), .ZN(n22) );
  INVD1 U7 ( .I(Reset), .ZN(n18) );
  INVD1 U8 ( .I(n21), .ZN(ReadAddr[0]) );
  INVD1 U9 ( .I(n24), .ZN(ReadAddr[1]) );
  INVD1 U10 ( .I(n28), .ZN(ReadAddr[3]) );
  INVD1 U11 ( .I(n26), .ZN(ReadAddr[2]) );
  INVD1 U12 ( .I(n30), .ZN(ReadAddr[4]) );
  INVD1 U13 ( .I(\add_308/carry[2] ), .ZN(n24) );
  INVD1 U14 ( .I(N169), .ZN(n21) );
  ND2D1 U15 ( .A1(CurState[1]), .A2(n110), .ZN(n36) );
  INVD1 U16 ( .I(n156), .ZN(n28) );
  CKXOR2D0 U17 ( .A1(ReadAddr[4]), .A2(\add_308/carry[4] ), .Z(N173) );
  AN2D0 U18 ( .A1(ReadAddr[3]), .A2(\add_308/carry[3] ), .Z(\add_308/carry[4] ) );
  CKXOR2D0 U19 ( .A1(\add_308/carry[3] ), .A2(ReadAddr[3]), .Z(N172) );
  AN2D0 U20 ( .A1(ReadAddr[2]), .A2(ReadAddr[1]), .Z(\add_308/carry[3] ) );
  CKXOR2D0 U21 ( .A1(ReadAddr[1]), .A2(ReadAddr[2]), .Z(N171) );
  CKXOR2D0 U22 ( .A1(WriteAddr[4]), .A2(\add_389/carry[4] ), .Z(N325) );
  AN2D0 U23 ( .A1(WriteAddr[3]), .A2(\add_389/carry[3] ), .Z(
        \add_389/carry[4] ) );
  CKXOR2D0 U24 ( .A1(\add_389/carry[3] ), .A2(WriteAddr[3]), .Z(N324) );
  AN2D0 U25 ( .A1(WriteAddr[2]), .A2(WriteAddr[1]), .Z(\add_389/carry[3] ) );
  CKXOR2D0 U26 ( .A1(WriteAddr[1]), .A2(WriteAddr[2]), .Z(N323) );
  MUX2ND0 U27 ( .I0(n82), .I1(n31), .S(n32), .ZN(n99) );
  MUX2ND0 U28 ( .I0(n81), .I1(n33), .S(n32), .ZN(n98) );
  MUX2ND0 U29 ( .I0(n80), .I1(n34), .S(n32), .ZN(n97) );
  MUX2ND0 U30 ( .I0(n79), .I1(n30), .S(n35), .ZN(n96) );
  MUX2ND0 U31 ( .I0(n78), .I1(n26), .S(n35), .ZN(n95) );
  MUX2ND0 U32 ( .I0(n77), .I1(n28), .S(n35), .ZN(n94) );
  OAI32D0 U33 ( .A1(n36), .A2(Reset), .A3(ReadReq), .B1(n76), .B2(n37), .ZN(
        n93) );
  AOI21D0 U34 ( .A1(n38), .A2(n39), .B(Reset), .ZN(n37) );
  MUX2ND0 U35 ( .I0(n75), .I1(n24), .S(n35), .ZN(n92) );
  OAI31D0 U36 ( .A1(n39), .A2(WriteReq), .A3(Reset), .B(n40), .ZN(n91) );
  OAI21D0 U37 ( .A1(Reset), .A2(n41), .B(EmptyFIFO), .ZN(n40) );
  MUX2ND0 U38 ( .I0(n73), .I1(n2), .S(n32), .ZN(n90) );
  MUX2ND0 U39 ( .I0(n89), .I1(n21), .S(n35), .ZN(n107) );
  INR3D0 U40 ( .A1(ReadReq), .B1(n42), .B2(n43), .ZN(n35) );
  MUX2ND0 U41 ( .I0(n44), .I1(n45), .S(n42), .ZN(n105) );
  NR2D0 U42 ( .A1(n46), .A2(n47), .ZN(n42) );
  CKND2D0 U43 ( .A1(n43), .A2(ReadReq), .ZN(n44) );
  AN3D0 U44 ( .A1(n48), .A2(n49), .A3(n50), .Z(n43) );
  NR3D0 U45 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n50) );
  CKXOR2D0 U46 ( .A1(n28), .A2(n77), .Z(n53) );
  CKXOR2D0 U47 ( .A1(n24), .A2(n75), .Z(n52) );
  CKXOR2D0 U48 ( .A1(n21), .A2(n89), .Z(n51) );
  CKXOR2D0 U49 ( .A1(n78), .A2(ReadAddr[2]), .Z(n49) );
  CKXOR2D0 U50 ( .A1(n79), .A2(ReadAddr[4]), .Z(n48) );
  MUX2ND0 U51 ( .I0(n87), .I1(n54), .S(n32), .ZN(n104) );
  NR3D0 U52 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n32) );
  MUX2ND0 U53 ( .I0(n58), .I1(n59), .S(n55), .ZN(n103) );
  NR2D0 U54 ( .A1(n46), .A2(n60), .ZN(n55) );
  CKND2D0 U55 ( .A1(n56), .A2(WriteReq), .ZN(n58) );
  AN3D0 U56 ( .A1(n61), .A2(n62), .A3(n63), .Z(n56) );
  NR3D0 U57 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n63) );
  CKXOR2D0 U58 ( .A1(n34), .A2(n80), .Z(n66) );
  CKXOR2D0 U59 ( .A1(n2), .A2(n73), .Z(n65) );
  CKXOR2D0 U60 ( .A1(n54), .A2(n87), .Z(n64) );
  CKXOR2D0 U61 ( .A1(n81), .A2(WriteAddr[2]), .Z(n62) );
  CKXOR2D0 U62 ( .A1(n82), .A2(WriteAddr[4]), .Z(n61) );
  MUX2ND0 U63 ( .I0(n67), .I1(n85), .S(n68), .ZN(n102) );
  NR2D0 U64 ( .A1(n60), .A2(n69), .ZN(n67) );
  MUX2ND0 U65 ( .I0(n70), .I1(n71), .S(CurState[1]), .ZN(n69) );
  OAI21D0 U66 ( .A1(n72), .A2(n74), .B(n86), .ZN(n71) );
  AOI31D0 U67 ( .A1(n88), .A2(n106), .A3(n108), .B(CurState[2]), .ZN(n86) );
  OAI21D0 U68 ( .A1(n108), .A2(n109), .B(n110), .ZN(n70) );
  CKND0 U69 ( .CLK(n111), .CN(n109) );
  AN3D0 U70 ( .A1(n112), .A2(n113), .A3(n114), .Z(n108) );
  NR3D0 U71 ( .A1(n115), .A2(n116), .A3(n117), .ZN(n114) );
  CKXOR2D0 U72 ( .A1(WriteAddr[3]), .A2(ReadAddr[3]), .Z(n117) );
  CKXOR2D0 U73 ( .A1(WriteAddr[1]), .A2(ReadAddr[1]), .Z(n116) );
  CKXOR2D0 U74 ( .A1(N321), .A2(ReadAddr[0]), .Z(n115) );
  CKXOR2D0 U75 ( .A1(ReadAddr[2]), .A2(n33), .Z(n113) );
  CKXOR2D0 U76 ( .A1(ReadAddr[4]), .A2(n31), .Z(n112) );
  MUX2ND0 U77 ( .I0(n118), .I1(n84), .S(n68), .ZN(n101) );
  AOI211D0 U78 ( .A1(n110), .A2(n111), .B(n47), .C(n119), .ZN(n118) );
  NR3D0 U79 ( .A1(n74), .A2(n120), .A3(n72), .ZN(n119) );
  ND3D0 U80 ( .A1(n121), .A2(n122), .A3(n123), .ZN(n74) );
  NR3D0 U81 ( .A1(n124), .A2(n125), .A3(n126), .ZN(n123) );
  CKXOR2D0 U82 ( .A1(ReadAddr[3]), .A2(N69), .Z(n126) );
  CKXOR2D0 U83 ( .A1(ReadAddr[1]), .A2(N67), .Z(n125) );
  CKXOR2D0 U84 ( .A1(ReadAddr[0]), .A2(N66), .Z(n124) );
  CKXOR2D0 U85 ( .A1(ReadAddr[2]), .A2(n127), .Z(n122) );
  CKXOR2D0 U86 ( .A1(ReadAddr[4]), .A2(n128), .Z(n121) );
  CKND0 U87 ( .CLK(n36), .CN(n47) );
  ND3D0 U88 ( .A1(n129), .A2(n130), .A3(n131), .ZN(n111) );
  NR3D0 U89 ( .A1(n132), .A2(n133), .A3(n134), .ZN(n131) );
  CKXOR2D0 U90 ( .A1(ReadAddr[3]), .A2(N324), .Z(n134) );
  CKXOR2D0 U91 ( .A1(ReadAddr[1]), .A2(n2), .Z(n133) );
  CKXOR2D0 U92 ( .A1(ReadAddr[0]), .A2(N321), .Z(n132) );
  CKXOR2D0 U93 ( .A1(N323), .A2(n26), .Z(n130) );
  CKXOR2D0 U94 ( .A1(N325), .A2(n30), .Z(n129) );
  MUX2ND0 U95 ( .I0(n135), .I1(n83), .S(n68), .ZN(n100) );
  OA211D0 U96 ( .A1(n57), .A2(n39), .B(n136), .C(n137), .Z(n68) );
  AOI21D0 U97 ( .A1(CurState[0]), .A2(n120), .B(n46), .ZN(n137) );
  MUX2ND0 U98 ( .I0(CurState[2]), .I1(n38), .S(n120), .ZN(n46) );
  CKND0 U99 ( .CLK(CurState[1]), .CN(n120) );
  OAI21D0 U100 ( .A1(ReadReq), .A2(n106), .B(CurState[2]), .ZN(n136) );
  CKND0 U101 ( .CLK(WriteReq), .CN(n57) );
  AOI21D0 U102 ( .A1(CurState[1]), .A2(n138), .B(n110), .ZN(n135) );
  OAI21D0 U103 ( .A1(n41), .A2(n88), .B(n72), .ZN(n138) );
  OAI31D0 U104 ( .A1(n139), .A2(n140), .A3(n141), .B(CurState[0]), .ZN(n72) );
  CKXOR2D0 U105 ( .A1(WriteAddr[4]), .A2(N47), .Z(n141) );
  CKXOR2D0 U106 ( .A1(WriteAddr[2]), .A2(N45), .Z(n140) );
  ND3D0 U107 ( .A1(n142), .A2(n143), .A3(n144), .ZN(n139) );
  CKXOR2D0 U108 ( .A1(N321), .A2(n22), .Z(n144) );
  CKXOR2D0 U109 ( .A1(WriteAddr[1]), .A2(n145), .Z(n143) );
  CKXOR2D0 U110 ( .A1(WriteAddr[3]), .A2(n146), .Z(n142) );
  ND3D0 U111 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n88) );
  NR3D0 U112 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n149) );
  CKXOR2D0 U113 ( .A1(WriteAddr[3]), .A2(N172), .Z(n152) );
  CKXOR2D0 U114 ( .A1(WriteAddr[1]), .A2(n24), .Z(n151) );
  CKXOR2D0 U115 ( .A1(N321), .A2(ReadAddr[0]), .Z(n150) );
  CKXOR2D0 U116 ( .A1(N171), .A2(n33), .Z(n148) );
  CKXOR2D0 U117 ( .A1(N173), .A2(n31), .Z(n147) );
  CKND2D0 U118 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  ND3D0 U119 ( .A1(n36), .A2(n39), .A3(n59), .ZN(N76) );
  OAI22D0 U120 ( .A1(n30), .A2(n36), .B1(n59), .B2(n128), .ZN(N75) );
  CKND0 U121 ( .CLK(N70), .CN(n128) );
  OAI22D0 U122 ( .A1(n28), .A2(n36), .B1(n59), .B2(n153), .ZN(N74) );
  CKND0 U123 ( .CLK(N69), .CN(n153) );
  OAI22D0 U124 ( .A1(n26), .A2(n36), .B1(n59), .B2(n127), .ZN(N73) );
  CKND0 U125 ( .CLK(N68), .CN(n127) );
  OAI22D0 U126 ( .A1(n24), .A2(n36), .B1(n59), .B2(n154), .ZN(N72) );
  CKND0 U127 ( .CLK(N67), .CN(n154) );
  OAI22D0 U128 ( .A1(n21), .A2(n36), .B1(n59), .B2(n155), .ZN(N71) );
  CKND0 U129 ( .CLK(N66), .CN(n155) );
  CKND2D0 U130 ( .A1(WriteCmd), .A2(n36), .ZN(n59) );
  CKND0 U131 ( .CLK(n38), .CN(n110) );
  CKND2D0 U132 ( .A1(CurState[2]), .A2(CurState[0]), .ZN(n38) );
  INR2D0 U133 ( .A1(N47), .B1(n45), .ZN(N53) );
  CKND2D0 U134 ( .A1(n39), .A2(n45), .ZN(N52) );
  NR2D0 U135 ( .A1(n45), .A2(n146), .ZN(N51) );
  CKND0 U136 ( .CLK(N46), .CN(n146) );
  INR2D0 U137 ( .A1(N45), .B1(n45), .ZN(N50) );
  NR2D0 U138 ( .A1(n45), .A2(n145), .ZN(N49) );
  CKND0 U139 ( .CLK(N44), .CN(n145) );
  NR2D0 U140 ( .A1(n45), .A2(n22), .ZN(N48) );
  CKND2D0 U141 ( .A1(ReadCmd), .A2(n39), .ZN(n45) );
  CKND0 U142 ( .CLK(n60), .CN(n39) );
  NR2D0 U143 ( .A1(n41), .A2(CurState[1]), .ZN(n60) );
  IND2D0 U144 ( .A1(CurState[2]), .B1(n106), .ZN(n41) );
  CKND0 U145 ( .CLK(CurState[0]), .CN(n106) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, ClockR, ClockW, Dreadyr, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N85, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n107,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  BUFTD1 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD1 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD1 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD1 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD1 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD1 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD1 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD1 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD1 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD1 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD1 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD1 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD1 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD1 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD1 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD1 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD1 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD1 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD1 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD1 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD1 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD1 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD1 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD1 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD1 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD1 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD1 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD1 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD1 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD1 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD1 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD1 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  XNR4D1 U18 ( .A1(n992), .A2(n989), .A3(n998), .A4(n995), .ZN(n84) );
  XOR4D1 U19 ( .A1(n1004), .A2(n1001), .A3(n1010), .A4(n1007), .Z(n83) );
  XOR4D1 U20 ( .A1(n980), .A2(n977), .A3(n986), .A4(n983), .Z(n80) );
  XOR4D1 U21 ( .A1(n959), .A2(n956), .A3(n965), .A4(n962), .Z(n77) );
  XNR4D1 U22 ( .A1(n938), .A2(n935), .A3(n944), .A4(n941), .ZN(n74) );
  XOR4D1 U27 ( .A1(n90), .A2(N72), .A3(n91), .A4(N75), .Z(n89) );
  XNR4D1 U28 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n91) );
  XNR4D1 U33 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n97) );
  XOR4D1 U34 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n96) );
  XNR4D1 U35 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .ZN(n93) );
  XNR4D1 U36 ( .A1(N80), .A2(N78), .A3(N82), .A4(N81), .ZN(n87) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(n718), .E(n663), .CP(n751), .CDN(n614), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(n1010), .E(n663), .CP(n751), .CDN(n613), 
        .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(n1008), .E(n662), .CP(n751), .CDN(n613), 
        .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(n1005), .E(n663), .CP(n751), .CDN(n613), 
        .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(n1001), .E(n662), .CP(n751), .CDN(n613), 
        .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(n998), .E(n663), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(n996), .E(n662), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(n993), .E(n663), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(n989), .E(n662), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(n986), .E(n663), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n984), .E(n662), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(n981), .E(n662), .CP(n752), .CDN(n613), 
        .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(n977), .E(n662), .CP(n752), .CDN(n612), 
        .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(n975), .E(n662), .CP(n752), .CDN(n612), 
        .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(n972), .E(n662), .CP(n752), .CDN(n612), 
        .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(n969), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(n965), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n963), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n960), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(n956), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n954), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(n951), .E(n662), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(n948), .E(n663), .CP(n753), .CDN(n612), 
        .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n944), .E(n663), .CP(n753), .CDN(n636), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(n942), .E(n663), .CP(n753), .CDN(n611), 
        .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n939), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n935), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n933), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n930), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(n927), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n924), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(n921), .E(n663), .CP(n754), .CDN(n612), 
        .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n918), .E(n663), .CP(n754), .CDN(n611), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(n718), .E(n667), .CP(n758), .CDN(n609), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(n1011), .E(n667), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(n1008), .E(n666), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(n1005), .E(n667), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(n1002), .E(n666), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(n999), .E(n667), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(n996), .E(n666), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(n993), .E(n667), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(n990), .E(n666), .CP(n758), .CDN(n608), 
        .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(n987), .E(n667), .CP(n759), .CDN(n608), 
        .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n984), .E(n666), .CP(n759), .CDN(n608), 
        .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(n981), .E(n666), .CP(n759), .CDN(n608), 
        .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(n978), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(n975), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(n972), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(n969), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(n966), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n963), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n960), .E(n666), .CP(n759), .CDN(n607), 
        .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(n957), .E(n666), .CP(n760), .CDN(n607), 
        .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n954), .E(n666), .CP(n760), .CDN(n607), 
        .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(n951), .E(n666), .CP(n760), .CDN(n607), 
        .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(n948), .E(n667), .CP(n760), .CDN(n607), 
        .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n945), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(n942), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n939), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n936), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n933), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n930), .E(n667), .CP(n760), .CDN(n606), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(n927), .E(n667), .CP(n761), .CDN(n606), 
        .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n924), .E(n667), .CP(n761), .CDN(n606), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(n921), .E(n667), .CP(n761), .CDN(n606), 
        .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n918), .E(n667), .CP(n761), .CDN(n606), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(n718), .E(n655), .CP(n738), .CDN(n624), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(n1011), .E(n655), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(n1008), .E(n654), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(n1005), .E(n655), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(n1002), .E(n654), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(n999), .E(n655), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(n990), .E(n654), .CP(n739), .CDN(n623), 
        .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(n987), .E(n655), .CP(n739), .CDN(n623), 
        .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(n984), .E(n654), .CP(n739), .CDN(n623), 
        .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(n981), .E(n654), .CP(n739), .CDN(n623), 
        .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(n978), .E(n654), .CP(n739), .CDN(n622), 
        .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(n975), .E(n654), .CP(n739), .CDN(n622), 
        .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(n972), .E(n654), .CP(n739), .CDN(n622), 
        .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(n969), .E(n654), .CP(n739), .CDN(n622), 
        .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(n966), .E(n654), .CP(n739), .CDN(n622), 
        .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(n963), .E(n654), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(n960), .E(n654), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(n957), .E(n654), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(n954), .E(n654), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(n951), .E(n654), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(n948), .E(n655), .CP(n740), .CDN(n622), 
        .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(n945), .E(n655), .CP(n740), .CDN(n635), 
        .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(n942), .E(n655), .CP(n740), .CDN(n630), 
        .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(n939), .E(n655), .CP(n740), .CDN(n621), 
        .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n936), .E(n655), .CP(n740), .CDN(n634), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(n933), .E(n655), .CP(n741), .CDN(n650), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(n930), .E(n655), .CP(n741), .CDN(n641), 
        .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(n927), .E(n655), .CP(n741), .CDN(n630), 
        .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(n924), .E(n655), .CP(n741), .CDN(n650), 
        .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(n921), .E(n655), .CP(n741), .CDN(n621), 
        .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(n918), .E(n655), .CP(n741), .CDN(n630), 
        .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n718), .E(n657), .CP(n741), .CDN(n580), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(n1011), .E(n657), .CP(n741), .CDN(n622), 
        .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(n1008), .E(n656), .CP(n741), .CDN(n641), 
        .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(n1005), .E(n657), .CP(n741), .CDN(n622), 
        .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(n1002), .E(n656), .CP(n742), .CDN(n622), 
        .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(n999), .E(n657), .CP(n742), .CDN(n622), 
        .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(n990), .E(n656), .CP(n742), .CDN(n622), 
        .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(n987), .E(n657), .CP(n742), .CDN(n622), 
        .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(n984), .E(n656), .CP(n742), .CDN(n621), 
        .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(n981), .E(n656), .CP(n742), .CDN(n622), 
        .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(n978), .E(n656), .CP(n742), .CDN(n621), 
        .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(n975), .E(n656), .CP(n742), .CDN(n621), 
        .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(n972), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(n969), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(n966), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(n963), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(n960), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(n957), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(n954), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(n951), .E(n656), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(n948), .E(n657), .CP(n743), .CDN(n621), 
        .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(n945), .E(n657), .CP(n743), .CDN(n620), 
        .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(n942), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(n939), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(n936), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(n933), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(n930), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(n927), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(n924), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(n921), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(n918), .E(n657), .CP(n744), .CDN(n620), 
        .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(n718), .E(n659), .CP(n744), .CDN(n620), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(n1011), .E(n659), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(n1008), .E(n658), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(n1005), .E(n659), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(n1002), .E(n658), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(n990), .E(n659), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(n987), .E(n658), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n984), .E(n659), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(n981), .E(n658), .CP(n746), .CDN(n619), 
        .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(n978), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(n975), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(n972), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(n969), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(n966), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(n963), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(n960), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(n957), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n954), .E(n658), .CP(n746), .CDN(n618), 
        .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(n951), .E(n658), .CP(n747), .CDN(n618), 
        .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(n948), .E(n659), .CP(n747), .CDN(n618), 
        .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n945), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(n942), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(n939), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n936), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n933), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n930), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(n927), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n924), .E(n659), .CP(n747), .CDN(n617), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(n921), .E(n659), .CP(n748), .CDN(n617), 
        .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n918), .E(n659), .CP(n748), .CDN(n617), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n718), .E(n661), .CP(n748), .CDN(n617), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(n1011), .E(n661), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(n1008), .E(n660), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(n1005), .E(n661), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(n1002), .E(n660), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(n999), .E(n661), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(n996), .E(n660), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(n993), .E(n661), .CP(n748), .CDN(n616), 
        .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(n990), .E(n660), .CP(n749), .CDN(n616), 
        .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(n987), .E(n661), .CP(n749), .CDN(n616), 
        .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n984), .E(n660), .CP(n749), .CDN(n616), 
        .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(n981), .E(n660), .CP(n749), .CDN(n616), 
        .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(n978), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(n975), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(n972), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(n969), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(n966), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n963), .E(n660), .CP(n749), .CDN(n615), 
        .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n960), .E(n660), .CP(n750), .CDN(n615), 
        .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(n957), .E(n660), .CP(n750), .CDN(n615), 
        .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n954), .E(n660), .CP(n750), .CDN(n615), 
        .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(n951), .E(n660), .CP(n750), .CDN(n615), 
        .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(n948), .E(n661), .CP(n750), .CDN(n615), 
        .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n945), .E(n661), .CP(n750), .CDN(n614), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(n942), .E(n661), .CP(n750), .CDN(n614), 
        .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n939), .E(n661), .CP(n750), .CDN(n614), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n936), .E(n661), .CP(n750), .CDN(n614), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n933), .E(n661), .CP(n750), .CDN(n614), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n930), .E(n661), .CP(n751), .CDN(n614), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(n927), .E(n661), .CP(n751), .CDN(n614), 
        .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n924), .E(n661), .CP(n751), .CDN(n614), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(n921), .E(n661), .CP(n751), .CDN(n614), 
        .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n918), .E(n661), .CP(n751), .CDN(n614), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n718), .E(n665), .CP(n754), .CDN(n610), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(n1011), .E(n665), .CP(n754), .CDN(n611), 
        .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(n1008), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(n1005), .E(n665), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(n1002), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(n999), .E(n665), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(n996), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(n993), .E(n665), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(n990), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(n987), .E(n665), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n984), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(n981), .E(n664), .CP(n755), .CDN(n611), 
        .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(n978), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(n975), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(n972), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(n969), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(n966), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(n963), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(n960), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(n957), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n954), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(n951), .E(n664), .CP(n756), .CDN(n610), 
        .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(n948), .E(n665), .CP(n757), .CDN(n610), 
        .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n945), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(n942), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(n939), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n936), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n933), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n930), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(n927), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n924), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(n921), .E(n665), .CP(n757), .CDN(n609), 
        .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n918), .E(n665), .CP(n758), .CDN(n609), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(n718), .E(n671), .CP(n764), .CDN(n604), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n1011), .E(n671), .CP(n764), .CDN(n603), 
        .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n1008), .E(n670), .CP(n764), .CDN(n603), 
        .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(n1005), .E(n671), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(n1002), .E(n670), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(n999), .E(n671), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n996), .E(n670), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(n993), .E(n671), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(n990), .E(n670), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(n987), .E(n671), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(n984), .E(n670), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(n981), .E(n670), .CP(n765), .CDN(n603), 
        .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(n978), .E(n670), .CP(n765), .CDN(n626), 
        .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(n975), .E(n670), .CP(n766), .CDN(n600), 
        .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(n972), .E(n670), .CP(n766), .CDN(n601), 
        .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n969), .E(n670), .CP(n766), .CDN(n602), 
        .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(n966), .E(n670), .CP(n766), .CDN(n635), 
        .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(n963), .E(n670), .CP(n766), .CDN(n618), 
        .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(n960), .E(n670), .CP(n766), .CDN(n617), 
        .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n957), .E(n670), .CP(n766), .CDN(n575), 
        .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(n954), .E(n670), .CP(n766), .CDN(n623), 
        .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(n951), .E(n670), .CP(n766), .CDN(n624), 
        .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(n948), .E(n671), .CP(n766), .CDN(n625), 
        .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(n945), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(n942), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(n939), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n936), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n933), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(n930), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(n927), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(n924), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(n921), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n918), .E(n671), .CP(n767), .CDN(n602), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(n719), .E(n673), .CP(n768), .CDN(n602), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n1011), .E(n673), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n1008), .E(n672), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n1005), .E(n673), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n1002), .E(n672), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(n999), .E(n673), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n996), .E(n672), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n993), .E(n673), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n990), .E(n672), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(n987), .E(n673), .CP(n768), .CDN(n601), 
        .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n984), .E(n672), .CP(n769), .CDN(n601), 
        .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n981), .E(n672), .CP(n769), .CDN(n601), 
        .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n978), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n974), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(n972), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n969), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n966), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n963), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n960), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n957), .E(n672), .CP(n769), .CDN(n600), 
        .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n953), .E(n672), .CP(n770), .CDN(n600), 
        .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n951), .E(n672), .CP(n770), .CDN(n600), 
        .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n948), .E(n673), .CP(n770), .CDN(n600), 
        .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n945), .E(n673), .CP(n770), .CDN(n630), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n942), .E(n673), .CP(n770), .CDN(n636), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n939), .E(n673), .CP(n770), .CDN(n639), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n936), .E(n673), .CP(n770), .CDN(n630), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n932), .E(n673), .CP(n770), .CDN(n638), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n930), .E(n673), .CP(n770), .CDN(n631), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(n927), .E(n673), .CP(n770), .CDN(n632), 
        .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n923), .E(n673), .CP(n771), .CDN(n636), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n921), .E(n673), .CP(n771), .CDN(n651), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n917), .E(n673), .CP(n771), .CDN(n630), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(n719), .E(n679), .CP(n777), .CDN(n596), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(n1011), .E(n679), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(n1008), .E(n678), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(n1005), .E(n679), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(n1002), .E(n678), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(n999), .E(n679), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(n996), .E(n678), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(n993), .E(n679), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(n990), .E(n678), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(n987), .E(n679), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n984), .E(n678), .CP(n778), .CDN(n595), 
        .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(n981), .E(n678), .CP(n779), .CDN(n595), 
        .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(n978), .E(n678), .CP(n779), .CDN(n622), 
        .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(n974), .E(n678), .CP(n779), .CDN(n592), 
        .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(n972), .E(n678), .CP(n779), .CDN(n593), 
        .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(n969), .E(n678), .CP(n779), .CDN(n594), 
        .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(n966), .E(n678), .CP(n779), .CDN(n637), 
        .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(n963), .E(n678), .CP(n779), .CDN(n549), 
        .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(n960), .E(n678), .CP(n779), .CDN(n644), 
        .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n957), .E(n678), .CP(n779), .CDN(n643), 
        .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n953), .E(n678), .CP(n779), .CDN(n647), 
        .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(n951), .E(n678), .CP(n780), .CDN(n613), 
        .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(n948), .E(n679), .CP(n780), .CDN(n614), 
        .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n945), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(n942), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(n939), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n936), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n932), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n930), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(n927), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n923), .E(n679), .CP(n780), .CDN(n594), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(n921), .E(n679), .CP(n781), .CDN(n594), 
        .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n917), .E(n679), .CP(n781), .CDN(n594), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n719), .E(n681), .CP(n781), .CDN(n594), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n1011), .E(n681), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n1008), .E(n680), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(n1005), .E(n681), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(n1002), .E(n680), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n999), .E(n681), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n996), .E(n680), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(n993), .E(n681), .CP(n781), .CDN(n593), 
        .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(n990), .E(n680), .CP(n782), .CDN(n593), 
        .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n987), .E(n681), .CP(n782), .CDN(n593), 
        .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n984), .E(n680), .CP(n782), .CDN(n593), 
        .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(n981), .E(n680), .CP(n782), .CDN(n593), 
        .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(n978), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(n974), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n972), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n969), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(n966), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(n963), .E(n680), .CP(n782), .CDN(n592), 
        .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(n960), .E(n680), .CP(n783), .CDN(n592), 
        .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n957), .E(n680), .CP(n783), .CDN(n592), 
        .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n953), .E(n680), .CP(n783), .CDN(n592), 
        .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(n951), .E(n680), .CP(n783), .CDN(n592), 
        .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(n948), .E(n681), .CP(n783), .CDN(n592), 
        .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n945), .E(n681), .CP(n783), .CDN(n572), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(n942), .E(n681), .CP(n783), .CDN(n639), 
        .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(n939), .E(n681), .CP(n783), .CDN(n573), 
        .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n936), .E(n681), .CP(n783), .CDN(n626), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n932), .E(n681), .CP(n783), .CDN(n627), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n930), .E(n681), .CP(n784), .CDN(n574), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n927), .E(n681), .CP(n784), .CDN(n650), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n923), .E(n681), .CP(n784), .CDN(n599), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(n921), .E(n681), .CP(n784), .CDN(n575), 
        .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n917), .E(n681), .CP(n784), .CDN(n615), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n719), .E(n687), .CP(n791), .CDN(n590), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n1011), .E(n687), .CP(n791), .CDN(n587), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n1008), .E(n686), .CP(n791), .CDN(n581), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n1005), .E(n687), .CP(n791), .CDN(n587), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n1002), .E(n686), .CP(n791), .CDN(n581), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n999), .E(n687), .CP(n791), .CDN(n587), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n996), .E(n686), .CP(n791), .CDN(n581), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n993), .E(n687), .CP(n791), .CDN(n587), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n990), .E(n686), .CP(n791), .CDN(n581), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n987), .E(n687), .CP(n792), .CDN(n587), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n984), .E(n686), .CP(n792), .CDN(n581), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n981), .E(n686), .CP(n792), .CDN(n587), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n978), .E(n686), .CP(n792), .CDN(n574), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n974), .E(n686), .CP(n792), .CDN(n581), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n972), .E(n686), .CP(n792), .CDN(n589), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n969), .E(n686), .CP(n792), .CDN(n587), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n966), .E(n686), .CP(n792), .CDN(n572), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n963), .E(n686), .CP(n792), .CDN(n627), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n960), .E(n686), .CP(n792), .CDN(n624), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n957), .E(n686), .CP(n793), .CDN(n625), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n953), .E(n686), .CP(n793), .CDN(n626), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n951), .E(n686), .CP(n793), .CDN(n623), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n948), .E(n687), .CP(n793), .CDN(n580), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n945), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n942), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n939), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n936), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n932), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n930), .E(n687), .CP(n793), .CDN(n589), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n927), .E(n687), .CP(n794), .CDN(n589), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n923), .E(n687), .CP(n794), .CDN(n589), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n921), .E(n687), .CP(n794), .CDN(n589), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n917), .E(n687), .CP(n794), .CDN(n589), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n719), .E(n689), .CP(n794), .CDN(n589), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n1011), .E(n689), .CP(n794), .CDN(n588), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n1008), .E(n688), .CP(n794), .CDN(n588), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n1005), .E(n689), .CP(n794), .CDN(n588), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n1002), .E(n688), .CP(n794), .CDN(n588), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n999), .E(n689), .CP(n794), .CDN(n588), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n996), .E(n688), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n993), .E(n689), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n990), .E(n688), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n987), .E(n689), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n984), .E(n688), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n981), .E(n688), .CP(n795), .CDN(n588), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n978), .E(n688), .CP(n795), .CDN(n587), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n974), .E(n688), .CP(n795), .CDN(n587), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n972), .E(n688), .CP(n795), .CDN(n587), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n969), .E(n688), .CP(n795), .CDN(n587), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n966), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n963), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n960), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n957), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n953), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n951), .E(n688), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n948), .E(n689), .CP(n796), .CDN(n587), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n945), .E(n689), .CP(n796), .CDN(n586), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n942), .E(n689), .CP(n796), .CDN(n586), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n939), .E(n689), .CP(n796), .CDN(n586), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n936), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n932), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n930), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n927), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n923), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n921), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n917), .E(n689), .CP(n797), .CDN(n586), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(n720), .E(n695), .CP(n804), .CDN(n581), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n1010), .E(n695), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n1007), .E(n694), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n1004), .E(n695), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n1001), .E(n694), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n998), .E(n695), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n995), .E(n694), .CP(n804), .CDN(n580), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n992), .E(n695), .CP(n805), .CDN(n580), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n989), .E(n694), .CP(n805), .CDN(n580), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n986), .E(n695), .CP(n805), .CDN(n580), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n983), .E(n694), .CP(n805), .CDN(n580), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n980), .E(n694), .CP(n805), .CDN(n580), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n977), .E(n694), .CP(n805), .CDN(n579), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n974), .E(n694), .CP(n805), .CDN(n579), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n971), .E(n694), .CP(n805), .CDN(n579), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n968), .E(n694), .CP(n805), .CDN(n579), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n965), .E(n694), .CP(n805), .CDN(n579), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n962), .E(n694), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n959), .E(n694), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n956), .E(n694), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n953), .E(n694), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n950), .E(n694), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n947), .E(n695), .CP(n806), .CDN(n579), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n944), .E(n695), .CP(n806), .CDN(n578), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n941), .E(n695), .CP(n806), .CDN(n578), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n938), .E(n695), .CP(n806), .CDN(n578), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n935), .E(n695), .CP(n806), .CDN(n578), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n932), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n929), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n926), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n923), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n920), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n917), .E(n695), .CP(n807), .CDN(n578), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n720), .E(n697), .CP(n807), .CDN(n578), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n1010), .E(n697), .CP(n807), .CDN(n577), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n1007), .E(n696), .CP(n807), .CDN(n577), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n1004), .E(n697), .CP(n807), .CDN(n577), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n1001), .E(n696), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n998), .E(n697), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n995), .E(n696), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n992), .E(n697), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n989), .E(n696), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n986), .E(n697), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n983), .E(n696), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n980), .E(n696), .CP(n808), .CDN(n577), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n977), .E(n696), .CP(n808), .CDN(n576), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n974), .E(n696), .CP(n808), .CDN(n576), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n971), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n968), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n965), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n962), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n959), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n956), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n953), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n950), .E(n696), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n947), .E(n697), .CP(n809), .CDN(n576), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n944), .E(n697), .CP(n809), .CDN(n575), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n941), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n938), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n935), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n933), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n929), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n926), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n923), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n920), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n917), .E(n697), .CP(n810), .CDN(n575), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n720), .E(n703), .CP(n817), .CDN(n569), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n1010), .E(n703), .CP(n817), .CDN(n568), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n1007), .E(n702), .CP(n817), .CDN(n568), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n1004), .E(n703), .CP(n817), .CDN(n568), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n1001), .E(n702), .CP(n817), .CDN(n568), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n998), .E(n703), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n995), .E(n702), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n992), .E(n703), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n989), .E(n702), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n986), .E(n703), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n983), .E(n702), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n980), .E(n702), .CP(n818), .CDN(n568), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n977), .E(n702), .CP(n818), .CDN(n567), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n975), .E(n702), .CP(n818), .CDN(n567), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n971), .E(n702), .CP(n818), .CDN(n567), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n968), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n965), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n962), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n959), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n956), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n954), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n950), .E(n702), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n947), .E(n703), .CP(n819), .CDN(n567), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n944), .E(n703), .CP(n819), .CDN(n566), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n941), .E(n703), .CP(n819), .CDN(n566), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n938), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n935), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n932), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n929), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n926), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n924), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n920), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n918), .E(n703), .CP(n820), .CDN(n566), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n720), .E(n705), .CP(n820), .CDN(n566), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n1010), .E(n705), .CP(n820), .CDN(n565), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n1007), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n1004), .E(n705), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n1001), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n998), .E(n705), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n995), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n992), .E(n705), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n989), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n986), .E(n705), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n983), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n980), .E(n704), .CP(n821), .CDN(n565), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n977), .E(n704), .CP(n822), .CDN(n633), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n974), .E(n704), .CP(n822), .CDN(n621), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n971), .E(n704), .CP(n822), .CDN(n646), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n968), .E(n704), .CP(n822), .CDN(n568), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n965), .E(n704), .CP(n822), .CDN(n570), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n962), .E(n704), .CP(n822), .CDN(n569), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n959), .E(n704), .CP(n822), .CDN(n571), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n956), .E(n704), .CP(n822), .CDN(n606), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n953), .E(n704), .CP(n822), .CDN(n607), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n950), .E(n704), .CP(n822), .CDN(n608), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n947), .E(n705), .CP(n823), .CDN(n609), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n944), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n941), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n938), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n935), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n932), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n929), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n926), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n923), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n920), .E(n705), .CP(n823), .CDN(n564), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n917), .E(n705), .CP(n824), .CDN(n564), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(n720), .E(n711), .CP(n830), .CDN(n558), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n1010), .E(n711), .CP(n830), .CDN(n557), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n1007), .E(n710), .CP(n830), .CDN(n557), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n1004), .E(n711), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n1001), .E(n710), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n998), .E(n711), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n995), .E(n710), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n992), .E(n711), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n989), .E(n710), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n986), .E(n711), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n983), .E(n710), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n980), .E(n710), .CP(n831), .CDN(n557), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n977), .E(n710), .CP(n831), .CDN(n556), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n974), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n971), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n968), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n965), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n962), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n959), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n956), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n953), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n950), .E(n710), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n947), .E(n711), .CP(n832), .CDN(n556), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n944), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n941), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n938), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n935), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n933), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n929), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n926), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n923), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n920), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n917), .E(n711), .CP(n833), .CDN(n555), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n720), .E(n712), .CP(n834), .CDN(n555), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n1010), .E(n712), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n1007), .E(n713), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n1004), .E(n712), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n1001), .E(n713), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n998), .E(n712), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n995), .E(n713), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n992), .E(n712), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n989), .E(n713), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n986), .E(n712), .CP(n834), .CDN(n554), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n983), .E(n713), .CP(n835), .CDN(n554), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n980), .E(n712), .CP(n835), .CDN(n554), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n977), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n975), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n971), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n968), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n965), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n962), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n959), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n956), .E(n712), .CP(n835), .CDN(n553), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n954), .E(n712), .CP(n836), .CDN(n553), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n950), .E(n712), .CP(n836), .CDN(n553), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n947), .E(n713), .CP(n836), .CDN(n553), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n944), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n941), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n938), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n935), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n932), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n929), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n926), .E(n713), .CP(n836), .CDN(n552), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n923), .E(n713), .CP(n837), .CDN(n552), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n920), .E(n713), .CP(n837), .CDN(n552), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n917), .E(n713), .CP(n837), .CDN(n552), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n718), .E(n669), .CP(n761), .CDN(n606), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(n1011), .E(n669), .CP(n761), .CDN(n605), 
        .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(n1008), .E(n668), .CP(n761), .CDN(n605), 
        .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(n1005), .E(n669), .CP(n761), .CDN(n605), 
        .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(n1002), .E(n668), .CP(n761), .CDN(n605), 
        .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(n999), .E(n669), .CP(n761), .CDN(n605), 
        .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(n996), .E(n668), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(n993), .E(n669), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(n990), .E(n668), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(n987), .E(n669), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n984), .E(n668), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(n981), .E(n668), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(n978), .E(n668), .CP(n762), .CDN(n621), 
        .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(n975), .E(n668), .CP(n762), .CDN(n605), 
        .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(n972), .E(n668), .CP(n762), .CDN(n603), 
        .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(n969), .E(n668), .CP(n762), .CDN(n604), 
        .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(n966), .E(n668), .CP(n763), .CDN(n634), 
        .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(n963), .E(n668), .CP(n763), .CDN(n565), 
        .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(n960), .E(n668), .CP(n763), .CDN(n624), 
        .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n957), .E(n668), .CP(n763), .CDN(n619), 
        .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n954), .E(n668), .CP(n763), .CDN(n620), 
        .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(n951), .E(n668), .CP(n763), .CDN(n621), 
        .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(n948), .E(n669), .CP(n763), .CDN(n624), 
        .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n945), .E(n669), .CP(n763), .CDN(n604), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(n942), .E(n669), .CP(n763), .CDN(n604), 
        .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(n939), .E(n669), .CP(n763), .CDN(n604), 
        .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n936), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n933), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n930), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(n927), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n924), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(n921), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n918), .E(n669), .CP(n764), .CDN(n604), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(n719), .E(n675), .CP(n771), .CDN(n651), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(n1011), .E(n675), .CP(n771), .CDN(n586), 
        .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(n1008), .E(n674), .CP(n771), .CDN(n621), 
        .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(n1005), .E(n675), .CP(n771), .CDN(n599), 
        .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(n1002), .E(n674), .CP(n771), .CDN(n630), 
        .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(n999), .E(n675), .CP(n771), .CDN(n582), 
        .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(n996), .E(n674), .CP(n771), .CDN(n591), 
        .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(n993), .E(n675), .CP(n772), .CDN(n621), 
        .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(n990), .E(n674), .CP(n772), .CDN(n588), 
        .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(n987), .E(n675), .CP(n772), .CDN(n631), 
        .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n984), .E(n674), .CP(n772), .CDN(n583), 
        .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(n981), .E(n674), .CP(n772), .CDN(n584), 
        .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(n978), .E(n674), .CP(n772), .CDN(n599), 
        .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(n974), .E(n674), .CP(n772), .CDN(n599), 
        .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(n972), .E(n674), .CP(n772), .CDN(n599), 
        .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(n969), .E(n674), .CP(n772), .CDN(n599), 
        .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(n966), .E(n674), .CP(n772), .CDN(n599), 
        .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(n963), .E(n674), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(n960), .E(n674), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(n957), .E(n674), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n953), .E(n674), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(n951), .E(n674), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(n948), .E(n675), .CP(n773), .CDN(n599), 
        .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n945), .E(n675), .CP(n773), .CDN(n581), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(n942), .E(n675), .CP(n773), .CDN(n631), 
        .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(n939), .E(n675), .CP(n773), .CDN(n632), 
        .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n936), .E(n675), .CP(n773), .CDN(n636), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n932), .E(n675), .CP(n774), .CDN(n638), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n930), .E(n675), .CP(n774), .CDN(n651), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(n927), .E(n675), .CP(n774), .CDN(n590), 
        .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n923), .E(n675), .CP(n774), .CDN(n651), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(n921), .E(n675), .CP(n774), .CDN(n587), 
        .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n917), .E(n675), .CP(n774), .CDN(n581), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(n719), .E(n677), .CP(n774), .CDN(n639), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(n1011), .E(n677), .CP(n774), .CDN(n598), 
        .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(n1008), .E(n676), .CP(n774), .CDN(n598), 
        .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(n1005), .E(n677), .CP(n774), .CDN(n598), 
        .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(n1002), .E(n676), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(n999), .E(n677), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(n996), .E(n676), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(n993), .E(n677), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(n990), .E(n676), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(n987), .E(n677), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n984), .E(n676), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(n981), .E(n676), .CP(n775), .CDN(n598), 
        .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(n978), .E(n676), .CP(n775), .CDN(n597), 
        .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(n974), .E(n676), .CP(n775), .CDN(n597), 
        .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(n972), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(n969), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(n966), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(n963), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(n960), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(n957), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n953), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(n951), .E(n676), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(n948), .E(n677), .CP(n776), .CDN(n597), 
        .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n945), .E(n677), .CP(n776), .CDN(n596), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(n942), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(n939), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n936), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n932), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n930), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(n927), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n923), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(n921), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n917), .E(n677), .CP(n777), .CDN(n596), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(n719), .E(n683), .CP(n784), .CDN(n589), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(n1011), .E(n683), .CP(n784), .CDN(n646), 
        .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(n1008), .E(n682), .CP(n784), .CDN(n648), 
        .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(n1005), .E(n683), .CP(n784), .CDN(n650), 
        .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(n1002), .E(n682), .CP(n784), .CDN(n616), 
        .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(n999), .E(n683), .CP(n785), .CDN(n567), 
        .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(n996), .E(n682), .CP(n785), .CDN(n623), 
        .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(n993), .E(n683), .CP(n785), .CDN(n650), 
        .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(n990), .E(n682), .CP(n785), .CDN(n566), 
        .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(n987), .E(n683), .CP(n785), .CDN(n580), 
        .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n984), .E(n682), .CP(n785), .CDN(n650), 
        .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(n981), .E(n682), .CP(n785), .CDN(n640), 
        .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(n978), .E(n682), .CP(n785), .CDN(n642), 
        .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(n974), .E(n682), .CP(n785), .CDN(n644), 
        .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(n972), .E(n682), .CP(n785), .CDN(n641), 
        .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(n969), .E(n682), .CP(n786), .CDN(n626), 
        .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(n966), .E(n682), .CP(n786), .CDN(n643), 
        .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(n963), .E(n682), .CP(n786), .CDN(n599), 
        .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(n960), .E(n682), .CP(n786), .CDN(n647), 
        .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(n957), .E(n682), .CP(n786), .CDN(n635), 
        .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n953), .E(n682), .CP(n786), .CDN(n634), 
        .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(n951), .E(n682), .CP(n786), .CDN(n650), 
        .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(n948), .E(n683), .CP(n786), .CDN(n588), 
        .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n945), .E(n683), .CP(n786), .CDN(n630), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(n942), .E(n683), .CP(n786), .CDN(n633), 
        .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(n939), .E(n683), .CP(n787), .CDN(n645), 
        .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n936), .E(n683), .CP(n787), .CDN(n640), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n932), .E(n683), .CP(n787), .CDN(n642), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n930), .E(n683), .CP(n787), .CDN(n645), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(n927), .E(n683), .CP(n787), .CDN(n633), 
        .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n923), .E(n683), .CP(n787), .CDN(n576), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(n921), .E(n683), .CP(n787), .CDN(n577), 
        .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n917), .E(n683), .CP(n787), .CDN(n578), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n719), .E(n685), .CP(n787), .CDN(n579), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n1011), .E(n685), .CP(n787), .CDN(n591), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n1008), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n1005), .E(n685), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n1002), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n999), .E(n685), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n996), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n993), .E(n685), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n990), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n987), .E(n685), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n984), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n981), .E(n684), .CP(n788), .CDN(n591), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n978), .E(n684), .CP(n789), .CDN(n621), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n974), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n972), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n969), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n966), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n963), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n960), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n957), .E(n684), .CP(n789), .CDN(n591), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n953), .E(n684), .CP(n789), .CDN(n581), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n951), .E(n684), .CP(n789), .CDN(n587), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n948), .E(n685), .CP(n790), .CDN(n591), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n945), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n942), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n939), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n936), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n932), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n930), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n927), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n923), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n921), .E(n685), .CP(n790), .CDN(n590), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n917), .E(n685), .CP(n791), .CDN(n590), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(n719), .E(n691), .CP(n797), .CDN(n586), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n1011), .E(n691), .CP(n797), .CDN(n585), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n1007), .E(n690), .CP(n797), .CDN(n585), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n1004), .E(n691), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n1002), .E(n690), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n999), .E(n691), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n995), .E(n690), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n992), .E(n691), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n990), .E(n690), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n987), .E(n691), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n983), .E(n690), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n980), .E(n690), .CP(n798), .CDN(n585), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n978), .E(n690), .CP(n798), .CDN(n584), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n974), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n971), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n968), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n966), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n962), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n959), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n957), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n953), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n950), .E(n690), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n947), .E(n691), .CP(n799), .CDN(n584), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n945), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n941), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n938), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n936), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n932), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n929), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n926), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n923), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n920), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n917), .E(n691), .CP(n800), .CDN(n583), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n720), .E(n693), .CP(n801), .CDN(n583), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n1011), .E(n693), .CP(n801), .CDN(n651), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n1007), .E(n692), .CP(n801), .CDN(n622), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n1004), .E(n693), .CP(n801), .CDN(n599), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n1002), .E(n692), .CP(n801), .CDN(n573), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n999), .E(n693), .CP(n801), .CDN(n589), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n995), .E(n692), .CP(n801), .CDN(n585), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n992), .E(n693), .CP(n801), .CDN(n636), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n990), .E(n692), .CP(n801), .CDN(n638), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n987), .E(n693), .CP(n801), .CDN(n580), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n983), .E(n692), .CP(n802), .CDN(n651), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n980), .E(n692), .CP(n802), .CDN(n632), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n978), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n974), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n971), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n968), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n966), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n962), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n959), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n957), .E(n692), .CP(n802), .CDN(n582), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n953), .E(n692), .CP(n803), .CDN(n582), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n950), .E(n692), .CP(n803), .CDN(n582), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n947), .E(n693), .CP(n803), .CDN(n582), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n945), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n941), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n938), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n936), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n932), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n929), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n926), .E(n693), .CP(n803), .CDN(n581), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n923), .E(n693), .CP(n804), .CDN(n581), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n920), .E(n693), .CP(n804), .CDN(n581), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n917), .E(n693), .CP(n804), .CDN(n581), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(n720), .E(n699), .CP(n810), .CDN(n575), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n1010), .E(n699), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n1007), .E(n698), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n1004), .E(n699), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n1001), .E(n698), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n998), .E(n699), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n995), .E(n698), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n992), .E(n699), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n989), .E(n698), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n986), .E(n699), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n983), .E(n698), .CP(n811), .CDN(n574), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n980), .E(n698), .CP(n812), .CDN(n574), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n977), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n974), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n971), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n968), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n965), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n962), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n959), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n956), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n953), .E(n698), .CP(n812), .CDN(n573), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n950), .E(n698), .CP(n813), .CDN(n573), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n947), .E(n699), .CP(n813), .CDN(n573), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n944), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n941), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n938), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n935), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n932), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n929), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n926), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n923), .E(n699), .CP(n813), .CDN(n572), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n920), .E(n699), .CP(n814), .CDN(n572), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n917), .E(n699), .CP(n814), .CDN(n572), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n720), .E(n701), .CP(n814), .CDN(n572), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n1010), .E(n701), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n1007), .E(n700), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n1004), .E(n701), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n1001), .E(n700), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n998), .E(n701), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n995), .E(n700), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n992), .E(n701), .CP(n814), .CDN(n571), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n989), .E(n700), .CP(n815), .CDN(n571), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n986), .E(n701), .CP(n815), .CDN(n571), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n983), .E(n700), .CP(n815), .CDN(n571), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n980), .E(n700), .CP(n815), .CDN(n571), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n977), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n975), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n971), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n968), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n965), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n962), .E(n700), .CP(n815), .CDN(n570), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n959), .E(n700), .CP(n816), .CDN(n570), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n956), .E(n700), .CP(n816), .CDN(n570), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n954), .E(n700), .CP(n816), .CDN(n570), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n950), .E(n700), .CP(n816), .CDN(n570), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n947), .E(n701), .CP(n816), .CDN(n570), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n944), .E(n701), .CP(n816), .CDN(n569), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n941), .E(n701), .CP(n816), .CDN(n569), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n938), .E(n701), .CP(n816), .CDN(n569), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n935), .E(n701), .CP(n816), .CDN(n569), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n932), .E(n701), .CP(n816), .CDN(n569), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n929), .E(n701), .CP(n817), .CDN(n569), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n926), .E(n701), .CP(n817), .CDN(n569), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n924), .E(n701), .CP(n817), .CDN(n569), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n920), .E(n701), .CP(n817), .CDN(n569), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n918), .E(n701), .CP(n817), .CDN(n569), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(n720), .E(n707), .CP(n824), .CDN(n564), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n1010), .E(n707), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n1007), .E(n706), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n1004), .E(n707), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n1001), .E(n706), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n998), .E(n707), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n995), .E(n706), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n992), .E(n707), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n989), .E(n706), .CP(n824), .CDN(n563), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n986), .E(n707), .CP(n825), .CDN(n563), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n983), .E(n706), .CP(n825), .CDN(n563), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n980), .E(n706), .CP(n825), .CDN(n563), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n977), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n975), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n971), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n968), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n965), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n962), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n959), .E(n706), .CP(n825), .CDN(n562), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n956), .E(n706), .CP(n826), .CDN(n562), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n954), .E(n706), .CP(n826), .CDN(n562), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n950), .E(n706), .CP(n826), .CDN(n562), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n947), .E(n707), .CP(n826), .CDN(n562), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n944), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n941), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n938), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n935), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n932), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n929), .E(n707), .CP(n826), .CDN(n561), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n926), .E(n707), .CP(n827), .CDN(n561), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n924), .E(n707), .CP(n827), .CDN(n561), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n920), .E(n707), .CP(n827), .CDN(n561), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n918), .E(n707), .CP(n827), .CDN(n561), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n720), .E(n709), .CP(n827), .CDN(n561), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n1010), .E(n709), .CP(n827), .CDN(n560), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n1007), .E(n708), .CP(n827), .CDN(n560), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n1004), .E(n709), .CP(n827), .CDN(n560), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n1001), .E(n708), .CP(n827), .CDN(n560), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n998), .E(n709), .CP(n827), .CDN(n560), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n995), .E(n708), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n992), .E(n709), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n989), .E(n708), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n986), .E(n709), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n983), .E(n708), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n980), .E(n708), .CP(n828), .CDN(n560), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n977), .E(n708), .CP(n828), .CDN(n559), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n974), .E(n708), .CP(n828), .CDN(n559), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n971), .E(n708), .CP(n828), .CDN(n559), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n968), .E(n708), .CP(n828), .CDN(n559), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n965), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n962), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n959), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n956), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n953), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n950), .E(n708), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n947), .E(n709), .CP(n829), .CDN(n559), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n944), .E(n709), .CP(n829), .CDN(n558), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n941), .E(n709), .CP(n829), .CDN(n558), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n938), .E(n709), .CP(n829), .CDN(n558), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n935), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n933), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n929), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n926), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n923), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n920), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n917), .E(n709), .CP(n830), .CDN(n558), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(n720), .E(n714), .CP(n837), .CDN(n552), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n1010), .E(n714), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n1007), .E(n714), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n1004), .E(n714), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n1001), .E(n715), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n998), .E(n714), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n995), .E(n715), .CP(n837), .CDN(n551), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n992), .E(n714), .CP(n838), .CDN(n551), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n989), .E(n715), .CP(n838), .CDN(n551), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n986), .E(n714), .CP(n838), .CDN(n551), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n983), .E(n715), .CP(n838), .CDN(n551), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n980), .E(n714), .CP(n838), .CDN(n551), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n977), .E(n714), .CP(n838), .CDN(n550), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n975), .E(n714), .CP(n838), .CDN(n550), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n971), .E(n714), .CP(n838), .CDN(n550), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n968), .E(n714), .CP(n838), .CDN(n550), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n965), .E(n714), .CP(n838), .CDN(n550), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n962), .E(n714), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n959), .E(n714), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n956), .E(n714), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n954), .E(n714), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n950), .E(n714), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n947), .E(n715), .CP(n839), .CDN(n550), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n944), .E(n715), .CP(n839), .CDN(n549), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n941), .E(n715), .CP(n839), .CDN(n549), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n938), .E(n715), .CP(n839), .CDN(n549), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n935), .E(n715), .CP(n839), .CDN(n549), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n933), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n929), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n926), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n924), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n920), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n918), .E(n715), .CP(n840), .CDN(n549), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n718), .E(n653), .CP(n735), .CDN(n627), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(n1011), .E(n653), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(n1008), .E(n652), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(n1005), .E(n653), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(n1002), .E(n652), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(n999), .E(n653), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(n993), .E(n652), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(n990), .E(n653), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(n987), .E(n652), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(n984), .E(n653), .CP(n736), .CDN(n626), 
        .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(n981), .E(n652), .CP(n736), .CDN(n626), 
        .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(n978), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(n975), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(n972), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(n969), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(n966), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(n963), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(n960), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(n957), .E(n652), .CP(n736), .CDN(n625), 
        .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(n954), .E(n652), .CP(n737), .CDN(n625), 
        .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(n951), .E(n652), .CP(n737), .CDN(n625), 
        .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(n948), .E(n653), .CP(n737), .CDN(n625), 
        .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(n945), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(n942), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(n939), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n936), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(n933), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(n930), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(n927), .E(n653), .CP(n737), .CDN(n624), 
        .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(n924), .E(n653), .CP(n738), .CDN(n624), 
        .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(n921), .E(n653), .CP(n738), .CDN(n624), 
        .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(n918), .E(n653), .CP(n738), .CDN(n624), 
        .Q(\Storage[31][0] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(n996), .E(n655), .CP(n738), .CDN(n623), 
        .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(n993), .E(n654), .CP(n739), .CDN(n623), 
        .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(n996), .E(n657), .CP(n742), .CDN(n625), 
        .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(n993), .E(n656), .CP(n742), .CDN(n627), 
        .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(n999), .E(n658), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(n996), .E(n659), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(n993), .E(n658), .CP(n745), .CDN(n619), 
        .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(n996), .E(n652), .CP(n735), .CDN(n626), 
        .Q(\Storage[31][26] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N51), .E(Read), .CP(n912), .CDN(n628), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N52), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N53), .E(Read), .CP(ClockR), .CDN(n629), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N54), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N55), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N56), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N57), .E(Read), .CP(n912), .CDN(n629), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N58), .E(n915), .CP(ClockR), .CDN(n629), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N59), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N60), .E(Read), .CP(n912), .CDN(n629), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N61), .E(Read), .CP(n912), .CDN(n629), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N62), .E(n914), .CP(ClockR), .CDN(n629), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N63), .E(Read), .CP(n912), .CDN(n628), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N64), .E(n914), .CP(ClockR), .CDN(n628), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N65), .E(n915), .CP(n912), .CDN(n628), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N66), .E(n914), .CP(ClockR), .CDN(n628), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N67), .E(n914), .CP(n912), .CDN(n628), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N68), .E(n914), .CP(ClockR), .CDN(n628), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N69), .E(n914), .CP(n912), .CDN(n628), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N70), .E(n914), .CP(ClockR), .CDN(n628), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N71), .E(n914), .CP(n912), .CDN(n628), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N72), .E(Read), .CP(n912), .CDN(n628), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N73), .E(Read), .CP(n912), .CDN(n628), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N74), .E(n915), .CP(n912), .CDN(n627), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N75), .E(n915), .CP(n912), .CDN(n627), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N76), .E(Read), .CP(n912), .CDN(n627), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N77), .E(n915), .CP(n912), .CDN(n627), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N78), .E(n915), .CP(n912), .CDN(n627), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N79), .E(n915), .CP(n912), .CDN(n627), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N80), .E(Read), .CP(n912), .CDN(n627), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N81), .E(n915), .CP(ClockR), .CDN(n627), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N82), .E(n915), .CP(ClockR), .CDN(n627), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N83), .E(n915), .CP(ClockR), .CDN(n627), .Q(
        ParityErr) );
  EDFCNQD1 Dreadyr_reg ( .D(n1), .E(n915), .CP(ClockR), .CDN(n108), .Q(Dreadyr) );
  TIEH U3 ( .Z(n1) );
  CKBD0 U4 ( .CLK(Read), .C(n914) );
  CKBD0 U5 ( .CLK(Read), .C(n915) );
  CKBD0 U6 ( .CLK(N46), .C(n916) );
  CKBD0 U7 ( .CLK(N45), .C(n518) );
  CKBD0 U8 ( .CLK(N45), .C(n517) );
  BUFFD0 U9 ( .I(n518), .Z(n519) );
  CKBD0 U10 ( .CLK(N45), .C(n516) );
  BUFFD0 U11 ( .I(n518), .Z(n530) );
  BUFFD0 U12 ( .I(n531), .Z(n532) );
  CKBD0 U13 ( .CLK(N44), .C(n531) );
  INVD0 U14 ( .I(n716), .ZN(n721) );
  CKND0 U15 ( .CLK(n721), .CN(n720) );
  INVD0 U16 ( .I(DataI[23]), .ZN(n988) );
  CKNXD0 U17 ( .I(n988), .ZN(n986) );
  INVD0 U23 ( .I(DataI[24]), .ZN(n991) );
  CKNXD0 U24 ( .I(n991), .ZN(n989) );
  INVD0 U25 ( .I(DataI[27]), .ZN(n1000) );
  CKNXD0 U26 ( .I(n1000), .ZN(n998) );
  INVD0 U29 ( .I(DataI[28]), .ZN(n1003) );
  CKNXD0 U30 ( .I(n1003), .ZN(n1001) );
  INVD0 U31 ( .I(DataI[31]), .ZN(n1012) );
  CKNXD0 U32 ( .I(n1012), .ZN(n1010) );
  INVD0 U37 ( .I(DataI[26]), .ZN(n997) );
  INVD0 U38 ( .I(DataI[25]), .ZN(n994) );
  INVD0 U39 ( .I(DataI[22]), .ZN(n985) );
  INVD0 U40 ( .I(DataI[29]), .ZN(n1006) );
  INVD0 U41 ( .I(DataI[30]), .ZN(n1009) );
  INVD0 U42 ( .I(DataI[0]), .ZN(n919) );
  INVD0 U43 ( .I(n919), .ZN(n918) );
  CKNXD0 U44 ( .I(n919), .ZN(n917) );
  INVD0 U45 ( .I(DataI[2]), .ZN(n925) );
  INVD0 U46 ( .I(n925), .ZN(n924) );
  CKNXD0 U47 ( .I(n925), .ZN(n923) );
  INVD0 U48 ( .I(DataI[5]), .ZN(n934) );
  INVD0 U49 ( .I(n934), .ZN(n933) );
  CKNXD0 U50 ( .I(n934), .ZN(n932) );
  INVD0 U51 ( .I(DataI[12]), .ZN(n955) );
  INVD0 U52 ( .I(n955), .ZN(n954) );
  CKND0 U53 ( .CLK(n955), .CN(n953) );
  INVD0 U54 ( .I(DataI[19]), .ZN(n976) );
  INVD0 U55 ( .I(n976), .ZN(n975) );
  CKND0 U56 ( .CLK(n976), .CN(n974) );
  INVD0 U57 ( .I(DataI[6]), .ZN(n937) );
  CKNXD0 U58 ( .I(n937), .ZN(n935) );
  INVD0 U59 ( .I(DataI[9]), .ZN(n946) );
  CKNXD0 U60 ( .I(n946), .ZN(n944) );
  INVD0 U61 ( .I(DataI[13]), .ZN(n958) );
  CKNXD0 U62 ( .I(n958), .ZN(n956) );
  INVD0 U63 ( .I(DataI[16]), .ZN(n967) );
  CKNXD0 U64 ( .I(n967), .ZN(n965) );
  INVD0 U65 ( .I(DataI[20]), .ZN(n979) );
  CKNXD0 U66 ( .I(n979), .ZN(n977) );
  INVD0 U67 ( .I(DataI[1]), .ZN(n922) );
  INVD0 U68 ( .I(DataI[3]), .ZN(n928) );
  INVD0 U69 ( .I(DataI[4]), .ZN(n931) );
  INVD0 U70 ( .I(DataI[10]), .ZN(n949) );
  INVD0 U71 ( .I(DataI[11]), .ZN(n952) );
  INVD0 U72 ( .I(DataI[17]), .ZN(n970) );
  INVD0 U73 ( .I(DataI[18]), .ZN(n973) );
  INVD0 U74 ( .I(DataI[7]), .ZN(n940) );
  INVD0 U75 ( .I(DataI[8]), .ZN(n943) );
  INVD0 U76 ( .I(DataI[14]), .ZN(n961) );
  INVD0 U77 ( .I(DataI[15]), .ZN(n964) );
  INVD0 U78 ( .I(DataI[21]), .ZN(n982) );
  CKAN2D0 U79 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U80 ( .I(N48), .ZN(n505) );
  BUFFD1 U81 ( .I(n640), .Z(n572) );
  BUFFD1 U82 ( .I(n640), .Z(n573) );
  BUFFD1 U83 ( .I(n640), .Z(n574) );
  BUFFD1 U84 ( .I(n640), .Z(n575) );
  BUFFD1 U85 ( .I(n639), .Z(n576) );
  BUFFD1 U86 ( .I(n639), .Z(n577) );
  BUFFD1 U87 ( .I(n639), .Z(n578) );
  BUFFD1 U88 ( .I(n639), .Z(n579) );
  BUFFD1 U89 ( .I(n630), .Z(n580) );
  BUFFD1 U90 ( .I(n651), .Z(n581) );
  BUFFD1 U91 ( .I(n638), .Z(n582) );
  BUFFD1 U92 ( .I(n638), .Z(n583) );
  BUFFD1 U93 ( .I(n638), .Z(n584) );
  BUFFD1 U94 ( .I(n638), .Z(n585) );
  BUFFD1 U95 ( .I(n638), .Z(n586) );
  BUFFD1 U96 ( .I(n651), .Z(n587) );
  BUFFD1 U97 ( .I(n640), .Z(n588) );
  BUFFD1 U98 ( .I(n630), .Z(n589) );
  BUFFD1 U99 ( .I(n632), .Z(n590) );
  BUFFD1 U100 ( .I(n651), .Z(n591) );
  BUFFD1 U101 ( .I(n637), .Z(n592) );
  BUFFD1 U102 ( .I(n637), .Z(n593) );
  BUFFD1 U103 ( .I(n637), .Z(n594) );
  BUFFD1 U104 ( .I(n636), .Z(n595) );
  BUFFD1 U105 ( .I(n636), .Z(n596) );
  BUFFD1 U106 ( .I(n636), .Z(n597) );
  BUFFD1 U107 ( .I(n636), .Z(n598) );
  BUFFD1 U108 ( .I(n630), .Z(n599) );
  BUFFD1 U109 ( .I(n635), .Z(n600) );
  BUFFD1 U110 ( .I(n635), .Z(n601) );
  BUFFD1 U111 ( .I(n635), .Z(n602) );
  BUFFD1 U112 ( .I(n634), .Z(n603) );
  BUFFD1 U113 ( .I(n634), .Z(n604) );
  BUFFD1 U114 ( .I(n634), .Z(n605) );
  BUFFD1 U115 ( .I(n633), .Z(n606) );
  BUFFD1 U116 ( .I(n633), .Z(n607) );
  BUFFD1 U117 ( .I(n633), .Z(n608) );
  BUFFD1 U118 ( .I(n633), .Z(n609) );
  BUFFD1 U119 ( .I(n631), .Z(n610) );
  BUFFD1 U120 ( .I(n646), .Z(n611) );
  BUFFD1 U121 ( .I(n637), .Z(n612) );
  BUFFD1 U122 ( .I(n632), .Z(n613) );
  BUFFD1 U123 ( .I(n632), .Z(n614) );
  BUFFD1 U124 ( .I(n632), .Z(n615) );
  BUFFD1 U125 ( .I(n632), .Z(n616) );
  BUFFD1 U126 ( .I(n631), .Z(n617) );
  BUFFD1 U127 ( .I(n631), .Z(n618) );
  BUFFD1 U128 ( .I(n631), .Z(n619) );
  BUFFD1 U129 ( .I(n631), .Z(n620) );
  BUFFD1 U130 ( .I(n649), .Z(n621) );
  BUFFD1 U131 ( .I(n108), .Z(n622) );
  BUFFD1 U132 ( .I(n630), .Z(n623) );
  BUFFD1 U133 ( .I(n630), .Z(n624) );
  BUFFD1 U134 ( .I(n630), .Z(n625) );
  BUFFD1 U135 ( .I(n630), .Z(n626) );
  BUFFD1 U136 ( .I(n642), .Z(n549) );
  BUFFD1 U137 ( .I(n639), .Z(n550) );
  BUFFD1 U138 ( .I(n645), .Z(n551) );
  BUFFD1 U139 ( .I(n645), .Z(n552) );
  BUFFD1 U140 ( .I(n645), .Z(n553) );
  BUFFD1 U141 ( .I(n645), .Z(n554) );
  BUFFD1 U142 ( .I(n645), .Z(n555) );
  BUFFD1 U143 ( .I(n645), .Z(n556) );
  BUFFD1 U144 ( .I(n644), .Z(n557) );
  BUFFD1 U145 ( .I(n644), .Z(n558) );
  BUFFD1 U146 ( .I(n644), .Z(n559) );
  BUFFD1 U147 ( .I(n644), .Z(n560) );
  BUFFD1 U148 ( .I(n643), .Z(n561) );
  BUFFD1 U149 ( .I(n643), .Z(n562) );
  BUFFD1 U150 ( .I(n643), .Z(n563) );
  BUFFD1 U151 ( .I(n643), .Z(n564) );
  BUFFD1 U152 ( .I(n642), .Z(n565) );
  BUFFD1 U153 ( .I(n642), .Z(n566) );
  BUFFD1 U154 ( .I(n642), .Z(n567) );
  BUFFD1 U155 ( .I(n641), .Z(n568) );
  BUFFD1 U156 ( .I(n641), .Z(n569) );
  BUFFD1 U157 ( .I(n641), .Z(n570) );
  BUFFD1 U158 ( .I(n641), .Z(n571) );
  BUFFD1 U159 ( .I(n649), .Z(n640) );
  BUFFD1 U160 ( .I(n649), .Z(n639) );
  BUFFD1 U161 ( .I(n651), .Z(n638) );
  BUFFD1 U162 ( .I(n647), .Z(n637) );
  BUFFD1 U163 ( .I(n651), .Z(n636) );
  BUFFD1 U164 ( .I(n650), .Z(n635) );
  BUFFD1 U165 ( .I(n650), .Z(n634) );
  BUFFD1 U166 ( .I(n648), .Z(n633) );
  BUFFD1 U167 ( .I(n651), .Z(n632) );
  BUFFD1 U168 ( .I(n651), .Z(n631) );
  BUFFD1 U169 ( .I(n548), .Z(n630) );
  BUFFD1 U170 ( .I(n841), .Z(n839) );
  BUFFD1 U171 ( .I(n842), .Z(n838) );
  BUFFD1 U172 ( .I(n842), .Z(n837) );
  BUFFD1 U173 ( .I(n843), .Z(n836) );
  BUFFD1 U174 ( .I(n843), .Z(n835) );
  BUFFD1 U175 ( .I(n844), .Z(n834) );
  BUFFD1 U176 ( .I(n844), .Z(n833) );
  BUFFD1 U177 ( .I(n845), .Z(n832) );
  BUFFD1 U178 ( .I(n845), .Z(n831) );
  BUFFD1 U179 ( .I(n846), .Z(n830) );
  BUFFD1 U180 ( .I(n846), .Z(n829) );
  BUFFD1 U181 ( .I(n847), .Z(n828) );
  BUFFD1 U182 ( .I(n847), .Z(n827) );
  BUFFD1 U183 ( .I(n848), .Z(n826) );
  BUFFD1 U184 ( .I(n848), .Z(n825) );
  BUFFD1 U185 ( .I(n849), .Z(n824) );
  BUFFD1 U186 ( .I(n849), .Z(n823) );
  BUFFD1 U187 ( .I(n850), .Z(n822) );
  BUFFD1 U188 ( .I(n850), .Z(n821) );
  BUFFD1 U189 ( .I(n851), .Z(n820) );
  BUFFD1 U190 ( .I(n851), .Z(n819) );
  BUFFD1 U191 ( .I(n852), .Z(n818) );
  BUFFD1 U192 ( .I(n852), .Z(n817) );
  BUFFD1 U193 ( .I(n853), .Z(n816) );
  BUFFD1 U194 ( .I(n853), .Z(n815) );
  BUFFD1 U195 ( .I(n854), .Z(n814) );
  BUFFD1 U196 ( .I(n854), .Z(n813) );
  BUFFD1 U197 ( .I(n855), .Z(n812) );
  BUFFD1 U198 ( .I(n855), .Z(n811) );
  BUFFD1 U199 ( .I(n856), .Z(n810) );
  BUFFD1 U200 ( .I(n856), .Z(n809) );
  BUFFD1 U201 ( .I(n857), .Z(n808) );
  BUFFD1 U202 ( .I(n857), .Z(n807) );
  BUFFD1 U203 ( .I(n858), .Z(n806) );
  BUFFD1 U204 ( .I(n858), .Z(n805) );
  BUFFD1 U205 ( .I(n859), .Z(n804) );
  BUFFD1 U206 ( .I(n859), .Z(n803) );
  BUFFD1 U207 ( .I(n860), .Z(n802) );
  BUFFD1 U208 ( .I(n860), .Z(n801) );
  BUFFD1 U209 ( .I(n861), .Z(n800) );
  BUFFD1 U210 ( .I(n861), .Z(n799) );
  BUFFD1 U211 ( .I(n862), .Z(n798) );
  BUFFD1 U212 ( .I(n862), .Z(n797) );
  BUFFD1 U213 ( .I(n863), .Z(n796) );
  BUFFD1 U214 ( .I(n863), .Z(n795) );
  BUFFD1 U215 ( .I(n864), .Z(n794) );
  BUFFD1 U216 ( .I(n864), .Z(n793) );
  BUFFD1 U217 ( .I(n865), .Z(n792) );
  BUFFD1 U218 ( .I(n865), .Z(n791) );
  BUFFD1 U219 ( .I(n866), .Z(n790) );
  BUFFD1 U220 ( .I(n866), .Z(n789) );
  BUFFD1 U221 ( .I(n867), .Z(n788) );
  BUFFD1 U222 ( .I(n867), .Z(n787) );
  BUFFD1 U223 ( .I(n868), .Z(n786) );
  BUFFD1 U224 ( .I(n868), .Z(n785) );
  BUFFD1 U225 ( .I(n869), .Z(n784) );
  BUFFD1 U226 ( .I(n869), .Z(n783) );
  BUFFD1 U227 ( .I(n870), .Z(n782) );
  BUFFD1 U228 ( .I(n870), .Z(n781) );
  BUFFD1 U229 ( .I(n871), .Z(n780) );
  BUFFD1 U230 ( .I(n871), .Z(n779) );
  BUFFD1 U231 ( .I(n872), .Z(n778) );
  BUFFD1 U232 ( .I(n872), .Z(n777) );
  BUFFD1 U233 ( .I(n873), .Z(n776) );
  BUFFD1 U234 ( .I(n873), .Z(n775) );
  BUFFD1 U235 ( .I(n874), .Z(n774) );
  BUFFD1 U236 ( .I(n874), .Z(n773) );
  BUFFD1 U237 ( .I(n875), .Z(n772) );
  BUFFD1 U238 ( .I(n875), .Z(n771) );
  BUFFD1 U239 ( .I(n876), .Z(n770) );
  BUFFD1 U240 ( .I(n876), .Z(n769) );
  BUFFD1 U241 ( .I(n877), .Z(n768) );
  BUFFD1 U242 ( .I(n877), .Z(n767) );
  BUFFD1 U243 ( .I(n878), .Z(n766) );
  BUFFD1 U244 ( .I(n878), .Z(n765) );
  BUFFD1 U245 ( .I(n879), .Z(n764) );
  BUFFD1 U246 ( .I(n879), .Z(n763) );
  BUFFD1 U247 ( .I(n880), .Z(n762) );
  BUFFD1 U248 ( .I(n880), .Z(n761) );
  BUFFD1 U249 ( .I(n881), .Z(n760) );
  BUFFD1 U250 ( .I(n881), .Z(n759) );
  BUFFD1 U251 ( .I(n882), .Z(n758) );
  BUFFD1 U252 ( .I(n882), .Z(n757) );
  BUFFD1 U253 ( .I(n883), .Z(n756) );
  BUFFD1 U254 ( .I(n883), .Z(n755) );
  BUFFD1 U255 ( .I(n884), .Z(n754) );
  BUFFD1 U256 ( .I(n884), .Z(n753) );
  BUFFD1 U257 ( .I(n885), .Z(n752) );
  BUFFD1 U258 ( .I(n885), .Z(n751) );
  BUFFD1 U259 ( .I(n886), .Z(n750) );
  BUFFD1 U260 ( .I(n886), .Z(n749) );
  BUFFD1 U261 ( .I(n887), .Z(n748) );
  BUFFD1 U262 ( .I(n887), .Z(n747) );
  BUFFD1 U263 ( .I(n888), .Z(n746) );
  BUFFD1 U264 ( .I(n888), .Z(n745) );
  BUFFD1 U265 ( .I(n889), .Z(n744) );
  BUFFD1 U266 ( .I(n889), .Z(n743) );
  BUFFD1 U267 ( .I(n890), .Z(n742) );
  BUFFD1 U268 ( .I(n890), .Z(n741) );
  BUFFD1 U269 ( .I(n891), .Z(n740) );
  BUFFD1 U270 ( .I(n891), .Z(n739) );
  BUFFD1 U271 ( .I(n892), .Z(n738) );
  BUFFD1 U272 ( .I(n892), .Z(n737) );
  BUFFD1 U273 ( .I(n893), .Z(n736) );
  BUFFD1 U274 ( .I(n893), .Z(n735) );
  BUFFD1 U275 ( .I(n841), .Z(n840) );
  BUFFD1 U276 ( .I(n535), .Z(n537) );
  BUFFD1 U277 ( .I(n517), .Z(n525) );
  BUFFD1 U278 ( .I(n535), .Z(n538) );
  BUFFD1 U279 ( .I(n534), .Z(n539) );
  BUFFD1 U280 ( .I(n534), .Z(n540) );
  BUFFD1 U281 ( .I(n534), .Z(n541) );
  BUFFD1 U282 ( .I(n533), .Z(n542) );
  BUFFD1 U283 ( .I(n533), .Z(n543) );
  BUFFD1 U284 ( .I(n533), .Z(n544) );
  BUFFD1 U285 ( .I(n532), .Z(n545) );
  BUFFD1 U286 ( .I(n532), .Z(n546) );
  BUFFD1 U287 ( .I(n520), .Z(n527) );
  BUFFD1 U288 ( .I(n520), .Z(n528) );
  BUFFD1 U289 ( .I(n519), .Z(n529) );
  BUFFD1 U290 ( .I(n521), .Z(n523) );
  BUFFD1 U291 ( .I(n521), .Z(n524) );
  BUFFD1 U292 ( .I(n520), .Z(n526) );
  BUFFD1 U293 ( .I(n521), .Z(n522) );
  BUFFD1 U294 ( .I(n535), .Z(n536) );
  INVD1 U295 ( .I(n722), .ZN(n719) );
  INVD1 U296 ( .I(n722), .ZN(n718) );
  BUFFD1 U297 ( .I(n630), .Z(n627) );
  BUFFD1 U298 ( .I(n646), .Z(n645) );
  BUFFD1 U299 ( .I(n647), .Z(n644) );
  BUFFD1 U300 ( .I(n647), .Z(n643) );
  BUFFD1 U301 ( .I(n648), .Z(n642) );
  BUFFD1 U302 ( .I(n648), .Z(n641) );
  BUFFD1 U303 ( .I(n547), .Z(n649) );
  BUFFD1 U304 ( .I(n548), .Z(n650) );
  BUFFD1 U305 ( .I(n108), .Z(n651) );
  BUFFD1 U306 ( .I(n910), .Z(n843) );
  BUFFD1 U307 ( .I(n910), .Z(n844) );
  BUFFD1 U308 ( .I(n910), .Z(n845) );
  BUFFD1 U309 ( .I(n909), .Z(n846) );
  BUFFD1 U310 ( .I(n909), .Z(n847) );
  BUFFD1 U311 ( .I(n909), .Z(n848) );
  BUFFD1 U312 ( .I(n908), .Z(n849) );
  BUFFD1 U313 ( .I(n908), .Z(n850) );
  BUFFD1 U314 ( .I(n908), .Z(n851) );
  BUFFD1 U315 ( .I(n907), .Z(n852) );
  BUFFD1 U316 ( .I(n907), .Z(n853) );
  BUFFD1 U317 ( .I(n907), .Z(n854) );
  BUFFD1 U318 ( .I(n906), .Z(n855) );
  BUFFD1 U319 ( .I(n906), .Z(n856) );
  BUFFD1 U320 ( .I(n906), .Z(n857) );
  BUFFD1 U321 ( .I(n905), .Z(n858) );
  BUFFD1 U322 ( .I(n905), .Z(n859) );
  BUFFD1 U323 ( .I(n905), .Z(n860) );
  BUFFD1 U324 ( .I(n904), .Z(n861) );
  BUFFD1 U325 ( .I(n904), .Z(n862) );
  BUFFD1 U326 ( .I(n904), .Z(n863) );
  BUFFD1 U327 ( .I(n903), .Z(n864) );
  BUFFD1 U328 ( .I(n903), .Z(n865) );
  BUFFD1 U329 ( .I(n903), .Z(n866) );
  BUFFD1 U330 ( .I(n902), .Z(n867) );
  BUFFD1 U331 ( .I(n902), .Z(n868) );
  BUFFD1 U332 ( .I(n902), .Z(n869) );
  BUFFD1 U333 ( .I(n901), .Z(n870) );
  BUFFD1 U334 ( .I(n901), .Z(n871) );
  BUFFD1 U335 ( .I(n901), .Z(n872) );
  BUFFD1 U336 ( .I(n900), .Z(n873) );
  BUFFD1 U337 ( .I(n900), .Z(n874) );
  BUFFD1 U338 ( .I(n900), .Z(n875) );
  BUFFD1 U339 ( .I(n899), .Z(n876) );
  BUFFD1 U340 ( .I(n899), .Z(n877) );
  BUFFD1 U341 ( .I(n899), .Z(n878) );
  BUFFD1 U342 ( .I(n898), .Z(n879) );
  BUFFD1 U343 ( .I(n898), .Z(n880) );
  BUFFD1 U344 ( .I(n898), .Z(n881) );
  BUFFD1 U345 ( .I(n897), .Z(n882) );
  BUFFD1 U346 ( .I(n897), .Z(n883) );
  BUFFD1 U347 ( .I(n897), .Z(n884) );
  BUFFD1 U348 ( .I(n896), .Z(n885) );
  BUFFD1 U349 ( .I(n896), .Z(n886) );
  BUFFD1 U350 ( .I(n896), .Z(n887) );
  BUFFD1 U351 ( .I(n895), .Z(n888) );
  BUFFD1 U352 ( .I(n895), .Z(n889) );
  BUFFD1 U353 ( .I(n895), .Z(n890) );
  BUFFD1 U354 ( .I(n894), .Z(n891) );
  BUFFD1 U355 ( .I(n894), .Z(n892) );
  BUFFD1 U356 ( .I(n894), .Z(n893) );
  BUFFD1 U357 ( .I(n911), .Z(n841) );
  BUFFD1 U358 ( .I(n911), .Z(n842) );
  BUFFD1 U359 ( .I(N44), .Z(n535) );
  BUFFD1 U360 ( .I(n507), .Z(n509) );
  BUFFD1 U361 ( .I(N47), .Z(n508) );
  BUFFD1 U362 ( .I(n510), .Z(n514) );
  BUFFD1 U363 ( .I(n510), .Z(n515) );
  BUFFD1 U364 ( .I(N46), .Z(n512) );
  BUFFD1 U365 ( .I(N46), .Z(n513) );
  BUFFD1 U366 ( .I(N47), .Z(n507) );
  BUFFD1 U367 ( .I(n531), .Z(n534) );
  BUFFD1 U368 ( .I(n531), .Z(n533) );
  BUFFD1 U369 ( .I(n517), .Z(n521) );
  BUFFD1 U370 ( .I(n517), .Z(n520) );
  BUFFD1 U371 ( .I(N46), .Z(n511) );
  BUFFD1 U372 ( .I(n642), .Z(n628) );
  BUFFD1 U373 ( .I(n628), .Z(n629) );
  INVD1 U374 ( .I(n716), .ZN(n722) );
  BUFFD1 U375 ( .I(n547), .Z(n647) );
  BUFFD1 U376 ( .I(n547), .Z(n648) );
  BUFFD1 U377 ( .I(n547), .Z(n646) );
  BUFFD1 U378 ( .I(n731), .Z(n910) );
  BUFFD1 U379 ( .I(n730), .Z(n909) );
  BUFFD1 U380 ( .I(n730), .Z(n908) );
  BUFFD1 U381 ( .I(n729), .Z(n907) );
  BUFFD1 U382 ( .I(n729), .Z(n906) );
  BUFFD1 U383 ( .I(n728), .Z(n905) );
  BUFFD1 U384 ( .I(n728), .Z(n904) );
  BUFFD1 U385 ( .I(n727), .Z(n903) );
  BUFFD1 U386 ( .I(n727), .Z(n902) );
  BUFFD1 U387 ( .I(n726), .Z(n901) );
  BUFFD1 U388 ( .I(n726), .Z(n900) );
  BUFFD1 U389 ( .I(n725), .Z(n899) );
  BUFFD1 U390 ( .I(n725), .Z(n898) );
  BUFFD1 U391 ( .I(n724), .Z(n897) );
  BUFFD1 U392 ( .I(n724), .Z(n896) );
  BUFFD1 U393 ( .I(n723), .Z(n895) );
  BUFFD1 U394 ( .I(n723), .Z(n894) );
  BUFFD1 U395 ( .I(n731), .Z(n911) );
  BUFFD1 U396 ( .I(n916), .Z(n510) );
  INVD1 U397 ( .I(n505), .ZN(n506) );
  XOR3D1 U398 ( .A1(n80), .A2(n947), .A3(n81), .Z(n79) );
  XOR3D1 U399 ( .A1(DataI[19]), .A2(n971), .A3(n82), .Z(n81) );
  XOR3D1 U400 ( .A1(n83), .A2(n968), .A3(n84), .Z(n82) );
  XOR3D1 U401 ( .A1(DataI[5]), .A2(n929), .A3(n76), .Z(n75) );
  XOR3D1 U402 ( .A1(n77), .A2(n926), .A3(n78), .Z(n76) );
  XOR3D1 U403 ( .A1(DataI[12]), .A2(n950), .A3(n79), .Z(n78) );
  INVD1 U404 ( .I(n717), .ZN(n716) );
  INVD1 U405 ( .I(N85), .ZN(n717) );
  XOR3D1 U406 ( .A1(DataI[2]), .A2(n920), .A3(n73), .Z(N85) );
  XOR3D1 U407 ( .A1(DataI[0]), .A2(n74), .A3(n75), .Z(n73) );
  BUFFD1 U408 ( .I(n732), .Z(n731) );
  BUFFD1 U409 ( .I(n732), .Z(n730) );
  BUFFD1 U410 ( .I(n732), .Z(n729) );
  BUFFD1 U411 ( .I(n733), .Z(n728) );
  BUFFD1 U412 ( .I(n733), .Z(n727) );
  BUFFD1 U413 ( .I(n733), .Z(n726) );
  BUFFD1 U414 ( .I(n734), .Z(n725) );
  BUFFD1 U415 ( .I(n734), .Z(n724) );
  BUFFD1 U416 ( .I(n734), .Z(n723) );
  BUFFD1 U417 ( .I(n548), .Z(n547) );
  BUFFD1 U418 ( .I(n108), .Z(n548) );
  XOR3D1 U419 ( .A1(N67), .A2(N66), .A3(n92), .Z(n90) );
  XOR3D1 U420 ( .A1(N65), .A2(n93), .A3(n94), .Z(n92) );
  XOR3D1 U421 ( .A1(N60), .A2(N59), .A3(n95), .Z(n94) );
  XOR3D1 U422 ( .A1(n96), .A2(N58), .A3(n97), .Z(n95) );
  XOR3D1 U423 ( .A1(N79), .A2(N74), .A3(n86), .Z(N83) );
  XOR3D1 U424 ( .A1(N73), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D1 U425 ( .A1(N77), .A2(N76), .A3(n89), .Z(n88) );
  INVD1 U426 ( .I(n5), .ZN(n677) );
  INVD1 U427 ( .I(n5), .ZN(n676) );
  INVD1 U428 ( .I(n6), .ZN(n675) );
  INVD1 U429 ( .I(n6), .ZN(n674) );
  INVD1 U430 ( .I(n7), .ZN(n673) );
  INVD1 U431 ( .I(n7), .ZN(n672) );
  INVD1 U432 ( .I(n8), .ZN(n671) );
  INVD1 U433 ( .I(n8), .ZN(n670) );
  INVD1 U434 ( .I(n9), .ZN(n669) );
  INVD1 U435 ( .I(n9), .ZN(n668) );
  INVD1 U436 ( .I(n10), .ZN(n667) );
  INVD1 U437 ( .I(n10), .ZN(n666) );
  INVD1 U438 ( .I(n11), .ZN(n665) );
  INVD1 U439 ( .I(n11), .ZN(n664) );
  INVD1 U440 ( .I(n12), .ZN(n663) );
  INVD1 U441 ( .I(n12), .ZN(n662) );
  INVD1 U442 ( .I(n13), .ZN(n661) );
  INVD1 U443 ( .I(n13), .ZN(n660) );
  INVD1 U444 ( .I(n14), .ZN(n659) );
  INVD1 U445 ( .I(n14), .ZN(n658) );
  INVD1 U446 ( .I(n15), .ZN(n657) );
  INVD1 U447 ( .I(n15), .ZN(n656) );
  INVD1 U448 ( .I(n16), .ZN(n655) );
  INVD1 U449 ( .I(n16), .ZN(n654) );
  INVD1 U450 ( .I(n17), .ZN(n653) );
  INVD1 U451 ( .I(n17), .ZN(n652) );
  INVD1 U452 ( .I(n18), .ZN(n715) );
  INVD1 U453 ( .I(n18), .ZN(n714) );
  INVD1 U454 ( .I(n19), .ZN(n713) );
  INVD1 U455 ( .I(n19), .ZN(n712) );
  INVD1 U456 ( .I(n20), .ZN(n711) );
  INVD1 U457 ( .I(n20), .ZN(n710) );
  INVD1 U458 ( .I(n21), .ZN(n709) );
  INVD1 U459 ( .I(n21), .ZN(n708) );
  INVD1 U460 ( .I(n22), .ZN(n707) );
  INVD1 U461 ( .I(n22), .ZN(n706) );
  INVD1 U462 ( .I(n23), .ZN(n705) );
  INVD1 U463 ( .I(n23), .ZN(n704) );
  INVD1 U464 ( .I(n24), .ZN(n703) );
  INVD1 U465 ( .I(n24), .ZN(n702) );
  INVD1 U466 ( .I(n25), .ZN(n701) );
  INVD1 U467 ( .I(n25), .ZN(n700) );
  INVD1 U468 ( .I(n26), .ZN(n699) );
  INVD1 U469 ( .I(n26), .ZN(n698) );
  INVD1 U470 ( .I(n27), .ZN(n697) );
  INVD1 U471 ( .I(n27), .ZN(n696) );
  INVD1 U472 ( .I(n28), .ZN(n695) );
  INVD1 U473 ( .I(n28), .ZN(n694) );
  INVD1 U474 ( .I(n29), .ZN(n693) );
  INVD1 U475 ( .I(n29), .ZN(n692) );
  INVD1 U476 ( .I(n30), .ZN(n691) );
  INVD1 U477 ( .I(n30), .ZN(n690) );
  INVD1 U478 ( .I(n31), .ZN(n689) );
  INVD1 U479 ( .I(n31), .ZN(n688) );
  INVD1 U480 ( .I(n32), .ZN(n687) );
  INVD1 U481 ( .I(n32), .ZN(n686) );
  INVD1 U482 ( .I(n33), .ZN(n685) );
  INVD1 U483 ( .I(n33), .ZN(n684) );
  INVD1 U484 ( .I(n2), .ZN(n683) );
  INVD1 U485 ( .I(n2), .ZN(n682) );
  INVD1 U486 ( .I(n3), .ZN(n681) );
  INVD1 U487 ( .I(n3), .ZN(n680) );
  INVD1 U488 ( .I(n4), .ZN(n679) );
  INVD1 U489 ( .I(n4), .ZN(n678) );
  INVD1 U490 ( .I(n913), .ZN(n912) );
  INVD1 U491 ( .I(n1009), .ZN(n1007) );
  INVD1 U492 ( .I(n940), .ZN(n938) );
  INVD1 U493 ( .I(n943), .ZN(n941) );
  INVD1 U494 ( .I(n961), .ZN(n959) );
  INVD1 U495 ( .I(n964), .ZN(n962) );
  INVD1 U496 ( .I(n982), .ZN(n980) );
  INVD1 U497 ( .I(n985), .ZN(n983) );
  INVD1 U498 ( .I(n994), .ZN(n992) );
  INVD1 U499 ( .I(n997), .ZN(n995) );
  INVD1 U500 ( .I(n1006), .ZN(n1004) );
  INVD1 U501 ( .I(n922), .ZN(n920) );
  INVD1 U502 ( .I(n928), .ZN(n926) );
  INVD1 U503 ( .I(n931), .ZN(n929) );
  INVD1 U504 ( .I(n949), .ZN(n947) );
  INVD1 U505 ( .I(n952), .ZN(n950) );
  INVD1 U506 ( .I(n970), .ZN(n968) );
  INVD1 U507 ( .I(n973), .ZN(n971) );
  INVD1 U508 ( .I(n940), .ZN(n939) );
  INVD1 U509 ( .I(n943), .ZN(n942) );
  INVD1 U510 ( .I(n961), .ZN(n960) );
  INVD1 U511 ( .I(n964), .ZN(n963) );
  INVD1 U512 ( .I(n982), .ZN(n981) );
  INVD1 U513 ( .I(n985), .ZN(n984) );
  INVD1 U514 ( .I(n994), .ZN(n993) );
  INVD1 U515 ( .I(n997), .ZN(n996) );
  INVD1 U516 ( .I(n1006), .ZN(n1005) );
  INVD1 U517 ( .I(n1009), .ZN(n1008) );
  INVD1 U518 ( .I(n922), .ZN(n921) );
  INVD1 U519 ( .I(n928), .ZN(n927) );
  INVD1 U520 ( .I(n931), .ZN(n930) );
  INVD1 U521 ( .I(n949), .ZN(n948) );
  INVD1 U522 ( .I(n952), .ZN(n951) );
  INVD1 U523 ( .I(n970), .ZN(n969) );
  INVD1 U524 ( .I(n973), .ZN(n972) );
  INVD1 U525 ( .I(n937), .ZN(n936) );
  INVD1 U526 ( .I(n946), .ZN(n945) );
  INVD1 U527 ( .I(n958), .ZN(n957) );
  INVD1 U528 ( .I(n967), .ZN(n966) );
  INVD1 U529 ( .I(n979), .ZN(n978) );
  INVD1 U530 ( .I(n988), .ZN(n987) );
  INVD1 U531 ( .I(n991), .ZN(n990) );
  INVD1 U532 ( .I(n1000), .ZN(n999) );
  INVD1 U533 ( .I(n1003), .ZN(n1002) );
  INVD1 U534 ( .I(n1012), .ZN(n1011) );
  INVD1 U535 ( .I(Reset), .ZN(n108) );
  BUFFD1 U536 ( .I(ClockW), .Z(n732) );
  BUFFD1 U537 ( .I(ClockW), .Z(n733) );
  BUFFD1 U538 ( .I(ClockW), .Z(n734) );
  OR2D1 U539 ( .A1(n69), .A2(n70), .Z(n2) );
  OR2D1 U540 ( .A1(n68), .A2(n70), .Z(n3) );
  OR2D1 U541 ( .A1(n67), .A2(n70), .Z(n4) );
  ND3D1 U542 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  ND3D1 U543 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U544 ( .I(AddrW[1]), .ZN(n106) );
  OR2D1 U545 ( .A1(n70), .A2(n99), .Z(n5) );
  OR2D1 U546 ( .A1(n70), .A2(n98), .Z(n6) );
  OR2D1 U547 ( .A1(n70), .A2(n85), .Z(n7) );
  OR2D1 U548 ( .A1(n70), .A2(n72), .Z(n8) );
  OR2D1 U549 ( .A1(n70), .A2(n71), .Z(n9) );
  OR2D1 U550 ( .A1(n66), .A2(n69), .Z(n10) );
  OR2D1 U551 ( .A1(n66), .A2(n68), .Z(n11) );
  OR2D1 U552 ( .A1(n66), .A2(n67), .Z(n12) );
  OR2D1 U553 ( .A1(n66), .A2(n99), .Z(n13) );
  OR2D1 U554 ( .A1(n66), .A2(n98), .Z(n14) );
  OR2D1 U555 ( .A1(n66), .A2(n85), .Z(n15) );
  OR2D1 U556 ( .A1(n66), .A2(n72), .Z(n16) );
  OR2D1 U557 ( .A1(n66), .A2(n71), .Z(n17) );
  OR2D1 U558 ( .A1(n69), .A2(n103), .Z(n18) );
  OR2D1 U559 ( .A1(n68), .A2(n103), .Z(n19) );
  OR2D1 U560 ( .A1(n67), .A2(n103), .Z(n20) );
  OR2D1 U561 ( .A1(n99), .A2(n103), .Z(n21) );
  OR2D1 U562 ( .A1(n98), .A2(n103), .Z(n22) );
  OR2D1 U563 ( .A1(n85), .A2(n103), .Z(n23) );
  OR2D1 U564 ( .A1(n72), .A2(n103), .Z(n24) );
  OR2D1 U565 ( .A1(n71), .A2(n103), .Z(n25) );
  OR2D1 U566 ( .A1(n69), .A2(n101), .Z(n26) );
  OR2D1 U567 ( .A1(n68), .A2(n101), .Z(n27) );
  OR2D1 U568 ( .A1(n67), .A2(n101), .Z(n28) );
  OR2D1 U569 ( .A1(n99), .A2(n101), .Z(n29) );
  OR2D1 U570 ( .A1(n98), .A2(n101), .Z(n30) );
  OR2D1 U571 ( .A1(n85), .A2(n101), .Z(n31) );
  OR2D1 U572 ( .A1(n72), .A2(n101), .Z(n32) );
  OR2D1 U573 ( .A1(n71), .A2(n101), .Z(n33) );
  INVD1 U574 ( .I(ClockR), .ZN(n913) );
  CKAN2D0 U575 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX4D0 U576 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n532), .S1(n519), .Z(
        n405) );
  MUX4D0 U577 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n534), .S1(N45), .Z(
        n418) );
  MUX4D0 U578 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n536), .S1(N45), .Z(
        n431) );
  MUX4D0 U579 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n531), .S1(n525), .Z(
        n444) );
  MUX4D0 U580 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n536), .S1(n525), .Z(
        n470) );
  MUX4D0 U581 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n536), .S1(n517), .Z(
        n409) );
  MUX4D0 U582 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n536), .S1(N45), .Z(
        n407) );
  MUX4D0 U583 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n532), .S1(n520), .Z(
        n420) );
  MUX4D0 U584 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n532), .S1(n520), .Z(
        n422) );
  MUX4D0 U585 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n536), .S1(n517), .Z(
        n433) );
  MUX4D0 U586 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n534), .S1(n518), .Z(
        n435) );
  MUX4D0 U587 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n536), .S1(n525), .Z(
        n448) );
  MUX4D0 U588 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n532), .S1(n525), .Z(
        n446) );
  MUX4D0 U589 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n536), .S1(n525), .Z(
        n461) );
  MUX4D0 U590 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n533), .S1(n525), .Z(
        n459) );
  MUX4D0 U591 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n535), .S1(n526), .Z(
        n472) );
  MUX4D0 U592 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n535), .S1(n526), .Z(
        n474) );
  MUX4D0 U593 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n535), .S1(n526), .Z(
        n485) );
  MUX4D0 U594 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n535), .S1(n526), .Z(
        n487) );
  MUX4D0 U595 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n535), .S1(N45), .Z(
        n406) );
  MUX4D0 U596 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n534), .S1(n518), .Z(
        n419) );
  MUX4D0 U597 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n531), .S1(N45), .Z(
        n432) );
  MUX4D0 U598 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n534), .S1(n525), .Z(
        n445) );
  MUX4D0 U599 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n534), .S1(n525), .Z(
        n458) );
  MUX4D0 U600 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n535), .S1(n526), .Z(
        n471) );
  MUX4D0 U601 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n535), .S1(n526), .Z(
        n484) );
  MUX4D0 U602 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n535), .S1(n518), .Z(
        n410) );
  MUX4D0 U603 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n534), .S1(N45), .Z(
        n408) );
  MUX4D0 U604 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n533), .S1(n520), .Z(
        n421) );
  MUX4D0 U605 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n533), .S1(n518), .Z(
        n423) );
  MUX4D0 U606 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n533), .S1(n520), .Z(
        n434) );
  MUX4D0 U607 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n532), .S1(n520), .Z(
        n436) );
  MUX4D0 U608 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n534), .S1(n525), .Z(
        n449) );
  MUX4D0 U609 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n534), .S1(n525), .Z(
        n447) );
  MUX4D0 U610 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n536), .S1(n525), .Z(
        n462) );
  MUX4D0 U611 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n536), .S1(n525), .Z(
        n460) );
  MUX4D0 U612 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n535), .S1(n526), .Z(
        n473) );
  MUX4D0 U613 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n535), .S1(n526), .Z(
        n475) );
  MUX4D0 U614 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n535), .S1(n526), .Z(
        n486) );
  MUX4D0 U615 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n535), .S1(n526), .Z(
        n488) );
  MUX4ND0 U616 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(N44), .S1(n526), .ZN(
        n495) );
  MUX4ND0 U617 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n531), .S1(n516), .ZN(
        n404) );
  MUX4ND0 U618 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n535), .S1(n516), .ZN(
        n417) );
  MUX4ND0 U619 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n532), .S1(n516), .ZN(
        n430) );
  MUX4ND0 U620 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n531), .S1(n516), .ZN(
        n443) );
  MUX4ND0 U621 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n534), .S1(n519), .ZN(
        n456) );
  MUX4ND0 U622 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(N44), .S1(n519), .ZN(
        n469) );
  MUX4ND0 U623 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n531), .S1(n520), .ZN(
        n482) );
  MUX4D0 U624 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n533), .S1(n526), .Z(
        n496) );
  MUX4D0 U625 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n540), .S1(n522), .Z(n38) );
  MUX4D0 U626 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n539), .S1(n527), .Z(n51) );
  MUX4D0 U627 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n534), .S1(n528), .Z(n64) );
  MUX4D0 U628 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n533), .S1(n528), .Z(
        n119) );
  MUX4D0 U629 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n534), .S1(n529), .Z(
        n132) );
  MUX4D0 U630 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n545), .S1(n529), .Z(
        n145) );
  MUX4D0 U631 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n545), .S1(N45), .Z(n158) );
  MUX4D0 U632 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n540), .S1(n521), .Z(
        n171) );
  MUX4D0 U633 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n532), .S1(N45), .Z(n184) );
  MUX4D0 U634 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n539), .S1(n516), .Z(
        n197) );
  MUX4D0 U635 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n539), .S1(n518), .Z(
        n210) );
  MUX4D0 U636 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n540), .S1(n530), .Z(
        n223) );
  MUX4D0 U637 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n540), .S1(n524), .Z(
        n236) );
  MUX4D0 U638 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n541), .S1(n520), .Z(
        n249) );
  MUX4D0 U639 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n541), .S1(n520), .Z(
        n262) );
  MUX4D0 U640 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n542), .S1(n519), .Z(
        n275) );
  MUX4D0 U641 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n542), .S1(n525), .Z(
        n288) );
  MUX4D0 U642 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n543), .S1(n526), .Z(
        n301) );
  MUX4D0 U643 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n543), .S1(n522), .Z(
        n314) );
  MUX4D0 U644 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n544), .S1(n522), .Z(
        n327) );
  MUX4D0 U645 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n544), .S1(n523), .Z(
        n340) );
  MUX4D0 U646 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n545), .S1(n523), .Z(
        n353) );
  MUX4D0 U647 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n545), .S1(n524), .Z(
        n366) );
  MUX4D0 U648 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n546), .S1(n524), .Z(
        n379) );
  MUX4D0 U649 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n546), .S1(n519), .Z(
        n392) );
  MUX4D0 U650 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(N44), .S1(n525), .Z(
        n457) );
  MUX4D0 U651 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n535), .S1(n526), .Z(
        n483) );
  MUX4D0 U652 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n536), .S1(n527), .Z(
        n498) );
  MUX4D0 U653 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n536), .S1(n527), .Z(
        n500) );
  MUX4D0 U654 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n540), .S1(n527), .Z(n42)
         );
  MUX4D0 U655 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n539), .S1(n527), .Z(n40) );
  MUX4D0 U656 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n539), .S1(n527), .Z(n53) );
  MUX4D0 U657 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n533), .S1(n528), .Z(n55)
         );
  MUX4D0 U658 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n533), .S1(n528), .Z(
        n107) );
  MUX4D0 U659 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n542), .S1(n528), .Z(n110)
         );
  MUX4D0 U660 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(N44), .S1(n528), .Z(n123)
         );
  MUX4D0 U661 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n534), .S1(n528), .Z(
        n121) );
  MUX4D0 U662 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n533), .S1(n529), .Z(n136)
         );
  MUX4D0 U663 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(N44), .S1(n529), .Z(n134) );
  MUX4D0 U664 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n540), .S1(n529), .Z(n149)
         );
  MUX4D0 U665 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n540), .S1(n529), .Z(
        n147) );
  MUX4D0 U666 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n541), .S1(N45), .Z(n160) );
  MUX4D0 U667 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n541), .S1(n516), .Z(n162)
         );
  MUX4D0 U668 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n539), .S1(n518), .Z(
        n173) );
  MUX4D0 U669 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n539), .S1(n520), .Z(n175)
         );
  MUX4D0 U670 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n539), .S1(n520), .Z(
        n186) );
  MUX4D0 U671 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n542), .S1(n518), .Z(n188)
         );
  MUX4D0 U672 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n539), .S1(n521), .Z(n201)
         );
  MUX4D0 U673 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n539), .S1(n526), .Z(
        n199) );
  MUX4D0 U674 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n539), .S1(n530), .Z(
        n214) );
  MUX4D0 U675 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n539), .S1(n530), .Z(
        n212) );
  MUX4D0 U676 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n540), .S1(n530), .Z(
        n227) );
  MUX4D0 U677 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n540), .S1(n530), .Z(
        n225) );
  MUX4D0 U678 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n540), .S1(n523), .Z(
        n238) );
  MUX4D0 U679 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n540), .S1(n525), .Z(
        n240) );
  MUX4D0 U680 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n541), .S1(n519), .Z(
        n251) );
  MUX4D0 U681 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n541), .S1(n521), .Z(
        n253) );
  MUX4D0 U682 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n541), .S1(n521), .Z(
        n266) );
  MUX4D0 U683 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n541), .S1(n518), .Z(
        n264) );
  MUX4D0 U684 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n542), .S1(n520), .Z(
        n279) );
  MUX4D0 U685 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n542), .S1(n521), .Z(
        n277) );
  MUX4D0 U686 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n542), .S1(n516), .Z(
        n290) );
  MUX4D0 U687 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n542), .S1(n523), .Z(
        n292) );
  MUX4D0 U688 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n543), .S1(n518), .Z(
        n305) );
  MUX4D0 U689 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n543), .S1(n524), .Z(
        n303) );
  MUX4D0 U690 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n543), .S1(n522), .Z(
        n318) );
  MUX4D0 U691 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n543), .S1(n522), .Z(
        n316) );
  MUX4D0 U692 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n544), .S1(n522), .Z(
        n329) );
  MUX4D0 U693 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n544), .S1(n523), .Z(
        n331) );
  MUX4D0 U694 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n544), .S1(n523), .Z(
        n342) );
  MUX4D0 U695 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n544), .S1(n523), .Z(
        n344) );
  MUX4D0 U696 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n545), .S1(n524), .Z(
        n357) );
  MUX4D0 U697 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n545), .S1(n523), .Z(
        n355) );
  MUX4D0 U698 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n545), .S1(n524), .Z(
        n370) );
  MUX4D0 U699 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n545), .S1(n524), .Z(
        n368) );
  MUX4D0 U700 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n546), .S1(n524), .Z(
        n381) );
  MUX4D0 U701 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n546), .S1(n524), .Z(
        n383) );
  MUX4D0 U702 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(N44), .S1(n517), .Z(n396) );
  MUX4D0 U703 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n546), .S1(n519), .Z(
        n394) );
  MUX4D0 U704 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(N44), .S1(n526), .Z(
        n497) );
  MUX4D0 U705 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n546), .S1(n527), .Z(n39) );
  MUX4D0 U706 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n541), .S1(n527), .Z(n52) );
  MUX4D0 U707 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n539), .S1(n528), .Z(n65) );
  MUX4D0 U708 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(N44), .S1(n528), .Z(n120) );
  MUX4D0 U709 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n536), .S1(n529), .Z(
        n133) );
  MUX4D0 U710 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n540), .S1(n529), .Z(
        n146) );
  MUX4D0 U711 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n541), .S1(N45), .Z(n159) );
  MUX4D0 U712 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n542), .S1(n525), .Z(
        n172) );
  MUX4D0 U713 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n542), .S1(n521), .Z(
        n185) );
  MUX4D0 U714 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n539), .S1(n518), .Z(
        n198) );
  MUX4D0 U715 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n539), .S1(n521), .Z(
        n211) );
  MUX4D0 U716 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n540), .S1(n530), .Z(
        n224) );
  MUX4D0 U717 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n540), .S1(n530), .Z(
        n237) );
  MUX4D0 U718 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n541), .S1(n525), .Z(
        n250) );
  MUX4D0 U719 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n541), .S1(n530), .Z(
        n263) );
  MUX4D0 U720 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n542), .S1(n524), .Z(
        n276) );
  MUX4D0 U721 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n542), .S1(n521), .Z(
        n289) );
  MUX4D0 U722 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n543), .S1(n522), .Z(
        n302) );
  MUX4D0 U723 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n543), .S1(n522), .Z(
        n315) );
  MUX4D0 U724 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n544), .S1(n522), .Z(
        n328) );
  MUX4D0 U725 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n544), .S1(n523), .Z(
        n341) );
  MUX4D0 U726 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n545), .S1(n523), .Z(
        n354) );
  MUX4D0 U727 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n545), .S1(n524), .Z(
        n367) );
  MUX4D0 U728 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n546), .S1(n524), .Z(
        n380) );
  MUX4D0 U729 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n546), .S1(n517), .Z(
        n393) );
  MUX4D0 U730 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n534), .S1(n527), .Z(
        n499) );
  MUX4D0 U731 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n536), .S1(n527), .Z(
        n501) );
  MUX4D0 U732 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n539), .S1(n527), .Z(n43)
         );
  MUX4D0 U733 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n541), .S1(n527), .Z(n41) );
  MUX4D0 U734 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n540), .S1(n527), .Z(n54) );
  MUX4D0 U735 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n543), .S1(n528), .Z(n56)
         );
  MUX4D0 U736 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n542), .S1(n528), .Z(
        n109) );
  MUX4D0 U737 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n541), .S1(n528), .Z(n111)
         );
  MUX4D0 U738 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n532), .S1(n529), .Z(n124)
         );
  MUX4D0 U739 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n536), .S1(n528), .Z(
        n122) );
  MUX4D0 U740 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n545), .S1(n529), .Z(n137)
         );
  MUX4D0 U741 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n534), .S1(n529), .Z(
        n135) );
  MUX4D0 U742 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n542), .S1(n529), .Z(n150)
         );
  MUX4D0 U743 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n540), .S1(n529), .Z(
        n148) );
  MUX4D0 U744 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n541), .S1(n518), .Z(
        n161) );
  MUX4D0 U745 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n540), .S1(n520), .Z(n163)
         );
  MUX4D0 U746 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n542), .S1(n522), .Z(
        n174) );
  MUX4D0 U747 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n542), .S1(n523), .Z(n176)
         );
  MUX4D0 U748 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n533), .S1(n516), .Z(
        n187) );
  MUX4D0 U749 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n541), .S1(n520), .Z(n189)
         );
  MUX4D0 U750 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n539), .S1(n527), .Z(n202)
         );
  MUX4D0 U751 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n539), .S1(n520), .Z(
        n200) );
  MUX4D0 U752 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n539), .S1(n530), .Z(
        n215) );
  MUX4D0 U753 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n539), .S1(n530), .Z(
        n213) );
  MUX4D0 U754 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n540), .S1(n530), .Z(
        n228) );
  MUX4D0 U755 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n540), .S1(n530), .Z(
        n226) );
  MUX4D0 U756 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n540), .S1(n520), .Z(
        n239) );
  MUX4D0 U757 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n541), .S1(n522), .Z(
        n241) );
  MUX4D0 U758 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n541), .S1(n522), .Z(
        n252) );
  MUX4D0 U759 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n541), .S1(n524), .Z(
        n254) );
  MUX4D0 U760 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n542), .S1(n520), .Z(
        n267) );
  MUX4D0 U761 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n541), .S1(n525), .Z(
        n265) );
  MUX4D0 U762 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n542), .S1(n522), .Z(
        n280) );
  MUX4D0 U763 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n542), .S1(n527), .Z(
        n278) );
  MUX4D0 U764 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n542), .S1(n521), .Z(
        n291) );
  MUX4D0 U765 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n543), .S1(n518), .Z(
        n293) );
  MUX4D0 U766 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n543), .S1(n522), .Z(
        n306) );
  MUX4D0 U767 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n543), .S1(n530), .Z(
        n304) );
  MUX4D0 U768 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n544), .S1(n522), .Z(
        n319) );
  MUX4D0 U769 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n543), .S1(n522), .Z(
        n317) );
  MUX4D0 U770 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n544), .S1(n523), .Z(
        n330) );
  MUX4D0 U771 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n544), .S1(n523), .Z(
        n332) );
  MUX4D0 U772 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n544), .S1(n523), .Z(
        n343) );
  MUX4D0 U773 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n545), .S1(n523), .Z(
        n345) );
  MUX4D0 U774 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n545), .S1(n524), .Z(
        n358) );
  MUX4D0 U775 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n545), .S1(n523), .Z(
        n356) );
  MUX4D0 U776 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n546), .S1(n524), .Z(
        n371) );
  MUX4D0 U777 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n545), .S1(n524), .Z(
        n369) );
  MUX4D0 U778 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n546), .S1(n524), .Z(
        n382) );
  MUX4D0 U779 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n546), .S1(n519), .Z(
        n384) );
  MUX4D0 U780 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(N44), .S1(n527), .Z(n397) );
  MUX4D0 U781 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n546), .S1(n517), .Z(
        n395) );
  MUX4ND0 U782 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n532), .S1(n522), .ZN(
        n37) );
  MUX4ND0 U783 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n536), .S1(n522), .ZN(
        n50) );
  MUX4ND0 U784 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n534), .S1(n522), .ZN(
        n63) );
  MUX4ND0 U785 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n546), .S1(n529), .ZN(
        n118) );
  MUX4ND0 U786 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n533), .S1(n528), .ZN(
        n131) );
  MUX4ND0 U787 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n533), .S1(n518), .ZN(
        n144) );
  MUX4ND0 U788 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n545), .S1(n529), .ZN(
        n157) );
  MUX4ND0 U789 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n544), .S1(n529), .ZN(
        n170) );
  MUX4ND0 U790 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n533), .S1(n528), .ZN(
        n183) );
  MUX4ND0 U791 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n534), .S1(N45), .ZN(
        n196) );
  MUX4ND0 U792 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n531), .S1(n529), .ZN(
        n209) );
  MUX4ND0 U793 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n535), .S1(n523), .ZN(
        n222) );
  MUX4ND0 U794 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n544), .S1(n528), .ZN(
        n235) );
  MUX4ND0 U795 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n546), .S1(n528), .ZN(
        n248) );
  MUX4ND0 U796 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n545), .S1(n523), .ZN(
        n261) );
  MUX4ND0 U797 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n531), .S1(n529), .ZN(
        n274) );
  MUX4ND0 U798 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n544), .S1(n521), .ZN(
        n287) );
  MUX4ND0 U799 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n543), .S1(n530), .ZN(
        n300) );
  MUX4ND0 U800 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n546), .S1(n528), .ZN(
        n313) );
  MUX4ND0 U801 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(N44), .S1(n516), .ZN(
        n326) );
  MUX4ND0 U802 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(N44), .S1(n516), .ZN(
        n339) );
  MUX4ND0 U803 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(N44), .S1(n527), .ZN(
        n352) );
  MUX4ND0 U804 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n544), .S1(n519), .ZN(
        n365) );
  MUX4ND0 U805 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n543), .S1(n523), .ZN(
        n378) );
  MUX4ND0 U806 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(N44), .S1(n516), .ZN(
        n391) );
  ND3D1 U807 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U808 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U809 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U810 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U811 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U812 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U813 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U814 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U815 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U816 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  INVD1 U817 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U818 ( .I(AddrW[2]), .ZN(n105) );
  INVD1 U819 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U820 ( .I(AddrW[4]), .ZN(n102) );
  CKAN2D0 U821 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U822 ( .I0(n35), .I1(n36), .I2(n37), .S0(n517), .S1(n511), .ZN(n34)
         );
  MUX3ND0 U823 ( .I0(n44), .I1(n45), .I2(n46), .S0(n509), .S1(n506), .ZN(N82)
         );
  MUX3ND0 U824 ( .I0(n48), .I1(n49), .I2(n50), .S0(n517), .S1(n511), .ZN(n47)
         );
  MUX3ND0 U825 ( .I0(n57), .I1(n58), .I2(n59), .S0(n509), .S1(n506), .ZN(N81)
         );
  MUX3ND0 U826 ( .I0(n61), .I1(n62), .I2(n63), .S0(n529), .S1(n512), .ZN(n60)
         );
  MUX3ND0 U827 ( .I0(n112), .I1(n113), .I2(n114), .S0(n509), .S1(n506), .ZN(
        N80) );
  MUX3ND0 U828 ( .I0(n116), .I1(n117), .I2(n118), .S0(n521), .S1(n512), .ZN(
        n115) );
  MUX3ND0 U829 ( .I0(n125), .I1(n126), .I2(n127), .S0(n509), .S1(n506), .ZN(
        N79) );
  MUX3ND0 U830 ( .I0(n129), .I1(n130), .I2(n131), .S0(n524), .S1(n512), .ZN(
        n128) );
  MUX3ND0 U831 ( .I0(n138), .I1(n139), .I2(n140), .S0(n509), .S1(n506), .ZN(
        N78) );
  MUX3ND0 U832 ( .I0(n142), .I1(n143), .I2(n144), .S0(n519), .S1(n512), .ZN(
        n141) );
  MUX3ND0 U833 ( .I0(n151), .I1(n152), .I2(n153), .S0(n509), .S1(n506), .ZN(
        N77) );
  MUX3ND0 U834 ( .I0(n155), .I1(n156), .I2(n157), .S0(n522), .S1(n512), .ZN(
        n154) );
  MUX3ND0 U835 ( .I0(n164), .I1(n165), .I2(n166), .S0(n509), .S1(n506), .ZN(
        N76) );
  MUX3ND0 U836 ( .I0(n168), .I1(n169), .I2(n170), .S0(n524), .S1(n512), .ZN(
        n167) );
  MUX3ND0 U837 ( .I0(n177), .I1(n178), .I2(n179), .S0(n509), .S1(n506), .ZN(
        N75) );
  MUX3ND0 U838 ( .I0(n181), .I1(n182), .I2(n183), .S0(n527), .S1(n512), .ZN(
        n180) );
  MUX3ND0 U839 ( .I0(n190), .I1(n191), .I2(n192), .S0(n509), .S1(n506), .ZN(
        N74) );
  MUX3ND0 U840 ( .I0(n194), .I1(n195), .I2(n196), .S0(n521), .S1(n512), .ZN(
        n193) );
  MUX3ND0 U841 ( .I0(n203), .I1(n204), .I2(n205), .S0(n509), .S1(n506), .ZN(
        N73) );
  MUX3ND0 U842 ( .I0(n207), .I1(n208), .I2(n209), .S0(n525), .S1(n512), .ZN(
        n206) );
  MUX3ND0 U843 ( .I0(n216), .I1(n217), .I2(n218), .S0(n509), .S1(n506), .ZN(
        N72) );
  MUX3ND0 U844 ( .I0(n220), .I1(n221), .I2(n222), .S0(n527), .S1(n512), .ZN(
        n219) );
  MUX3ND0 U845 ( .I0(n229), .I1(n230), .I2(n231), .S0(n509), .S1(n506), .ZN(
        N71) );
  MUX3ND0 U846 ( .I0(n233), .I1(n234), .I2(n235), .S0(n518), .S1(n512), .ZN(
        n232) );
  MUX3ND0 U847 ( .I0(n242), .I1(n243), .I2(n244), .S0(n509), .S1(n506), .ZN(
        N70) );
  MUX3ND0 U848 ( .I0(n246), .I1(n247), .I2(n248), .S0(n529), .S1(n512), .ZN(
        n245) );
  MUX3ND0 U849 ( .I0(n255), .I1(n256), .I2(n257), .S0(n508), .S1(n506), .ZN(
        N69) );
  MUX3ND0 U850 ( .I0(n259), .I1(n260), .I2(n261), .S0(n520), .S1(n512), .ZN(
        n258) );
  MUX3ND0 U851 ( .I0(n268), .I1(n269), .I2(n270), .S0(n508), .S1(n506), .ZN(
        N68) );
  MUX3ND0 U852 ( .I0(n272), .I1(n273), .I2(n274), .S0(n526), .S1(n513), .ZN(
        n271) );
  MUX3ND0 U853 ( .I0(n281), .I1(n282), .I2(n283), .S0(n508), .S1(n506), .ZN(
        N67) );
  MUX3ND0 U854 ( .I0(n285), .I1(n286), .I2(n287), .S0(n516), .S1(n513), .ZN(
        n284) );
  MUX3ND0 U855 ( .I0(n294), .I1(n295), .I2(n296), .S0(n508), .S1(n506), .ZN(
        N66) );
  MUX3ND0 U856 ( .I0(n298), .I1(n299), .I2(n300), .S0(n519), .S1(n513), .ZN(
        n297) );
  MUX3ND0 U857 ( .I0(n307), .I1(n308), .I2(n309), .S0(n508), .S1(n506), .ZN(
        N65) );
  MUX3ND0 U858 ( .I0(n311), .I1(n312), .I2(n313), .S0(n525), .S1(n513), .ZN(
        n310) );
  MUX3ND0 U859 ( .I0(n320), .I1(n321), .I2(n322), .S0(n508), .S1(n506), .ZN(
        N64) );
  MUX3ND0 U860 ( .I0(n324), .I1(n325), .I2(n326), .S0(n516), .S1(n513), .ZN(
        n323) );
  MUX3ND0 U861 ( .I0(n333), .I1(n334), .I2(n335), .S0(n508), .S1(n506), .ZN(
        N63) );
  MUX3ND0 U862 ( .I0(n337), .I1(n338), .I2(n339), .S0(n524), .S1(n513), .ZN(
        n336) );
  MUX3ND0 U863 ( .I0(n346), .I1(n347), .I2(n348), .S0(n508), .S1(N48), .ZN(N62) );
  MUX3ND0 U864 ( .I0(n350), .I1(n351), .I2(n352), .S0(n528), .S1(n513), .ZN(
        n349) );
  MUX3ND0 U865 ( .I0(n359), .I1(n360), .I2(n361), .S0(n508), .S1(N48), .ZN(N61) );
  MUX3ND0 U866 ( .I0(n363), .I1(n364), .I2(n365), .S0(n527), .S1(n513), .ZN(
        n362) );
  MUX3ND0 U867 ( .I0(n372), .I1(n373), .I2(n374), .S0(n508), .S1(N48), .ZN(N60) );
  MUX3ND0 U868 ( .I0(n376), .I1(n377), .I2(n378), .S0(n523), .S1(n513), .ZN(
        n375) );
  MUX3ND0 U869 ( .I0(n385), .I1(n386), .I2(n387), .S0(n508), .S1(N48), .ZN(N59) );
  MUX3ND0 U870 ( .I0(n389), .I1(n390), .I2(n391), .S0(n528), .S1(n513), .ZN(
        n388) );
  MUX3ND0 U871 ( .I0(n398), .I1(n399), .I2(n400), .S0(n508), .S1(N48), .ZN(N58) );
  MUX3ND0 U872 ( .I0(n402), .I1(n403), .I2(n404), .S0(n519), .S1(n513), .ZN(
        n401) );
  MUX3ND0 U873 ( .I0(n411), .I1(n412), .I2(n413), .S0(n508), .S1(N48), .ZN(N57) );
  MUX3ND0 U874 ( .I0(n415), .I1(n416), .I2(n417), .S0(n521), .S1(n513), .ZN(
        n414) );
  MUX3ND0 U875 ( .I0(n424), .I1(n425), .I2(n426), .S0(n508), .S1(N48), .ZN(N56) );
  MUX3ND0 U876 ( .I0(n428), .I1(n429), .I2(n430), .S0(n521), .S1(n513), .ZN(
        n427) );
  MUX3ND0 U877 ( .I0(n437), .I1(n438), .I2(n439), .S0(n508), .S1(N48), .ZN(N55) );
  MUX3ND0 U878 ( .I0(n441), .I1(n442), .I2(n443), .S0(n521), .S1(n511), .ZN(
        n440) );
  MUX3ND0 U879 ( .I0(n450), .I1(n451), .I2(n452), .S0(n508), .S1(N48), .ZN(N54) );
  MUX3ND0 U880 ( .I0(n454), .I1(n455), .I2(n456), .S0(n516), .S1(n511), .ZN(
        n453) );
  MUX3ND0 U881 ( .I0(n463), .I1(n464), .I2(n465), .S0(N47), .S1(N48), .ZN(N53)
         );
  MUX3ND0 U882 ( .I0(n467), .I1(n468), .I2(n469), .S0(n521), .S1(n511), .ZN(
        n466) );
  MUX3ND0 U883 ( .I0(n476), .I1(n477), .I2(n478), .S0(n508), .S1(N48), .ZN(N52) );
  MUX3ND0 U884 ( .I0(n480), .I1(n481), .I2(n482), .S0(n516), .S1(n916), .ZN(
        n479) );
  MUX3ND0 U885 ( .I0(n489), .I1(n490), .I2(n491), .S0(N47), .S1(N48), .ZN(N51)
         );
  MUX3ND0 U886 ( .I0(n493), .I1(n494), .I2(n495), .S0(n521), .S1(n512), .ZN(
        n492) );
  MUX3ND0 U887 ( .I0(n502), .I1(n503), .I2(n504), .S0(n507), .S1(N48), .ZN(N50) );
  MUX2ND0 U888 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n536), .ZN(
        n36) );
  MUX2ND0 U889 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n536), .ZN(
        n35) );
  MUX3ND0 U890 ( .I0(n39), .I1(n38), .I2(n34), .S0(n515), .S1(n509), .ZN(n46)
         );
  MUX2ND0 U891 ( .I0(n41), .I1(n40), .S(n510), .ZN(n45) );
  MUX2ND0 U892 ( .I0(n43), .I1(n42), .S(N46), .ZN(n44) );
  MUX2ND0 U893 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n537), .ZN(
        n49) );
  MUX2ND0 U894 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n537), .ZN(
        n48) );
  MUX3ND0 U895 ( .I0(n52), .I1(n51), .I2(n47), .S0(n515), .S1(n509), .ZN(n59)
         );
  MUX2ND0 U896 ( .I0(n54), .I1(n53), .S(n510), .ZN(n58) );
  MUX2ND0 U897 ( .I0(n56), .I1(n55), .S(n514), .ZN(n57) );
  MUX2ND0 U898 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n537), .ZN(
        n62) );
  MUX2ND0 U899 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n537), .ZN(
        n61) );
  MUX3ND0 U900 ( .I0(n65), .I1(n64), .I2(n60), .S0(n515), .S1(n509), .ZN(n114)
         );
  MUX2ND0 U901 ( .I0(n109), .I1(n107), .S(n510), .ZN(n113) );
  MUX2ND0 U902 ( .I0(n111), .I1(n110), .S(n916), .ZN(n112) );
  MUX2ND0 U903 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n537), .ZN(
        n117) );
  MUX2ND0 U904 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n538), .ZN(
        n116) );
  MUX3ND0 U905 ( .I0(n120), .I1(n119), .I2(n115), .S0(n515), .S1(n509), .ZN(
        n127) );
  MUX2ND0 U906 ( .I0(n122), .I1(n121), .S(n916), .ZN(n126) );
  MUX2ND0 U907 ( .I0(n124), .I1(n123), .S(N46), .ZN(n125) );
  MUX2ND0 U908 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n538), .ZN(
        n130) );
  MUX2ND0 U909 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n538), .ZN(
        n129) );
  MUX3ND0 U910 ( .I0(n133), .I1(n132), .I2(n128), .S0(n515), .S1(n509), .ZN(
        n140) );
  MUX2ND0 U911 ( .I0(n135), .I1(n134), .S(n916), .ZN(n139) );
  MUX2ND0 U912 ( .I0(n137), .I1(n136), .S(n916), .ZN(n138) );
  MUX2ND0 U913 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n538), .ZN(
        n143) );
  MUX2ND0 U914 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n543), .ZN(
        n142) );
  MUX3ND0 U915 ( .I0(n146), .I1(n145), .I2(n141), .S0(n514), .S1(n509), .ZN(
        n153) );
  MUX2ND0 U916 ( .I0(n148), .I1(n147), .S(N46), .ZN(n152) );
  MUX2ND0 U917 ( .I0(n150), .I1(n149), .S(N46), .ZN(n151) );
  MUX2ND0 U918 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n544), .ZN(
        n156) );
  MUX2ND0 U919 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n543), .ZN(
        n155) );
  MUX3ND0 U920 ( .I0(n159), .I1(n158), .I2(n154), .S0(n514), .S1(n507), .ZN(
        n166) );
  MUX2ND0 U921 ( .I0(n161), .I1(n160), .S(N46), .ZN(n165) );
  MUX2ND0 U922 ( .I0(n163), .I1(n162), .S(N46), .ZN(n164) );
  MUX2ND0 U923 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n531), .ZN(
        n169) );
  MUX2ND0 U924 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n533), .ZN(
        n168) );
  MUX3ND0 U925 ( .I0(n172), .I1(n171), .I2(n167), .S0(n510), .S1(n507), .ZN(
        n179) );
  MUX2ND0 U926 ( .I0(n174), .I1(n173), .S(n515), .ZN(n178) );
  MUX2ND0 U927 ( .I0(n176), .I1(n175), .S(n512), .ZN(n177) );
  MUX2ND0 U928 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n544), .ZN(
        n182) );
  MUX2ND0 U929 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n546), .ZN(
        n181) );
  MUX3ND0 U930 ( .I0(n185), .I1(n184), .I2(n180), .S0(n515), .S1(n507), .ZN(
        n192) );
  MUX2ND0 U931 ( .I0(n187), .I1(n186), .S(N46), .ZN(n191) );
  MUX2ND0 U932 ( .I0(n189), .I1(n188), .S(N46), .ZN(n190) );
  MUX2ND0 U933 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n544), .ZN(
        n195) );
  MUX2ND0 U934 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n543), .ZN(
        n194) );
  MUX3ND0 U935 ( .I0(n198), .I1(n197), .I2(n193), .S0(n514), .S1(n507), .ZN(
        n205) );
  MUX2ND0 U936 ( .I0(n200), .I1(n199), .S(N46), .ZN(n204) );
  MUX2ND0 U937 ( .I0(n202), .I1(n201), .S(n511), .ZN(n203) );
  MUX2ND0 U938 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n546), 
        .ZN(n208) );
  MUX2ND0 U939 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n533), 
        .ZN(n207) );
  MUX3ND0 U940 ( .I0(n211), .I1(n210), .I2(n206), .S0(n510), .S1(n507), .ZN(
        n218) );
  MUX2ND0 U941 ( .I0(n213), .I1(n212), .S(n512), .ZN(n217) );
  MUX2ND0 U942 ( .I0(n215), .I1(n214), .S(n510), .ZN(n216) );
  MUX2ND0 U943 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n536), 
        .ZN(n221) );
  MUX2ND0 U944 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n536), 
        .ZN(n220) );
  MUX3ND0 U945 ( .I0(n224), .I1(n223), .I2(n219), .S0(n510), .S1(n507), .ZN(
        n231) );
  MUX2ND0 U946 ( .I0(n226), .I1(n225), .S(n510), .ZN(n230) );
  MUX2ND0 U947 ( .I0(n228), .I1(n227), .S(n514), .ZN(n229) );
  MUX2ND0 U948 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n545), 
        .ZN(n234) );
  MUX2ND0 U949 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n543), 
        .ZN(n233) );
  MUX3ND0 U950 ( .I0(n237), .I1(n236), .I2(n232), .S0(n514), .S1(n507), .ZN(
        n244) );
  MUX2ND0 U951 ( .I0(n239), .I1(n238), .S(n512), .ZN(n243) );
  MUX2ND0 U952 ( .I0(n241), .I1(n240), .S(n510), .ZN(n242) );
  MUX2ND0 U953 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n535), 
        .ZN(n247) );
  MUX2ND0 U954 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n544), 
        .ZN(n246) );
  MUX3ND0 U955 ( .I0(n250), .I1(n249), .I2(n245), .S0(n514), .S1(n507), .ZN(
        n257) );
  MUX2ND0 U956 ( .I0(n252), .I1(n251), .S(n510), .ZN(n256) );
  MUX2ND0 U957 ( .I0(n254), .I1(n253), .S(n515), .ZN(n255) );
  MUX2ND0 U958 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n533), 
        .ZN(n260) );
  MUX2ND0 U959 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n533), 
        .ZN(n259) );
  MUX3ND0 U960 ( .I0(n263), .I1(n262), .I2(n258), .S0(n510), .S1(n507), .ZN(
        n270) );
  MUX2ND0 U961 ( .I0(n265), .I1(n264), .S(n510), .ZN(n269) );
  MUX2ND0 U962 ( .I0(n267), .I1(n266), .S(n511), .ZN(n268) );
  MUX2ND0 U963 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n543), 
        .ZN(n273) );
  MUX2ND0 U964 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n531), 
        .ZN(n272) );
  MUX3ND0 U965 ( .I0(n276), .I1(n275), .I2(n271), .S0(n510), .S1(n507), .ZN(
        n283) );
  MUX2ND0 U966 ( .I0(n278), .I1(n277), .S(n511), .ZN(n282) );
  MUX2ND0 U967 ( .I0(n280), .I1(n279), .S(n916), .ZN(n281) );
  MUX2ND0 U968 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n535), 
        .ZN(n286) );
  MUX2ND0 U969 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n538), 
        .ZN(n285) );
  MUX3ND0 U970 ( .I0(n289), .I1(n288), .I2(n284), .S0(n514), .S1(n507), .ZN(
        n296) );
  MUX2ND0 U971 ( .I0(n291), .I1(n290), .S(n916), .ZN(n295) );
  MUX2ND0 U972 ( .I0(n293), .I1(n292), .S(N46), .ZN(n294) );
  MUX2ND0 U973 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n538), 
        .ZN(n299) );
  MUX2ND0 U974 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n538), 
        .ZN(n298) );
  MUX3ND0 U975 ( .I0(n302), .I1(n301), .I2(n297), .S0(n514), .S1(n507), .ZN(
        n309) );
  MUX2ND0 U976 ( .I0(n304), .I1(n303), .S(n510), .ZN(n308) );
  MUX2ND0 U977 ( .I0(n306), .I1(n305), .S(n514), .ZN(n307) );
  MUX2ND0 U978 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n538), 
        .ZN(n312) );
  MUX2ND0 U979 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n538), 
        .ZN(n311) );
  MUX3ND0 U980 ( .I0(n315), .I1(n314), .I2(n310), .S0(n514), .S1(n507), .ZN(
        n322) );
  MUX2ND0 U981 ( .I0(n317), .I1(n316), .S(n513), .ZN(n321) );
  MUX2ND0 U982 ( .I0(n319), .I1(n318), .S(n513), .ZN(n320) );
  MUX2ND0 U983 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n538), 
        .ZN(n325) );
  MUX2ND0 U984 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n538), 
        .ZN(n324) );
  MUX3ND0 U985 ( .I0(n328), .I1(n327), .I2(n323), .S0(n916), .S1(n508), .ZN(
        n335) );
  MUX2ND0 U986 ( .I0(n330), .I1(n329), .S(n511), .ZN(n334) );
  MUX2ND0 U987 ( .I0(n332), .I1(n331), .S(n511), .ZN(n333) );
  MUX2ND0 U988 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n538), 
        .ZN(n338) );
  MUX2ND0 U989 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n538), 
        .ZN(n337) );
  MUX3ND0 U990 ( .I0(n341), .I1(n340), .I2(n336), .S0(n514), .S1(N47), .ZN(
        n348) );
  MUX2ND0 U991 ( .I0(n343), .I1(n342), .S(n513), .ZN(n347) );
  MUX2ND0 U992 ( .I0(n345), .I1(n344), .S(n513), .ZN(n346) );
  MUX2ND0 U993 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n538), 
        .ZN(n351) );
  MUX2ND0 U994 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n538), 
        .ZN(n350) );
  MUX3ND0 U995 ( .I0(n354), .I1(n353), .I2(n349), .S0(n515), .S1(N47), .ZN(
        n361) );
  MUX2ND0 U996 ( .I0(n356), .I1(n355), .S(n511), .ZN(n360) );
  MUX2ND0 U997 ( .I0(n358), .I1(n357), .S(n511), .ZN(n359) );
  MUX2ND0 U998 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n538), 
        .ZN(n364) );
  MUX2ND0 U999 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n538), 
        .ZN(n363) );
  MUX3ND0 U1000 ( .I0(n367), .I1(n366), .I2(n362), .S0(n515), .S1(N47), .ZN(
        n374) );
  MUX2ND0 U1001 ( .I0(n369), .I1(n368), .S(n510), .ZN(n373) );
  MUX2ND0 U1002 ( .I0(n371), .I1(n370), .S(n513), .ZN(n372) );
  MUX2ND0 U1003 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n538), 
        .ZN(n377) );
  MUX2ND0 U1004 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n538), 
        .ZN(n376) );
  MUX3ND0 U1005 ( .I0(n380), .I1(n379), .I2(n375), .S0(n514), .S1(N47), .ZN(
        n387) );
  MUX2ND0 U1006 ( .I0(n382), .I1(n381), .S(n512), .ZN(n386) );
  MUX2ND0 U1007 ( .I0(n384), .I1(n383), .S(n510), .ZN(n385) );
  MUX2ND0 U1008 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n538), 
        .ZN(n390) );
  MUX2ND0 U1009 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n537), 
        .ZN(n389) );
  MUX3ND0 U1010 ( .I0(n393), .I1(n392), .I2(n388), .S0(n514), .S1(N47), .ZN(
        n400) );
  MUX2ND0 U1011 ( .I0(n395), .I1(n394), .S(n916), .ZN(n399) );
  MUX2ND0 U1012 ( .I0(n397), .I1(n396), .S(n916), .ZN(n398) );
  MUX2ND0 U1013 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n537), 
        .ZN(n403) );
  MUX2ND0 U1014 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n537), 
        .ZN(n402) );
  MUX3ND0 U1015 ( .I0(n406), .I1(n405), .I2(n401), .S0(n514), .S1(n508), .ZN(
        n413) );
  MUX2ND0 U1016 ( .I0(n408), .I1(n407), .S(n511), .ZN(n412) );
  MUX2ND0 U1017 ( .I0(n410), .I1(n409), .S(n511), .ZN(n411) );
  MUX2ND0 U1018 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n537), 
        .ZN(n416) );
  MUX2ND0 U1019 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n537), 
        .ZN(n415) );
  MUX3ND0 U1020 ( .I0(n419), .I1(n418), .I2(n414), .S0(n515), .S1(n508), .ZN(
        n426) );
  MUX2ND0 U1021 ( .I0(n421), .I1(n420), .S(n510), .ZN(n425) );
  MUX2ND0 U1022 ( .I0(n423), .I1(n422), .S(n513), .ZN(n424) );
  MUX2ND0 U1023 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n537), 
        .ZN(n429) );
  MUX2ND0 U1024 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n537), 
        .ZN(n428) );
  MUX3ND0 U1025 ( .I0(n432), .I1(n431), .I2(n427), .S0(n514), .S1(N47), .ZN(
        n439) );
  MUX2ND0 U1026 ( .I0(n434), .I1(n433), .S(n511), .ZN(n438) );
  MUX2ND0 U1027 ( .I0(n436), .I1(n435), .S(n511), .ZN(n437) );
  MUX2ND0 U1028 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n537), 
        .ZN(n442) );
  MUX2ND0 U1029 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n537), 
        .ZN(n441) );
  MUX3ND0 U1030 ( .I0(n445), .I1(n444), .I2(n440), .S0(n515), .S1(N47), .ZN(
        n452) );
  MUX2ND0 U1031 ( .I0(n447), .I1(n446), .S(n916), .ZN(n451) );
  MUX2ND0 U1032 ( .I0(n449), .I1(n448), .S(n511), .ZN(n450) );
  MUX2ND0 U1033 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n537), 
        .ZN(n455) );
  MUX2ND0 U1034 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n537), 
        .ZN(n454) );
  MUX3ND0 U1035 ( .I0(n458), .I1(n457), .I2(n453), .S0(n515), .S1(N47), .ZN(
        n465) );
  MUX2ND0 U1036 ( .I0(n460), .I1(n459), .S(n916), .ZN(n464) );
  MUX2ND0 U1037 ( .I0(n462), .I1(n461), .S(n916), .ZN(n463) );
  MUX2ND0 U1038 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n537), 
        .ZN(n468) );
  MUX2ND0 U1039 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n537), 
        .ZN(n467) );
  MUX3ND0 U1040 ( .I0(n471), .I1(n470), .I2(n466), .S0(n515), .S1(N47), .ZN(
        n478) );
  MUX2ND0 U1041 ( .I0(n473), .I1(n472), .S(n513), .ZN(n477) );
  MUX2ND0 U1042 ( .I0(n475), .I1(n474), .S(n511), .ZN(n476) );
  MUX2ND0 U1043 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n537), 
        .ZN(n481) );
  MUX2ND0 U1044 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n537), 
        .ZN(n480) );
  MUX3ND0 U1045 ( .I0(n484), .I1(n483), .I2(n479), .S0(n515), .S1(N47), .ZN(
        n491) );
  MUX2ND0 U1046 ( .I0(n486), .I1(n485), .S(n511), .ZN(n490) );
  MUX2ND0 U1047 ( .I0(n488), .I1(n487), .S(n511), .ZN(n489) );
  MUX2ND0 U1048 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n536), 
        .ZN(n494) );
  MUX2ND0 U1049 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n534), 
        .ZN(n493) );
  MUX3ND0 U1050 ( .I0(n497), .I1(n496), .I2(n492), .S0(n515), .S1(n507), .ZN(
        n504) );
  MUX2ND0 U1051 ( .I0(n499), .I1(n498), .S(n512), .ZN(n503) );
  MUX2ND0 U1052 ( .I0(n501), .I1(n500), .S(n512), .ZN(n502) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] , n1;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(n1), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  INVD0 U1 ( .I(SUM[0]), .ZN(n1) );
  INVD0 U2 ( .I(A[0]), .ZN(SUM[0]) );
  CKXOR2D0 U3 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
endmodule

