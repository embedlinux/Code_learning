
`ifndef RKV_I2C_USER_ELEMENT_SEQUENCES_SVH
`define RKV_I2C_USER_ELEMENT_SEQUENCES_SVH


`endif // RKV_I2C_USER_ELEMENT_SEQUENCES_SVH

