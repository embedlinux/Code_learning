
module FullDup ( OutParDataA, OutParDataB, InParDataA, InParDataB, InParValidA, 
        InParValidB, ClockA, ClockB, Reset, tms, tdi, tdo );
  output [31:0] OutParDataA;
  output [31:0] OutParDataB;
  input [31:0] InParDataA;
  input [31:0] InParDataB;
  input InParValidA, InParValidB, ClockA, ClockB, Reset, tms, tdi;
  output tdo;
  wire   n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, \SerDes_U1/Rx_ParClk ,
         \SerDes_U1/Tx_SerClk , \SerDes_U1/Tx_F_Full , \SerDes_U1/Tx_F_Empty ,
         \SerDes_U1/SerLineValid , \SerDes_U1/Des_U1/SerRxToDecode ,
         \SerDes_U1/Des_U1/SerialClk , \SerDes_U1/Des_U1/ParValidDecode ,
         \SerDes_U2/Rx_ParClk , \SerDes_U2/Tx_SerClk , \SerDes_U2/Tx_F_Full ,
         \SerDes_U2/Tx_F_Empty , \SerDes_U2/SerLineValid ,
         \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ,
         \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N84 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N82 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N80 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N78 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N76 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N74 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N72 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N70 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N68 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N66 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N64 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N62 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N60 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N58 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N56 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N54 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N28 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N26 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N24 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N83 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N81 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N79 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N77 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N75 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N73 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N71 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N69 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N67 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N65 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N63 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N61 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N59 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N57 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N55 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N53 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N29 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N27 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N25 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N24 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N23 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 , \SerDes_U2/Des_U1/SerRxToDecode ,
         \SerDes_U2/Des_U1/SerialClk , \SerDes_U2/Des_U1/ParValidDecode ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ,
         \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ,
         \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N79 , \SerDes_U1/Des_U1/DesDec_Rx1/N47 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N43 , \SerDes_U1/Des_U1/DesDec_Rx1/N42 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N41 , \SerDes_U1/Des_U1/DesDec_Rx1/N40 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N39 , \SerDes_U1/Des_U1/DesDec_Rx1/N38 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N37 , \SerDes_U1/Des_U1/DesDec_Rx1/N34 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N33 , \SerDes_U1/Des_U1/DesDec_Rx1/N32 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N31 , \SerDes_U1/Des_U1/DesDec_Rx1/N30 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[63] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ,
         \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[0] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[1] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[2] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[3] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N79 , \SerDes_U2/Des_U1/DesDec_Rx1/N47 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N43 , \SerDes_U2/Des_U1/DesDec_Rx1/N42 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N41 , \SerDes_U2/Des_U1/DesDec_Rx1/N40 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N39 , \SerDes_U2/Des_U1/DesDec_Rx1/N38 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N37 , \SerDes_U2/Des_U1/DesDec_Rx1/N34 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N33 , \SerDes_U2/Des_U1/DesDec_Rx1/N32 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N31 , \SerDes_U2/Des_U1/DesDec_Rx1/N30 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[63] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ,
         \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[0] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[1] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[2] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[3] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 , n712, n713, n714,
         n715, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n837, n841,
         n842, n849, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n985, n989,
         n990, n997, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1030, n1031,
         n1032, n1033, n1035, n1036, n1048, n1050, n1052, n1310, n1312, n1314,
         n1319, n1324, n1327, n1394, n1397, n1399, n1401, n1403, n1417, n1419,
         n1421, n1423, n1425, n1427, n1429, n1431, n1433, n1435, n1437, n1439,
         n1441, n1443, n1445, n1447, n1449, n1451, n1453, n1455, n1457, n1459,
         n1461, n1463, n1465, n1467, n1469, n1471, n1473, n1475, n1477, n1479,
         n1481, n1483, n1485, n1487, n1491, n1493, n1495, n1497, n1499, n1501,
         n1503, n1505, n1507, n1509, n1511, n1513, n1515, n1517, n1519, n1521,
         n1523, n1525, n1527, n1529, n1531, n1533, n1535, n1537, n1539, n1541,
         n1543, n1545, n1547, n1549, n1551, n1553, n1619, n1623, n1625, n1646,
         n1650, n1652, n1655, n1672, n1674, n1676, n1678, n2192, n2194, n2196,
         n2198, n2204, n2207, n2213, n2280, n2283, n2285, n2287, n2289, n2303,
         n2305, n2307, n2309, n2311, n2313, n2315, n2317, n2319, n2321, n2323,
         n2325, n2327, n2329, n2331, n2333, n2335, n2337, n2339, n2341, n2343,
         n2345, n2347, n2349, n2351, n2353, n2355, n2357, n2359, n2361, n2363,
         n2365, n2367, n2369, n2371, n2373, n2377, n2379, n2381, n2383, n2385,
         n2387, n2389, n2391, n2393, n2395, n2397, n2399, n2401, n2403, n2405,
         n2407, n2409, n2411, n2413, n2415, n2417, n2419, n2421, n2423, n2425,
         n2427, n2429, n2431, n2433, n2435, n2437, n2439, n2505, n2509, n2511,
         n2532, n2536, n2538, n2541, n2549, n2553, n2876, n2878, n2880, n2882,
         n2884, n2886, n2888, n2893, n2896, n2901, n2904, n2906, n2909, n2945,
         n2947, n2949, n2951, n2953, n3467, n3469, n3471, n3473, n3479, n3482,
         n3485, n3523, n3526, n3528, n3530, n1037, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3594,
         n3595, n3597, n3598, n3600, n3601, n3603, n3604, n3606, n3607, n3609,
         n3610, n3612, n3613, n3615, n3616, n3618, n3619, n3621, n3622, n3624,
         n3625, n3627, n3628, n3630, n3631, n3633, n3634, n3636, n3637, n3639,
         n3640, n3642, n3643, n3645, n3646, n3648, n3649, n3651, n3652, n3654,
         n3655, n3657, n3658, n3660, n3661, n3663, n3664, n3666, n3667, n3669,
         n3670, n3672, n3673, n3675, n3676, n3678, n3679, n3681, n3682, n3684,
         n3685, n3687, n3688, n3690, n3692, n3694, n3696, n3698, n3700, n3702,
         n3704, n3706, n3708, n3710, n3712, n3714, n3716, n3718, n3720, n3722,
         n3724, n3726, n3728, n3730, n3732, n3734, n3736, n3738, n3740, n3742,
         n3744, n3746, n3748, n3750, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124;
  wire   [31:0] \SerDes_U1/Des_U1/DecodeToFIFO ;
  wire   [3:0] \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr ;
  wire   [3:0] \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState ;
  wire   [2:0] \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState ;
  wire   [31:0] \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr ;
  wire   [31:0] \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr ;
  wire   [31:0] \SerDes_U2/Des_U1/DecodeToFIFO ;
  wire   [2:0] \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState ;
  wire   [2:0] \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState ;
  wire   [31:0] \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr ;
  wire   [31:0] \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr ;
  wire   [31:0] \SerDes_U1/Des_U1/DesDec_Rx1/Decoder ;
  wire   [31:0] \SerDes_U2/Des_U1/DesDec_Rx1/Decoder ;
  wire   [1:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq ;
  wire   [1:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq ;
  wire   [1:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq ;
  wire   [1:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq ;
  wire   [5:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD ;
  wire   [3:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr ;

  DEL005 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleDelay1  ( .I(ClockA), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleDelay1  ( .I(
        \SerDes_U1/Rx_ParClk ), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleDelay1  ( .I(ClockB), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleDelay1  ( .I(
        \SerDes_U2/Rx_ParClk ), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]) );
  CKND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/I_2  ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/I_2  ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/I_2  ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/I_2  ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]) );
  FullDup_DW01_inc_0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/add_16  ( .A(
        {\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/add_16  ( .A(
        {\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_2 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/add_16  ( .A(
        {\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_3 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/add_16  ( .A(
        {\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 }) );
  FullDup_DW01_dec_0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 }) );
  FullDup_DW01_inc_4 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 }) );
  FullDup_DW01_inc_5 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 }) );
  FullDup_DW01_dec_1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 }) );
  FullDup_DW01_inc_6 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 }) );
  FullDup_DW01_inc_7 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 }) );
  FullDup_DW01_dec_2 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 }) );
  FullDup_DW01_inc_8 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 }) );
  FullDup_DW01_inc_9 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 }) );
  FullDup_DW01_dec_3 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 }) );
  FullDup_DW01_inc_10 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 }) );
  FullDup_DW01_inc_11 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 }) );
  FullDup_DW01_inc_12 \SerDes_U2/Des_U1/DesDec_Rx1/ClkGen/add_206  ( .A({
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] }), .SUM({
        \SerDes_U2/Des_U1/DesDec_Rx1/N34 , \SerDes_U2/Des_U1/DesDec_Rx1/N33 , 
        \SerDes_U2/Des_U1/DesDec_Rx1/N32 , \SerDes_U2/Des_U1/DesDec_Rx1/N31 , 
        \SerDes_U2/Des_U1/DesDec_Rx1/N30 }) );
  FullDup_DW01_inc_13 \SerDes_U1/Des_U1/DesDec_Rx1/ClkGen/add_206  ( .A({
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] }), .SUM({
        \SerDes_U1/Des_U1/DesDec_Rx1/N34 , \SerDes_U1/Des_U1/DesDec_Rx1/N33 , 
        \SerDes_U1/Des_U1/DesDec_Rx1/N32 , \SerDes_U1/Des_U1/DesDec_Rx1/N31 , 
        \SerDes_U1/Des_U1/DesDec_Rx1/N30 }) );
  FullDup_DW01_dec_4 \SerDes_U2/Ser_U1/SerEnc_Tx1/ShifterBlock/sub_132  ( .A({
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 }), .SUM({
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 })
         );
  FullDup_DW01_dec_5 \SerDes_U1/Ser_U1/SerEnc_Tx1/ShifterBlock/sub_132  ( .A({
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 }), .SUM({
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 })
         );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[31]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]), .SI(n3684), .SE(
        n1037), .CP(ClockA), .CDN(n4415), .Q(n5125) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[30]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]), .SI(n3678), .SE(
        n1037), .CP(ClockA), .CDN(n4390), .Q(n5126) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[29]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]), .SI(n3672), .SE(
        n1037), .CP(ClockA), .CDN(n4442), .Q(n5127) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[28]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]), .SI(n3666), .SE(
        n1037), .CP(ClockA), .CDN(n3530), .Q(n5128) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[27]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]), .SI(n3660), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(n5129) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[26]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]), .SI(n3654), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(n5130) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[25]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]), .SI(n3648), .SE(
        n1037), .CP(ClockA), .CDN(n4389), .Q(n5131) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[24]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]), .SI(n3642), .SE(
        n1037), .CP(ClockA), .CDN(n4452), .Q(n5132) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[23]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]), .SI(n3636), .SE(
        n1037), .CP(ClockA), .CDN(n4427), .Q(n5133) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[22]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]), .SI(n3630), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(n5134) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[21]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]), .SI(n3624), .SE(
        n1037), .CP(ClockA), .CDN(n4457), .Q(n5135) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[20]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]), .SI(n3618), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(n5136) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[19]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]), .SI(n3612), .SE(
        n1037), .CP(ClockA), .CDN(n4374), .Q(n5137) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[18]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]), .SI(n3606), .SE(
        n1037), .CP(ClockA), .CDN(n4374), .Q(n5138) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[17]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]), .SI(n3600), .SE(
        n1037), .CP(ClockA), .CDN(n4376), .Q(n5139) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[16]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]), .SI(n3594), .SE(
        n1037), .CP(ClockA), .CDN(n4383), .Q(n5140) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[15]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]), .SI(n3597), .SE(
        n1037), .CP(ClockA), .CDN(n4414), .Q(n5141) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[14]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]), .SI(n3603), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(n5142) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[13]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]), .SI(n3609), .SE(
        n1037), .CP(ClockA), .CDN(n4457), .Q(n5143) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[12]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]), .SI(n3615), .SE(
        n1037), .CP(ClockA), .CDN(n4420), .Q(n5144) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[11]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]), .SI(n3621), .SE(
        n1037), .CP(ClockA), .CDN(n4429), .Q(n5145) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[10]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]), .SI(n3627), .SE(
        n1037), .CP(ClockA), .CDN(n4374), .Q(n5146) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[9]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]), .SI(n3633), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(n5147) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[8]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]), .SI(n3639), .SE(
        n1037), .CP(ClockA), .CDN(n4385), .Q(n5148) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[7]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]), .SI(n3645), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(n5149) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[6]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]), .SI(n3651), .SE(
        n1037), .CP(ClockA), .CDN(n4419), .Q(n5150) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[5]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]), .SI(n3657), .SE(
        n1037), .CP(ClockA), .CDN(n4379), .Q(n5151) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[4]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]), .SI(n3663), .SE(
        n1037), .CP(ClockA), .CDN(n4442), .Q(n5152) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[3]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]), .SI(n3669), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(n5153) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]), .SI(n3675), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(n5154) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]), .SI(n3681), .SE(
        n1037), .CP(ClockA), .CDN(n4447), .Q(n5155) );
  SDFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]), .SI(n3687), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(n5156) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[31]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]), .SI(n5157), .SE(
        n1037), .CP(ClockB), .CDN(n4416), .Q(n5157) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[30]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]), .SI(n5158), .SE(
        n1037), .CP(ClockB), .CDN(n4412), .Q(n5158) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[29]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]), .SI(n5159), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(n5159) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[28]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]), .SI(n5160), .SE(
        n1037), .CP(ClockB), .CDN(n4446), .Q(n5160) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[27]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]), .SI(n5161), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(n5161) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[26]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]), .SI(n5162), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(n5162) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[25]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]), .SI(n5163), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(n5163) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[24]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]), .SI(n5164), .SE(
        n1037), .CP(ClockB), .CDN(n4411), .Q(n5164) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[23]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]), .SI(n5165), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(n5165) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[22]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]), .SI(n5166), .SE(
        n1037), .CP(ClockB), .CDN(n4464), .Q(n5166) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[21]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]), .SI(n5167), .SE(
        n1037), .CP(ClockB), .CDN(n4422), .Q(n5167) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[20]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]), .SI(n5168), .SE(
        n1037), .CP(ClockB), .CDN(n4453), .Q(n5168) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[19]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]), .SI(n5169), .SE(
        n1037), .CP(ClockB), .CDN(n4423), .Q(n5169) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[18]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]), .SI(n5170), .SE(
        n1037), .CP(ClockB), .CDN(n4383), .Q(n5170) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[17]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]), .SI(n5171), .SE(
        n1037), .CP(ClockB), .CDN(n4453), .Q(n5171) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[16]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]), .SI(n5172), .SE(
        n1037), .CP(ClockB), .CDN(n4401), .Q(n5172) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[15]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]), .SI(n5173), .SE(
        n1037), .CP(ClockB), .CDN(n4420), .Q(n5173) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[14]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]), .SI(n5174), .SE(
        n1037), .CP(ClockB), .CDN(n4379), .Q(n5174) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[13]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]), .SI(n5175), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(n5175) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[12]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]), .SI(n5176), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(n5176) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[11]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]), .SI(n5177), .SE(
        n1037), .CP(ClockB), .CDN(n4437), .Q(n5177) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[10]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]), .SI(n5178), .SE(
        n1037), .CP(ClockB), .CDN(n4456), .Q(n5178) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[9]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]), .SI(n5179), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(n5179) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[8]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]), .SI(n5180), .SE(
        n1037), .CP(ClockB), .CDN(n4382), .Q(n5180) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[7]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]), .SI(n5181), .SE(
        n1037), .CP(ClockB), .CDN(n4447), .Q(n5181) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[6]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]), .SI(n5182), .SE(
        n1037), .CP(ClockB), .CDN(n4392), .Q(n5182) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[5]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]), .SI(n5183), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(n5183) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[4]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]), .SI(n5184), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(n5184) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]), .SI(n5185), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(n5185) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]), .SI(n5186), .SE(
        n1037), .CP(ClockB), .CDN(n4454), .Q(n5186) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]), .SI(n5187), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(n5187) );
  SDFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]), .SI(n5188), .SE(
        n1037), .CP(ClockB), .CDN(n4455), .Q(n5188) );
  SDFND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/FullFIFOr_reg  ( .D(n3528), .SI(
        \SerDes_U2/Tx_F_Full ), .SE(n1037), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(
        \SerDes_U2/Tx_F_Full ) );
  SDFND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/EmptyFIFOr_reg  ( .D(n2945), .SI(
        \SerDes_U2/Tx_F_Empty ), .SE(n1037), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(
        \SerDes_U2/Tx_F_Empty ), .QN(n1036) );
  SDFND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/EmptyFIFOr_reg  ( .D(n2909), .SI(
        \SerDes_U1/Tx_F_Empty ), .SE(n1037), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(
        \SerDes_U1/Tx_F_Empty ), .QN(n1035) );
  SDFND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/FullFIFOr_reg  ( .D(n2906), .SI(
        \SerDes_U1/Tx_F_Full ), .SE(n1037), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(
        \SerDes_U1/Tx_F_Full ), .QN(n1017) );
  SDFCND0 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ), .SE(
        n1037), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(
        n2553), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ), .QN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ) );
  SDFCND0 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ), .SE(
        n1037), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(
        n2553), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ), .QN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ) );
  SDFCND0 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ), .SE(
        n1037), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(
        n2511), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ), .QN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ) );
  SDFCND0 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ), .SE(
        n1037), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(
        n2511), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ), .QN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ) );
  SDFCND0 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ), .SE(
        n1037), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(
        n2549), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[0] ), .QN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ) );
  SDFCND0 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ), .SE(
        n1037), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(
        n2549), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN[1] ), .QN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ) );
  SDFCND0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ), .SE(
        n1037), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(
        n1625), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[1] ), .QN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ) );
  SDFCND0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ), .SE(
        n1037), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(
        n1625), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN[0] ), .QN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ) );
  SDFCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4382), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .QN(n722) );
  SDFCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4391), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .QN(n870) );
  SDFCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .QN(n1031) );
  SDFCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .QN(n1033) );
  SDFCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .QN(n1032) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteCmdr_reg  ( .D(n3482), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .SE(n1037), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4415), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .QN(n1023) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[3]  ( .D(n3473), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[3] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4416), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[3] ), .QN(n1022) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n3471), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4416), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ), .QN(n1020) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n3469), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4416), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ), .QN(n1019) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n3467), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4416), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ), .QN(n1021) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[3]  ( .D(n2953), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[3] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4440), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[3] ), .QN(n1028) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n2951), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4440), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ), .QN(n1026) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n2949), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4440), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ), .QN(n1025) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n2947), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ), .QN(n1027) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteCmdr_reg  ( .D(n2207), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .QN(n863) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[3]  ( .D(n2198), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[3] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4420), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[3] ), .QN(n862) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n2196), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4420), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ), .QN(n860) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n2194), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4417), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ), .QN(n859) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n2192), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4416), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ), .QN(n861) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[3]  ( .D(n1678), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[3] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[3] ), .QN(n868) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1676), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ), .QN(n866) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1674), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ), .QN(n865) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1672), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ), .QN(n867) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteCmdr_reg  ( .D(n2893), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .SE(n1037), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .QN(n1010) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n2888), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[2] ), .QN(n1007) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n2886), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[0] ), .QN(n1008) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n2884), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr[1] ), .QN(n1009) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n2880), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[2] ), .QN(n1012) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n2878), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[0] ), .QN(n1013) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n2876), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr[1] ), .QN(n1014) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteCmdr_reg  ( .D(n1319), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .QN(n715) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n1314), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[2] ), .QN(n712) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n1312), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[0] ), .QN(n713) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n1310), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr[1] ), .QN(n714) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1052), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4412), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[2] ), .QN(n718) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1050), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4413), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[0] ), .QN(n719) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1048), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4411), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr[1] ), .QN(n720) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[63]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[63] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[63] ), .QN(n1004)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[31]  ( .D(n2439), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [31]), .SE(n1037), .CPN(n4477), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [31]), .QN(n1005)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[30]  ( .D(n2437), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [30]), .SE(n1037), .CPN(n4474), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [30]), .QN(n971)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[29]  ( .D(n2435), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [29]), .SE(n1037), .CPN(n4477), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [29]), .QN(n969)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[28]  ( .D(n2433), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [28]), .SE(n1037), .CPN(n4475), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [28]), .QN(n967)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[27]  ( .D(n2431), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [27]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4419), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [27]), .QN(n965) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[26]  ( .D(n2429), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [26]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4419), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [26]), .QN(n963) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[25]  ( .D(n2427), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [25]), .SE(n1037), .CPN(n4474), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [25]), .QN(n961)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[24]  ( .D(n2425), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [24]), .SE(n1037), .CPN(n4476), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [24]), .QN(n959)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[23]  ( .D(n2423), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [23]), .SE(n1037), .CPN(n4476), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [23]), .QN(n957)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[22]  ( .D(n2421), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [22]), .SE(n1037), .CPN(n4475), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [22]), .QN(n955)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[21]  ( .D(n2419), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [21]), .SE(n1037), .CPN(n4476), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [21]), .QN(n953)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[20]  ( .D(n2417), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [20]), .SE(n1037), .CPN(n4477), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [20]), .QN(n951)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[19]  ( .D(n2415), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [19]), .SE(n1037), .CPN(n4475), 
        .CDN(n4419), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [19]), .QN(n949)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[18]  ( .D(n2413), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [18]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [18]), .QN(n947) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[17]  ( .D(n2411), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [17]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [17]), .QN(n945) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[16]  ( .D(n2409), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [16]), .SE(n1037), .CPN(n4475), 
        .CDN(n4418), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [16]), .QN(n943)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[15]  ( .D(n2407), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [15]), .SE(n1037), .CPN(n4474), 
        .CDN(n4418), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [15]), .QN(n941)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[14]  ( .D(n2405), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [14]), .SE(n1037), .CPN(n4475), 
        .CDN(n4418), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [14]), .QN(n939)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[13]  ( .D(n2403), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [13]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [13]), .QN(n937) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[12]  ( .D(n2401), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [12]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [12]), .QN(n935) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[11]  ( .D(n2399), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [11]), .SE(n1037), .CPN(n4474), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [11]), .QN(n933)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[10]  ( .D(n2397), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [10]), .SE(n1037), .CPN(n4475), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [10]), .QN(n931)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[9]  ( .D(n2395), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [9]), .SE(n1037), .CPN(n4477), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [9]), .QN(n929)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[8]  ( .D(n2393), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [8]), .SE(n1037), .CPN(n4476), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [8]), .QN(n927)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[7]  ( .D(n2391), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [7]), .SE(n1037), .CPN(n4474), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [7]), .QN(n925)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[6]  ( .D(n2389), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [6]), .SE(n1037), .CPN(n4477), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [6]), .QN(n923)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[5]  ( .D(n2387), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [5]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4417), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [5]), .QN(n921) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[4]  ( .D(n2385), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [4]), .SE(n1037), .CPN(n4476), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [4]), .QN(n919)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[3]  ( .D(n2383), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [3]), .SE(n1037), .CPN(n4477), 
        .CDN(n4425), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [3]), .QN(n917)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[2]  ( .D(n2381), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [2]), .SE(n1037), .CPN(n4476), 
        .CDN(n4412), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [2]), .QN(n915)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[1]  ( .D(n2379), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [1]), .SE(n1037), .CPN(n4476), 
        .CDN(n4411), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [1]), .QN(n913)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[0]  ( .D(n2377), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Decoder [0]), .SE(n1037), .CPN(n4474), 
        .CDN(n4411), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Decoder [0]), .QN(n911)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/doParSync_reg  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N47 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .SE(n1037), .CPN(n4477), 
        .CDN(n4412), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/doParSync ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad_reg  ( .D(n4478), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .QN(n909) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[0]  ( .D(n2309), 
        .SI(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[0] ), .SE(n1037), .CPN(
        n4474), .CDN(n4415), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[0] ), .QN(n876) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[1]  ( .D(n2307), 
        .SI(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[1] ), .SE(n1037), .CPN(
        n4474), .CDN(n4415), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[1] ), .QN(n874) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[2]  ( .D(n2305), 
        .SI(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[2] ), .SE(n1037), .CPN(
        n4474), .CDN(n4416), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[2] ), .QN(n873) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[3]  ( .D(n2303), 
        .SI(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[3] ), .SE(n1037), .CPN(
        n4474), .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer[3] ), .QN(n875) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidr_reg  ( .D(n2285), .SI(
        \SerDes_U1/Des_U1/ParValidDecode ), .SE(n1037), .CPN(n4475), .CDN(
        n4418), .Q(\SerDes_U1/Des_U1/ParValidDecode ), .QN(n872) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[63]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[63] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[63] ), .QN(n856) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[31]  ( .D(n1553), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [31]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [31]), .QN(n857) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[30]  ( .D(n1551), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [30]), .SE(n1037), .CPN(n4470), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [30]), .QN(n823)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[29]  ( .D(n1549), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [29]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [29]), .QN(n821) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[28]  ( .D(n1547), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [28]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [28]), .QN(n819) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[27]  ( .D(n1545), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [27]), .SE(n1037), .CPN(n4467), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [27]), .QN(n817)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[26]  ( .D(n1543), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [26]), .SE(n1037), .CPN(n4467), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [26]), .QN(n815)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[25]  ( .D(n1541), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [25]), .SE(n1037), .CPN(n4470), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [25]), .QN(n813)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[24]  ( .D(n1539), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [24]), .SE(n1037), .CPN(n4468), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [24]), .QN(n811)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[23]  ( .D(n1537), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [23]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4432), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [23]), .QN(n809) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[22]  ( .D(n1535), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [22]), .SE(n1037), .CPN(n4469), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [22]), .QN(n807)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[21]  ( .D(n1533), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [21]), .SE(n1037), .CPN(n4469), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [21]), .QN(n805)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[20]  ( .D(n1531), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [20]), .SE(n1037), .CPN(n4469), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [20]), .QN(n803)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[19]  ( .D(n1529), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [19]), .SE(n1037), .CPN(n4468), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [19]), .QN(n801)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[18]  ( .D(n1527), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [18]), .SE(n1037), .CPN(n4471), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [18]), .QN(n799)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[17]  ( .D(n1525), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [17]), .SE(n1037), .CPN(n4470), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [17]), .QN(n797)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[16]  ( .D(n1523), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [16]), .SE(n1037), .CPN(n4471), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [16]), .QN(n795)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[15]  ( .D(n1521), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [15]), .SE(n1037), .CPN(n4467), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [15]), .QN(n793)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[14]  ( .D(n1519), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [14]), .SE(n1037), .CPN(n4471), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [14]), .QN(n791)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[13]  ( .D(n1517), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [13]), .SE(n1037), .CPN(n4467), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [13]), .QN(n789)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[12]  ( .D(n1515), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [12]), .SE(n1037), .CPN(n4471), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [12]), .QN(n787)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[11]  ( .D(n1513), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [11]), .SE(n1037), .CPN(n4470), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [11]), .QN(n785)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[10]  ( .D(n1511), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [10]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [10]), .QN(n783) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[9]  ( .D(n1509), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [9]), .SE(n1037), .CPN(n4468), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [9]), .QN(n781)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[8]  ( .D(n1507), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [8]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [8]), .QN(n779) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[7]  ( .D(n1505), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [7]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [7]), .QN(n777) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[6]  ( .D(n1503), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [6]), .SE(n1037), .CPN(n4471), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [6]), .QN(n775)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[5]  ( .D(n1501), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [5]), .SE(n1037), .CPN(n4471), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [5]), .QN(n773)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[4]  ( .D(n1499), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [4]), .SE(n1037), .CPN(n4468), 
        .CDN(n4433), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [4]), .QN(n771)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[3]  ( .D(n1497), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [3]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [3]), .QN(n769) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[2]  ( .D(n1495), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [2]), .SE(n1037), .CPN(n4470), 
        .CDN(n4434), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [2]), .QN(n767)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[1]  ( .D(n1493), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [1]), .SE(n1037), .CPN(n4470), 
        .CDN(n4434), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [1]), .QN(n765)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[0]  ( .D(n1491), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Decoder [0]), .SE(n1037), .CPN(n4467), 
        .CDN(n4434), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Decoder [0]), .QN(n763)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/doParSync_reg  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N47 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .SE(n1037), .CPN(n4471), 
        .CDN(n4434), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/doParSync ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad_reg  ( .D(n4472), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .SE(n1037), .CPN(n4468), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .QN(n761) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[0]  ( .D(n1423), 
        .SI(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[0] ), .SE(n1037), .CPN(
        n4469), .CDN(n4437), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[0] ), .QN(n728) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[1]  ( .D(n1421), 
        .SI(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[1] ), .SE(n1037), .CPN(
        n4469), .CDN(n4437), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[1] ), .QN(n726) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[2]  ( .D(n1419), 
        .SI(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[2] ), .SE(n1037), .CPN(
        n4469), .CDN(n4437), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[2] ), .QN(n725) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[3]  ( .D(n1417), 
        .SI(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[3] ), .SE(n1037), .CPN(
        n4469), .CDN(n4437), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer[3] ), .QN(n727) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidr_reg  ( .D(n1399), .SI(
        \SerDes_U2/Des_U1/ParValidDecode ), .SE(n1037), .CPN(n4470), .CDN(
        n4437), .Q(\SerDes_U2/Des_U1/ParValidDecode ), .QN(n724) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4420), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4432), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4428), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4415), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), .E(n4487), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4434), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4428), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4415), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), .E(n4483), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[30]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N83 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4460), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[29]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4452), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[26]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N79 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4451), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[25]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ), .SE(n1037), .CP(n4520), 
        .CDN(n4435), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[22]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N75 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ), .SE(n1037), .CP(n4520), 
        .CDN(n4400), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[21]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[18]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N71 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4399), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[17]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4397), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[14]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N67 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ), .SE(n1037), .CP(n4520), 
        .CDN(n4434), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[13]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4404), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[10]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N63 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ), .SE(n1037), .CP(n4520), 
        .CDN(n4446), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[9]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ), .SE(n1037), .CP(n4520), .CDN(
        n4392), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[6]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N59 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ), .SE(n1037), .CP(n4520), .CDN(
        n4400), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ), .SE(n1037), .CP(n4520), .CDN(
        n4438), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N55 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ), .SE(n1037), .CP(n4520), .CDN(
        n4435), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ), .SE(n1037), .CP(n4520), .CDN(
        n4433), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N54 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4462), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N58 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ), .SE(n1037), .CP(n4522), .CDN(
        n4437), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[6]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ), .SE(n1037), .CP(n4522), .CDN(
        n4376), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[9]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N62 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ), .SE(n1037), .CP(n4522), .CDN(
        n4453), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[10]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ), .SE(n1037), .CP(n4522), 
        .CDN(n4375), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[13]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N66 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ), .SE(n1037), .CP(n4522), 
        .CDN(n4431), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[14]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ), .SE(n1037), .CP(n4522), 
        .CDN(n4435), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[17]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N70 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4424), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[18]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4451), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[21]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N74 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ), .SE(n1037), .CP(n4522), 
        .CDN(n4374), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[22]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ), .SE(n1037), .CP(n4522), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[25]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N78 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[26]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ), .SE(n1037), .CP(n4522), 
        .CDN(n4395), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[29]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N82 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4406), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[30]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ), .SE(n1037), .CP(n4522), 
        .CDN(n4402), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[31]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[28]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N81 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4444), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[27]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4443), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[24]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N77 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ), .SE(n1037), .CP(n4520), 
        .CDN(n4403), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[23]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4401), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[20]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N73 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ), .SE(n1037), .CP(n4520), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[19]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ), .SE(n1037), .CP(n4520), 
        .CDN(n4407), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[16]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N69 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[15]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ), .SE(n1037), .CP(n4520), 
        .CDN(n4405), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[12]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N65 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4434), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[11]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ), .SE(n1037), .CP(n4520), 
        .CDN(n4383), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[8]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N61 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ), .SE(n1037), .CP(n4520), .CDN(
        n4449), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[7]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ), .SE(n1037), .CP(n4520), .CDN(
        n4393), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N57 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ), .SE(n1037), .CP(n4520), .CDN(
        n4436), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ), .SE(n1037), .CP(n4520), .CDN(
        n4418), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N53 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4419), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4462), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N56 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4387), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4379), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[7]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N60 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ), .SE(n1037), .CP(n4522), .CDN(
        n4378), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[8]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ), .SE(n1037), .CP(n4522), .CDN(
        n4377), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[11]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N64 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ), .SE(n1037), .CP(n4522), 
        .CDN(n4376), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[12]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ), .SE(n1037), .CP(n4522), 
        .CDN(n4400), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[15]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N68 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ), .SE(n1037), .CP(n4522), 
        .CDN(n4449), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[16]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[19]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N72 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ), .SE(n1037), .CP(n4522), 
        .CDN(n4420), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[20]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4458), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[23]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N76 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[24]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ), .SE(n1037), .CP(n4522), 
        .CDN(n4397), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[27]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N80 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4408), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[28]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ), .SE(n1037), .CP(n4522), 
        .CDN(n4407), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[31]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N84 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4392), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4435), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4436), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .E(n4495), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4393), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4411), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4392), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4418), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4384), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .E(n4493), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4408), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4425), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), .E(n4491), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4382), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .E(n4489), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4420), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4430), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .E(n4485), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4430), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4428), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4433), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4436), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .E(n4497), .SE(
        n1037), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ) );
  SDFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SDN(n4410), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]) );
  SDFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SDN(n4409), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]) );
  SDFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SDN(n4410), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]) );
  SDFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SDN(n4410), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4391), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4425), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ), .E(n4592), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ), .E(n4592), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4420), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4375), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4432), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4432), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ), .E(n4590), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4375), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ), .E(n4590), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4388), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4435), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4375), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ), .E(n4584), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4415), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ), .E(n4584), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4437), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4427), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4434), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4411), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4425), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ), .E(n4582), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4432), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4408), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .E(n4576), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4408), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4401), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4388), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4401), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4382), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4420), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .E(n4574), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4391), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4392), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4377), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4375), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4420), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4430), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4400), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), .E(n4568), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4437), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4433), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4393), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4434), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4411), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4400), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .E(n4566), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4382), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4410), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4431), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ), .E(n4594), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ), .E(n4594), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4430), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4437), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4375), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4415), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ), .E(n4588), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4408), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4389), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ), .E(n4588), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4383), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4392), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4448), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4379), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ), .E(n4586), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4437), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4432), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4392), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ), .E(n4586), 
        .SE(n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4428), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4436), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4419), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4453), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4438), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4400), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ), .E(n4580), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4454), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4455), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4415), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4465), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4417), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4376), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4404), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .E(n4578), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4436), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4381), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4417), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4426), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4451), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4449), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4443), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4446), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), .E(n4572), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4464), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4396), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4427), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4444), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4378), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4409), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4437), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4406), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4407), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4408), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4399), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4429), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4393), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4388), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4385), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4401), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .E(n4570), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4403), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4386), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4436), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4439), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4434), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n3530), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4425), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4466), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4458), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4460), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4456), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4397), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4398), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4440), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4463), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4442), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), .E(n4564), .SE(
        n1037), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4434), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n4394), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4413), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4403), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]), .E(n4519), .SE(n1037), .CP(ClockA), .CDN(n4431), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4388), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4446), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4422), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4430), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4396), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4439), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4436), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4419), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4408), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4418), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4449), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4374), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4427), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4433), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4428), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4465), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4460), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4422), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4463), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4423), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4425), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4426), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4459), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4414), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4411), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4435), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]), .E(n4519), .SE(
        n1037), .CP(ClockA), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4404), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4404), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4404), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4404), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4404), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), .E(n4502), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4395), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), .E(n4506), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4436), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4384), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4439), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4382), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4442), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4378), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4386), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4448), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4391), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4412), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4441), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4455), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4440), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4441), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4408), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4375), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4380), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4458), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4402), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4419), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4429), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4463), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4425), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4415), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4419), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4427), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4428), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .E(n4514), .SE(
        n1037), .CP(ClockA), .CDN(n4432), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4465), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4417), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4419), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4426), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4423), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4422), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4425), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4418), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4414), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4416), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4415), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4444), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4448), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4442), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4391), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4462), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4441), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4457), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4445), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4406), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4418), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4440), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4375), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4389), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4391), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4410), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4442), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4456), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4438), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4437), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), .E(n4510), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4463), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4457), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4460), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4386), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4378), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4464), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4447), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4389), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4428), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4377), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4411), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4434), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4409), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4417), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4420), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4435), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4463), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4466), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4456), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4439), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4436), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4421), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4424), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4431), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4430), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4429), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4392), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4415), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4446), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4427), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .E(n4512), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4375), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4442), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4401), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4401), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4399), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .E(n4504), .SE(
        n1037), .CP(ClockA), .CDN(n4398), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4394), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4394), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4395), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4396), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4409), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4409), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4410), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4464), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4426), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4428), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4423), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4430), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4431), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4415), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4413), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4383), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4412), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4432), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .E(n4508), .SE(
        n1037), .CP(ClockA), .CDN(n4388), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4392), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4464), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        InParDataA[0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4400), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        InParDataA[1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4393), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        InParDataA[2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4459), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        InParDataA[3]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4386), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        InParDataA[4]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4374), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        InParDataA[5]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4410), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        InParDataA[6]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4390), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        InParDataA[7]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4391), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        InParDataA[8]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4440), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        InParDataA[9]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4447), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        InParDataA[10]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4413), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        InParDataA[11]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4410), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        InParDataA[12]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4414), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        InParDataA[13]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4434), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        InParDataA[14]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4378), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        InParDataA[15]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4397), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        InParDataA[16]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4455), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        InParDataA[17]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4437), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        InParDataA[18]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4417), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        InParDataA[19]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4424), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        InParDataA[20]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4386), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        InParDataA[21]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4416), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        InParDataA[22]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4382), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        InParDataA[23]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4451), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        InParDataA[24]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4385), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        InParDataA[25]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4409), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        InParDataA[26]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4392), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        InParDataA[27]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4408), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        InParDataA[28]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4407), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        InParDataA[29]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .E(n4516), .SE(
        n1037), .CP(ClockA), .CDN(n4420), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ) );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        InParDataA[30]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4415), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] )
         );
  SEDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        InParDataA[31]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .SE(n1037), .CP(ClockA), 
        .CDN(n4461), .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] )
         );
  SEDFCNQHD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[4]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N42 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ), .E(\SerDes_U1/SerLineValid ), .SE(n1037), .CP(n4475), .CDN(n4391), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[4]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N42 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ), .E(\SerDes_U2/SerLineValid ), .SE(n1037), .CP(n4470), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), .SE(n1037), 
        .CP(\SerDes_U2/Rx_ParClk ), .CDN(n1625), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]), .E(n3582), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]), .E(n4596), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4383), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4383), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4383), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]), .E(n4596), .SE(n1037), .CP(ClockB), .CDN(n4383), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4403), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4401), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4376), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n4393), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n4402), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n4414), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4446), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4374), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n4402), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), .SE(n1037), 
        .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2511), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4396), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4466), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4464), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4411), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4401), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4445), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4400), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4427), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4443), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4374), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ), .E(n4556), .SE(
        n1037), .CP(ClockB), .CDN(n4448), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4410), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ), .E(n4556), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4379), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4379), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4379), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4379), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4378), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4378), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ), .E(n4554), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4377), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n3530), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4418), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4400), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ), .E(n4554), 
        .SE(n1037), .CP(ClockB), .CDN(n4451), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4462), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4411), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4392), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4391), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4391), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ), .E(n4548), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4390), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ), .E(n4548), 
        .SE(n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4389), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4389), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4386), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4445), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4418), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4438), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4465), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ), .E(n4546), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4383), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4412), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4443), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4444), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4452), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4451), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4450), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4449), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4401), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4465), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4417), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4448), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4447), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4441), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4454), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4453), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4455), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4394), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4375), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4426), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4448), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4425), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4410), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4456), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4396), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .E(n4540), .SE(
        n1037), .CP(ClockB), .CDN(n4386), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4429), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4399), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4397), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4407), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4402), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4403), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4388), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4387), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4457), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4418), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4436), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4446), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .E(n4538), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4376), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4376), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4417), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4424), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4395), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4430), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4459), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4440), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4454), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4400), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4404), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4448), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4397), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4454), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4453), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4455), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4418), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4396), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4394), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4413), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), .E(n4532), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4402), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4403), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4401), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4387), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4378), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4439), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4456), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4399), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4436), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4431), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4420), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4446), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4434), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4422), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4402), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .E(n4530), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4382), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4382), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4382), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4381), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n3530), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ), .E(n4558), .SE(
        n1037), .CP(ClockB), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n3530), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4411), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4401), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4400), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4427), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ), .E(n4558), 
        .SE(n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4460), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4401), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4409), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4437), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4461), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4433), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4417), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4421), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4439), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4436), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4449), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4403), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4389), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4457), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4453), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4454), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ), .E(n4552), .SE(
        n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4388), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4385), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4403), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4437), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ), .E(n4552), 
        .SE(n1037), .CP(ClockB), .CDN(n4412), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4382), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4430), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4415), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4413), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4449), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4424), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4429), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4411), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4464), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4400), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4405), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4423), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4414), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4416), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4425), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4466), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4461), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4459), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4463), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ), .E(n4550), .SE(
        n1037), .CP(ClockB), .CDN(n4402), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4460), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4458), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4410), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ), .E(n4550), 
        .SE(n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4392), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4392), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4416), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4415), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4413), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4424), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4463), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4437), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4434), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4436), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4417), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4420), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4393), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4419), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4464), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4423), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4422), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4425), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4426), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4427), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4429), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4458), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4448), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4397), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4455), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ), .E(n4544), .SE(
        n1037), .CP(ClockB), .CDN(n4465), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4380), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4420), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n3530), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4411), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4413), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4374), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4434), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4387), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4457), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4407), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4417), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4444), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4430), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4464), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4430), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4461), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4455), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4394), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4438), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4421), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4427), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .E(n4542), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4440), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4396), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4375), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4375), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4375), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4444), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4456), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4391), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4442), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4396), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4440), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4410), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4441), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4424), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4385), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4447), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4394), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4397), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4399), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4398), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4384), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4425), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), .E(n4536), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4376), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4449), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4379), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4412), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4439), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4375), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4454), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4413), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4436), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4421), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4419), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4377), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4376), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4375), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4380), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4445), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4430), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4466), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4450), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4465), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4435), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4450), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4374), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4458), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4409), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4431), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4445), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4429), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4438), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .E(n4534), .SE(
        n1037), .CP(ClockB), .CDN(n4466), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4440), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4394), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        InParDataB[31]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        InParDataB[29]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        InParDataB[27]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        InParDataB[25]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4408), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        InParDataB[23]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        InParDataB[21]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        InParDataB[19]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        InParDataB[17]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4408), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        InParDataB[15]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        InParDataB[13]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        InParDataB[11]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4407), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        InParDataB[9]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        InParDataB[7]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        InParDataB[5]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        InParDataB[3]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        InParDataB[1]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        InParDataB[0]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        InParDataB[2]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4407), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        InParDataB[4]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        InParDataB[6]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        InParDataB[8]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        InParDataB[10]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        InParDataB[12]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        InParDataB[14]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        InParDataB[16]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        InParDataB[18]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        InParDataB[20]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        InParDataB[22]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4406), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        InParDataB[24]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4390), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        InParDataB[26]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), .E(n4528), .SE(
        n1037), .CP(ClockB), .CDN(n4405), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ) );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        InParDataB[28]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4405), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] )
         );
  SEDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        InParDataB[30]), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .SE(n1037), .CP(ClockB), 
        .CDN(n4405), .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] )
         );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4441), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n4380), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4451), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n4400), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), .SE(n1037), 
        .CP(ClockA), .CDN(n2553), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4382), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4417), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4461), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4452), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ) );
  SDFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[1]  ( 
        .D(n1650), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .SE(n1037), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ) );
  SDFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[1]  ( 
        .D(n2536), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .SE(n1037), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ) );
  SDFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[1]  ( 
        .D(n1403), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .SE(n1037), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ) );
  SDFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[1]  ( 
        .D(n2289), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .SE(n1037), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4411), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ) );
  SDFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[4]  ( 
        .D(n1655), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .SE(n1037), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ) );
  SDFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[4]  ( 
        .D(n2541), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .SE(n1037), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4409), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ) );
  SDFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[4]  ( 
        .D(n1623), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .SE(n1037), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ) );
  SDFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[4]  ( 
        .D(n2509), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .SE(n1037), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4409), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .SE(n1037), 
        .CP(\SerDes_U2/Rx_ParClk ), .CDN(n1625), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), .SE(n1037), 
        .CP(ClockB), .CDN(n2549), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[1]  ( .D(n3526), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4411), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .QN(n1030) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[0]  ( .D(n3485), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4415), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .QN(n1024) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[2]  ( .D(n3479), 
        .SI(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .SE(n1037), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4415), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .QN(n1018) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[1]  ( .D(n2283), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4418), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .QN(n871) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[0]  ( .D(n2213), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4425), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .QN(n864) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[2]  ( .D(n2204), 
        .SI(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .SE(n1037), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4423), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .QN(n858) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[1]  ( .D(n2904), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .QN(n1016) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[0]  ( .D(n2896), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .QN(n1011) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[2]  ( .D(n2882), 
        .SI(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .SE(n1037), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .QN(n1006) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[1]  ( .D(n1397), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4437), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .QN(n723) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[0]  ( .D(n1327), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .QN(n717) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[8]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4416), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ), .QN(n910)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[9]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ), .QN(n912)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[10]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ), .QN(n914)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[11]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ), .QN(n916)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[12]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ), .QN(n918)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[13]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ), .QN(n920)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[14]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ), .QN(n922) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[15]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4425), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ), .QN(n924)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[18]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4425), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ), .QN(n997)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[19]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4425), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ), .QN(n1003) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[23]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ), .QN(n4615)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[24]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ), .QN(n926)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[25]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ), .QN(n928) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[26]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ), .QN(n930)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[27]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ), .QN(n932)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[28]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ), .QN(n934)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[29]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ), .QN(n936)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[30]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ), .QN(n938)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[31]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ), .QN(n940)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[32]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ), .QN(n4614)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[34]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ), .QN(n989)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[35]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ), .QN(n990)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[37]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ), .QN(n4613)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[40]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ), .QN(n942)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[41]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ), .QN(n944)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[42]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ), .QN(n946)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[43]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ), .QN(n948)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[44]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ), .QN(n950) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[45]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ), .QN(n952)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[46]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4422), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ), .QN(n954) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[47]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ), .QN(n956)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[48]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ), .QN(n985)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[54]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ), .QN(n4612)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[55]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ), .QN(n4611)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[56]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ), .QN(n958)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[57]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ), .QN(n960)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[58]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4420), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ), .QN(n962) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[59]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ), .QN(n964)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[60]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ), .QN(n966)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[61]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ), .QN(n968)
         );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[62]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4420), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ), .QN(n970)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[8]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ), .QN(n762)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[9]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ), .QN(n764)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[10]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ), .QN(n766)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[11]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ), .QN(n768)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[12]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ), .QN(n770)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[13]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ), .QN(n772)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[14]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ), .QN(n774)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[15]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ), .QN(n776)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[18]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ), .QN(n849)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[19]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ), .QN(n855)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[23]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ), .QN(n4610)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[24]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ), .QN(n778) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[25]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ), .QN(n780) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[26]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ), .QN(n782)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[27]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ), .QN(n784)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[28]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ), .QN(n786)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[29]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ), .QN(n788)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[30]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ), .QN(n790)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[31]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ), .QN(n792)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[32]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ), .QN(n4609)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[34]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ), .QN(n841)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[35]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4428), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ), .QN(n842) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[37]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ), .QN(n4608)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[40]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ), .QN(n794)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[41]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4429), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ), .QN(n796) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[42]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ), .QN(n798)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[43]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ), .QN(n800)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[44]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ), .QN(n802)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[45]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ), .QN(n804)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[46]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4429), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ), .QN(n806) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[47]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ), .QN(n808)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[48]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ), .QN(n837)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[54]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ), .QN(n4607)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[55]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ), .QN(n4606)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[56]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4430), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ), .QN(n810) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[57]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ), .QN(n812)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[58]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ), .QN(n814)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[59]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4430), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ), .QN(n816) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[60]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ), .QN(n818)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[61]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ), .QN(n820)
         );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[62]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4431), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ), .QN(n822)
         );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .SE(n1037), 
        .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2511), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[1]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N39 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ), .E(\SerDes_U1/SerLineValid ), .SE(n1037), .CP(n4475), .CDN(n4387), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[1]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N39 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ), .E(\SerDes_U2/SerLineValid ), .SE(n1037), .CP(n4470), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ) );
  SDFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[0]  ( 
        .D(n1652), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .SE(n1037), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ) );
  SDFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[0]  ( 
        .D(n2538), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .SE(n1037), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ) );
  SDFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[0]  ( 
        .D(n1401), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .SE(n1037), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4410), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ) );
  SDFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[0]  ( 
        .D(n2287), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .SE(n1037), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(n4411), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4443), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4437), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4443), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4450), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[2]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N40 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ), .E(\SerDes_U1/SerLineValid ), .SE(n1037), .CP(n4475), .CDN(n4389), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[3]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N41 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ), .E(\SerDes_U1/SerLineValid ), .SE(n1037), .CP(n4475), .CDN(n4390), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[2]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N40 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ), .E(\SerDes_U2/SerLineValid ), .SE(n1037), .CP(n4470), .CDN(n4450), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[3]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N41 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ), .E(\SerDes_U2/SerLineValid ), .SE(n1037), .CP(n4470), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .SE(n1037), 
        .CP(ClockA), .CDN(n2553), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[0]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N38 ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ), .E(\SerDes_U1/SerLineValid ), .SE(n1037), .CP(n4474), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[0]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N38 ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ), .E(\SerDes_U2/SerLineValid ), .SE(n1037), .CP(n4469), .CDN(n4405), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4446), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4435), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4454), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4392), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4393), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4465), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .SE(n1037), 
        .CP(ClockB), .CDN(n2549), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n4438), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n4432), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n4386), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4421), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4424), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4382), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4410), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4425), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4433), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4416), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4385), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4449), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4444), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4417), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), .SE(n1037), 
        .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4406), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), .SE(n1037), 
        .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4414), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), .SE(n1037), 
        .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4417), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), .SE(n1037), 
        .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4443), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[0]  ( .D(n1487), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .SE(n1037), .CPN(n4467), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [0]), .QN(n760) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[1]  ( .D(n1485), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .SE(n1037), .CPN(n4469), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [1]), .QN(n759) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[2]  ( .D(n1483), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .SE(n1037), .CPN(n4469), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [2]), .QN(n758) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[3]  ( .D(n1481), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4434), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .QN(n757) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[4]  ( .D(n1479), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .SE(n1037), .CPN(n4471), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [4]), .QN(n756) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[5]  ( .D(n1477), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .SE(n1037), .CPN(n4470), .CDN(
        n4434), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [5]), .QN(n755) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[6]  ( .D(n1475), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4435), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .QN(n754) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[7]  ( .D(n1473), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .SE(n1037), .CPN(n4469), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [7]), .QN(n753) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[8]  ( .D(n1471), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .SE(n1037), .CPN(n4468), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [8]), .QN(n752) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[9]  ( .D(n1469), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .SE(n1037), .CPN(n4471), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [9]), .QN(n751) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[10]  ( .D(n1467), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [10]), .QN(n750) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[11]  ( .D(n1465), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [11]), .QN(n749) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[12]  ( .D(n1463), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [12]), .QN(n748) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[13]  ( .D(n1461), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [13]), .QN(n747) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[14]  ( .D(n1459), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [14]), .QN(n746) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[15]  ( .D(n1457), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [15]), .QN(n745) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[16]  ( .D(n1455), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .SE(n1037), .CPN(n4467), .CDN(
        n4435), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [16]), .QN(n744) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[17]  ( .D(n1453), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .SE(n1037), .CPN(n4467), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [17]), .QN(n743) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[18]  ( .D(n1451), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .SE(n1037), .CPN(n4467), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [18]), .QN(n742) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[19]  ( .D(n1449), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [19]), .QN(n741) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[20]  ( .D(n1447), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [20]), .QN(n740) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[21]  ( .D(n1445), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [21]), .QN(n739) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[22]  ( .D(n1443), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [22]), .QN(n738) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[23]  ( .D(n1441), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [23]), .QN(n737) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[24]  ( .D(n1439), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [24]), .QN(n736) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[25]  ( .D(n1437), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [25]), .QN(n735) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[26]  ( .D(n1435), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [26]), .QN(n734) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[27]  ( .D(n1433), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .SE(n1037), .CPN(n4468), .CDN(
        n4436), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [27]), .QN(n733) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[28]  ( .D(n1431), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .SE(n1037), .CPN(n4469), .CDN(
        n4437), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [28]), .QN(n732) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[29]  ( .D(n1429), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .SE(n1037), .CPN(n4469), .CDN(
        n4437), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [29]), .QN(n731) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[30]  ( .D(n1427), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .SE(n1037), .CPN(n4469), .CDN(
        n4437), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [30]), .QN(n730) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[31]  ( .D(n1425), .SI(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .SE(n1037), .CPN(n4469), .CDN(
        n4437), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [31]), .QN(n729) );
  SDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4423), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[36]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4423), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[52]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[36]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[52]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ) );
  SDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4434), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[2]  ( .D(n1324), 
        .SI(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .SE(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4438), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[51]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[51]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRxToDecode ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4415), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[1]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4415), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[2]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4415), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[4]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4417), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[5]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4416), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[6]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4416), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[16]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4411), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[17]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4425), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[20]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ), .SE(n1037), .CPN(n4474), 
        .CDN(n4425), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[21]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4424), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[22]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4424), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[33]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[38]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4423), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[39]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ), .SE(n1037), .CPN(n4476), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[49]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[50]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ), .SE(n1037), .CPN(n4475), 
        .CDN(n4421), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[53]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4421), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRxToDecode ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4411), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[1]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4432), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[2]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4425), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[4]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4425), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[5]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4425), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[6]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[16]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[17]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[20]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[21]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4427), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[22]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4427), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[33]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ), .SE(n1037), .CPN(n4469), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[38]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4428), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[39]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ), .SE(n1037), .CPN(n4471), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[49]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ), .SE(n1037), .CPN(n4467), 
        .CDN(n4429), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[50]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ), .SE(n1037), .CPN(n4468), 
        .CDN(n4430), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[53]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4430), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4451), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[3]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4416), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[7]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ), .SI(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ), .SE(n1037), .CPN(n4477), 
        .CDN(n4416), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[3]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4425), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ) );
  SDFNCND0 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[7]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ), .SI(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ), .SE(n1037), .CPN(n4470), 
        .CDN(n4426), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4420), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n4430), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4430), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4417), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4428), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4457), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4453), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ) );
  SDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4384), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4404), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]) );
  SDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutReg_reg  ( .D(
        n2505), .SI(\SerDes_U1/Des_U1/SerialClk ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4446), 
        .Q(\SerDes_U1/Des_U1/SerialClk ) );
  SDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutReg_reg  ( .D(
        n1619), .SI(\SerDes_U2/Des_U1/SerialClk ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n4440), 
        .Q(\SerDes_U2/Des_U1/SerialClk ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutReg_reg  ( .D(
        n2532), .SI(\SerDes_U1/Tx_SerClk ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4425), 
        .Q(\SerDes_U1/Tx_SerClk ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutReg_reg  ( .D(
        n1646), .SI(\SerDes_U2/Tx_SerClk ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n4434), 
        .Q(\SerDes_U2/Tx_SerClk ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4427), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n4454), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n4400), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]) );
  SDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[0]  ( .D(n2373), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .SE(n1037), .CPN(n4476), .CDN(
        n4412), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [0]), .QN(n908) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[1]  ( .D(n2371), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .QN(n907) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[2]  ( .D(n2369), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .SE(n1037), .CPN(n4476), .CDN(
        n4412), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [2]), .QN(n906) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[3]  ( .D(n2367), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .SE(n1037), .CPN(n4474), .CDN(
        n4412), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [3]), .QN(n905) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[4]  ( .D(n2365), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .QN(n904) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[5]  ( .D(n2363), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .QN(n903) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[6]  ( .D(n2361), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .QN(n902) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[7]  ( .D(n2359), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .SE(n1037), .CPN(n4476), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [7]), .QN(n901) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[8]  ( .D(n2357), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .SE(n1037), .CPN(n4477), .CDN(
        n4412), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [8]), .QN(n900) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[9]  ( .D(n2355), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .QN(n899) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[10]  ( .D(n2353), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .QN(n898) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[11]  ( .D(n2351), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .SE(n1037), .CPN(n4476), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [11]), .QN(n897) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[12]  ( .D(n2349), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .SE(n1037), .CPN(n4477), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [12]), .QN(n896) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[13]  ( .D(n2347), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4413), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .QN(n895) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[14]  ( .D(n2345), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .SE(n1037), .CPN(n4477), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [14]), .QN(n894) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[15]  ( .D(n2343), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .SE(n1037), .CPN(n4477), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [15]), .QN(n893) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[16]  ( .D(n2341), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .SE(n1037), .CPN(n4476), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [16]), .QN(n892) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[17]  ( .D(n2339), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .SE(n1037), .CPN(n4476), .CDN(
        n4413), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [17]), .QN(n891) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[18]  ( .D(n2337), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4415), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .QN(n890) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[19]  ( .D(n2335), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .SE(n1037), .CPN(n4475), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [19]), .QN(n889) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[20]  ( .D(n2333), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .SE(n1037), .CPN(n4477), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [20]), .QN(n888) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[21]  ( .D(n2331), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .SE(n1037), .CPN(n4477), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [21]), .QN(n887) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[22]  ( .D(n2329), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .SE(n1037), .CPN(n4475), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [22]), .QN(n886) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[23]  ( .D(n2327), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .SE(n1037), .CPN(n4474), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [23]), .QN(n885) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[24]  ( .D(n2325), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .SE(n1037), .CPN(n4477), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [24]), .QN(n884) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[25]  ( .D(n2323), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n4415), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .QN(n883) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[26]  ( .D(n2321), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .SE(n1037), .CPN(n4474), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [26]), .QN(n882) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[27]  ( .D(n2319), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .SE(n1037), .CPN(n4476), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [27]), .QN(n881) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[28]  ( .D(n2317), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .SE(n1037), .CPN(n4474), .CDN(
        n4418), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [28]), .QN(n880) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[29]  ( .D(n2315), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .SE(n1037), .CPN(n4474), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [29]), .QN(n879) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[30]  ( .D(n2313), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .SE(n1037), .CPN(n4474), .CDN(
        n4414), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [30]), .QN(n878) );
  SDFNCND0 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[31]  ( .D(n2311), .SI(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .SE(n1037), .CPN(n4474), .CDN(
        n4415), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [31]), .QN(n877) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4382), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/SerValidr_reg  ( .D(n1036), .SI(
        \SerDes_U2/SerLineValid ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4445), .Q(
        \SerDes_U2/SerLineValid ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/SerValidr_reg  ( .D(n1035), .SI(
        \SerDes_U1/SerLineValid ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n4422), .Q(
        \SerDes_U1/SerLineValid ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4385), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4426), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4410), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4390), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4429), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4413), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4431), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ), .SI(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4383), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4405), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4445), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4374), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4441), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ) );
  SEDFCNQHD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .SE(n1037), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4409), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4457), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ) );
  SEDFCNQHD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .SE(n1037), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4377), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr_reg  ( .D(n4523), .SI(
        n4522), .SE(n1037), .CP(ClockA), .CDN(n4426), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr_reg  ( .D(n4521), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .SE(n1037), .CP(ClockB), 
        .CDN(n4439), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4449), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4427), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ) );
  SDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 ), .SI(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4393), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ) );
  SDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 ), .SI(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4411), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ) );
  SDFNCND0 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadCmdr_reg  ( .D(n3523), .SI(
        n3582), .SE(n1037), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4411), .Q(
        n3582), .QN(n3587) );
  SDFNCND0 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadCmdr_reg  ( .D(n2280), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CPN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4418), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .QN(n869) );
  SDFNCND0 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadCmdr_reg  ( .D(n2901), .SI(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .SE(n1037), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n4439), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .QN(n1015) );
  SDFNCND0 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadCmdr_reg  ( .D(n1394), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CPN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n4437), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .QN(n721) );
  SEDFCNQHD2 \SerDes_U2/Des_U1/DesDec_Rx1/ParClkr_reg  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N37 ), .SI(n1037), .E(
        \SerDes_U2/Des_U1/DesDec_Rx1/N43 ), .SE(n1037), .CP(n4470), .CDN(n4465), .Q(\SerDes_U2/Rx_ParClk ) );
  SEDFCNQHD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/SerOutr_reg  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 ), .SI(
        \SerDes_U1/Des_U1/SerRxToDecode ), .E(n5124), .SE(n1037), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n4393), .Q(
        \SerDes_U1/Des_U1/SerRxToDecode ) );
  SEDFCNQHD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/SerOutr_reg  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ), .SI(
        \SerDes_U2/Des_U1/SerRxToDecode ), .E(n5124), .SE(n1037), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n4448), .Q(
        \SerDes_U2/Des_U1/SerRxToDecode ) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4398), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4453), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4463), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4458), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4463), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4412), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4444), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4380), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4446), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4462), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4451), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4455), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4453), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4454), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4426), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4456), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4442), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4447), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4408), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4445), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]), .E(n4518), .SE(
        n1037), .CP(ClockA), .CDN(n4444), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4443), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4449), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4450), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockA), 
        .CDN(n4452), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4451), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4448), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4445), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n3530), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4402), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]) );
  SEDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ), .SI(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]), .E(n4518), .SE(n1037), .CP(ClockA), .CDN(n4391), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4415), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [31]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4425), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [30]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4395), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [29]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4422), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [28]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4432), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [27]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4464), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [26]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4381), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [25]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4440), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [24]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4447), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [23]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4455), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [22]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4411), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [21]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4433), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [20]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4452), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [19]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4446), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [18]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4447), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [17]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .SE(n1037), .CP(ClockB), 
        .CDN(n4449), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [16]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4412), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [15]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4450), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [14]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4459), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [13]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4462), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [12]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4461), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [11]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]), .E(n4597), .SE(
        n1037), .CP(ClockB), .CDN(n4392), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [10]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4466), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [9]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4399), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [8]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4377), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [7]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4395), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [6]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4448), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [5]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4460), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [4]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4466), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [3]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4438), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [2]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4450), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [1]) );
  SEDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ), .SI(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]), .E(n4597), .SE(n1037), .CP(ClockB), .CDN(n4441), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr [0]) );
  SDFSND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .SI(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ), .SE(n1037), 
        .CP(\SerDes_U2/Rx_ParClk ), .SDN(n4411), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ), .QN(n1625)
         );
  SDFSND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .SI(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ), .SE(n1037), 
        .CP(\SerDes_U1/Rx_ParClk ), .SDN(n4411), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters ), .QN(n2511)
         );
  SDFSND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .SI(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ), .SE(n1037), 
        .CP(ClockA), .SDN(n4409), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ), .QN(n2553)
         );
  SDFSND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .SI(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ), .SE(n1037), 
        .CP(ClockB), .SDN(n4409), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters ), .QN(n2549)
         );
  SEDF4CCNQXD4 \SerDes_U1/Des_U1/DesDec_Rx1/ParClkr_reg  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N37 ), .SI(n1037), .E(
        \SerDes_U1/Des_U1/DesDec_Rx1/N43 ), .SE(n1037), .CP(n4475), .CDN(n3530), .Q(\SerDes_U1/Rx_ParClk ) );
  INVD16 U3311 ( .I(n3649), .ZN(n3651) );
  INVD16 U3312 ( .I(n3655), .ZN(n3657) );
  INVD16 U3313 ( .I(n3661), .ZN(n3663) );
  INVD16 U3314 ( .I(n3643), .ZN(n3645) );
  INVD16 U3315 ( .I(n3646), .ZN(n3648) );
  INVD16 U3316 ( .I(n3652), .ZN(n3654) );
  INVD16 U3317 ( .I(n3667), .ZN(n3669) );
  INVD16 U3318 ( .I(n3637), .ZN(n3639) );
  INVD16 U3319 ( .I(n3640), .ZN(n3642) );
  INVD16 U3320 ( .I(n3658), .ZN(n3660) );
  INVD16 U3321 ( .I(n3673), .ZN(n3675) );
  INVD16 U3322 ( .I(n3631), .ZN(n3633) );
  INVD16 U3323 ( .I(n3634), .ZN(n3636) );
  INVD16 U3324 ( .I(n3664), .ZN(n3666) );
  INVD16 U3325 ( .I(n3679), .ZN(n3681) );
  INVD16 U3326 ( .I(n3625), .ZN(n3627) );
  INVD16 U3327 ( .I(n3628), .ZN(n3630) );
  INVD16 U3328 ( .I(n3670), .ZN(n3672) );
  INVD16 U3329 ( .I(n3685), .ZN(n3687) );
  INVD16 U3330 ( .I(n3619), .ZN(n3621) );
  INVD16 U3331 ( .I(n3622), .ZN(n3624) );
  INVD16 U3332 ( .I(n3676), .ZN(n3678) );
  INVD16 U3333 ( .I(n3604), .ZN(n3606) );
  INVD16 U3334 ( .I(n3613), .ZN(n3615) );
  INVD16 U3335 ( .I(n3616), .ZN(n3618) );
  INVD16 U3336 ( .I(n3682), .ZN(n3684) );
  INVD16 U3337 ( .I(n3607), .ZN(n3609) );
  INVD16 U3338 ( .I(n3598), .ZN(n3600) );
  INVD16 U3339 ( .I(n3610), .ZN(n3612) );
  INVD16 U3340 ( .I(n3595), .ZN(n3597) );
  INVD16 U3341 ( .I(n3592), .ZN(n3594) );
  INVD16 U3342 ( .I(n3601), .ZN(n3603) );
  AN2D1 U3343 ( .A1(\SerDes_U2/Des_U1/SerialClk ), .A2(
        \SerDes_U2/SerLineValid ), .Z(\SerDes_U2/Des_U1/DesDec_Rx1/SerClock )
         );
  AN2D1 U3344 ( .A1(\SerDes_U1/Des_U1/SerialClk ), .A2(
        \SerDes_U1/SerLineValid ), .Z(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock )
         );
  NR2D1P5 U3345 ( .A1(\SerDes_U1/Tx_F_Empty ), .A2(Reset), .ZN(n3580) );
  INVD1 U3346 ( .I(Reset), .ZN(n3530) );
  NR2D1 U3347 ( .A1(n4996), .A2(n4999), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ) );
  NR2D1 U3348 ( .A1(n1023), .A2(n4987), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ) );
  NR2D1 U3349 ( .A1(n4996), .A2(n4997), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ) );
  NR2D1 U3350 ( .A1(n4994), .A2(n4997), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ) );
  NR2D1 U3351 ( .A1(n4995), .A2(n4996), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ) );
  NR2D1 U3352 ( .A1(n4988), .A2(n4999), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ) );
  NR2D1 U3353 ( .A1(n4989), .A2(n4999), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ) );
  NR2D1 U3354 ( .A1(n4988), .A2(n4998), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ) );
  NR2D1 U3355 ( .A1(n4995), .A2(n4989), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ) );
  NR2D1 U3356 ( .A1(n4764), .A2(n5075), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ) );
  NR2D1 U3357 ( .A1(n863), .A2(n5095), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ) );
  NR2D1 U3358 ( .A1(n5106), .A2(n5107), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ) );
  NR2D1 U3359 ( .A1(n5104), .A2(n5107), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ) );
  NR2D1 U3360 ( .A1(n5096), .A2(n5109), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ) );
  NR2D1 U3361 ( .A1(n5097), .A2(n5109), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ) );
  NR2D1 U3362 ( .A1(n4943), .A2(n5018), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ) );
  NR2D1 U3363 ( .A1(n4944), .A2(n5018), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ) );
  NR2D1 U3364 ( .A1(n4994), .A2(n4999), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ) );
  NR2D1 U3365 ( .A1(n4996), .A2(n4998), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ) );
  NR2D1 U3366 ( .A1(n4994), .A2(n4995), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ) );
  NR2D1 U3367 ( .A1(n4989), .A2(n4998), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ) );
  NR2D1 U3368 ( .A1(n4988), .A2(n4997), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ) );
  NR2D1 U3369 ( .A1(n4989), .A2(n4997), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ) );
  NR2D1 U3370 ( .A1(n4995), .A2(n4988), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ) );
  NR2D1 U3371 ( .A1(n4764), .A2(n5069), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ) );
  NR2D1 U3372 ( .A1(n4747), .A2(n5069), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ) );
  NR2D1 U3373 ( .A1(n4747), .A2(n5075), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ) );
  NR2D1 U3374 ( .A1(n5106), .A2(n5109), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ) );
  NR2D1 U3375 ( .A1(n5104), .A2(n5109), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ) );
  NR2D1 U3376 ( .A1(n5106), .A2(n5108), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ) );
  NR2D1 U3377 ( .A1(n5105), .A2(n5106), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ) );
  NR2D1 U3378 ( .A1(n5104), .A2(n5105), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ) );
  NR2D1 U3379 ( .A1(n5096), .A2(n5108), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ) );
  NR2D1 U3380 ( .A1(n5097), .A2(n5108), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ) );
  NR2D1 U3381 ( .A1(n5096), .A2(n5107), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ) );
  NR2D1 U3382 ( .A1(n5097), .A2(n5107), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ) );
  NR2D1 U3383 ( .A1(n5105), .A2(n5096), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ) );
  NR2D1 U3384 ( .A1(n5105), .A2(n5097), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ) );
  NR2D1 U3385 ( .A1(n4944), .A2(n5021), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ) );
  NR2D1 U3386 ( .A1(n4943), .A2(n5021), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ) );
  INR2D1 U3387 ( .A1(n5110), .B1(n5111), .ZN(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ) );
  INR2D1 U3388 ( .A1(n5022), .B1(n5023), .ZN(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ) );
  OR2D1 U3389 ( .A1(\SerDes_U2/Tx_F_Empty ), .A2(Reset), .Z(n3581) );
  MUX2ND0 U3390 ( .I0(n3760), .I1(n3761), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3583) );
  MUX2ND0 U3391 ( .I0(n3764), .I1(n3765), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3584) );
  MUX2ND0 U3392 ( .I0(n3752), .I1(n3753), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3585) );
  MUX2ND0 U3393 ( .I0(n3756), .I1(n3757), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3586) );
  MUX2ND0 U3394 ( .I0(n3762), .I1(n3763), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3588) );
  MUX2ND0 U3395 ( .I0(n3766), .I1(n3767), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3589) );
  MUX2ND0 U3396 ( .I0(n3754), .I1(n3755), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3590) );
  MUX2ND0 U3397 ( .I0(n3758), .I1(n3759), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n3591) );
  CKBXD0 U3398 ( .I(n4355), .Z(n3592) );
  CKNXD16 U3399 ( .I(n3592), .ZN(OutParDataA[16]) );
  CKBXD0 U3400 ( .I(n4354), .Z(n3595) );
  CKNXD16 U3401 ( .I(n3595), .ZN(OutParDataA[15]) );
  CKBXD0 U3402 ( .I(n4356), .Z(n3598) );
  CKNXD16 U3403 ( .I(n3598), .ZN(OutParDataA[17]) );
  CKBXD0 U3404 ( .I(n4353), .Z(n3601) );
  CKNXD16 U3405 ( .I(n3601), .ZN(OutParDataA[14]) );
  CKBXD0 U3406 ( .I(n4357), .Z(n3604) );
  CKNXD16 U3407 ( .I(n3604), .ZN(OutParDataA[18]) );
  CKBXD0 U3408 ( .I(n4352), .Z(n3607) );
  CKNXD16 U3409 ( .I(n3607), .ZN(OutParDataA[13]) );
  CKBXD0 U3410 ( .I(n4358), .Z(n3610) );
  CKNXD16 U3411 ( .I(n3610), .ZN(OutParDataA[19]) );
  CKBXD0 U3412 ( .I(n4351), .Z(n3613) );
  CKNXD16 U3413 ( .I(n3613), .ZN(OutParDataA[12]) );
  CKBXD0 U3414 ( .I(n4359), .Z(n3616) );
  CKNXD16 U3415 ( .I(n3616), .ZN(OutParDataA[20]) );
  CKBXD0 U3416 ( .I(n4350), .Z(n3619) );
  CKNXD16 U3417 ( .I(n3619), .ZN(OutParDataA[11]) );
  CKBXD0 U3418 ( .I(n4360), .Z(n3622) );
  CKNXD16 U3419 ( .I(n3622), .ZN(OutParDataA[21]) );
  CKBXD0 U3420 ( .I(n4349), .Z(n3625) );
  CKNXD16 U3421 ( .I(n3625), .ZN(OutParDataA[10]) );
  CKBXD0 U3422 ( .I(n4361), .Z(n3628) );
  CKNXD16 U3423 ( .I(n3628), .ZN(OutParDataA[22]) );
  CKBXD0 U3424 ( .I(n4348), .Z(n3631) );
  CKNXD16 U3425 ( .I(n3631), .ZN(OutParDataA[9]) );
  CKBXD0 U3426 ( .I(n4362), .Z(n3634) );
  CKNXD16 U3427 ( .I(n3634), .ZN(OutParDataA[23]) );
  CKBXD0 U3428 ( .I(n4347), .Z(n3637) );
  CKNXD16 U3429 ( .I(n3637), .ZN(OutParDataA[8]) );
  CKBXD0 U3430 ( .I(n4363), .Z(n3640) );
  CKNXD16 U3431 ( .I(n3640), .ZN(OutParDataA[24]) );
  CKBXD0 U3432 ( .I(n4346), .Z(n3643) );
  CKNXD16 U3433 ( .I(n3643), .ZN(OutParDataA[7]) );
  CKBXD0 U3434 ( .I(n4364), .Z(n3646) );
  CKNXD16 U3435 ( .I(n3646), .ZN(OutParDataA[25]) );
  CKBXD0 U3436 ( .I(n4345), .Z(n3649) );
  CKNXD16 U3437 ( .I(n3649), .ZN(OutParDataA[6]) );
  CKBXD0 U3438 ( .I(n4365), .Z(n3652) );
  CKNXD16 U3439 ( .I(n3652), .ZN(OutParDataA[26]) );
  CKBXD0 U3440 ( .I(n4344), .Z(n3655) );
  CKNXD16 U3441 ( .I(n3655), .ZN(OutParDataA[5]) );
  CKBXD0 U3442 ( .I(n4366), .Z(n3658) );
  CKNXD16 U3443 ( .I(n3658), .ZN(OutParDataA[27]) );
  CKBXD0 U3444 ( .I(n4343), .Z(n3661) );
  CKNXD16 U3445 ( .I(n3661), .ZN(OutParDataA[4]) );
  CKBXD0 U3446 ( .I(n4367), .Z(n3664) );
  CKNXD16 U3447 ( .I(n3664), .ZN(OutParDataA[28]) );
  CKBXD0 U3448 ( .I(n4342), .Z(n3667) );
  CKNXD16 U3449 ( .I(n3667), .ZN(OutParDataA[3]) );
  CKBXD0 U3450 ( .I(n4368), .Z(n3670) );
  CKNXD16 U3451 ( .I(n3670), .ZN(OutParDataA[29]) );
  CKBXD0 U3452 ( .I(n4341), .Z(n3673) );
  CKNXD16 U3453 ( .I(n3673), .ZN(OutParDataA[2]) );
  CKBXD0 U3454 ( .I(n4369), .Z(n3676) );
  CKNXD16 U3455 ( .I(n3676), .ZN(OutParDataA[30]) );
  CKBXD0 U3456 ( .I(n4340), .Z(n3679) );
  CKNXD16 U3457 ( .I(n3679), .ZN(OutParDataA[1]) );
  CKBXD0 U3458 ( .I(n4370), .Z(n3682) );
  CKNXD16 U3459 ( .I(n3682), .ZN(OutParDataA[31]) );
  CKBXD0 U3460 ( .I(n4339), .Z(n3685) );
  CKNXD16 U3461 ( .I(n3685), .ZN(OutParDataA[0]) );
  CKBD0 U3462 ( .CLK(n4338), .C(n3688) );
  CKND16 U3463 ( .CLK(n3688), .CN(OutParDataB[31]) );
  CKBD0 U3464 ( .CLK(n4337), .C(n3690) );
  CKND16 U3465 ( .CLK(n3690), .CN(OutParDataB[30]) );
  CKBD0 U3466 ( .CLK(n4336), .C(n3692) );
  CKND16 U3467 ( .CLK(n3692), .CN(OutParDataB[29]) );
  CKBD0 U3468 ( .CLK(n4335), .C(n3694) );
  CKND16 U3469 ( .CLK(n3694), .CN(OutParDataB[28]) );
  CKBD0 U3470 ( .CLK(n4334), .C(n3696) );
  CKND16 U3471 ( .CLK(n3696), .CN(OutParDataB[27]) );
  CKBD0 U3472 ( .CLK(n4333), .C(n3698) );
  CKND16 U3473 ( .CLK(n3698), .CN(OutParDataB[26]) );
  CKBD0 U3474 ( .CLK(n4332), .C(n3700) );
  CKND16 U3475 ( .CLK(n3700), .CN(OutParDataB[25]) );
  CKBD0 U3476 ( .CLK(n4331), .C(n3702) );
  CKND16 U3477 ( .CLK(n3702), .CN(OutParDataB[24]) );
  CKBD0 U3478 ( .CLK(n4330), .C(n3704) );
  CKND16 U3479 ( .CLK(n3704), .CN(OutParDataB[23]) );
  CKBD0 U3480 ( .CLK(n4329), .C(n3706) );
  CKND16 U3481 ( .CLK(n3706), .CN(OutParDataB[22]) );
  CKBD0 U3482 ( .CLK(n4328), .C(n3708) );
  CKND16 U3483 ( .CLK(n3708), .CN(OutParDataB[21]) );
  CKBD0 U3484 ( .CLK(n4327), .C(n3710) );
  CKND16 U3485 ( .CLK(n3710), .CN(OutParDataB[20]) );
  CKBD0 U3486 ( .CLK(n4326), .C(n3712) );
  CKND16 U3487 ( .CLK(n3712), .CN(OutParDataB[19]) );
  CKBD0 U3488 ( .CLK(n4325), .C(n3714) );
  CKND16 U3489 ( .CLK(n3714), .CN(OutParDataB[18]) );
  CKBD0 U3490 ( .CLK(n4324), .C(n3716) );
  CKND16 U3491 ( .CLK(n3716), .CN(OutParDataB[17]) );
  CKBD0 U3492 ( .CLK(n4323), .C(n3718) );
  CKND16 U3493 ( .CLK(n3718), .CN(OutParDataB[16]) );
  CKBD0 U3494 ( .CLK(n4322), .C(n3720) );
  CKND16 U3495 ( .CLK(n3720), .CN(OutParDataB[15]) );
  CKBD0 U3496 ( .CLK(n4321), .C(n3722) );
  CKND16 U3497 ( .CLK(n3722), .CN(OutParDataB[14]) );
  CKBD0 U3498 ( .CLK(n4320), .C(n3724) );
  CKND16 U3499 ( .CLK(n3724), .CN(OutParDataB[13]) );
  CKBD0 U3500 ( .CLK(n4319), .C(n3726) );
  CKND16 U3501 ( .CLK(n3726), .CN(OutParDataB[12]) );
  CKBD0 U3502 ( .CLK(n4318), .C(n3728) );
  CKND16 U3503 ( .CLK(n3728), .CN(OutParDataB[11]) );
  CKBD0 U3504 ( .CLK(n4317), .C(n3730) );
  CKND16 U3505 ( .CLK(n3730), .CN(OutParDataB[10]) );
  CKBD0 U3506 ( .CLK(n4316), .C(n3732) );
  CKND16 U3507 ( .CLK(n3732), .CN(OutParDataB[9]) );
  CKBD0 U3508 ( .CLK(n4315), .C(n3734) );
  CKND16 U3509 ( .CLK(n3734), .CN(OutParDataB[8]) );
  CKBD0 U3510 ( .CLK(n4314), .C(n3736) );
  CKND16 U3511 ( .CLK(n3736), .CN(OutParDataB[7]) );
  CKBD0 U3512 ( .CLK(n4313), .C(n3738) );
  CKND16 U3513 ( .CLK(n3738), .CN(OutParDataB[6]) );
  CKBD0 U3514 ( .CLK(n4312), .C(n3740) );
  CKND16 U3515 ( .CLK(n3740), .CN(OutParDataB[5]) );
  CKBD0 U3516 ( .CLK(n4311), .C(n3742) );
  CKND16 U3517 ( .CLK(n3742), .CN(OutParDataB[4]) );
  CKBD0 U3518 ( .CLK(n4310), .C(n3744) );
  CKND16 U3519 ( .CLK(n3744), .CN(OutParDataB[3]) );
  CKBD0 U3520 ( .CLK(n4309), .C(n3746) );
  CKND16 U3521 ( .CLK(n3746), .CN(OutParDataB[2]) );
  CKBD0 U3522 ( .CLK(n4308), .C(n3748) );
  CKND16 U3523 ( .CLK(n3748), .CN(OutParDataB[1]) );
  CKBD0 U3524 ( .CLK(n4307), .C(n3750) );
  CKND16 U3525 ( .CLK(n3750), .CN(OutParDataB[0]) );
  BUFFD1 U3526 ( .I(n4442), .Z(n4436) );
  BUFFD1 U3527 ( .I(n4442), .Z(n4435) );
  BUFFD1 U3528 ( .I(n4447), .Z(n4414) );
  BUFFD1 U3529 ( .I(n4447), .Z(n4413) );
  BUFFD1 U3530 ( .I(n4448), .Z(n4412) );
  BUFFD1 U3531 ( .I(n4448), .Z(n4409) );
  BUFFD1 U3532 ( .I(n4442), .Z(n4434) );
  BUFFD1 U3533 ( .I(n4448), .Z(n4410) );
  BUFFD1 U3534 ( .I(n4441), .Z(n4437) );
  BUFFD1 U3535 ( .I(n4447), .Z(n4415) );
  BUFFD1 U3536 ( .I(n4448), .Z(n4411) );
  BUFFD1 U3537 ( .I(n4446), .Z(n4418) );
  BUFFD1 U3538 ( .I(n4442), .Z(n4433) );
  BUFFD1 U3539 ( .I(n4443), .Z(n4431) );
  BUFFD1 U3540 ( .I(n4443), .Z(n4430) );
  BUFFD1 U3541 ( .I(n4443), .Z(n4429) );
  BUFFD1 U3542 ( .I(n4444), .Z(n4428) );
  BUFFD1 U3543 ( .I(n4444), .Z(n4427) );
  BUFFD1 U3544 ( .I(n4444), .Z(n4426) );
  BUFFD1 U3545 ( .I(n4443), .Z(n4432) );
  BUFFD1 U3546 ( .I(n4446), .Z(n4419) );
  BUFFD1 U3547 ( .I(n4445), .Z(n4422) );
  BUFFD1 U3548 ( .I(n4445), .Z(n4423) );
  BUFFD1 U3549 ( .I(n4444), .Z(n4425) );
  BUFFD1 U3550 ( .I(n4445), .Z(n4424) );
  BUFFD1 U3551 ( .I(n4445), .Z(n4421) );
  BUFFD1 U3552 ( .I(n4446), .Z(n4420) );
  BUFFD1 U3553 ( .I(n4446), .Z(n4417) );
  BUFFD1 U3554 ( .I(n4441), .Z(n4438) );
  BUFFD1 U3555 ( .I(n4441), .Z(n4439) );
  BUFFD1 U3556 ( .I(n4447), .Z(n4416) );
  BUFFD1 U3557 ( .I(n4452), .Z(n4394) );
  BUFFD1 U3558 ( .I(n4452), .Z(n4395) );
  BUFFD1 U3559 ( .I(n4452), .Z(n4396) );
  BUFFD1 U3560 ( .I(n4451), .Z(n4397) );
  BUFFD1 U3561 ( .I(n4451), .Z(n4398) );
  BUFFD1 U3562 ( .I(n4451), .Z(n4399) );
  BUFFD1 U3563 ( .I(n4451), .Z(n4400) );
  BUFFD1 U3564 ( .I(n4450), .Z(n4401) );
  BUFFD1 U3565 ( .I(n4450), .Z(n4403) );
  BUFFD1 U3566 ( .I(n4450), .Z(n4404) );
  BUFFD1 U3567 ( .I(n4449), .Z(n4406) );
  BUFFD1 U3568 ( .I(n4449), .Z(n4407) );
  BUFFD1 U3569 ( .I(n4449), .Z(n4408) );
  BUFFD1 U3570 ( .I(n4450), .Z(n4402) );
  BUFFD1 U3571 ( .I(n4449), .Z(n4405) );
  BUFFD1 U3572 ( .I(n4437), .Z(n4375) );
  BUFFD1 U3573 ( .I(n4456), .Z(n4376) );
  BUFFD1 U3574 ( .I(n4452), .Z(n4393) );
  BUFFD1 U3575 ( .I(n4454), .Z(n4387) );
  BUFFD1 U3576 ( .I(n4454), .Z(n4388) );
  BUFFD1 U3577 ( .I(n4453), .Z(n4389) );
  BUFFD1 U3578 ( .I(n4453), .Z(n4390) );
  BUFFD1 U3579 ( .I(n4453), .Z(n4391) );
  BUFFD1 U3580 ( .I(n4453), .Z(n4392) );
  BUFFD1 U3581 ( .I(n4456), .Z(n4377) );
  BUFFD1 U3582 ( .I(n4456), .Z(n4378) );
  BUFFD1 U3583 ( .I(n4456), .Z(n4379) );
  BUFFD1 U3584 ( .I(n4421), .Z(n4380) );
  BUFFD1 U3585 ( .I(n4455), .Z(n4381) );
  BUFFD1 U3586 ( .I(n4455), .Z(n4382) );
  BUFFD1 U3587 ( .I(n4455), .Z(n4383) );
  BUFFD1 U3588 ( .I(n4455), .Z(n4384) );
  BUFFD1 U3589 ( .I(n4454), .Z(n4385) );
  BUFFD1 U3590 ( .I(n4454), .Z(n4386) );
  BUFFD1 U3591 ( .I(n4441), .Z(n4440) );
  BUFFD1 U3592 ( .I(n4463), .Z(n4442) );
  BUFFD1 U3593 ( .I(n4462), .Z(n4443) );
  BUFFD1 U3594 ( .I(n4462), .Z(n4444) );
  BUFFD1 U3595 ( .I(n4461), .Z(n4445) );
  BUFFD1 U3596 ( .I(n4461), .Z(n4446) );
  BUFFD1 U3597 ( .I(n4458), .Z(n4451) );
  BUFFD1 U3598 ( .I(n4463), .Z(n4441) );
  BUFFD1 U3599 ( .I(n4459), .Z(n4450) );
  BUFFD1 U3600 ( .I(n4459), .Z(n4449) );
  BUFFD1 U3601 ( .I(n4458), .Z(n4452) );
  BUFFD1 U3602 ( .I(n4457), .Z(n4453) );
  BUFFD1 U3603 ( .I(n4396), .Z(n4456) );
  BUFFD1 U3604 ( .I(n4460), .Z(n4447) );
  BUFFD1 U3605 ( .I(n4446), .Z(n4455) );
  BUFFD1 U3606 ( .I(n4457), .Z(n4454) );
  BUFFD1 U3607 ( .I(n4460), .Z(n4448) );
  BUFFD1 U3608 ( .I(n4464), .Z(n4462) );
  BUFFD1 U3609 ( .I(n4464), .Z(n4461) );
  BUFFD1 U3610 ( .I(n4464), .Z(n4463) );
  BUFFD1 U3611 ( .I(n4465), .Z(n4459) );
  BUFFD1 U3612 ( .I(n4465), .Z(n4458) );
  BUFFD1 U3613 ( .I(n4379), .Z(n4457) );
  BUFFD1 U3614 ( .I(n4465), .Z(n4460) );
  BUFFD1 U3615 ( .I(n4466), .Z(n4464) );
  BUFFD1 U3616 ( .I(n4466), .Z(n4465) );
  INVD1 U3617 ( .I(n4565), .ZN(n4564) );
  INVD1 U3618 ( .I(n4529), .ZN(n4528) );
  INVD1 U3619 ( .I(n4571), .ZN(n4570) );
  INVD1 U3620 ( .I(n4492), .ZN(n4491) );
  INVD1 U3621 ( .I(n4535), .ZN(n4534) );
  BUFFD1 U3622 ( .I(n4306), .Z(n4305) );
  BUFFD1 U3623 ( .I(n4306), .Z(n4304) );
  BUFFD1 U3624 ( .I(n4203), .Z(n4202) );
  BUFFD1 U3625 ( .I(n4203), .Z(n4201) );
  BUFFD1 U3626 ( .I(n3947), .Z(n3951) );
  BUFFD1 U3627 ( .I(n3948), .Z(n3952) );
  BUFFD1 U3628 ( .I(n4089), .Z(n4090) );
  BUFFD1 U3629 ( .I(n3948), .Z(n3949) );
  BUFFD1 U3630 ( .I(n3948), .Z(n3950) );
  BUFFD1 U3631 ( .I(n4088), .Z(n4089) );
  BUFFD1 U3632 ( .I(n4087), .Z(n4091) );
  BUFFD1 U3633 ( .I(n4087), .Z(n4092) );
  BUFFD1 U3634 ( .I(n4306), .Z(n4303) );
  BUFFD1 U3635 ( .I(n4203), .Z(n4200) );
  BUFFD1 U3636 ( .I(n4302), .Z(n4301) );
  BUFFD1 U3637 ( .I(n3943), .Z(n3945) );
  BUFFD1 U3638 ( .I(n3943), .Z(n3946) );
  BUFFD1 U3639 ( .I(n4083), .Z(n4085) );
  BUFFD1 U3640 ( .I(n4083), .Z(n4086) );
  INVD1 U3641 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .ZN(n4565) );
  INVD1 U3642 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .ZN(n4529) );
  INVD1 U3643 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .ZN(n4571) );
  INVD1 U3644 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .ZN(n4535) );
  INVD1 U3645 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .ZN(n4492) );
  BUFFD1 U3646 ( .I(n4199), .Z(n4198) );
  BUFFD1 U3647 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3944) );
  BUFFD1 U3648 ( .I(n4083), .Z(n4084) );
  BUFFD1 U3649 ( .I(n4471), .Z(n4468) );
  BUFFD1 U3650 ( .I(n4471), .Z(n4467) );
  BUFFD1 U3651 ( .I(n4471), .Z(n4469) );
  BUFFD1 U3652 ( .I(n4476), .Z(n4474) );
  BUFFD1 U3653 ( .I(n4374), .Z(n4466) );
  INVD1 U3654 ( .I(n4501), .ZN(n4197) );
  INVD1 U3655 ( .I(n4482), .ZN(n4300) );
  INVD1 U3656 ( .I(n4526), .ZN(n4082) );
  INVD1 U3657 ( .I(n4562), .ZN(n3942) );
  INVD1 U3658 ( .I(n4563), .ZN(n3941) );
  INVD1 U3659 ( .I(n4527), .ZN(n4081) );
  BUFFD1 U3660 ( .I(n4467), .Z(n4470) );
  BUFFD1 U3661 ( .I(n4476), .Z(n4475) );
  INVD1 U3662 ( .I(n4488), .ZN(n4487) );
  INVD1 U3663 ( .I(n4490), .ZN(n4489) );
  INVD1 U3664 ( .I(n4573), .ZN(n4572) );
  INVD1 U3665 ( .I(n4581), .ZN(n4580) );
  INVD1 U3666 ( .I(n4589), .ZN(n4588) );
  INVD1 U3667 ( .I(n4591), .ZN(n4590) );
  INVD1 U3668 ( .I(n4593), .ZN(n4592) );
  INVD1 U3669 ( .I(n4509), .ZN(n4508) );
  INVD1 U3670 ( .I(n4507), .ZN(n4506) );
  INVD1 U3671 ( .I(n4537), .ZN(n4536) );
  INVD1 U3672 ( .I(n4545), .ZN(n4544) );
  INVD1 U3673 ( .I(n4553), .ZN(n4552) );
  INVD1 U3674 ( .I(n4555), .ZN(n4554) );
  INVD1 U3675 ( .I(n4557), .ZN(n4556) );
  INVD1 U3676 ( .I(n4494), .ZN(n4493) );
  INVD1 U3677 ( .I(n4567), .ZN(n4566) );
  INVD1 U3678 ( .I(n4569), .ZN(n4568) );
  INVD1 U3679 ( .I(n4575), .ZN(n4574) );
  INVD1 U3680 ( .I(n4577), .ZN(n4576) );
  INVD1 U3681 ( .I(n4583), .ZN(n4582) );
  INVD1 U3682 ( .I(n4585), .ZN(n4584) );
  INVD1 U3683 ( .I(n4587), .ZN(n4586) );
  INVD1 U3684 ( .I(n4595), .ZN(n4594) );
  INVD1 U3685 ( .I(n4513), .ZN(n4512) );
  INVD1 U3686 ( .I(n4531), .ZN(n4530) );
  INVD1 U3687 ( .I(n4533), .ZN(n4532) );
  INVD1 U3688 ( .I(n4541), .ZN(n4540) );
  INVD1 U3689 ( .I(n4549), .ZN(n4548) );
  INVD1 U3690 ( .I(n4511), .ZN(n4510) );
  INVD1 U3691 ( .I(n4539), .ZN(n4538) );
  INVD1 U3692 ( .I(n4547), .ZN(n4546) );
  INVD1 U3693 ( .I(n4551), .ZN(n4550) );
  INVD1 U3694 ( .I(n4559), .ZN(n4558) );
  INVD1 U3695 ( .I(n4496), .ZN(n4495) );
  INVD1 U3696 ( .I(n4498), .ZN(n4497) );
  INVD1 U3697 ( .I(n4517), .ZN(n4516) );
  INVD1 U3698 ( .I(n4515), .ZN(n4514) );
  INVD1 U3699 ( .I(n3581), .ZN(n4371) );
  INVD1 U3700 ( .I(n4473), .ZN(n4472) );
  INVD1 U3701 ( .I(n4479), .ZN(n4478) );
  INVD1 U3702 ( .I(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), .ZN(n4473) );
  INVD1 U3703 ( .I(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), .ZN(n4479) );
  INVD1 U3704 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .ZN(n4488) );
  INVD1 U3705 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .ZN(n4490) );
  INVD1 U3706 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .ZN(n4573) );
  INVD1 U3707 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .ZN(n4581) );
  INVD1 U3708 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .ZN(n4589) );
  INVD1 U3709 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .ZN(n4591) );
  INVD1 U3710 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .ZN(n4593) );
  INVD1 U3711 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .ZN(n4509) );
  INVD1 U3712 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .ZN(n4507) );
  INVD1 U3713 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .ZN(n4537) );
  INVD1 U3714 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .ZN(n4545) );
  INVD1 U3715 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .ZN(n4553) );
  INVD1 U3716 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .ZN(n4555) );
  INVD1 U3717 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .ZN(n4557) );
  INVD1 U3718 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .ZN(n4567) );
  INVD1 U3719 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .ZN(n4569) );
  INVD1 U3720 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .ZN(n4575) );
  INVD1 U3721 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .ZN(n4577) );
  INVD1 U3722 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .ZN(n4583) );
  INVD1 U3723 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .ZN(n4585) );
  INVD1 U3724 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .ZN(n4513) );
  INVD1 U3725 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .ZN(n4531) );
  INVD1 U3726 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .ZN(n4533) );
  INVD1 U3727 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .ZN(n4539) );
  INVD1 U3728 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .ZN(n4541) );
  INVD1 U3729 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .ZN(n4547) );
  INVD1 U3730 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .ZN(n4549) );
  INVD1 U3731 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .ZN(n4494) );
  INVD1 U3732 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .ZN(n4587) );
  INVD1 U3733 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .ZN(n4595) );
  INVD1 U3734 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .ZN(n4551) );
  INVD1 U3735 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .ZN(n4559) );
  INVD1 U3736 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .ZN(n4511) );
  INVD1 U3737 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .ZN(n4517) );
  INVD1 U3738 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .ZN(n4515) );
  INVD1 U3739 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .ZN(n4496) );
  INVD1 U3740 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .ZN(n4498) );
  BUFFD1 U3741 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .Z(n4306) );
  BUFFD1 U3742 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .Z(n4203) );
  BUFFD1 U3743 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .Z(n4302) );
  BUFFD1 U3744 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .Z(n4199) );
  BUFFD1 U3745 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .Z(n4088) );
  BUFFD1 U3746 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .Z(n3948) );
  BUFFD1 U3747 ( .I(n3530), .Z(n4374) );
  BUFFD1 U3748 ( .I(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .Z(n4477) );
  BUFFD1 U3749 ( .I(\SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .Z(n4471) );
  BUFFD1 U3750 ( .I(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .Z(n4476) );
  BUFFD1 U3751 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .Z(n4087) );
  BUFFD1 U3752 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3943) );
  BUFFD1 U3753 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .Z(n3947) );
  BUFFD1 U3754 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4083) );
  INVD1 U3755 ( .I(n4579), .ZN(n4578) );
  INVD1 U3756 ( .I(n4543), .ZN(n4542) );
  INVD1 U3757 ( .I(n761), .ZN(n4373) );
  INVD1 U3758 ( .I(n909), .ZN(n4372) );
  INVD1 U3759 ( .I(n4484), .ZN(n4483) );
  INVD1 U3760 ( .I(n4486), .ZN(n4485) );
  INVD1 U3761 ( .I(n4505), .ZN(n4504) );
  INVD1 U3762 ( .I(n4503), .ZN(n4502) );
  INVD1 U3763 ( .I(n721), .ZN(n4518) );
  INVD1 U3764 ( .I(n869), .ZN(n4597) );
  INVD1 U3765 ( .I(n1015), .ZN(n4519) );
  INVD1 U3766 ( .I(n3587), .ZN(n4596) );
  INVD1 U3767 ( .I(n4521), .ZN(n4520) );
  INVD1 U3768 ( .I(n4523), .ZN(n4522) );
  INVD1 U3769 ( .I(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .ZN(n4521) );
  INVD1 U3770 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .ZN(n4579) );
  INVD1 U3771 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .ZN(n4543) );
  INVD1 U3772 ( .I(\SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .ZN(n4523) );
  INVD1 U3773 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .ZN(n4484) );
  INVD1 U3774 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .ZN(n4486) );
  INVD1 U3775 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .ZN(n4505) );
  INVD1 U3776 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .ZN(n4503) );
  INVD1 U3777 ( .I(n4605), .ZN(n4602) );
  INVD1 U3778 ( .I(n4601), .ZN(n4598) );
  MUX4ND0 U3779 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .S0(n4303), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4224) );
  MUX4ND0 U3780 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4227) );
  MUX4ND0 U3781 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .S0(n4306), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4230) );
  MUX4ND0 U3782 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4233) );
  MUX4ND0 U3783 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .S0(n4306), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4236) );
  MUX4ND0 U3784 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4239) );
  MUX4ND0 U3785 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .S0(n4306), 
        .S1(n4302), .ZN(n4242) );
  MUX4ND0 U3786 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4245) );
  MUX4ND0 U3787 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .S0(n4306), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4248) );
  MUX4ND0 U3788 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4251) );
  MUX4ND0 U3789 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .S0(n4306), 
        .S1(n4302), .ZN(n4254) );
  MUX4ND0 U3790 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4257) );
  MUX4ND0 U3791 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .S0(n4306), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4260) );
  MUX4ND0 U3792 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4263) );
  MUX4ND0 U3793 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .S0(n4306), 
        .S1(n4302), .ZN(n4266) );
  MUX4ND0 U3794 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4281) );
  MUX4ND0 U3795 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4284) );
  MUX4ND0 U3796 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .S0(n4303), 
        .S1(n4301), .ZN(n4287) );
  MUX4ND0 U3797 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .S0(n4305), 
        .S1(n4302), .ZN(n4290) );
  MUX4ND0 U3798 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .S0(n4203), 
        .S1(n4198), .ZN(n4187) );
  MUX4ND0 U3799 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .S0(n4200), 
        .S1(n4198), .ZN(n4184) );
  MUX4ND0 U3800 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4198), .ZN(n4181) );
  MUX4ND0 U3801 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4198), .ZN(n4178) );
  MUX4ND0 U3802 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .S0(n4203), 
        .S1(n4198), .ZN(n4163) );
  MUX4ND0 U3803 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4160) );
  MUX4ND0 U3804 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .S0(n4200), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4157) );
  MUX4ND0 U3805 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .S0(n4203), 
        .S1(n4199), .ZN(n4154) );
  MUX4ND0 U3806 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4151) );
  MUX4ND0 U3807 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .S0(n4203), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4148) );
  MUX4ND0 U3808 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .S0(n4203), 
        .S1(n4199), .ZN(n4145) );
  MUX4ND0 U3809 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .S0(n4203), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4142) );
  MUX4ND0 U3810 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4199), .ZN(n4139) );
  MUX4ND0 U3811 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4199), .ZN(n4136) );
  MUX4ND0 U3812 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .S0(n4203), 
        .S1(n4199), .ZN(n4133) );
  MUX4ND0 U3813 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .S0(n4203), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4130) );
  MUX4ND0 U3814 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4199), .ZN(n4127) );
  MUX4ND0 U3815 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .S0(n4203), .S1(
        n4199), .ZN(n4124) );
  MUX4ND0 U3816 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4121) );
  MUX4ND0 U3817 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4206) );
  MUX4ND0 U3818 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4209) );
  MUX4ND0 U3819 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .S0(n4306), .S1(
        n4302), .ZN(n4212) );
  MUX4ND0 U3820 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n4302), .ZN(n4215) );
  MUX4ND0 U3821 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .S0(n4306), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4218) );
  MUX4ND0 U3822 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .S0(n4303), .S1(
        n4301), .ZN(n4221) );
  MUX4ND0 U3823 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .S0(n4306), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4269) );
  MUX4ND0 U3824 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .S0(n4306), 
        .S1(n4302), .ZN(n4272) );
  MUX4ND0 U3825 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .S0(n4306), 
        .S1(n4302), .ZN(n4275) );
  MUX4ND0 U3826 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .S0(n4306), 
        .S1(n4302), .ZN(n4278) );
  MUX4ND0 U3827 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .S0(n4306), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4293) );
  MUX4ND0 U3828 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .S0(n4306), 
        .S1(n4302), .ZN(n4296) );
  MUX4ND0 U3829 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .S0(n4304), 
        .S1(n4302), .ZN(n4299) );
  MUX4ND0 U3830 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .S0(n4203), 
        .S1(n4198), .ZN(n4196) );
  MUX4ND0 U3831 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4198), .ZN(n4193) );
  MUX4ND0 U3832 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4198), .ZN(n4190) );
  MUX4ND0 U3833 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .S0(n4203), 
        .S1(n4198), .ZN(n4175) );
  MUX4ND0 U3834 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .S0(n4202), 
        .S1(n4198), .ZN(n4172) );
  MUX4ND0 U3835 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .S0(n4203), 
        .S1(n4198), .ZN(n4169) );
  MUX4ND0 U3836 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .S0(n4201), 
        .S1(n4198), .ZN(n4166) );
  MUX4ND0 U3837 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4199), .ZN(n4118) );
  MUX4ND0 U3838 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .S0(n4203), .S1(
        n4198), .ZN(n4115) );
  MUX4ND0 U3839 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .S0(n4200), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4112) );
  MUX4ND0 U3840 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n4199), .ZN(n4109) );
  MUX4ND0 U3841 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .S0(n4203), .S1(
        n4198), .ZN(n4106) );
  MUX4ND0 U3842 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .S0(n4203), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4103) );
  AN2D1 U3843 ( .A1(n4602), .A2(n4603), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N24 )
         );
  AN2D1 U3844 ( .A1(n4598), .A2(n4599), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N24 )
         );
  ND2D1 U3845 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .ZN(n4605) );
  ND2D1 U3846 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .ZN(n4601) );
  INVD1 U3847 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .ZN(n4562) );
  MUX4D0 U3848 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ), .S0(n3949), 
        .S1(n3945), .Z(n3821) );
  MUX4D0 U3849 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ), .S0(n3949), 
        .S1(n3945), .Z(n3825) );
  MUX4D0 U3850 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ), .S0(n3949), 
        .S1(n3945), .Z(n3829) );
  MUX4D0 U3851 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ), .S0(n3950), 
        .S1(n3946), .Z(n3833) );
  MUX4D0 U3852 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ), .S0(n3950), 
        .S1(n3946), .Z(n3837) );
  MUX4D0 U3853 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ), .S0(n3950), 
        .S1(n3946), .Z(n3841) );
  MUX4D0 U3854 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ), .S0(n3951), 
        .S1(n3944), .Z(n3845) );
  MUX4D0 U3855 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ), .S0(n3948), 
        .S1(n3944), .Z(n3849) );
  MUX4D0 U3856 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ), .S0(n3947), 
        .S1(n3944), .Z(n3853) );
  MUX4D0 U3857 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ), .S0(n3948), 
        .S1(n3943), .Z(n3857) );
  MUX4D0 U3858 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ), .S0(n3947), 
        .S1(n3946), .Z(n3861) );
  MUX4D0 U3859 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3865) );
  MUX4D0 U3860 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ), .S0(n3948), 
        .S1(n3945), .Z(n3869) );
  MUX4D0 U3861 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ), .S0(n3947), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3873) );
  MUX4D0 U3862 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ), .S0(n3947), 
        .S1(n3946), .Z(n3877) );
  MUX4D0 U3863 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ), .S0(n3951), 
        .S1(n3945), .Z(n3881) );
  MUX4D0 U3864 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ), .S0(n3951), 
        .S1(n3943), .Z(n3885) );
  MUX4D0 U3865 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ), .S0(n3951), 
        .S1(n3944), .Z(n3889) );
  MUX4D0 U3866 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ), .S0(n3952), 
        .S1(n3943), .Z(n3893) );
  MUX4D0 U3867 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ), .S0(n3949), 
        .S1(n3944), .Z(n3897) );
  MUX4D0 U3868 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ), .S0(n3950), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3901) );
  MUX4D0 U3869 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ), .S0(n3952), 
        .S1(n3943), .Z(n3905) );
  MUX4D0 U3870 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ), .S0(n3952), 
        .S1(n3943), .Z(n3909) );
  MUX4D0 U3871 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ), .S0(n3952), 
        .S1(n3943), .Z(n3913) );
  MUX4D0 U3872 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ), .S0(n3951), 
        .S1(n3944), .Z(n3917) );
  MUX4D0 U3873 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ), .S0(n3951), 
        .S1(n3946), .Z(n3921) );
  MUX4D0 U3874 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ), .S0(n3952), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3925) );
  MUX4D0 U3875 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ), .S0(n3950), 
        .S1(n3944), .Z(n3929) );
  MUX4D0 U3876 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ), .S0(n3947), 
        .S1(n3943), .Z(n3933) );
  MUX4D0 U3877 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ), .S0(n3947), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3937) );
  MUX4D0 U3878 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ), .S0(n4089), 
        .S1(n4085), .Z(n3961) );
  MUX4D0 U3879 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ), .S0(n4089), 
        .S1(n4083), .Z(n3965) );
  MUX4D0 U3880 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ), .S0(n4089), 
        .S1(n4083), .Z(n3969) );
  MUX4D0 U3881 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ), .S0(n4091), 
        .S1(n4085), .Z(n3973) );
  MUX4D0 U3882 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ), .S0(n4092), 
        .S1(n4085), .Z(n3977) );
  MUX4D0 U3883 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ), .S0(n4088), 
        .S1(n4085), .Z(n3981) );
  MUX4D0 U3884 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ), .S0(n4089), 
        .S1(n4084), .Z(n3985) );
  MUX4D0 U3885 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ), .S0(n4092), 
        .S1(n4085), .Z(n3989) );
  MUX4D0 U3886 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ), .S0(n4091), 
        .S1(n4086), .Z(n3993) );
  MUX4D0 U3887 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ), .S0(n4091), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n3997) );
  MUX4D0 U3888 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ), .S0(n4092), 
        .S1(n4084), .Z(n4001) );
  MUX4D0 U3889 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ), .S0(n4088), 
        .S1(n4085), .Z(n4005) );
  MUX4D0 U3890 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ), .S0(n4088), 
        .S1(n4083), .Z(n4009) );
  MUX4D0 U3891 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4013) );
  MUX4D0 U3892 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4017) );
  MUX4D0 U3893 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ), .S0(n4087), 
        .S1(n4085), .Z(n4021) );
  MUX4D0 U3894 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ), .S0(n4089), 
        .S1(n4086), .Z(n4025) );
  MUX4D0 U3895 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ), .S0(n4088), 
        .S1(n4083), .Z(n4029) );
  MUX4D0 U3896 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ), .S0(n4088), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4033) );
  MUX4D0 U3897 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ), .S0(n4087), 
        .S1(n4084), .Z(n4037) );
  MUX4D0 U3898 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ), .S0(n4087), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4041) );
  MUX4D0 U3899 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ), .S0(n4090), 
        .S1(n4084), .Z(n4045) );
  MUX4D0 U3900 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ), .S0(n4090), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4049) );
  MUX4D0 U3901 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ), .S0(n4090), 
        .S1(n4083), .Z(n4053) );
  MUX4D0 U3902 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ), .S0(n4091), 
        .S1(n4086), .Z(n4057) );
  MUX4D0 U3903 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ), .S0(n4091), 
        .S1(n4086), .Z(n4061) );
  MUX4D0 U3904 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ), .S0(n4091), 
        .S1(n4086), .Z(n4065) );
  MUX4D0 U3905 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ), .S0(n4092), 
        .S1(n4086), .Z(n4069) );
  MUX4D0 U3906 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ), .S0(n4092), 
        .S1(n4083), .Z(n4073) );
  MUX4D0 U3907 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ), .S0(n4092), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4077) );
  MUX4D0 U3908 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3813) );
  MUX4D0 U3909 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ), .S0(n3947), 
        .S1(n3944), .Z(n3817) );
  MUX4D0 U3910 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ), .S0(n4088), 
        .S1(n4084), .Z(n3953) );
  MUX4D0 U3911 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4084), .Z(n3957) );
  INVD1 U3912 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(n4482) );
  MUX4ND0 U3913 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3752) );
  MUX4ND0 U3914 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3753) );
  MUX4ND0 U3915 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3754) );
  MUX4ND0 U3916 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3755) );
  MUX4ND0 U3917 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3756) );
  MUX4ND0 U3918 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3757) );
  MUX4ND0 U3919 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3758) );
  MUX4ND0 U3920 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3759) );
  MUX4ND0 U3921 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3760) );
  MUX4ND0 U3922 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3761) );
  MUX4ND0 U3923 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3762) );
  MUX4ND0 U3924 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3763) );
  MUX4ND0 U3925 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3764) );
  MUX4ND0 U3926 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3765) );
  MUX4ND0 U3927 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3766) );
  MUX4ND0 U3928 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n3767) );
  INVD1 U3929 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .ZN(n4563) );
  INVD1 U3930 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .ZN(n4526) );
  INVD1 U3931 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .ZN(n4525) );
  INVD1 U3932 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .ZN(n4527) );
  INVD1 U3933 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n4481) );
  INVD1 U3934 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .ZN(n4561) );
  INVD1 U3935 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(n4501) );
  INVD1 U3936 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n4500) );
  INVD1 U3937 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .ZN(n4560) );
  INVD1 U3938 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .ZN(n4524) );
  MUX4D0 U3939 ( .I0(n3816), .I1(n3814), .I2(n3815), .I3(n3813), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ) );
  MUX4D0 U3940 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .S0(n3952), .S1(
        n3944), .Z(n3815) );
  MUX4D0 U3941 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ), .S0(n3951), 
        .S1(n3944), .Z(n3814) );
  MUX4D0 U3942 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .S0(n3948), .S1(
        n3944), .Z(n3816) );
  MUX4D0 U3943 ( .I0(n3820), .I1(n3818), .I2(n3819), .I3(n3817), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ) );
  MUX4D0 U3944 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3819) );
  MUX4D0 U3945 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ), .S0(n3950), 
        .S1(n3944), .Z(n3818) );
  MUX4D0 U3946 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .S0(n3949), .S1(
        n3944), .Z(n3820) );
  MUX4D0 U3947 ( .I0(n3824), .I1(n3822), .I2(n3823), .I3(n3821), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ) );
  MUX4D0 U3948 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .S0(n3949), .S1(
        n3945), .Z(n3823) );
  MUX4D0 U3949 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ), .S0(n3949), 
        .S1(n3945), .Z(n3822) );
  MUX4D0 U3950 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .S0(n3949), .S1(
        n3945), .Z(n3824) );
  MUX4D0 U3951 ( .I0(n3828), .I1(n3826), .I2(n3827), .I3(n3825), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ) );
  MUX4D0 U3952 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .S0(n3949), .S1(
        n3945), .Z(n3827) );
  MUX4D0 U3953 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ), .S0(n3949), 
        .S1(n3945), .Z(n3826) );
  MUX4D0 U3954 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .S0(n3949), .S1(
        n3945), .Z(n3828) );
  MUX4D0 U3955 ( .I0(n3832), .I1(n3830), .I2(n3831), .I3(n3829), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ) );
  MUX4D0 U3956 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .S0(n3949), .S1(
        n3945), .Z(n3831) );
  MUX4D0 U3957 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ), .S0(n3949), 
        .S1(n3945), .Z(n3830) );
  MUX4D0 U3958 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .S0(n3949), .S1(
        n3945), .Z(n3832) );
  MUX4D0 U3959 ( .I0(n3836), .I1(n3834), .I2(n3835), .I3(n3833), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ) );
  MUX4D0 U3960 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .S0(n3950), .S1(
        n3946), .Z(n3835) );
  MUX4D0 U3961 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ), .S0(n3950), 
        .S1(n3946), .Z(n3834) );
  MUX4D0 U3962 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .S0(n3950), .S1(
        n3946), .Z(n3836) );
  MUX4D0 U3963 ( .I0(n3840), .I1(n3838), .I2(n3839), .I3(n3837), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ) );
  MUX4D0 U3964 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .S0(n3950), .S1(
        n3946), .Z(n3839) );
  MUX4D0 U3965 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ), .S0(n3950), 
        .S1(n3946), .Z(n3838) );
  MUX4D0 U3966 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .S0(n3950), .S1(
        n3946), .Z(n3840) );
  MUX4D0 U3967 ( .I0(n3844), .I1(n3842), .I2(n3843), .I3(n3841), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ) );
  MUX4D0 U3968 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .S0(n3950), .S1(
        n3946), .Z(n3843) );
  MUX4D0 U3969 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ), .S0(n3950), 
        .S1(n3946), .Z(n3842) );
  MUX4D0 U3970 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .S0(n3950), .S1(
        n3946), .Z(n3844) );
  MUX4D0 U3971 ( .I0(n3848), .I1(n3846), .I2(n3847), .I3(n3845), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ) );
  MUX4D0 U3972 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .S0(n3952), .S1(
        n3944), .Z(n3847) );
  MUX4D0 U3973 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3846) );
  MUX4D0 U3974 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3943), .Z(n3848) );
  MUX4D0 U3975 ( .I0(n3852), .I1(n3850), .I2(n3851), .I3(n3849), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ) );
  MUX4D0 U3976 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3943), .Z(n3851) );
  MUX4D0 U3977 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ), .S0(n3947), 
        .S1(n3946), .Z(n3850) );
  MUX4D0 U3978 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .S0(n3948), .S1(
        n3945), .Z(n3852) );
  MUX4D0 U3979 ( .I0(n3856), .I1(n3854), .I2(n3855), .I3(n3853), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ) );
  MUX4D0 U3980 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .S0(n3947), 
        .S1(n3943), .Z(n3855) );
  MUX4D0 U3981 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ), .S0(n3949), 
        .S1(n3946), .Z(n3854) );
  MUX4D0 U3982 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .S0(n3947), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3856) );
  MUX4D0 U3983 ( .I0(n3860), .I1(n3858), .I2(n3859), .I3(n3857), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ) );
  MUX4D0 U3984 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .S0(n3947), 
        .S1(n3945), .Z(n3859) );
  MUX4D0 U3985 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ), .S0(n3948), 
        .S1(n3943), .Z(n3858) );
  MUX4D0 U3986 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3860) );
  MUX4D0 U3987 ( .I0(n3864), .I1(n3862), .I2(n3863), .I3(n3861), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ) );
  MUX4D0 U3988 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .S0(n3948), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3863) );
  MUX4D0 U3989 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ), .S0(n3950), 
        .S1(n3945), .Z(n3862) );
  MUX4D0 U3990 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3946), .Z(n3864) );
  MUX4D0 U3991 ( .I0(n3868), .I1(n3866), .I2(n3867), .I3(n3865), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ) );
  MUX4D0 U3992 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .S0(n3948), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3867) );
  MUX4D0 U3993 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ), .S0(n3947), 
        .S1(n3945), .Z(n3866) );
  MUX4D0 U3994 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .S0(n3947), 
        .S1(n3943), .Z(n3868) );
  MUX4D0 U3995 ( .I0(n3872), .I1(n3870), .I2(n3871), .I3(n3869), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ) );
  MUX4D0 U3996 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .S0(n3947), 
        .S1(n3944), .Z(n3871) );
  MUX4D0 U3997 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ), .S0(n3948), 
        .S1(n3945), .Z(n3870) );
  MUX4D0 U3998 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3946), .Z(n3872) );
  MUX4D0 U3999 ( .I0(n3876), .I1(n3874), .I2(n3875), .I3(n3873), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ) );
  MUX4D0 U4000 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .S0(n3947), 
        .S1(n3943), .Z(n3875) );
  MUX4D0 U4001 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ), .S0(n3948), 
        .S1(n3945), .Z(n3874) );
  MUX4D0 U4002 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .S0(n3949), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3876) );
  MUX4D0 U4003 ( .I0(n3880), .I1(n3878), .I2(n3879), .I3(n3877), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ) );
  MUX4D0 U4004 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3879) );
  MUX4D0 U4005 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ), .S0(n3948), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3878) );
  MUX4D0 U4006 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3880) );
  MUX4D0 U4007 ( .I0(n3884), .I1(n3882), .I2(n3883), .I3(n3881), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ) );
  MUX4D0 U4008 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .S0(n3951), 
        .S1(n3944), .Z(n3883) );
  MUX4D0 U4009 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ), .S0(n3951), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3882) );
  MUX4D0 U4010 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .S0(n3951), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3884) );
  MUX4D0 U4011 ( .I0(n3888), .I1(n3886), .I2(n3887), .I3(n3885), .S0(n3941), 
        .S1(n3942), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ) );
  MUX4D0 U4012 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .S0(n3951), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3887) );
  MUX4D0 U4013 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ), .S0(n3951), 
        .S1(n3944), .Z(n3886) );
  MUX4D0 U4014 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .S0(n3951), 
        .S1(n3943), .Z(n3888) );
  MUX4D0 U4015 ( .I0(n3892), .I1(n3890), .I2(n3891), .I3(n3889), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ) );
  MUX4D0 U4016 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .S0(n3951), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3891) );
  MUX4D0 U4017 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ), .S0(n3951), 
        .S1(n3943), .Z(n3890) );
  MUX4D0 U4018 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .S0(n3951), 
        .S1(n3946), .Z(n3892) );
  MUX4D0 U4019 ( .I0(n3896), .I1(n3894), .I2(n3895), .I3(n3893), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ) );
  MUX4D0 U4020 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .S0(n3948), 
        .S1(n3943), .Z(n3895) );
  MUX4D0 U4021 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ), .S0(n3951), 
        .S1(n3945), .Z(n3894) );
  MUX4D0 U4022 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .S0(n3948), 
        .S1(n3946), .Z(n3896) );
  MUX4D0 U4023 ( .I0(n3900), .I1(n3898), .I2(n3899), .I3(n3897), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ) );
  MUX4D0 U4024 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .S0(n3952), 
        .S1(n3946), .Z(n3899) );
  MUX4D0 U4025 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ), .S0(n3947), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3898) );
  MUX4D0 U4026 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3900) );
  MUX4D0 U4027 ( .I0(n3904), .I1(n3902), .I2(n3903), .I3(n3901), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ) );
  MUX4D0 U4028 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .S0(n3947), 
        .S1(n3944), .Z(n3903) );
  MUX4D0 U4029 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ), .S0(n3950), 
        .S1(n3946), .Z(n3902) );
  MUX4D0 U4030 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .S0(n3949), 
        .S1(n3943), .Z(n3904) );
  MUX4D0 U4031 ( .I0(n3908), .I1(n3906), .I2(n3907), .I3(n3905), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ) );
  MUX4D0 U4032 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .S0(n3952), 
        .S1(n3943), .Z(n3907) );
  MUX4D0 U4033 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ), .S0(n3952), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3906) );
  MUX4D0 U4034 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .S0(n3952), 
        .S1(n3945), .Z(n3908) );
  MUX4D0 U4035 ( .I0(n3912), .I1(n3910), .I2(n3911), .I3(n3909), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ) );
  MUX4D0 U4036 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .S0(n3952), 
        .S1(n3943), .Z(n3911) );
  MUX4D0 U4037 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ), .S0(n3952), 
        .S1(n3943), .Z(n3910) );
  MUX4D0 U4038 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .S0(n3952), 
        .S1(n3943), .Z(n3912) );
  MUX4D0 U4039 ( .I0(n3916), .I1(n3914), .I2(n3915), .I3(n3913), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ) );
  MUX4D0 U4040 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .S0(n3952), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3915) );
  MUX4D0 U4041 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ), .S0(n3952), 
        .S1(n3945), .Z(n3914) );
  MUX4D0 U4042 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .S0(n3952), 
        .S1(n3944), .Z(n3916) );
  MUX4D0 U4043 ( .I0(n3920), .I1(n3918), .I2(n3919), .I3(n3917), .S0(n3941), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ) );
  MUX4D0 U4044 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3945), .Z(n3919) );
  MUX4D0 U4045 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ), .S0(n3950), 
        .S1(n3944), .Z(n3918) );
  MUX4D0 U4046 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .S0(n3949), 
        .S1(n3943), .Z(n3920) );
  MUX4D0 U4047 ( .I0(n3924), .I1(n3922), .I2(n3923), .I3(n3921), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ) );
  MUX4D0 U4048 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .S0(n3947), 
        .S1(n3943), .Z(n3923) );
  MUX4D0 U4049 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ), .S0(n3948), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3922) );
  MUX4D0 U4050 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3946), .Z(n3924) );
  MUX4D0 U4051 ( .I0(n3928), .I1(n3926), .I2(n3927), .I3(n3925), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ) );
  MUX4D0 U4052 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .S0(n3948), 
        .S1(n3946), .Z(n3927) );
  MUX4D0 U4053 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3944), .Z(n3926) );
  MUX4D0 U4054 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .S0(n3951), 
        .S1(n3945), .Z(n3928) );
  MUX4D0 U4055 ( .I0(n3932), .I1(n3930), .I2(n3931), .I3(n3929), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ) );
  MUX4D0 U4056 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .S0(n3951), 
        .S1(n3945), .Z(n3931) );
  MUX4D0 U4057 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ), .S0(n3948), 
        .S1(n3946), .Z(n3930) );
  MUX4D0 U4058 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n3945), .Z(n3932) );
  MUX4D0 U4059 ( .I0(n3936), .I1(n3934), .I2(n3935), .I3(n3933), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ) );
  MUX4D0 U4060 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .S0(n3950), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3935) );
  MUX4D0 U4061 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ), .S0(n3949), 
        .S1(n3943), .Z(n3934) );
  MUX4D0 U4062 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .S0(n3952), 
        .S1(n3944), .Z(n3936) );
  MUX4D0 U4063 ( .I0(n3940), .I1(n3938), .I2(n3939), .I3(n3937), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n3942), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ) );
  MUX4D0 U4064 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .S0(n3952), 
        .S1(n3946), .Z(n3939) );
  MUX4D0 U4065 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ), .S0(n3947), 
        .S1(n3943), .Z(n3938) );
  MUX4D0 U4066 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .S0(n3948), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n3940) );
  MUX4D0 U4067 ( .I0(n3956), .I1(n3954), .I2(n3955), .I3(n3953), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ) );
  MUX4D0 U4068 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .S0(n4092), .S1(
        n4084), .Z(n3955) );
  MUX4D0 U4069 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ), .S0(n4091), 
        .S1(n4084), .Z(n3954) );
  MUX4D0 U4070 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .S0(n4090), .S1(
        n4084), .Z(n3956) );
  MUX4D0 U4071 ( .I0(n3960), .I1(n3958), .I2(n3959), .I3(n3957), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ) );
  MUX4D0 U4072 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .S0(n4088), .S1(
        n4084), .Z(n3959) );
  MUX4D0 U4073 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ), .S0(n4090), 
        .S1(n4084), .Z(n3958) );
  MUX4D0 U4074 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .S0(n4090), .S1(
        n4084), .Z(n3960) );
  MUX4D0 U4075 ( .I0(n3964), .I1(n3962), .I2(n3963), .I3(n3961), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ) );
  MUX4D0 U4076 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .S0(n4089), .S1(
        n4085), .Z(n3963) );
  MUX4D0 U4077 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ), .S0(n4089), 
        .S1(n4086), .Z(n3962) );
  MUX4D0 U4078 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .S0(n4089), .S1(
        n4085), .Z(n3964) );
  MUX4D0 U4079 ( .I0(n3968), .I1(n3966), .I2(n3967), .I3(n3965), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ) );
  MUX4D0 U4080 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .S0(n4089), .S1(
        n4083), .Z(n3967) );
  MUX4D0 U4081 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ), .S0(n4089), 
        .S1(n4083), .Z(n3966) );
  MUX4D0 U4082 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .S0(n4089), .S1(
        n4083), .Z(n3968) );
  MUX4D0 U4083 ( .I0(n3972), .I1(n3970), .I2(n3971), .I3(n3969), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ) );
  MUX4D0 U4084 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .S0(n4089), .S1(
        n4086), .Z(n3971) );
  MUX4D0 U4085 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ), .S0(n4089), 
        .S1(n4083), .Z(n3970) );
  MUX4D0 U4086 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .S0(n4089), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n3972) );
  MUX4D0 U4087 ( .I0(n3976), .I1(n3974), .I2(n3975), .I3(n3973), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ) );
  MUX4D0 U4088 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4085), .Z(n3975) );
  MUX4D0 U4089 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ), .S0(n4087), 
        .S1(n4085), .Z(n3974) );
  MUX4D0 U4090 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .S0(n4089), .S1(
        n4085), .Z(n3976) );
  MUX4D0 U4091 ( .I0(n3980), .I1(n3978), .I2(n3979), .I3(n3977), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ) );
  MUX4D0 U4092 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .S0(n4092), .S1(
        n4085), .Z(n3979) );
  MUX4D0 U4093 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ), .S0(n4091), 
        .S1(n4085), .Z(n3978) );
  MUX4D0 U4094 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .S0(n4090), .S1(
        n4085), .Z(n3980) );
  MUX4D0 U4095 ( .I0(n3984), .I1(n3982), .I2(n3983), .I3(n3981), .S0(n4081), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ) );
  MUX4D0 U4096 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .S0(n4087), .S1(
        n4085), .Z(n3983) );
  MUX4D0 U4097 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ), .S0(n4089), 
        .S1(n4085), .Z(n3982) );
  MUX4D0 U4098 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .S0(n4088), .S1(
        n4085), .Z(n3984) );
  MUX4D0 U4099 ( .I0(n3988), .I1(n3986), .I2(n3987), .I3(n3985), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ) );
  MUX4D0 U4100 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4083), .Z(n3987) );
  MUX4D0 U4101 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n3986) );
  MUX4D0 U4102 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .S0(n4088), .S1(
        n4085), .Z(n3988) );
  MUX4D0 U4103 ( .I0(n3992), .I1(n3990), .I2(n3991), .I3(n3989), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ) );
  MUX4D0 U4104 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4086), .Z(n3991) );
  MUX4D0 U4105 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ), .S0(n4090), 
        .S1(n4084), .Z(n3990) );
  MUX4D0 U4106 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .S0(n4087), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n3992) );
  MUX4D0 U4107 ( .I0(n3996), .I1(n3994), .I2(n3995), .I3(n3993), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ) );
  MUX4D0 U4108 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .S0(n4089), 
        .S1(n4086), .Z(n3995) );
  MUX4D0 U4109 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ), .S0(n4090), 
        .S1(n4085), .Z(n3994) );
  MUX4D0 U4110 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .S0(n4089), 
        .S1(n4086), .Z(n3996) );
  MUX4D0 U4111 ( .I0(n4000), .I1(n3998), .I2(n3999), .I3(n3997), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ) );
  MUX4D0 U4112 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .S0(n4087), 
        .S1(n4086), .Z(n3999) );
  MUX4D0 U4113 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ), .S0(n4088), 
        .S1(n4085), .Z(n3998) );
  MUX4D0 U4114 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4083), .Z(n4000) );
  MUX4D0 U4115 ( .I0(n4004), .I1(n4002), .I2(n4003), .I3(n4001), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ) );
  MUX4D0 U4116 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4003) );
  MUX4D0 U4117 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ), .S0(n4088), 
        .S1(n4083), .Z(n4002) );
  MUX4D0 U4118 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .S0(n4088), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4004) );
  MUX4D0 U4119 ( .I0(n4008), .I1(n4006), .I2(n4007), .I3(n4005), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ) );
  MUX4D0 U4120 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .S0(n4087), 
        .S1(n4085), .Z(n4007) );
  MUX4D0 U4121 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ), .S0(n4087), 
        .S1(n4084), .Z(n4006) );
  MUX4D0 U4122 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .S0(n4087), 
        .S1(n4084), .Z(n4008) );
  MUX4D0 U4123 ( .I0(n4012), .I1(n4010), .I2(n4011), .I3(n4009), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ) );
  MUX4D0 U4124 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .S0(n4088), 
        .S1(n4083), .Z(n4011) );
  MUX4D0 U4125 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ), .S0(n4091), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4010) );
  MUX4D0 U4126 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .S0(n4087), 
        .S1(n4084), .Z(n4012) );
  MUX4D0 U4127 ( .I0(n4016), .I1(n4014), .I2(n4015), .I3(n4013), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ) );
  MUX4D0 U4128 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .S0(n4087), 
        .S1(n4085), .Z(n4015) );
  MUX4D0 U4129 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4086), .Z(n4014) );
  MUX4D0 U4130 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .S0(n4091), 
        .S1(n4086), .Z(n4016) );
  MUX4D0 U4131 ( .I0(n4020), .I1(n4018), .I2(n4019), .I3(n4017), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ) );
  MUX4D0 U4132 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .S0(n4089), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4019) );
  MUX4D0 U4133 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ), .S0(n4092), 
        .S1(n4083), .Z(n4018) );
  MUX4D0 U4134 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .S0(n4092), 
        .S1(n4083), .Z(n4020) );
  MUX4D0 U4135 ( .I0(n4024), .I1(n4022), .I2(n4023), .I3(n4021), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ) );
  MUX4D0 U4136 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .S0(n4087), 
        .S1(n4083), .Z(n4023) );
  MUX4D0 U4137 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4022) );
  MUX4D0 U4138 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .S0(n4088), 
        .S1(n4085), .Z(n4024) );
  MUX4D0 U4139 ( .I0(n4028), .I1(n4026), .I2(n4027), .I3(n4025), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ) );
  MUX4D0 U4140 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4084), .Z(n4027) );
  MUX4D0 U4141 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ), .S0(n4088), 
        .S1(n4084), .Z(n4026) );
  MUX4D0 U4142 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .S0(n4087), 
        .S1(n4085), .Z(n4028) );
  MUX4D0 U4143 ( .I0(n4032), .I1(n4030), .I2(n4031), .I3(n4029), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ) );
  MUX4D0 U4144 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4086), .Z(n4031) );
  MUX4D0 U4145 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ), .S0(n4088), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4030) );
  MUX4D0 U4146 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .S0(n4087), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4032) );
  MUX4D0 U4147 ( .I0(n4036), .I1(n4034), .I2(n4035), .I3(n4033), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ) );
  MUX4D0 U4148 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .S0(n4087), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4035) );
  MUX4D0 U4149 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ), .S0(n4088), 
        .S1(n4083), .Z(n4034) );
  MUX4D0 U4150 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4084), .Z(n4036) );
  MUX4D0 U4151 ( .I0(n4040), .I1(n4038), .I2(n4039), .I3(n4037), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ) );
  MUX4D0 U4152 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .S0(n4088), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4039) );
  MUX4D0 U4153 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ), .S0(n4088), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4038) );
  MUX4D0 U4154 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .S0(n4087), 
        .S1(n4084), .Z(n4040) );
  MUX4D0 U4155 ( .I0(n4044), .I1(n4042), .I2(n4043), .I3(n4041), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ) );
  MUX4D0 U4156 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .S0(n4090), 
        .S1(n4083), .Z(n4043) );
  MUX4D0 U4157 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ), .S0(n4087), 
        .S1(n4086), .Z(n4042) );
  MUX4D0 U4158 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n4083), .Z(n4044) );
  MUX4D0 U4159 ( .I0(n4048), .I1(n4046), .I2(n4047), .I3(n4045), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ) );
  MUX4D0 U4160 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .S0(n4090), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4047) );
  MUX4D0 U4161 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ), .S0(n4090), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4046) );
  MUX4D0 U4162 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .S0(n4090), 
        .S1(n4083), .Z(n4048) );
  MUX4D0 U4163 ( .I0(n4052), .I1(n4050), .I2(n4051), .I3(n4049), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ) );
  MUX4D0 U4164 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .S0(n4090), 
        .S1(n4084), .Z(n4051) );
  MUX4D0 U4165 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ), .S0(n4090), 
        .S1(n4083), .Z(n4050) );
  MUX4D0 U4166 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .S0(n4090), 
        .S1(n4086), .Z(n4052) );
  MUX4D0 U4167 ( .I0(n4056), .I1(n4054), .I2(n4055), .I3(n4053), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ) );
  MUX4D0 U4168 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .S0(n4090), 
        .S1(n4083), .Z(n4055) );
  MUX4D0 U4169 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ), .S0(n4090), 
        .S1(n4085), .Z(n4054) );
  MUX4D0 U4170 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .S0(n4090), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n4056) );
  MUX4D0 U4171 ( .I0(n4060), .I1(n4058), .I2(n4059), .I3(n4057), .S0(n4081), 
        .S1(n4082), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ) );
  MUX4D0 U4172 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .S0(n4091), 
        .S1(n4086), .Z(n4059) );
  MUX4D0 U4173 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ), .S0(n4091), 
        .S1(n4086), .Z(n4058) );
  MUX4D0 U4174 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .S0(n4091), 
        .S1(n4086), .Z(n4060) );
  MUX4D0 U4175 ( .I0(n4064), .I1(n4062), .I2(n4063), .I3(n4061), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ) );
  MUX4D0 U4176 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .S0(n4091), 
        .S1(n4086), .Z(n4063) );
  MUX4D0 U4177 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ), .S0(n4091), 
        .S1(n4086), .Z(n4062) );
  MUX4D0 U4178 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .S0(n4091), 
        .S1(n4086), .Z(n4064) );
  MUX4D0 U4179 ( .I0(n4068), .I1(n4066), .I2(n4067), .I3(n4065), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ) );
  MUX4D0 U4180 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .S0(n4091), 
        .S1(n4086), .Z(n4067) );
  MUX4D0 U4181 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ), .S0(n4091), 
        .S1(n4086), .Z(n4066) );
  MUX4D0 U4182 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .S0(n4091), 
        .S1(n4086), .Z(n4068) );
  MUX4D0 U4183 ( .I0(n4072), .I1(n4070), .I2(n4071), .I3(n4069), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ) );
  MUX4D0 U4184 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .S0(n4092), 
        .S1(n4086), .Z(n4071) );
  MUX4D0 U4185 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ), .S0(n4092), 
        .S1(n4085), .Z(n4070) );
  MUX4D0 U4186 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .S0(n4092), 
        .S1(n4084), .Z(n4072) );
  MUX4D0 U4187 ( .I0(n4076), .I1(n4074), .I2(n4075), .I3(n4073), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n4082), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ) );
  MUX4D0 U4188 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .S0(n4092), 
        .S1(n4084), .Z(n4075) );
  MUX4D0 U4189 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ), .S0(n4092), 
        .S1(n4084), .Z(n4074) );
  MUX4D0 U4190 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .S0(n4092), 
        .S1(n4083), .Z(n4076) );
  MUX4D0 U4191 ( .I0(n4080), .I1(n4078), .I2(n4079), .I3(n4077), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ) );
  MUX4D0 U4192 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .S0(n4092), 
        .S1(n4084), .Z(n4079) );
  MUX4D0 U4193 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ), .S0(n4092), 
        .S1(n4084), .Z(n4078) );
  MUX4D0 U4194 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .S0(n4092), 
        .S1(n4084), .Z(n4080) );
  INVD1 U4195 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n4499) );
  INVD1 U4196 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n4480) );
  INVD1 U4197 ( .I(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), .ZN(n4603) );
  INVD1 U4198 ( .I(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), .ZN(n4599) );
  INR2D1 U4199 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), .B1(n4604), .ZN(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ) );
  INR2D1 U4200 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), .B1(n4600), .ZN(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N26 ) );
  TIEH U4201 ( .Z(n5124) );
  TIEL U4202 ( .ZN(n1037) );
  MUX2ND0 U4203 ( .I0(n4093), .I1(n4094), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ) );
  MUX2ND0 U4204 ( .I0(n4095), .I1(n4096), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ) );
  MUX2ND0 U4205 ( .I0(n4094), .I1(n4093), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ) );
  MUX2ND0 U4206 ( .I0(n4096), .I1(n4095), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ) );
  MUX2ND0 U4207 ( .I0(n3584), .I1(n3588), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4094) );
  MUX2ND0 U4208 ( .I0(n3583), .I1(n3589), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4093) );
  MUX2ND0 U4209 ( .I0(n3588), .I1(n3583), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4096) );
  MUX2ND0 U4210 ( .I0(n3589), .I1(n3584), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4095) );
  MUX2ND0 U4211 ( .I0(n4097), .I1(n4098), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N29 ) );
  MUX2ND0 U4212 ( .I0(n4099), .I1(n4100), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N27 ) );
  MUX2ND0 U4213 ( .I0(n4098), .I1(n4097), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N25 ) );
  MUX2ND0 U4214 ( .I0(n4100), .I1(n4099), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N23 ) );
  MUX2ND0 U4215 ( .I0(n3586), .I1(n3590), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4098) );
  MUX2ND0 U4216 ( .I0(n3585), .I1(n3591), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4097) );
  MUX2ND0 U4217 ( .I0(n3590), .I1(n3585), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4100) );
  MUX2ND0 U4218 ( .I0(n3591), .I1(n3586), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n4099) );
  MUX3ND0 U4219 ( .I0(n4101), .I1(n4102), .I2(n4103), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ) );
  MUX3ND0 U4220 ( .I0(n4104), .I1(n4105), .I2(n4106), .S0(n4199), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ) );
  MUX3ND0 U4221 ( .I0(n4107), .I1(n4108), .I2(n4109), .S0(n4198), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ) );
  MUX3ND0 U4222 ( .I0(n4110), .I1(n4111), .I2(n4112), .S0(n4198), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ) );
  MUX3ND0 U4223 ( .I0(n4113), .I1(n4114), .I2(n4115), .S0(n4199), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ) );
  MUX3ND0 U4224 ( .I0(n4116), .I1(n4117), .I2(n4118), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ) );
  MUX3ND0 U4225 ( .I0(n4119), .I1(n4120), .I2(n4121), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ) );
  MUX3ND0 U4226 ( .I0(n4122), .I1(n4123), .I2(n4124), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ) );
  MUX3ND0 U4227 ( .I0(n4125), .I1(n4126), .I2(n4127), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ) );
  MUX3ND0 U4228 ( .I0(n4128), .I1(n4129), .I2(n4130), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n4197), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ) );
  MUX3ND0 U4229 ( .I0(n4131), .I1(n4132), .I2(n4133), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ) );
  MUX3ND0 U4230 ( .I0(n4134), .I1(n4135), .I2(n4136), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ) );
  MUX3ND0 U4231 ( .I0(n4137), .I1(n4138), .I2(n4139), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ) );
  MUX3ND0 U4232 ( .I0(n4140), .I1(n4141), .I2(n4142), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n4197), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ) );
  MUX3ND0 U4233 ( .I0(n4143), .I1(n4144), .I2(n4145), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ) );
  MUX3ND0 U4234 ( .I0(n4146), .I1(n4147), .I2(n4148), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ) );
  MUX3ND0 U4235 ( .I0(n4149), .I1(n4150), .I2(n4151), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n4197), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ) );
  MUX3ND0 U4236 ( .I0(n4152), .I1(n4153), .I2(n4154), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ) );
  MUX3ND0 U4237 ( .I0(n4155), .I1(n4156), .I2(n4157), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ) );
  MUX3ND0 U4238 ( .I0(n4158), .I1(n4159), .I2(n4160), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ) );
  MUX3ND0 U4239 ( .I0(n4161), .I1(n4162), .I2(n4163), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ) );
  MUX3ND0 U4240 ( .I0(n4164), .I1(n4165), .I2(n4166), .S0(n4199), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ) );
  MUX3ND0 U4241 ( .I0(n4167), .I1(n4168), .I2(n4169), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n4197), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ) );
  MUX3ND0 U4242 ( .I0(n4170), .I1(n4171), .I2(n4172), .S0(n4198), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ) );
  MUX3ND0 U4243 ( .I0(n4173), .I1(n4174), .I2(n4175), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ) );
  MUX3ND0 U4244 ( .I0(n4176), .I1(n4177), .I2(n4178), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ) );
  MUX3ND0 U4245 ( .I0(n4179), .I1(n4180), .I2(n4181), .S0(n4199), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ) );
  MUX3ND0 U4246 ( .I0(n4182), .I1(n4183), .I2(n4184), .S0(n4199), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ) );
  MUX3ND0 U4247 ( .I0(n4185), .I1(n4186), .I2(n4187), .S0(n4198), .S1(n4197), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ) );
  MUX3ND0 U4248 ( .I0(n4188), .I1(n4189), .I2(n4190), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ) );
  MUX3ND0 U4249 ( .I0(n4191), .I1(n4192), .I2(n4193), .S0(n4199), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ) );
  MUX3ND0 U4250 ( .I0(n4194), .I1(n4195), .I2(n4196), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n4197), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ) );
  MUX2ND0 U4251 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .S(n4200), 
        .ZN(n4102) );
  MUX2ND0 U4252 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .S(n4200), 
        .ZN(n4101) );
  MUX2ND0 U4253 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .S(n4200), 
        .ZN(n4105) );
  MUX2ND0 U4254 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .S(n4200), 
        .ZN(n4104) );
  MUX2ND0 U4255 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .S(n4200), 
        .ZN(n4108) );
  MUX2ND0 U4256 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .S(n4200), 
        .ZN(n4107) );
  MUX2ND0 U4257 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .S(n4200), 
        .ZN(n4111) );
  MUX2ND0 U4258 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .S(n4200), 
        .ZN(n4110) );
  MUX2ND0 U4259 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .S(n4200), 
        .ZN(n4114) );
  MUX2ND0 U4260 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .S(n4200), 
        .ZN(n4113) );
  MUX2ND0 U4261 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .S(n4200), 
        .ZN(n4117) );
  MUX2ND0 U4262 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .S(n4200), 
        .ZN(n4116) );
  MUX2ND0 U4263 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .S(n4201), 
        .ZN(n4120) );
  MUX2ND0 U4264 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .S(n4201), 
        .ZN(n4119) );
  MUX2ND0 U4265 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .S(n4201), 
        .ZN(n4123) );
  MUX2ND0 U4266 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .S(n4201), 
        .ZN(n4122) );
  MUX2ND0 U4267 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .S(n4201), 
        .ZN(n4126) );
  MUX2ND0 U4268 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .S(n4201), 
        .ZN(n4125) );
  MUX2ND0 U4269 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .S(n4201), 
        .ZN(n4129) );
  MUX2ND0 U4270 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .S(n4201), 
        .ZN(n4128) );
  MUX2ND0 U4271 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .S(n4201), 
        .ZN(n4132) );
  MUX2ND0 U4272 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .S(n4201), 
        .ZN(n4131) );
  MUX2ND0 U4273 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .S(n4201), 
        .ZN(n4135) );
  MUX2ND0 U4274 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .S(n4201), 
        .ZN(n4134) );
  MUX2ND0 U4275 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .S(n4201), 
        .ZN(n4138) );
  MUX2ND0 U4276 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .S(n4201), 
        .ZN(n4137) );
  MUX2ND0 U4277 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .S(n4202), 
        .ZN(n4141) );
  MUX2ND0 U4278 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .S(n4202), 
        .ZN(n4140) );
  MUX2ND0 U4279 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .S(n4202), 
        .ZN(n4144) );
  MUX2ND0 U4280 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .S(n4202), 
        .ZN(n4143) );
  MUX2ND0 U4281 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .S(n4202), 
        .ZN(n4147) );
  MUX2ND0 U4282 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .S(n4202), 
        .ZN(n4146) );
  MUX2ND0 U4283 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .S(n4202), 
        .ZN(n4150) );
  MUX2ND0 U4284 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .S(n4202), 
        .ZN(n4149) );
  MUX2ND0 U4285 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .S(n4202), 
        .ZN(n4153) );
  MUX2ND0 U4286 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .S(n4202), 
        .ZN(n4152) );
  MUX2ND0 U4287 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .S(n4202), 
        .ZN(n4156) );
  MUX2ND0 U4288 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .S(n4201), 
        .ZN(n4155) );
  MUX2ND0 U4289 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .S(n4202), 
        .ZN(n4159) );
  MUX2ND0 U4290 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .S(n4202), 
        .ZN(n4158) );
  MUX2ND0 U4291 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .S(n4202), 
        .ZN(n4162) );
  MUX2ND0 U4292 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .S(n4202), 
        .ZN(n4161) );
  MUX2ND0 U4293 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .S(n4203), 
        .ZN(n4165) );
  MUX2ND0 U4294 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n4164) );
  MUX2ND0 U4295 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .S(n4200), 
        .ZN(n4168) );
  MUX2ND0 U4296 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .S(n4203), 
        .ZN(n4167) );
  MUX2ND0 U4297 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .S(n4202), 
        .ZN(n4171) );
  MUX2ND0 U4298 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n4170) );
  MUX2ND0 U4299 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .S(n4202), 
        .ZN(n4174) );
  MUX2ND0 U4300 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .S(n4201), 
        .ZN(n4173) );
  MUX2ND0 U4301 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .S(n4202), 
        .ZN(n4177) );
  MUX2ND0 U4302 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .S(n4202), 
        .ZN(n4176) );
  MUX2ND0 U4303 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .S(n4201), 
        .ZN(n4180) );
  MUX2ND0 U4304 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .S(n4202), 
        .ZN(n4179) );
  MUX2ND0 U4305 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .S(n4202), 
        .ZN(n4183) );
  MUX2ND0 U4306 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .S(n4201), 
        .ZN(n4182) );
  MUX2ND0 U4307 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .S(n4201), 
        .ZN(n4186) );
  MUX2ND0 U4308 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .S(n4201), 
        .ZN(n4185) );
  MUX2ND0 U4309 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .S(n4201), 
        .ZN(n4189) );
  MUX2ND0 U4310 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .S(n4200), 
        .ZN(n4188) );
  MUX2ND0 U4311 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .S(n4200), 
        .ZN(n4192) );
  MUX2ND0 U4312 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .S(n4200), 
        .ZN(n4191) );
  MUX2ND0 U4313 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .S(n4200), 
        .ZN(n4195) );
  MUX2ND0 U4314 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .S(n4200), 
        .ZN(n4194) );
  MUX3ND0 U4315 ( .I0(n4204), .I1(n4205), .I2(n4206), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ) );
  MUX3ND0 U4316 ( .I0(n4207), .I1(n4208), .I2(n4209), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ) );
  MUX3ND0 U4317 ( .I0(n4210), .I1(n4211), .I2(n4212), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ) );
  MUX3ND0 U4318 ( .I0(n4213), .I1(n4214), .I2(n4215), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ) );
  MUX3ND0 U4319 ( .I0(n4216), .I1(n4217), .I2(n4218), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ) );
  MUX3ND0 U4320 ( .I0(n4219), .I1(n4220), .I2(n4221), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ) );
  MUX3ND0 U4321 ( .I0(n4222), .I1(n4223), .I2(n4224), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ) );
  MUX3ND0 U4322 ( .I0(n4225), .I1(n4226), .I2(n4227), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ) );
  MUX3ND0 U4323 ( .I0(n4228), .I1(n4229), .I2(n4230), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ) );
  MUX3ND0 U4324 ( .I0(n4231), .I1(n4232), .I2(n4233), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ) );
  MUX3ND0 U4325 ( .I0(n4234), .I1(n4235), .I2(n4236), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ) );
  MUX3ND0 U4326 ( .I0(n4237), .I1(n4238), .I2(n4239), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ) );
  MUX3ND0 U4327 ( .I0(n4240), .I1(n4241), .I2(n4242), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ) );
  MUX3ND0 U4328 ( .I0(n4243), .I1(n4244), .I2(n4245), .S0(n4302), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ) );
  MUX3ND0 U4329 ( .I0(n4246), .I1(n4247), .I2(n4248), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ) );
  MUX3ND0 U4330 ( .I0(n4249), .I1(n4250), .I2(n4251), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ) );
  MUX3ND0 U4331 ( .I0(n4252), .I1(n4253), .I2(n4254), .S0(n4302), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ) );
  MUX3ND0 U4332 ( .I0(n4255), .I1(n4256), .I2(n4257), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n4300), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ) );
  MUX3ND0 U4333 ( .I0(n4258), .I1(n4259), .I2(n4260), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ) );
  MUX3ND0 U4334 ( .I0(n4261), .I1(n4262), .I2(n4263), .S0(n4302), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ) );
  MUX3ND0 U4335 ( .I0(n4264), .I1(n4265), .I2(n4266), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n4300), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ) );
  MUX3ND0 U4336 ( .I0(n4267), .I1(n4268), .I2(n4269), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ) );
  MUX3ND0 U4337 ( .I0(n4270), .I1(n4271), .I2(n4272), .S0(n4302), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ) );
  MUX3ND0 U4338 ( .I0(n4273), .I1(n4274), .I2(n4275), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ) );
  MUX3ND0 U4339 ( .I0(n4276), .I1(n4277), .I2(n4278), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ) );
  MUX3ND0 U4340 ( .I0(n4279), .I1(n4280), .I2(n4281), .S0(n4302), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ) );
  MUX3ND0 U4341 ( .I0(n4282), .I1(n4283), .I2(n4284), .S0(n4301), .S1(n4300), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ) );
  MUX3ND0 U4342 ( .I0(n4285), .I1(n4286), .I2(n4287), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ) );
  MUX3ND0 U4343 ( .I0(n4288), .I1(n4289), .I2(n4290), .S0(n4302), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ) );
  MUX3ND0 U4344 ( .I0(n4291), .I1(n4292), .I2(n4293), .S0(n4302), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ) );
  MUX3ND0 U4345 ( .I0(n4294), .I1(n4295), .I2(n4296), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ) );
  MUX3ND0 U4346 ( .I0(n4297), .I1(n4298), .I2(n4299), .S0(n4301), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ) );
  MUX2ND0 U4347 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .S(n4303), 
        .ZN(n4205) );
  MUX2ND0 U4348 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .S(n4303), 
        .ZN(n4204) );
  MUX2ND0 U4349 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .S(n4303), 
        .ZN(n4208) );
  MUX2ND0 U4350 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .S(n4303), 
        .ZN(n4207) );
  MUX2ND0 U4351 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .S(n4303), 
        .ZN(n4211) );
  MUX2ND0 U4352 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .S(n4303), 
        .ZN(n4210) );
  MUX2ND0 U4353 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .S(n4303), 
        .ZN(n4214) );
  MUX2ND0 U4354 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .S(n4303), 
        .ZN(n4213) );
  MUX2ND0 U4355 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .S(n4303), 
        .ZN(n4217) );
  MUX2ND0 U4356 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .S(n4303), 
        .ZN(n4216) );
  MUX2ND0 U4357 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .S(n4303), 
        .ZN(n4220) );
  MUX2ND0 U4358 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .S(n4303), 
        .ZN(n4219) );
  MUX2ND0 U4359 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .S(n4304), 
        .ZN(n4223) );
  MUX2ND0 U4360 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .S(n4304), 
        .ZN(n4222) );
  MUX2ND0 U4361 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .S(n4304), 
        .ZN(n4226) );
  MUX2ND0 U4362 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .S(n4304), 
        .ZN(n4225) );
  MUX2ND0 U4363 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .S(n4304), 
        .ZN(n4229) );
  MUX2ND0 U4364 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .S(n4304), 
        .ZN(n4228) );
  MUX2ND0 U4365 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .S(n4304), 
        .ZN(n4232) );
  MUX2ND0 U4366 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .S(n4304), 
        .ZN(n4231) );
  MUX2ND0 U4367 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .S(n4304), 
        .ZN(n4235) );
  MUX2ND0 U4368 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .S(n4304), 
        .ZN(n4234) );
  MUX2ND0 U4369 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .S(n4304), 
        .ZN(n4238) );
  MUX2ND0 U4370 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .S(n4304), 
        .ZN(n4237) );
  MUX2ND0 U4371 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .S(n4304), 
        .ZN(n4241) );
  MUX2ND0 U4372 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .S(n4304), 
        .ZN(n4240) );
  MUX2ND0 U4373 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .S(n4305), 
        .ZN(n4244) );
  MUX2ND0 U4374 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .S(n4305), 
        .ZN(n4243) );
  MUX2ND0 U4375 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .S(n4305), 
        .ZN(n4247) );
  MUX2ND0 U4376 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .S(n4305), 
        .ZN(n4246) );
  MUX2ND0 U4377 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .S(n4305), 
        .ZN(n4250) );
  MUX2ND0 U4378 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .S(n4305), 
        .ZN(n4249) );
  MUX2ND0 U4379 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .S(n4305), 
        .ZN(n4253) );
  MUX2ND0 U4380 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .S(n4305), 
        .ZN(n4252) );
  MUX2ND0 U4381 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .S(n4305), 
        .ZN(n4256) );
  MUX2ND0 U4382 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .S(n4305), 
        .ZN(n4255) );
  MUX2ND0 U4383 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .S(n4305), 
        .ZN(n4259) );
  MUX2ND0 U4384 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .S(n4304), 
        .ZN(n4258) );
  MUX2ND0 U4385 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .S(n4305), 
        .ZN(n4262) );
  MUX2ND0 U4386 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .S(n4305), 
        .ZN(n4261) );
  MUX2ND0 U4387 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n4265) );
  MUX2ND0 U4388 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .S(n4305), 
        .ZN(n4264) );
  MUX2ND0 U4389 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .S(n4306), 
        .ZN(n4268) );
  MUX2ND0 U4390 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n4267) );
  MUX2ND0 U4391 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .S(n4305), 
        .ZN(n4271) );
  MUX2ND0 U4392 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .S(n4303), 
        .ZN(n4270) );
  MUX2ND0 U4393 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .S(n4305), 
        .ZN(n4274) );
  MUX2ND0 U4394 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .S(n4304), 
        .ZN(n4273) );
  MUX2ND0 U4395 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .S(n4305), 
        .ZN(n4277) );
  MUX2ND0 U4396 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .S(n4306), 
        .ZN(n4276) );
  MUX2ND0 U4397 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .S(n4305), 
        .ZN(n4280) );
  MUX2ND0 U4398 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .S(n4305), 
        .ZN(n4279) );
  MUX2ND0 U4399 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .S(n4304), 
        .ZN(n4283) );
  MUX2ND0 U4400 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .S(n4305), 
        .ZN(n4282) );
  MUX2ND0 U4401 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .S(n4305), 
        .ZN(n4286) );
  MUX2ND0 U4402 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .S(n4304), 
        .ZN(n4285) );
  MUX2ND0 U4403 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .S(n4304), 
        .ZN(n4289) );
  MUX2ND0 U4404 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .S(n4304), 
        .ZN(n4288) );
  MUX2ND0 U4405 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .S(n4304), 
        .ZN(n4292) );
  MUX2ND0 U4406 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .S(n4303), 
        .ZN(n4291) );
  MUX2ND0 U4407 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .S(n4303), 
        .ZN(n4295) );
  MUX2ND0 U4408 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .S(n4303), 
        .ZN(n4294) );
  MUX2ND0 U4409 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .S(n4303), 
        .ZN(n4298) );
  MUX2ND0 U4410 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .S(n4303), 
        .ZN(n4297) );
  CKND0 U4411 ( .CLK(n5188), .CN(n4307) );
  CKND0 U4412 ( .CLK(n5187), .CN(n4308) );
  CKND0 U4413 ( .CLK(n5186), .CN(n4309) );
  CKND0 U4414 ( .CLK(n5185), .CN(n4310) );
  CKND0 U4415 ( .CLK(n5184), .CN(n4311) );
  CKND0 U4416 ( .CLK(n5183), .CN(n4312) );
  CKND0 U4417 ( .CLK(n5182), .CN(n4313) );
  CKND0 U4418 ( .CLK(n5181), .CN(n4314) );
  CKND0 U4419 ( .CLK(n5180), .CN(n4315) );
  CKND0 U4420 ( .CLK(n5179), .CN(n4316) );
  CKND0 U4421 ( .CLK(n5178), .CN(n4317) );
  CKND0 U4422 ( .CLK(n5177), .CN(n4318) );
  CKND0 U4423 ( .CLK(n5176), .CN(n4319) );
  CKND0 U4424 ( .CLK(n5175), .CN(n4320) );
  CKND0 U4425 ( .CLK(n5174), .CN(n4321) );
  CKND0 U4426 ( .CLK(n5173), .CN(n4322) );
  CKND0 U4427 ( .CLK(n5172), .CN(n4323) );
  CKND0 U4428 ( .CLK(n5171), .CN(n4324) );
  CKND0 U4429 ( .CLK(n5170), .CN(n4325) );
  CKND0 U4430 ( .CLK(n5169), .CN(n4326) );
  CKND0 U4431 ( .CLK(n5168), .CN(n4327) );
  CKND0 U4432 ( .CLK(n5167), .CN(n4328) );
  CKND0 U4433 ( .CLK(n5166), .CN(n4329) );
  CKND0 U4434 ( .CLK(n5165), .CN(n4330) );
  CKND0 U4435 ( .CLK(n5164), .CN(n4331) );
  CKND0 U4436 ( .CLK(n5163), .CN(n4332) );
  CKND0 U4437 ( .CLK(n5162), .CN(n4333) );
  CKND0 U4438 ( .CLK(n5161), .CN(n4334) );
  CKND0 U4439 ( .CLK(n5160), .CN(n4335) );
  CKND0 U4440 ( .CLK(n5159), .CN(n4336) );
  CKND0 U4441 ( .CLK(n5158), .CN(n4337) );
  CKND0 U4442 ( .CLK(n5157), .CN(n4338) );
  CKND0 U4443 ( .CLK(n5156), .CN(n4339) );
  CKND0 U4444 ( .CLK(n5155), .CN(n4340) );
  CKND0 U4445 ( .CLK(n5154), .CN(n4341) );
  CKND0 U4446 ( .CLK(n5153), .CN(n4342) );
  CKND0 U4447 ( .CLK(n5152), .CN(n4343) );
  CKND0 U4448 ( .CLK(n5151), .CN(n4344) );
  CKND0 U4449 ( .CLK(n5150), .CN(n4345) );
  CKND0 U4450 ( .CLK(n5149), .CN(n4346) );
  CKND0 U4451 ( .CLK(n5148), .CN(n4347) );
  CKND0 U4452 ( .CLK(n5147), .CN(n4348) );
  CKND0 U4453 ( .CLK(n5146), .CN(n4349) );
  CKND0 U4454 ( .CLK(n5145), .CN(n4350) );
  CKND0 U4455 ( .CLK(n5144), .CN(n4351) );
  CKND0 U4456 ( .CLK(n5143), .CN(n4352) );
  CKND0 U4457 ( .CLK(n5142), .CN(n4353) );
  CKND0 U4458 ( .CLK(n5141), .CN(n4354) );
  CKND0 U4459 ( .CLK(n5140), .CN(n4355) );
  CKND0 U4460 ( .CLK(n5139), .CN(n4356) );
  CKND0 U4461 ( .CLK(n5138), .CN(n4357) );
  CKND0 U4462 ( .CLK(n5137), .CN(n4358) );
  CKND0 U4463 ( .CLK(n5136), .CN(n4359) );
  CKND0 U4464 ( .CLK(n5135), .CN(n4360) );
  CKND0 U4465 ( .CLK(n5134), .CN(n4361) );
  CKND0 U4466 ( .CLK(n5133), .CN(n4362) );
  CKND0 U4467 ( .CLK(n5132), .CN(n4363) );
  CKND0 U4468 ( .CLK(n5131), .CN(n4364) );
  CKND0 U4469 ( .CLK(n5130), .CN(n4365) );
  CKND0 U4470 ( .CLK(n5129), .CN(n4366) );
  CKND0 U4471 ( .CLK(n5128), .CN(n4367) );
  CKND0 U4472 ( .CLK(n5127), .CN(n4368) );
  CKND0 U4473 ( .CLK(n5126), .CN(n4369) );
  CKND0 U4474 ( .CLK(n5125), .CN(n4370) );
  OR2D1 U4475 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .Z(n4600) );
  MUX2ND0 U4476 ( .I0(n4601), .I1(n4600), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N28 ) );
  OR2D1 U4477 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .Z(n4604) );
  MUX2ND0 U4478 ( .I0(n4605), .I1(n4604), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ) );
  OAI31D0 U4479 ( .A1(n4616), .A2(Reset), .A3(n4617), .B(n4618), .ZN(n3528) );
  OAI21D0 U4480 ( .A1(n4619), .A2(Reset), .B(\SerDes_U2/Tx_F_Full ), .ZN(n4618) );
  AOI21D0 U4481 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .B(n4620), .ZN(
        n4619) );
  NR3D0 U4482 ( .A1(\SerDes_U2/Tx_F_Empty ), .A2(n4521), .A3(n4621), .ZN(n4617) );
  MUX2ND0 U4483 ( .I0(n4622), .I1(n1030), .S(n4623), .ZN(n3526) );
  AOI211D0 U4484 ( .A1(n4624), .A2(n4625), .B(n4626), .C(n4620), .ZN(n4622) );
  AOI21D0 U4485 ( .A1(n4627), .A2(n4628), .B(n4629), .ZN(n4626) );
  MUX2D0 U4486 ( .I0(n4630), .I1(n4628), .S(n1033), .Z(n4624) );
  ND4D0 U4487 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n4628) );
  AOI211D0 U4488 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .A2(n4524), .B(n4635), .C(n4636), .ZN(n4634) );
  XNR2D0 U4489 ( .A1(n4637), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .ZN(n4636) );
  XNR2D0 U4490 ( .A1(n4638), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), 
        .ZN(n4635) );
  OAI33D0 U4491 ( .A1(n4639), .A2(n4640), .A3(n4641), .B1(n4642), .B2(n4643), 
        .B3(n4644), .ZN(n3523) );
  XNR2D0 U4492 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .A2(n1028), 
        .ZN(n4640) );
  ND3D0 U4493 ( .A1(n4645), .A2(n4646), .A3(n4647), .ZN(n4639) );
  XNR2D0 U4494 ( .A1(n1027), .A2(n4526), .ZN(n4647) );
  XNR2D0 U4495 ( .A1(n1026), .A2(n4525), .ZN(n4646) );
  XNR2D0 U4496 ( .A1(n1025), .A2(n4524), .ZN(n4645) );
  MUX2ND0 U4497 ( .I0(n4648), .I1(n1024), .S(n4623), .ZN(n3485) );
  AOI32D0 U4498 ( .A1(n4625), .A2(n4649), .A3(n4650), .B1(n4651), .B2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n4648) );
  OAI21D0 U4499 ( .A1(n1031), .A2(n4652), .B(n1032), .ZN(n4651) );
  NR4D0 U4500 ( .A1(n4650), .A2(n4653), .A3(n4654), .A4(n4655), .ZN(n4652) );
  XNR2D0 U4501 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n4656), 
        .ZN(n4655) );
  XNR2D0 U4502 ( .A1(n4657), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), 
        .ZN(n4654) );
  XNR2D0 U4503 ( .A1(n4658), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n4653) );
  OAI31D0 U4504 ( .A1(n4659), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), 
        .A3(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .B(n4660), .ZN(n4649) );
  MUX2ND0 U4505 ( .I0(n4661), .I1(n4662), .S(n4526), .ZN(n4660) );
  OAI32D0 U4506 ( .A1(n4663), .A2(n4527), .A3(n4631), .B1(n4632), .B2(n4664), 
        .ZN(n4662) );
  OAI32D0 U4507 ( .A1(n4663), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .A3(n4632), .B1(n4631), .B2(n4664), .ZN(n4661) );
  CKND2D0 U4508 ( .A1(n4665), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .ZN(n4664) );
  XNR2D0 U4509 ( .A1(n4637), .A2(n4527), .ZN(n4665) );
  MUX2ND0 U4510 ( .I0(n4666), .I1(n4667), .S(n4526), .ZN(n4659) );
  NR2D0 U4511 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .A2(n4631), 
        .ZN(n4667) );
  NR2D0 U4512 ( .A1(n4527), .A2(n4632), .ZN(n4666) );
  OAI33D0 U4513 ( .A1(n4668), .A2(n4669), .A3(n4670), .B1(n4671), .B2(n4620), 
        .B3(n4644), .ZN(n3482) );
  XNR2D0 U4514 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .A2(n1022), 
        .ZN(n4669) );
  ND3D0 U4515 ( .A1(n4672), .A2(n4673), .A3(n4674), .ZN(n4668) );
  XNR2D0 U4516 ( .A1(n1021), .A2(n4638), .ZN(n4674) );
  XNR2D0 U4517 ( .A1(n1020), .A2(n4675), .ZN(n4673) );
  XNR2D0 U4518 ( .A1(n1019), .A2(n4676), .ZN(n4672) );
  MUX2ND0 U4519 ( .I0(n4677), .I1(n1018), .S(n4623), .ZN(n3479) );
  OA211D0 U4520 ( .A1(n1033), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .B(n4678), .C(n4679), .Z(n4623) );
  AOI22D0 U4521 ( .A1(n4680), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .B1(n4620), .B2(
        n4681), .ZN(n4679) );
  AO31D0 U4522 ( .A1(n4371), .A2(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), 
        .A3(InParValidB), .B(n1033), .Z(n4680) );
  AOI21D0 U4523 ( .A1(n4682), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .B(n4643), .ZN(
        n4677) );
  IOA22D0 U4524 ( .B1(n1031), .B2(n4630), .A1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(n4627), .ZN(
        n4682) );
  ND4D0 U4525 ( .A1(n4683), .A2(n4650), .A3(n4684), .A4(n4658), .ZN(n4627) );
  CKND2D0 U4526 ( .A1(n4632), .A2(n4631), .ZN(n4658) );
  CKND2D0 U4527 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n4525), 
        .ZN(n4631) );
  CKND2D0 U4528 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .A2(n4675), 
        .ZN(n4632) );
  XNR2D0 U4529 ( .A1(n4685), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .ZN(n4684) );
  CKND2D0 U4530 ( .A1(n4686), .A2(n4663), .ZN(n4685) );
  MUX2ND0 U4531 ( .I0(n4675), .I1(n4687), .S(n4637), .ZN(n4686) );
  NR2D0 U4532 ( .A1(n4675), .A2(n4638), .ZN(n4687) );
  CKND0 U4533 ( .CLK(n4688), .CN(n4650) );
  XNR3D0 U4534 ( .A1(n4638), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), 
        .A3(n4526), .ZN(n4683) );
  ND4D0 U4535 ( .A1(n4689), .A2(n4690), .A3(n4691), .A4(n4688), .ZN(n4630) );
  OAI21D0 U4536 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .A2(n4676), 
        .B(n4633), .ZN(n4688) );
  CKND2D0 U4537 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .A2(n4676), 
        .ZN(n4633) );
  XNR2D0 U4538 ( .A1(n4692), .A2(n4525), .ZN(n4691) );
  XNR2D0 U4539 ( .A1(n4527), .A2(n4693), .ZN(n4690) );
  XNR2D0 U4540 ( .A1(n4694), .A2(n4526), .ZN(n4689) );
  MUX2ND0 U4541 ( .I0(n4637), .I1(n1022), .S(n4670), .ZN(n3473) );
  MUX2ND0 U4542 ( .I0(n4675), .I1(n1020), .S(n4670), .ZN(n3471) );
  MUX2ND0 U4543 ( .I0(n4676), .I1(n1019), .S(n4670), .ZN(n3469) );
  MUX2ND0 U4544 ( .I0(n4638), .I1(n1021), .S(n4670), .ZN(n3467) );
  OAI21D0 U4545 ( .A1(n4620), .A2(n4644), .B(n4681), .ZN(n4670) );
  CKND0 U4546 ( .CLK(n4678), .CN(n4644) );
  MUX2ND0 U4547 ( .I0(n4527), .I1(n1028), .S(n4641), .ZN(n2953) );
  MUX2ND0 U4548 ( .I0(n4525), .I1(n1026), .S(n4641), .ZN(n2951) );
  MUX2ND0 U4549 ( .I0(n4524), .I1(n1025), .S(n4641), .ZN(n2949) );
  MUX2ND0 U4550 ( .I0(n4526), .I1(n1027), .S(n4641), .ZN(n2947) );
  ND3D0 U4551 ( .A1(n4371), .A2(InParValidB), .A3(n4695), .ZN(n4641) );
  AOI21D0 U4552 ( .A1(n4678), .A2(n4616), .B(n4521), .ZN(n4695) );
  INR2D0 U4553 ( .A1(n4629), .B1(n4625), .ZN(n4678) );
  ND3D0 U4554 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .A3(n1031), .ZN(
        n4629) );
  OAI31D0 U4555 ( .A1(n4696), .A2(Reset), .A3(n4681), .B(n4697), .ZN(n2945) );
  OAI21D0 U4556 ( .A1(n4698), .A2(Reset), .B(\SerDes_U2/Tx_F_Empty ), .ZN(
        n4697) );
  AOI21D0 U4557 ( .A1(n4625), .A2(n1033), .B(n4620), .ZN(n4698) );
  NR2D0 U4558 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        n1031), .ZN(n4625) );
  NR2D0 U4559 ( .A1(\SerDes_U2/Tx_F_Full ), .A2(n4621), .ZN(n4681) );
  CKND0 U4560 ( .CLK(InParValidB), .CN(n4621) );
  OAI31D0 U4561 ( .A1(n4699), .A2(Reset), .A3(n4700), .B(n4701), .ZN(n2909) );
  OAI21D0 U4562 ( .A1(Reset), .A2(n4702), .B(\SerDes_U1/Tx_F_Empty ), .ZN(
        n4701) );
  OAI22D0 U4563 ( .A1(n1017), .A2(n4703), .B1(n4704), .B2(n4705), .ZN(n2906)
         );
  AO31D0 U4564 ( .A1(n1035), .A2(\SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), 
        .A3(InParValidA), .B(Reset), .Z(n4705) );
  AOI21D0 U4565 ( .A1(n4699), .A2(n4706), .B(Reset), .ZN(n4703) );
  CKND0 U4566 ( .CLK(n4707), .CN(n4706) );
  MUX2ND0 U4567 ( .I0(n4708), .I1(n1016), .S(n4709), .ZN(n2904) );
  NR2D0 U4568 ( .A1(n4710), .A2(n4711), .ZN(n4708) );
  MUX2ND0 U4569 ( .I0(n4712), .I1(n4713), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .ZN(n4711) );
  OAI21D0 U4570 ( .A1(n4714), .A2(n4715), .B(n4716), .ZN(n4713) );
  MUX2ND0 U4571 ( .I0(n4717), .I1(n4718), .S(n4719), .ZN(n4715) );
  NR2D0 U4572 ( .A1(n4720), .A2(n4721), .ZN(n4714) );
  OAI21D0 U4573 ( .A1(n4722), .A2(n4718), .B(n4707), .ZN(n4712) );
  OA211D0 U4574 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n4723), 
        .B(n4721), .C(n4724), .Z(n4718) );
  NR2D0 U4575 ( .A1(n4725), .A2(n4726), .ZN(n4724) );
  CKND0 U4576 ( .CLK(n4727), .CN(n4722) );
  MUX2ND0 U4577 ( .I0(n4728), .I1(n4729), .S(n4730), .ZN(n2901) );
  IND4D0 U4578 ( .A1(n4731), .B1(n4732), .B2(n4733), .B3(n4734), .ZN(n4729) );
  XNR2D0 U4579 ( .A1(n1013), .A2(n4499), .ZN(n4734) );
  XNR2D0 U4580 ( .A1(n1014), .A2(n4500), .ZN(n4733) );
  XNR2D0 U4581 ( .A1(n1012), .A2(n4501), .ZN(n4732) );
  MUX2ND0 U4582 ( .I0(n4735), .I1(n1011), .S(n4709), .ZN(n2896) );
  AOI21D0 U4583 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A2(
        n4736), .B(n4707), .ZN(n4735) );
  OAI31D0 U4584 ( .A1(n4737), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A3(n4726), .B(
        n4738), .ZN(n4736) );
  OAI31D0 U4585 ( .A1(n4739), .A2(n4740), .A3(n4741), .B(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n4738) );
  XNR2D0 U4586 ( .A1(n4742), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .ZN(n4739) );
  MUX2ND0 U4587 ( .I0(n4743), .I1(n4744), .S(n4500), .ZN(n4737) );
  NR2D0 U4588 ( .A1(n4745), .A2(n4746), .ZN(n4744) );
  XNR2D0 U4589 ( .A1(n4723), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), 
        .ZN(n4746) );
  OAI22D0 U4590 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n4747), 
        .B1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .B2(n4721), .ZN(
        n4743) );
  OAI33D0 U4591 ( .A1(n4748), .A2(n4749), .A3(n4750), .B1(n4730), .B2(n1010), 
        .B3(n4710), .ZN(n2893) );
  XNR2D0 U4592 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n1007), 
        .ZN(n4749) );
  OAI211D0 U4593 ( .A1(n4710), .A2(n4751), .B(n4752), .C(n4753), .ZN(n4748) );
  XNR2D0 U4594 ( .A1(n1009), .A2(n4745), .ZN(n4753) );
  XNR2D0 U4595 ( .A1(n1008), .A2(n4754), .ZN(n4752) );
  CKND0 U4596 ( .CLK(n4755), .CN(n4751) );
  MUX2ND0 U4597 ( .I0(n1007), .I1(n4723), .S(n4756), .ZN(n2888) );
  MUX2ND0 U4598 ( .I0(n1008), .I1(n4754), .S(n4756), .ZN(n2886) );
  MUX2ND0 U4599 ( .I0(n1009), .I1(n4745), .S(n4756), .ZN(n2884) );
  AOI21D0 U4600 ( .A1(n4699), .A2(n4755), .B(n4750), .ZN(n4756) );
  MUX2ND0 U4601 ( .I0(n4757), .I1(n1006), .S(n4709), .ZN(n2882) );
  OA211D0 U4602 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A2(
        n4719), .B(n4755), .C(n4758), .Z(n4709) );
  AOI22D0 U4603 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        n4759), .B1(n4700), .B2(n4710), .ZN(n4758) );
  CKND0 U4604 ( .CLK(n4750), .CN(n4700) );
  CKND2D0 U4605 ( .A1(n1017), .A2(InParValidA), .ZN(n4750) );
  CKND2D0 U4606 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .A2(
        n4731), .ZN(n4759) );
  OAI221D0 U4607 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        n4760), .B1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .B2(
        n4727), .C(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(
        n4757) );
  OAI211D0 U4608 ( .A1(n4761), .A2(n4762), .B(n4725), .C(n4740), .ZN(n4727) );
  CKND0 U4609 ( .CLK(n4726), .CN(n4740) );
  MUX2ND0 U4610 ( .I0(n4747), .I1(n4763), .S(n4501), .ZN(n4762) );
  CKND2D0 U4611 ( .A1(n4764), .A2(n4747), .ZN(n4763) );
  NR2D0 U4612 ( .A1(n4745), .A2(n4721), .ZN(n4761) );
  OA211D0 U4613 ( .A1(n4721), .A2(n4720), .B(n4717), .C(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .Z(n4760) );
  AN3D0 U4614 ( .A1(n4741), .A2(n4726), .A3(n4765), .Z(n4717) );
  MUX2ND0 U4615 ( .I0(n4766), .I1(n4767), .S(n4501), .ZN(n4765) );
  OAI21D0 U4616 ( .A1(n4723), .A2(n4499), .B(n4768), .ZN(n4767) );
  NR2D0 U4617 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .A2(n4720), 
        .ZN(n4766) );
  XNR2D0 U4618 ( .A1(n4754), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(n4726) );
  XNR2D0 U4619 ( .A1(n4725), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n4741) );
  XNR2D0 U4620 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n4500), 
        .ZN(n4725) );
  CKND2D0 U4621 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n4723), 
        .ZN(n4721) );
  MUX2ND0 U4622 ( .I0(n1012), .I1(n4501), .S(n4769), .ZN(n2880) );
  MUX2ND0 U4623 ( .I0(n1013), .I1(n4499), .S(n4769), .ZN(n2878) );
  MUX2ND0 U4624 ( .I0(n1014), .I1(n4500), .S(n4769), .ZN(n2876) );
  INR2D0 U4625 ( .A1(n4730), .B1(n4731), .ZN(n4769) );
  ND3D0 U4626 ( .A1(InParValidA), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .A3(n3580), .ZN(n4731) );
  CKND2D0 U4627 ( .A1(n4755), .A2(n4704), .ZN(n4730) );
  MUX2ND0 U4628 ( .I0(n4707), .I1(n4716), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .ZN(n4755) );
  AO222D0 U4629 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ), .A2(
        n4770), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ), .B2(n4771), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .C2(n4772), 
        .Z(n2541) );
  AO222D0 U4630 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ), .A2(
        n4770), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ), .B2(n4771), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .C2(n4772), 
        .Z(n2538) );
  AO222D0 U4631 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ), .A2(
        n4770), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ), .B2(n4771), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .C2(n4772), 
        .Z(n2536) );
  CKND0 U4632 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CN(
        n4772) );
  AN2D0 U4633 ( .A1(n4773), .A2(n4774), .Z(n4771) );
  AN3D0 U4634 ( .A1(n4775), .A2(n4776), .A3(n4777), .Z(n4770) );
  CKXOR2D0 U4635 ( .A1(\SerDes_U1/Tx_SerClk ), .A2(n4778), .Z(n2532) );
  AO222D0 U4636 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ), .A2(
        n4779), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ), .B2(n4780), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .C2(n4781), 
        .Z(n2509) );
  XNR2D0 U4637 ( .A1(n4782), .A2(\SerDes_U1/Des_U1/SerialClk ), .ZN(n2505) );
  MUX2ND0 U4638 ( .I0(n1005), .I1(n1004), .S(n4478), .ZN(n2439) );
  MUX2ND0 U4639 ( .I0(n971), .I1(n970), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2437) );
  MUX2ND0 U4640 ( .I0(n969), .I1(n968), .S(n4478), .ZN(n2435) );
  MUX2ND0 U4641 ( .I0(n967), .I1(n966), .S(n4478), .ZN(n2433) );
  MUX2ND0 U4642 ( .I0(n965), .I1(n964), .S(n4478), .ZN(n2431) );
  MUX2ND0 U4643 ( .I0(n963), .I1(n962), .S(n4478), .ZN(n2429) );
  MUX2ND0 U4644 ( .I0(n961), .I1(n960), .S(n4478), .ZN(n2427) );
  MUX2ND0 U4645 ( .I0(n959), .I1(n958), .S(n4478), .ZN(n2425) );
  MUX2ND0 U4646 ( .I0(n957), .I1(n956), .S(n4478), .ZN(n2423) );
  MUX2ND0 U4647 ( .I0(n955), .I1(n954), .S(n4478), .ZN(n2421) );
  MUX2ND0 U4648 ( .I0(n953), .I1(n952), .S(n4478), .ZN(n2419) );
  MUX2ND0 U4649 ( .I0(n951), .I1(n950), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2417) );
  MUX2ND0 U4650 ( .I0(n949), .I1(n948), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2415) );
  MUX2ND0 U4651 ( .I0(n947), .I1(n946), .S(n4478), .ZN(n2413) );
  MUX2ND0 U4652 ( .I0(n945), .I1(n944), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2411) );
  MUX2ND0 U4653 ( .I0(n943), .I1(n942), .S(n4478), .ZN(n2409) );
  MUX2ND0 U4654 ( .I0(n941), .I1(n940), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2407) );
  MUX2ND0 U4655 ( .I0(n939), .I1(n938), .S(n4478), .ZN(n2405) );
  MUX2ND0 U4656 ( .I0(n937), .I1(n936), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2403) );
  MUX2ND0 U4657 ( .I0(n935), .I1(n934), .S(n4478), .ZN(n2401) );
  MUX2ND0 U4658 ( .I0(n933), .I1(n932), .S(n4478), .ZN(n2399) );
  MUX2ND0 U4659 ( .I0(n931), .I1(n930), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2397) );
  MUX2ND0 U4660 ( .I0(n929), .I1(n928), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2395) );
  MUX2ND0 U4661 ( .I0(n927), .I1(n926), .S(n4478), .ZN(n2393) );
  MUX2ND0 U4662 ( .I0(n925), .I1(n924), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2391) );
  MUX2ND0 U4663 ( .I0(n923), .I1(n922), .S(n4478), .ZN(n2389) );
  MUX2ND0 U4664 ( .I0(n921), .I1(n920), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2387) );
  MUX2ND0 U4665 ( .I0(n919), .I1(n918), .S(n4478), .ZN(n2385) );
  MUX2ND0 U4666 ( .I0(n917), .I1(n916), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n2383) );
  MUX2ND0 U4667 ( .I0(n915), .I1(n914), .S(n4478), .ZN(n2381) );
  MUX2ND0 U4668 ( .I0(n913), .I1(n912), .S(n4478), .ZN(n2379) );
  MUX2ND0 U4669 ( .I0(n911), .I1(n910), .S(n4478), .ZN(n2377) );
  MUX2ND0 U4670 ( .I0(n908), .I1(n911), .S(n4372), .ZN(n2373) );
  MUX2ND0 U4671 ( .I0(n907), .I1(n913), .S(n4372), .ZN(n2371) );
  MUX2ND0 U4672 ( .I0(n906), .I1(n915), .S(n4372), .ZN(n2369) );
  MUX2ND0 U4673 ( .I0(n905), .I1(n917), .S(n4372), .ZN(n2367) );
  MUX2ND0 U4674 ( .I0(n904), .I1(n919), .S(n4372), .ZN(n2365) );
  MUX2ND0 U4675 ( .I0(n903), .I1(n921), .S(n4372), .ZN(n2363) );
  MUX2ND0 U4676 ( .I0(n902), .I1(n923), .S(n4372), .ZN(n2361) );
  MUX2ND0 U4677 ( .I0(n901), .I1(n925), .S(n4372), .ZN(n2359) );
  MUX2ND0 U4678 ( .I0(n900), .I1(n927), .S(n4372), .ZN(n2357) );
  MUX2ND0 U4679 ( .I0(n899), .I1(n929), .S(n4372), .ZN(n2355) );
  MUX2ND0 U4680 ( .I0(n898), .I1(n931), .S(n4372), .ZN(n2353) );
  MUX2ND0 U4681 ( .I0(n897), .I1(n933), .S(n4372), .ZN(n2351) );
  MUX2ND0 U4682 ( .I0(n896), .I1(n935), .S(n4372), .ZN(n2349) );
  MUX2ND0 U4683 ( .I0(n895), .I1(n937), .S(n4372), .ZN(n2347) );
  MUX2ND0 U4684 ( .I0(n894), .I1(n939), .S(n4372), .ZN(n2345) );
  MUX2ND0 U4685 ( .I0(n893), .I1(n941), .S(n4372), .ZN(n2343) );
  MUX2ND0 U4686 ( .I0(n892), .I1(n943), .S(n4372), .ZN(n2341) );
  MUX2ND0 U4687 ( .I0(n891), .I1(n945), .S(n4372), .ZN(n2339) );
  MUX2ND0 U4688 ( .I0(n890), .I1(n947), .S(n4372), .ZN(n2337) );
  MUX2ND0 U4689 ( .I0(n889), .I1(n949), .S(n4372), .ZN(n2335) );
  MUX2ND0 U4690 ( .I0(n888), .I1(n951), .S(n4372), .ZN(n2333) );
  MUX2ND0 U4691 ( .I0(n887), .I1(n953), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2331) );
  MUX2ND0 U4692 ( .I0(n886), .I1(n955), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2329) );
  MUX2ND0 U4693 ( .I0(n885), .I1(n957), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2327) );
  MUX2ND0 U4694 ( .I0(n884), .I1(n959), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2325) );
  MUX2ND0 U4695 ( .I0(n883), .I1(n961), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2323) );
  MUX2ND0 U4696 ( .I0(n882), .I1(n963), .S(n4372), .ZN(n2321) );
  MUX2ND0 U4697 ( .I0(n881), .I1(n965), .S(n4372), .ZN(n2319) );
  MUX2ND0 U4698 ( .I0(n880), .I1(n967), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2317) );
  MUX2ND0 U4699 ( .I0(n879), .I1(n969), .S(n4372), .ZN(n2315) );
  MUX2ND0 U4700 ( .I0(n878), .I1(n971), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2313) );
  MUX2ND0 U4701 ( .I0(n877), .I1(n1005), .S(
        \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n2311) );
  NR2D0 U4702 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4783), .ZN(
        n2309) );
  CKXOR2D0 U4703 ( .A1(n876), .A2(n875), .Z(n4783) );
  NR2D0 U4704 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4784), .ZN(
        n2307) );
  XNR2D0 U4705 ( .A1(n4785), .A2(n874), .ZN(n4784) );
  NR2D0 U4706 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4786), .ZN(
        n2305) );
  CKXOR2D0 U4707 ( .A1(n873), .A2(n4787), .Z(n4786) );
  NR2D0 U4708 ( .A1(n874), .A2(n4785), .ZN(n4787) );
  IND2D0 U4709 ( .A1(n876), .B1(n875), .ZN(n4785) );
  NR2D0 U4710 ( .A1(n4788), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/UnLoad ), .ZN(
        n2303) );
  OA31D0 U4711 ( .A1(n874), .A2(n876), .A3(n873), .B(n875), .Z(n4788) );
  AO222D0 U4712 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ), .A2(
        n4779), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ), .B2(n4780), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .C2(n4781), 
        .Z(n2289) );
  AO222D0 U4713 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ), .A2(
        n4779), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ), .B2(n4780), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .C2(n4781), 
        .Z(n2287) );
  CKND0 U4714 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CN(
        n4781) );
  AN2D0 U4715 ( .A1(n4789), .A2(n4790), .Z(n4780) );
  AN3D0 U4716 ( .A1(n4791), .A2(n4792), .A3(n4793), .Z(n4779) );
  OAI21D0 U4717 ( .A1(n872), .A2(n4794), .B(n909), .ZN(n2285) );
  NR2D0 U4718 ( .A1(\SerDes_U1/Rx_ParClk ), .A2(n875), .ZN(n4794) );
  MUX2ND0 U4719 ( .I0(n871), .I1(n4795), .S(n4796), .ZN(n2283) );
  AOI211D0 U4720 ( .A1(n4797), .A2(n870), .B(n4798), .C(n4799), .ZN(n4795) );
  AOI211D0 U4721 ( .A1(n4800), .A2(n4801), .B(n4802), .C(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .ZN(n4798) );
  ND4D0 U4722 ( .A1(n4803), .A2(n4804), .A3(n4805), .A4(n4806), .ZN(n4801) );
  MUX2ND0 U4723 ( .I0(n4807), .I1(n4808), .S(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(n4797) );
  CKND2D0 U4724 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n4809), .ZN(n4808) );
  AN4D0 U4725 ( .A1(n4806), .A2(n4805), .A3(n4804), .A4(n4803), .Z(n4807) );
  OA211D0 U4726 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n4562), 
        .B(n4810), .C(n4811), .Z(n4803) );
  AOI21D0 U4727 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .A2(n4812), 
        .B(n4813), .ZN(n4811) );
  AOI22D0 U4728 ( .A1(n4563), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), 
        .B1(n4562), .B2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .ZN(
        n4804) );
  OAI33D0 U4729 ( .A1(n4814), .A2(n869), .A3(n4815), .B1(n4816), .B2(n4817), 
        .B3(n4818), .ZN(n2280) );
  XNR2D0 U4730 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .A2(n868), 
        .ZN(n4818) );
  XNR2D0 U4731 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .A2(n866), 
        .ZN(n4817) );
  IND3D0 U4732 ( .A1(n4819), .B1(n4820), .B2(n4821), .ZN(n4816) );
  XNR2D0 U4733 ( .A1(n867), .A2(n4562), .ZN(n4821) );
  XNR2D0 U4734 ( .A1(n865), .A2(n4560), .ZN(n4820) );
  OAI211D0 U4735 ( .A1(n864), .A2(n4796), .B(n4822), .C(n4823), .ZN(n2213) );
  AOI31D0 U4736 ( .A1(n4824), .A2(n4825), .A3(n4826), .B(n4827), .ZN(n4823) );
  OAI31D0 U4737 ( .A1(n4828), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), 
        .A3(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .B(n4829), .ZN(n4825) );
  MUX2ND0 U4738 ( .I0(n4830), .I1(n4831), .S(n4562), .ZN(n4829) );
  OAI32D0 U4739 ( .A1(n4832), .A2(n4563), .A3(n4806), .B1(n4810), .B2(n4833), 
        .ZN(n4831) );
  OAI32D0 U4740 ( .A1(n4832), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), 
        .A3(n4810), .B1(n4806), .B2(n4833), .ZN(n4830) );
  CKND2D0 U4741 ( .A1(n4834), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n4833) );
  XNR2D0 U4742 ( .A1(n4812), .A2(n4563), .ZN(n4834) );
  MUX2ND0 U4743 ( .I0(n4835), .I1(n4836), .S(n4562), .ZN(n4828) );
  NR2D0 U4744 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .A2(n4806), 
        .ZN(n4836) );
  NR2D0 U4745 ( .A1(n4563), .A2(n4810), .ZN(n4835) );
  ND3D0 U4746 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n4837), .A3(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(
        n4822) );
  ND4D0 U4747 ( .A1(n4838), .A2(n4839), .A3(n4840), .A4(n4841), .ZN(n4837) );
  XNR2D0 U4748 ( .A1(n4842), .A2(n4843), .ZN(n4840) );
  XNR2D0 U4749 ( .A1(n4812), .A2(n4844), .ZN(n4839) );
  XNR2D0 U4750 ( .A1(n4845), .A2(n4846), .ZN(n4838) );
  OAI32D0 U4751 ( .A1(n4847), .A2(n4848), .A3(n4849), .B1(n4814), .B2(n4850), 
        .ZN(n2207) );
  XNR2D0 U4752 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .A2(n862), 
        .ZN(n4848) );
  ND3D0 U4753 ( .A1(n4851), .A2(n4852), .A3(n4853), .ZN(n4847) );
  XNR2D0 U4754 ( .A1(n861), .A2(n4846), .ZN(n4853) );
  XNR2D0 U4755 ( .A1(n860), .A2(n4854), .ZN(n4852) );
  XNR2D0 U4756 ( .A1(n859), .A2(n4842), .ZN(n4851) );
  OAI221D0 U4757 ( .A1(n4855), .A2(n4802), .B1(n858), .B2(n4796), .C(n4856), 
        .ZN(n2204) );
  AOI31D0 U4758 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A3(n4857), .B(
        n4815), .ZN(n4856) );
  CKND0 U4759 ( .CLK(n4858), .CN(n4815) );
  CKND0 U4760 ( .CLK(n4809), .CN(n4857) );
  ND4D0 U4761 ( .A1(n4859), .A2(n4860), .A3(n4861), .A4(n4841), .ZN(n4809) );
  XNR2D0 U4762 ( .A1(n4563), .A2(n4862), .ZN(n4861) );
  XNR2D0 U4763 ( .A1(n4863), .A2(n4561), .ZN(n4860) );
  XNR2D0 U4764 ( .A1(n4864), .A2(n4562), .ZN(n4859) );
  CKND2D0 U4765 ( .A1(n872), .A2(n4799), .ZN(n4796) );
  CKND0 U4766 ( .CLK(n4800), .CN(n4855) );
  ND4D0 U4767 ( .A1(n4865), .A2(n4824), .A3(n4866), .A4(n4843), .ZN(n4800) );
  CKND2D0 U4768 ( .A1(n4810), .A2(n4806), .ZN(n4843) );
  CKND2D0 U4769 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n4561), 
        .ZN(n4806) );
  CKND2D0 U4770 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .A2(n4854), 
        .ZN(n4810) );
  XNR2D0 U4771 ( .A1(n4867), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), 
        .ZN(n4866) );
  CKND2D0 U4772 ( .A1(n4868), .A2(n4832), .ZN(n4867) );
  MUX2ND0 U4773 ( .I0(n4854), .I1(n4869), .S(n4812), .ZN(n4868) );
  NR2D0 U4774 ( .A1(n4854), .A2(n4846), .ZN(n4869) );
  CKND0 U4775 ( .CLK(n4841), .CN(n4824) );
  IND2D0 U4776 ( .A1(n4813), .B1(n4805), .ZN(n4841) );
  CKND2D0 U4777 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .A2(n4560), 
        .ZN(n4805) );
  NR2D0 U4778 ( .A1(n4560), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), 
        .ZN(n4813) );
  XNR3D0 U4779 ( .A1(n4846), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), 
        .A3(n4562), .ZN(n4865) );
  MUX2ND0 U4780 ( .I0(n4812), .I1(n862), .S(n4849), .ZN(n2198) );
  MUX2ND0 U4781 ( .I0(n4854), .I1(n860), .S(n4849), .ZN(n2196) );
  MUX2ND0 U4782 ( .I0(n4842), .I1(n859), .S(n4849), .ZN(n2194) );
  MUX2ND0 U4783 ( .I0(n4846), .I1(n861), .S(n4849), .ZN(n2192) );
  IND2D0 U4784 ( .A1(n872), .B1(n4814), .ZN(n4849) );
  OAI221D0 U4785 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n4802), .B1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .B2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .C(n4870), .ZN(
        n4814) );
  MUX2ND0 U4786 ( .I0(n4563), .I1(n868), .S(n4819), .ZN(n1678) );
  MUX2ND0 U4787 ( .I0(n4561), .I1(n866), .S(n4819), .ZN(n1676) );
  MUX2ND0 U4788 ( .I0(n4560), .I1(n865), .S(n4819), .ZN(n1674) );
  MUX2ND0 U4789 ( .I0(n4562), .I1(n867), .S(n4819), .ZN(n1672) );
  NR2D0 U4790 ( .A1(n4827), .A2(n4826), .ZN(n4819) );
  CKND0 U4791 ( .CLK(n4870), .CN(n4826) );
  CKND2D0 U4792 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n870), .ZN(n4870) );
  AO222D0 U4793 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ), .A2(
        n4871), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ), .B2(n4872), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .C2(n4873), 
        .Z(n1655) );
  AO222D0 U4794 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ), .A2(
        n4871), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ), .B2(n4872), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .C2(n4873), 
        .Z(n1652) );
  AO222D0 U4795 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ), .A2(
        n4871), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ), .B2(n4872), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .C2(n4873), 
        .Z(n1650) );
  CKND0 U4796 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CN(
        n4873) );
  AN2D0 U4797 ( .A1(n4874), .A2(n4875), .Z(n4872) );
  AN3D0 U4798 ( .A1(n4876), .A2(n4877), .A3(n4878), .Z(n4871) );
  CKXOR2D0 U4799 ( .A1(\SerDes_U2/Tx_SerClk ), .A2(n4879), .Z(n1646) );
  AO222D0 U4800 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ), .A2(
        n4880), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ), .B2(n4881), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .C2(n4882), 
        .Z(n1623) );
  XNR2D0 U4801 ( .A1(n4883), .A2(\SerDes_U2/Des_U1/SerialClk ), .ZN(n1619) );
  MUX2ND0 U4802 ( .I0(n857), .I1(n856), .S(n4472), .ZN(n1553) );
  MUX2ND0 U4803 ( .I0(n823), .I1(n822), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1551) );
  MUX2ND0 U4804 ( .I0(n821), .I1(n820), .S(n4472), .ZN(n1549) );
  MUX2ND0 U4805 ( .I0(n819), .I1(n818), .S(n4472), .ZN(n1547) );
  MUX2ND0 U4806 ( .I0(n817), .I1(n816), .S(n4472), .ZN(n1545) );
  MUX2ND0 U4807 ( .I0(n815), .I1(n814), .S(n4472), .ZN(n1543) );
  MUX2ND0 U4808 ( .I0(n813), .I1(n812), .S(n4472), .ZN(n1541) );
  MUX2ND0 U4809 ( .I0(n811), .I1(n810), .S(n4472), .ZN(n1539) );
  MUX2ND0 U4810 ( .I0(n809), .I1(n808), .S(n4472), .ZN(n1537) );
  MUX2ND0 U4811 ( .I0(n807), .I1(n806), .S(n4472), .ZN(n1535) );
  MUX2ND0 U4812 ( .I0(n805), .I1(n804), .S(n4472), .ZN(n1533) );
  MUX2ND0 U4813 ( .I0(n803), .I1(n802), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1531) );
  MUX2ND0 U4814 ( .I0(n801), .I1(n800), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1529) );
  MUX2ND0 U4815 ( .I0(n799), .I1(n798), .S(n4472), .ZN(n1527) );
  MUX2ND0 U4816 ( .I0(n797), .I1(n796), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1525) );
  MUX2ND0 U4817 ( .I0(n795), .I1(n794), .S(n4472), .ZN(n1523) );
  MUX2ND0 U4818 ( .I0(n793), .I1(n792), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1521) );
  MUX2ND0 U4819 ( .I0(n791), .I1(n790), .S(n4472), .ZN(n1519) );
  MUX2ND0 U4820 ( .I0(n789), .I1(n788), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1517) );
  MUX2ND0 U4821 ( .I0(n787), .I1(n786), .S(n4472), .ZN(n1515) );
  MUX2ND0 U4822 ( .I0(n785), .I1(n784), .S(n4472), .ZN(n1513) );
  MUX2ND0 U4823 ( .I0(n783), .I1(n782), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1511) );
  MUX2ND0 U4824 ( .I0(n781), .I1(n780), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1509) );
  MUX2ND0 U4825 ( .I0(n779), .I1(n778), .S(n4472), .ZN(n1507) );
  MUX2ND0 U4826 ( .I0(n777), .I1(n776), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1505) );
  MUX2ND0 U4827 ( .I0(n775), .I1(n774), .S(n4472), .ZN(n1503) );
  MUX2ND0 U4828 ( .I0(n773), .I1(n772), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1501) );
  MUX2ND0 U4829 ( .I0(n771), .I1(n770), .S(n4472), .ZN(n1499) );
  MUX2ND0 U4830 ( .I0(n769), .I1(n768), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1497) );
  MUX2ND0 U4831 ( .I0(n767), .I1(n766), .S(n4472), .ZN(n1495) );
  MUX2ND0 U4832 ( .I0(n765), .I1(n764), .S(n4472), .ZN(n1493) );
  MUX2ND0 U4833 ( .I0(n763), .I1(n762), .S(n4472), .ZN(n1491) );
  MUX2ND0 U4834 ( .I0(n760), .I1(n763), .S(n4373), .ZN(n1487) );
  MUX2ND0 U4835 ( .I0(n759), .I1(n765), .S(n4373), .ZN(n1485) );
  MUX2ND0 U4836 ( .I0(n758), .I1(n767), .S(n4373), .ZN(n1483) );
  MUX2ND0 U4837 ( .I0(n757), .I1(n769), .S(n4373), .ZN(n1481) );
  MUX2ND0 U4838 ( .I0(n756), .I1(n771), .S(n4373), .ZN(n1479) );
  MUX2ND0 U4839 ( .I0(n755), .I1(n773), .S(n4373), .ZN(n1477) );
  MUX2ND0 U4840 ( .I0(n754), .I1(n775), .S(n4373), .ZN(n1475) );
  MUX2ND0 U4841 ( .I0(n753), .I1(n777), .S(n4373), .ZN(n1473) );
  MUX2ND0 U4842 ( .I0(n752), .I1(n779), .S(n4373), .ZN(n1471) );
  MUX2ND0 U4843 ( .I0(n751), .I1(n781), .S(n4373), .ZN(n1469) );
  MUX2ND0 U4844 ( .I0(n750), .I1(n783), .S(n4373), .ZN(n1467) );
  MUX2ND0 U4845 ( .I0(n749), .I1(n785), .S(n4373), .ZN(n1465) );
  MUX2ND0 U4846 ( .I0(n748), .I1(n787), .S(n4373), .ZN(n1463) );
  MUX2ND0 U4847 ( .I0(n747), .I1(n789), .S(n4373), .ZN(n1461) );
  MUX2ND0 U4848 ( .I0(n746), .I1(n791), .S(n4373), .ZN(n1459) );
  MUX2ND0 U4849 ( .I0(n745), .I1(n793), .S(n4373), .ZN(n1457) );
  MUX2ND0 U4850 ( .I0(n744), .I1(n795), .S(n4373), .ZN(n1455) );
  MUX2ND0 U4851 ( .I0(n743), .I1(n797), .S(n4373), .ZN(n1453) );
  MUX2ND0 U4852 ( .I0(n742), .I1(n799), .S(n4373), .ZN(n1451) );
  MUX2ND0 U4853 ( .I0(n741), .I1(n801), .S(n4373), .ZN(n1449) );
  MUX2ND0 U4854 ( .I0(n740), .I1(n803), .S(n4373), .ZN(n1447) );
  MUX2ND0 U4855 ( .I0(n739), .I1(n805), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1445) );
  MUX2ND0 U4856 ( .I0(n738), .I1(n807), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1443) );
  MUX2ND0 U4857 ( .I0(n737), .I1(n809), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1441) );
  MUX2ND0 U4858 ( .I0(n736), .I1(n811), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1439) );
  MUX2ND0 U4859 ( .I0(n735), .I1(n813), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1437) );
  MUX2ND0 U4860 ( .I0(n734), .I1(n815), .S(n4373), .ZN(n1435) );
  MUX2ND0 U4861 ( .I0(n733), .I1(n817), .S(n4373), .ZN(n1433) );
  MUX2ND0 U4862 ( .I0(n732), .I1(n819), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1431) );
  MUX2ND0 U4863 ( .I0(n731), .I1(n821), .S(n4373), .ZN(n1429) );
  MUX2ND0 U4864 ( .I0(n730), .I1(n823), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1427) );
  MUX2ND0 U4865 ( .I0(n729), .I1(n857), .S(
        \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(n1425) );
  NR2D0 U4866 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4884), .ZN(
        n1423) );
  CKXOR2D0 U4867 ( .A1(n728), .A2(n727), .Z(n4884) );
  NR2D0 U4868 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4885), .ZN(
        n1421) );
  XNR2D0 U4869 ( .A1(n4886), .A2(n726), .ZN(n4885) );
  NR2D0 U4870 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .A2(n4887), .ZN(
        n1419) );
  CKXOR2D0 U4871 ( .A1(n725), .A2(n4888), .Z(n4887) );
  NR2D0 U4872 ( .A1(n726), .A2(n4886), .ZN(n4888) );
  IND2D0 U4873 ( .A1(n728), .B1(n727), .ZN(n4886) );
  NR2D0 U4874 ( .A1(n4889), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/UnLoad ), .ZN(
        n1417) );
  OA31D0 U4875 ( .A1(n726), .A2(n728), .A3(n725), .B(n727), .Z(n4889) );
  AO222D0 U4876 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ), .A2(
        n4880), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ), .B2(n4881), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .C2(n4882), 
        .Z(n1403) );
  AO222D0 U4877 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ), .A2(
        n4880), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ), .B2(n4881), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .C2(n4882), 
        .Z(n1401) );
  CKND0 U4878 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CN(
        n4882) );
  AN2D0 U4879 ( .A1(n4890), .A2(n4891), .Z(n4881) );
  AN3D0 U4880 ( .A1(n4892), .A2(n4893), .A3(n4894), .Z(n4880) );
  OAI21D0 U4881 ( .A1(n724), .A2(n4895), .B(n761), .ZN(n1399) );
  NR2D0 U4882 ( .A1(\SerDes_U2/Rx_ParClk ), .A2(n727), .ZN(n4895) );
  MUX2ND0 U4883 ( .I0(n723), .I1(n4896), .S(n4897), .ZN(n1397) );
  AOI32D0 U4884 ( .A1(n4898), .A2(n4899), .A3(n4900), .B1(n722), .B2(n4901), 
        .ZN(n4896) );
  IOA22D0 U4885 ( .B1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .B2(
        n4902), .A1(n4903), .A2(n4904), .ZN(n4901) );
  NR4D0 U4886 ( .A1(n4905), .A2(n4906), .A3(n4907), .A4(n4899), .ZN(n4902) );
  OAI32D0 U4887 ( .A1(n4907), .A2(n4905), .A3(n4906), .B1(n4908), .B2(n4909), 
        .ZN(n4898) );
  CKND0 U4888 ( .CLK(n4910), .CN(n4909) );
  OA22D0 U4889 ( .A1(n4911), .A2(n4912), .B1(n4913), .B2(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .Z(n4908) );
  OAI221D0 U4890 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .A2(n4914), 
        .B1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .B2(n4915), .C(n4911), 
        .ZN(n4906) );
  OAI22D0 U4891 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n4481), 
        .B1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .B2(n4480), .ZN(
        n4907) );
  OAI31D0 U4892 ( .A1(n4916), .A2(n721), .A3(n4917), .B(n4918), .ZN(n1394) );
  IND4D0 U4893 ( .A1(n4919), .B1(n4920), .B2(n4921), .B3(n4922), .ZN(n4918) );
  XNR2D0 U4894 ( .A1(n719), .A2(n4480), .ZN(n4922) );
  XNR2D0 U4895 ( .A1(n720), .A2(n4481), .ZN(n4921) );
  XNR2D0 U4896 ( .A1(n718), .A2(n4482), .ZN(n4920) );
  OAI211D0 U4897 ( .A1(n717), .A2(n4897), .B(n4923), .C(n4924), .ZN(n1327) );
  AOI31D0 U4898 ( .A1(n722), .A2(n4925), .A3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .B(n4900), .ZN(
        n4924) );
  OAI32D0 U4899 ( .A1(n4926), .A2(n4911), .A3(n4912), .B1(n4927), .B2(n4913), 
        .ZN(n4925) );
  CKND2D0 U4900 ( .A1(n4928), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), 
        .ZN(n4913) );
  AOI22D0 U4901 ( .A1(n4905), .A2(n4929), .B1(n4930), .B2(n4482), .ZN(n4927)
         );
  NR2D0 U4902 ( .A1(n4482), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n4905) );
  CKND2D0 U4903 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n4481), 
        .ZN(n4911) );
  XNR2D0 U4904 ( .A1(n4915), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), 
        .ZN(n4926) );
  OAI31D0 U4905 ( .A1(n4931), .A2(n4928), .A3(n4932), .B(n4904), .ZN(n4923) );
  XNR2D0 U4906 ( .A1(n4929), .A2(n4933), .ZN(n4932) );
  XNR2D0 U4907 ( .A1(n4934), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n4931) );
  CKND0 U4908 ( .CLK(n4935), .CN(n4897) );
  OAI211D0 U4909 ( .A1(n4936), .A2(n4903), .B(n4937), .C(n4938), .ZN(n1324) );
  AOI21D0 U4910 ( .A1(n4935), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .B(n4939), .ZN(
        n4938) );
  AOI31D0 U4911 ( .A1(n4940), .A2(n4910), .A3(n4928), .B(n4941), .ZN(n4939) );
  CKND0 U4912 ( .CLK(n4912), .CN(n4928) );
  CKXOR2D0 U4913 ( .A1(n4482), .A2(n4942), .Z(n4910) );
  CKND2D0 U4914 ( .A1(n4943), .A2(n4944), .ZN(n4942) );
  XNR2D0 U4915 ( .A1(n4929), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), 
        .ZN(n4940) );
  NR2D0 U4916 ( .A1(\SerDes_U2/Des_U1/ParValidDecode ), .A2(n4945), .ZN(n4935)
         );
  ND3D0 U4917 ( .A1(n4946), .A2(n4912), .A3(n4947), .ZN(n4903) );
  XNR2D0 U4918 ( .A1(n4948), .A2(n4481), .ZN(n4947) );
  XNR2D0 U4919 ( .A1(n4914), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), 
        .ZN(n4912) );
  XNR2D0 U4920 ( .A1(n4482), .A2(n4949), .ZN(n4946) );
  CKND0 U4921 ( .CLK(n4904), .CN(n4936) );
  NR2D0 U4922 ( .A1(n4899), .A2(n4950), .ZN(n4904) );
  MUX2ND0 U4923 ( .I0(n4951), .I1(n4952), .S(n4916), .ZN(n1319) );
  ND4D0 U4924 ( .A1(n4953), .A2(n4954), .A3(n4955), .A4(
        \SerDes_U2/Des_U1/ParValidDecode ), .ZN(n4952) );
  XNR2D0 U4925 ( .A1(n713), .A2(n4914), .ZN(n4955) );
  XNR2D0 U4926 ( .A1(n714), .A2(n4929), .ZN(n4954) );
  XNR2D0 U4927 ( .A1(n712), .A2(n4915), .ZN(n4953) );
  MUX2ND0 U4928 ( .I0(n712), .I1(n4915), .S(n4956), .ZN(n1314) );
  MUX2ND0 U4929 ( .I0(n713), .I1(n4914), .S(n4956), .ZN(n1312) );
  MUX2ND0 U4930 ( .I0(n714), .I1(n4929), .S(n4956), .ZN(n1310) );
  AN2D0 U4931 ( .A1(n4916), .A2(\SerDes_U2/Des_U1/ParValidDecode ), .Z(n4956)
         );
  OAI22D0 U4932 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n4941), .B1(n4957), .B2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .ZN(n4916) );
  NR2D0 U4933 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n4950), .ZN(n4957) );
  MUX2ND0 U4934 ( .I0(n4482), .I1(n718), .S(n4919), .ZN(n1052) );
  MUX2ND0 U4935 ( .I0(n4480), .I1(n719), .S(n4919), .ZN(n1050) );
  MUX2ND0 U4936 ( .I0(n4481), .I1(n720), .S(n4919), .ZN(n1048) );
  AOI21D0 U4937 ( .A1(n722), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .B(n4900), .ZN(
        n4919) );
  AO22D0 U4938 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ), .A2(
        n4878), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ), .B2(n4874), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ) );
  MUX2ND0 U4939 ( .I0(n4958), .I1(n4959), .S(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .ZN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ) );
  CKND2D0 U4940 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        n4875), .ZN(n4959) );
  ND3D0 U4941 ( .A1(n4960), .A2(n4877), .A3(n4961), .ZN(n4875) );
  ND4D0 U4942 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .ZN(n4961) );
  IND3D0 U4943 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .B1(
        n4877), .B2(n4876), .ZN(n4958) );
  CKND2D0 U4944 ( .A1(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .ZN(n4876) );
  AO22D0 U4945 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ), .A2(
        n4878), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ), .B2(n4874), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ) );
  AO22D0 U4946 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ), .A2(
        n4878), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ), .B2(n4874), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ) );
  AN2D0 U4947 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .Z(n4874) );
  NR2D0 U4948 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .ZN(n4878) );
  INR2D0 U4949 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ), .B1(
        n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ) );
  INR2D0 U4950 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ), .B1(
        n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ) );
  INR2D0 U4951 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ), .B1(
        n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ) );
  INR2D0 U4952 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ), .B1(
        n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ) );
  INR2D0 U4953 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ), .B1(
        n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ) );
  INR2D0 U4954 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ), .B1(n4879), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ) );
  OA21D0 U4955 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), 
        .A2(n4877), .B(n4962), .Z(n4879) );
  IOA22D0 U4956 ( .B1(n4963), .B2(n4964), .A1(n4877), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .ZN(n4962)
         );
  AOI221D0 U4957 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .A2(n4960), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .B2(n4965), .C(n4966), .ZN(n4964) );
  AOI221D0 U4958 ( .A1(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(n4967), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B2(n4968), 
        .C(n4969), .ZN(n4966) );
  IAO21D0 U4959 ( .A1(n4968), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .ZN(n4969)
         );
  OAI32D0 U4960 ( .A1(n4970), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .A3(n4971), 
        .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .B2(
        n4972), .ZN(n4968) );
  AN2D0 U4961 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), 
        .A2(n4972), .Z(n4971) );
  CKND0 U4962 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .CN(n4972) );
  CKND0 U4963 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .CN(n4970) );
  CKND0 U4964 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .CN(n4967) );
  CKND0 U4965 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .CN(n4965) );
  NR2D0 U4966 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), 
        .A2(n4960), .ZN(n4963) );
  CKND0 U4967 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .CN(n4960) );
  CKND0 U4968 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .CN(n4877) );
  AN2D0 U4969 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]), .A2(
        n4440), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ) );
  CKXOR2D0 U4970 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ) );
  XNR2D0 U4971 ( .A1(n4973), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ) );
  AO221D0 U4972 ( .A1(n4974), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .B1(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), .B2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .C(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ) );
  NR2D0 U4973 ( .A1(n4973), .A2(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ) );
  CKND0 U4974 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ) );
  IOA21D0 U4975 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .B(n4973), 
        .ZN(n4974) );
  CKND0 U4976 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .CN(n4973) );
  AN2D0 U4977 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ) );
  AN2D0 U4978 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N83 ) );
  AN2D0 U4979 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ) );
  AN2D0 U4980 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N81 ) );
  AN2D0 U4981 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ) );
  AN2D0 U4982 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N79 ) );
  AN2D0 U4983 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ) );
  AN2D0 U4984 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N77 ) );
  AN2D0 U4985 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ) );
  AN2D0 U4986 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N75 ) );
  AN2D0 U4987 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ) );
  AN2D0 U4988 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N73 ) );
  AN2D0 U4989 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ) );
  AN2D0 U4990 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N71 ) );
  AN2D0 U4991 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ) );
  AN2D0 U4992 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N69 ) );
  AN2D0 U4993 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ) );
  AN2D0 U4994 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N67 ) );
  AN2D0 U4995 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ) );
  AN2D0 U4996 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N65 ) );
  AN2D0 U4997 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ) );
  AN2D0 U4998 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N63 ) );
  AN2D0 U4999 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ) );
  AN2D0 U5000 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N61 ) );
  AN2D0 U5001 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ) );
  AN2D0 U5002 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N59 ) );
  AN2D0 U5003 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ) );
  AN2D0 U5004 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N57 ) );
  AN2D0 U5005 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ) );
  AN2D0 U5006 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N55 ) );
  AN2D0 U5007 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ) );
  AN2D0 U5008 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]), .A2(
        n4371), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N53 ) );
  OAI31D0 U5009 ( .A1(n4975), .A2(n4976), .A3(n4977), .B(n4978), .ZN(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ) );
  OAI21D0 U5010 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N23 ), .A2(n4979), .B(n4980), .ZN(n4978) );
  MUX2ND0 U5011 ( .I0(n4981), .I1(n4982), .S(n4979), .ZN(n4980) );
  MUX3ND0 U5012 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/N25 ), .I1(n4983), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N24 ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .S1(n4984), .ZN(n4982) );
  NR2D0 U5013 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .ZN(n4984) );
  MUX2D0 U5014 ( .I0(n4985), .I1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ), .S(n4976), 
        .Z(n4983) );
  AN2D0 U5015 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N27 ), .A2(n4977), .Z(n4985)
         );
  IND2D0 U5016 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .B1(n4977), .ZN(
        n4979) );
  CKND0 U5017 ( .CLK(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), .CN(n4977) );
  OAI21D0 U5018 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .B(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .ZN(n4976) );
  MUX2ND0 U5019 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/N29 ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ), .S(n4981), .ZN(n4975) );
  CKND0 U5020 ( .CLK(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .CN(n4981) );
  CKND0 U5021 ( .CLK(ClockB), .CN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U5022 ( .A1(n4696), .A2(n4616), .A3(n4671), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ) );
  OAI22D0 U5023 ( .A1(n4616), .A2(n4527), .B1(n4693), .B2(n4671), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ) );
  OA211D0 U5024 ( .A1(n4986), .A2(n4637), .B(n4987), .C(n4663), .Z(n4693) );
  OAI22D0 U5025 ( .A1(n4616), .A2(n4526), .B1(n4694), .B2(n4671), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ) );
  XNR2D0 U5026 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n4986), 
        .ZN(n4694) );
  OAI22D0 U5027 ( .A1(n4616), .A2(n4525), .B1(n4692), .B2(n4671), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ) );
  AN2D0 U5028 ( .A1(n4988), .A2(n4989), .Z(n4692) );
  OAI22D0 U5029 ( .A1(n4616), .A2(n4524), .B1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .B2(n4671), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ) );
  CKND2D0 U5030 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .A2(n4616), 
        .ZN(n4671) );
  CKND0 U5031 ( .CLK(n4643), .CN(n4616) );
  NR3D0 U5032 ( .A1(n1032), .A2(n1033), .A3(n1031), .ZN(n4643) );
  NR2D0 U5033 ( .A1(n4657), .A2(n4642), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ) );
  XNR2D0 U5034 ( .A1(n4990), .A2(n4527), .ZN(n4657) );
  CKND2D0 U5035 ( .A1(n4696), .A2(n4642), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ) );
  NR2D0 U5036 ( .A1(n4642), .A2(n4656), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ) );
  OAI21D0 U5037 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .A2(n4991), 
        .B(n4990), .ZN(n4656) );
  CKND2D0 U5038 ( .A1(n4991), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), 
        .ZN(n4990) );
  NR2D0 U5039 ( .A1(n4525), .A2(n4524), .ZN(n4991) );
  MUX2ND0 U5040 ( .I0(n4992), .I1(n4993), .S(n4525), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ) );
  OR2D0 U5041 ( .A1(n4642), .A2(n4524), .Z(n4993) );
  CKND0 U5042 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .CN(n4992) );
  NR2D0 U5043 ( .A1(n4642), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), 
        .ZN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ) );
  CKND2D0 U5044 ( .A1(n3582), .A2(n4696), .ZN(n4642) );
  CKND0 U5045 ( .CLK(n4620), .CN(n4696) );
  NR3D0 U5046 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n4620) );
  ND3D0 U5047 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), .A3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .ZN(n4995) );
  OR2D0 U5048 ( .A1(n4663), .A2(n1023), .Z(n4997) );
  CKND2D0 U5049 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .A2(n4638), 
        .ZN(n4663) );
  ND3D0 U5050 ( .A1(n4986), .A2(n4637), .A3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .ZN(n4987) );
  ND3D0 U5051 ( .A1(n4637), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), 
        .A3(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .ZN(n4998) );
  CKND0 U5052 ( .CLK(n4986), .CN(n4994) );
  NR2D0 U5053 ( .A1(n4675), .A2(n4676), .ZN(n4986) );
  CKND2D0 U5054 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n4676), 
        .ZN(n4989) );
  CKND2D0 U5055 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .A2(n4675), 
        .ZN(n4988) );
  ND3D0 U5056 ( .A1(n4637), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_MemWriteCmd ), 
        .A3(n4638), .ZN(n4999) );
  CKND0 U5057 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .CN(n4638)
         );
  CKND0 U5058 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .CN(n4637)
         );
  CKND2D0 U5059 ( .A1(n4676), .A2(n4675), .ZN(n4996) );
  CKND0 U5060 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .CN(n4675)
         );
  CKND0 U5061 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .CN(n4676)
         );
  AO22D0 U5062 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ), .A2(
        n4894), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ), .B2(n4890), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ) );
  MUX2ND0 U5063 ( .I0(n5000), .I1(n5001), .S(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .ZN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ) );
  CKND2D0 U5064 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        n4891), .ZN(n5001) );
  ND3D0 U5065 ( .A1(n5002), .A2(n4893), .A3(n5003), .ZN(n4891) );
  ND4D0 U5066 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .ZN(n5003) );
  IND3D0 U5067 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .B1(
        n4893), .B2(n4892), .ZN(n5000) );
  CKND2D0 U5068 ( .A1(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n4892) );
  AO22D0 U5069 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ), .A2(
        n4894), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ), .B2(n4890), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ) );
  AO22D0 U5070 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ), .A2(
        n4894), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ), .B2(n4890), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ) );
  AN2D0 U5071 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .Z(n4890) );
  NR2D0 U5072 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .ZN(n4894) );
  AN2D0 U5073 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ), .A2(n4883), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ) );
  AN2D0 U5074 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ), .A2(n4883), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ) );
  AN2D0 U5075 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ), .A2(n4883), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ) );
  AN2D0 U5076 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ), .A2(n4883), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ) );
  AN2D0 U5077 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ), .A2(n4883), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ) );
  AN2D0 U5078 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ), .A2(n4883), 
        .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ) );
  OAI21D0 U5079 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), 
        .A2(n4893), .B(n5004), .ZN(n4883) );
  IOA22D0 U5080 ( .B1(n5005), .B2(n5006), .A1(n4893), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .ZN(n5004)
         );
  AOI221D0 U5081 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .A2(n5002), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .B2(n5007), .C(n5008), .ZN(n5006) );
  AOI221D0 U5082 ( .A1(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(n5009), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B2(n5010), 
        .C(n5011), .ZN(n5008) );
  IAO21D0 U5083 ( .A1(n5010), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .ZN(n5011)
         );
  OAI32D0 U5084 ( .A1(n5012), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .A3(n5013), 
        .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .B2(
        n5014), .ZN(n5010) );
  AN2D0 U5085 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), 
        .A2(n5014), .Z(n5013) );
  CKND0 U5086 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .CN(n5014) );
  CKND0 U5087 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .CN(n5012) );
  CKND0 U5088 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .CN(n5009) );
  CKND0 U5089 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .CN(n5007) );
  NR2D0 U5090 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), 
        .A2(n5002), .ZN(n5005) );
  CKND0 U5091 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .CN(n5002) );
  CKND0 U5092 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .CN(n4893) );
  AN2D0 U5093 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]), .A2(
        n4440), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ) );
  CKXOR2D0 U5094 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ) );
  XNR2D0 U5095 ( .A1(n5015), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ) );
  AO221D0 U5096 ( .A1(n5016), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .B1(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), .B2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .C(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ) );
  NR2D0 U5097 ( .A1(n5015), .A2(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .ZN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ) );
  CKND0 U5098 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ) );
  IOA21D0 U5099 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .B(n5015), 
        .ZN(n5016) );
  CKND0 U5100 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .CN(n5015) );
  CKND2D0 U5101 ( .A1(\SerDes_U2/Rx_ParClk ), .A2(ClockA), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U5102 ( .A1(n4945), .A2(n4937), .A3(n715), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ) );
  OAI22D0 U5103 ( .A1(n4482), .A2(n4937), .B1(n4949), .B2(n4951), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ) );
  AN2D0 U5104 ( .A1(n5017), .A2(n4943), .Z(n4949) );
  MUX2D0 U5105 ( .I0(n4915), .I1(n4944), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .Z(n5017) );
  OAI22D0 U5106 ( .A1(n4481), .A2(n4937), .B1(n4948), .B2(n4951), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ) );
  CKND2D0 U5107 ( .A1(n4937), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), 
        .ZN(n4951) );
  XNR2D0 U5108 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .ZN(n4948) );
  MUX2ND0 U5109 ( .I0(n4480), .I1(n5018), .S(n4937), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ) );
  CKND0 U5110 ( .CLK(n4917), .CN(n4937) );
  NR2D0 U5111 ( .A1(n4899), .A2(n4941), .ZN(n4917) );
  CKND0 U5112 ( .CLK(n4900), .CN(n4941) );
  NR2D0 U5113 ( .A1(n4950), .A2(n722), .ZN(n4900) );
  NR2D0 U5114 ( .A1(n4934), .A2(n5019), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ) );
  XNR2D0 U5115 ( .A1(n4482), .A2(n5020), .ZN(n4934) );
  CKND2D0 U5116 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n5020) );
  CKND2D0 U5117 ( .A1(n721), .A2(n4945), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ) );
  INR2D0 U5118 ( .A1(n4933), .B1(n5019), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ) );
  XNR2D0 U5119 ( .A1(n4481), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), 
        .ZN(n4933) );
  NR2D0 U5120 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .A2(n5019), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ) );
  IND2D0 U5121 ( .A1(n721), .B1(n4945), .ZN(n5019) );
  ND3D0 U5122 ( .A1(n4950), .A2(n4899), .A3(n722), .ZN(n4945) );
  CKND0 U5123 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .CN(
        n4899) );
  CKND0 U5124 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .CN(
        n4950) );
  NR3D0 U5125 ( .A1(n5018), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ) );
  NR3D0 U5126 ( .A1(n5021), .A2(n4929), .A3(n4915), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ) );
  NR3D0 U5127 ( .A1(n5018), .A2(n4929), .A3(n4915), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ) );
  CKND0 U5128 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .CN(n4929)
         );
  CKND0 U5129 ( .CLK(n4930), .CN(n4943) );
  NR2D0 U5130 ( .A1(n4915), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), 
        .ZN(n4930) );
  CKND2D0 U5131 ( .A1(n4914), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), 
        .ZN(n5018) );
  CKND0 U5132 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .CN(n4914)
         );
  CKND2D0 U5133 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n4915), 
        .ZN(n4944) );
  CKND0 U5134 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .CN(n4915)
         );
  NR3D0 U5135 ( .A1(n5021), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ) );
  CKND2D0 U5136 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .ZN(n5021) );
  NR2D0 U5137 ( .A1(n5022), .A2(n5023), .ZN(\SerDes_U2/Des_U1/DesDec_Rx1/N47 )
         );
  CKND2D0 U5138 ( .A1(n5024), .A2(n5025), .ZN(n5023) );
  NR4D0 U5139 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ), .ZN(n5025) );
  NR4D0 U5140 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ), .ZN(n5024) );
  AN4D0 U5141 ( .A1(n5026), .A2(n5027), .A3(n5028), .A4(n5029), .Z(n5022) );
  NR4D0 U5142 ( .A1(n5030), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ), 
        .A3(n855), .A4(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ), .ZN(n5029)
         );
  ND3D0 U5143 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ), .ZN(n5030) );
  NR4D0 U5144 ( .A1(n5031), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ), .ZN(n5028) );
  ND3D0 U5145 ( .A1(n841), .A2(n837), .A3(n842), .ZN(n5031) );
  NR4D0 U5146 ( .A1(n5032), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ), .ZN(n5027) );
  ND3D0 U5147 ( .A1(n4606), .A2(n849), .A3(n4607), .ZN(n5032) );
  NR4D0 U5148 ( .A1(n5033), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ), .ZN(n5026) );
  ND3D0 U5149 ( .A1(n4609), .A2(n4608), .A3(n4610), .ZN(n5033) );
  OA21D0 U5150 ( .A1(n5034), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .B(
        \SerDes_U2/SerLineValid ), .Z(\SerDes_U2/Des_U1/DesDec_Rx1/N43 ) );
  NR4D0 U5151 ( .A1(n5035), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ), .ZN(n5034) );
  OR2D0 U5152 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ), .Z(n5035) );
  INR2D0 U5153 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N34 ), .B1(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N42 ) );
  INR2D0 U5154 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N33 ), .B1(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N41 ) );
  INR2D0 U5155 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N32 ), .B1(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N40 ) );
  INR2D0 U5156 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N31 ), .B1(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N39 ) );
  INR2D0 U5157 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N30 ), .B1(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N38 ) );
  NR2D0 U5158 ( .A1(\SerDes_U2/Rx_ParClk ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N37 ) );
  AO22D0 U5159 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ), .A2(
        n4777), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ), .B2(n4773), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ) );
  MUX2ND0 U5160 ( .I0(n5036), .I1(n5037), .S(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .ZN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ) );
  CKND2D0 U5161 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        n4774), .ZN(n5037) );
  ND3D0 U5162 ( .A1(n5038), .A2(n4776), .A3(n5039), .ZN(n4774) );
  ND4D0 U5163 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .ZN(n5039) );
  IND3D0 U5164 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .B1(
        n4776), .B2(n4775), .ZN(n5036) );
  CKND2D0 U5165 ( .A1(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .ZN(n4775) );
  AO22D0 U5166 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ), .A2(
        n4777), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ), .B2(n4773), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ) );
  AO22D0 U5167 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ), .A2(
        n4777), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ), .B2(n4773), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ) );
  AN2D0 U5168 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .Z(n4773) );
  NR2D0 U5169 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .ZN(n4777) );
  INR2D0 U5170 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ), .B1(
        n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ) );
  INR2D0 U5171 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ), .B1(
        n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ) );
  INR2D0 U5172 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ), .B1(
        n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ) );
  INR2D0 U5173 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ), .B1(
        n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ) );
  INR2D0 U5174 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ), .B1(
        n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ) );
  INR2D0 U5175 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ), .B1(n4778), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ) );
  OA21D0 U5176 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), 
        .A2(n4776), .B(n5040), .Z(n4778) );
  IOA22D0 U5177 ( .B1(n5041), .B2(n5042), .A1(n4776), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .ZN(n5040)
         );
  AOI221D0 U5178 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .A2(n5038), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .B2(n5043), .C(n5044), .ZN(n5042) );
  AOI221D0 U5179 ( .A1(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(n5045), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B2(n5046), 
        .C(n5047), .ZN(n5044) );
  IAO21D0 U5180 ( .A1(n5046), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .ZN(n5047)
         );
  OAI32D0 U5181 ( .A1(n5048), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .A3(n5049), 
        .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .B2(
        n5050), .ZN(n5046) );
  AN2D0 U5182 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), 
        .A2(n5050), .Z(n5049) );
  CKND0 U5183 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .CN(n5050) );
  CKND0 U5184 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .CN(n5048) );
  CKND0 U5185 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .CN(n5045) );
  CKND0 U5186 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .CN(n5043) );
  NR2D0 U5187 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), 
        .A2(n5038), .ZN(n5041) );
  CKND0 U5188 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .CN(n5038) );
  CKND0 U5189 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .CN(n4776) );
  AN2D0 U5190 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]), .A2(
        n4440), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ) );
  CKXOR2D0 U5191 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ) );
  XNR2D0 U5192 ( .A1(n5051), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ) );
  AO221D0 U5193 ( .A1(n5052), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .B1(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), .B2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .C(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ) );
  NR2D0 U5194 ( .A1(n5051), .A2(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ) );
  CKND0 U5195 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ) );
  IOA21D0 U5196 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .B(n5051), 
        .ZN(n5052) );
  CKND0 U5197 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .CN(n5051) );
  AN2D0 U5198 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [31]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N84 ) );
  AN2D0 U5199 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [30]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ) );
  AN2D0 U5200 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [29]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N82 ) );
  AN2D0 U5201 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [28]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ) );
  AN2D0 U5202 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [27]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N80 ) );
  AN2D0 U5203 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [26]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ) );
  AN2D0 U5204 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [25]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N78 ) );
  AN2D0 U5205 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [24]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ) );
  AN2D0 U5206 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [23]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N76 ) );
  AN2D0 U5207 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [22]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ) );
  AN2D0 U5208 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [21]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N74 ) );
  AN2D0 U5209 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [20]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ) );
  AN2D0 U5210 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [19]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N72 ) );
  AN2D0 U5211 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [18]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ) );
  AN2D0 U5212 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [17]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N70 ) );
  AN2D0 U5213 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [16]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ) );
  AN2D0 U5214 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [15]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N68 ) );
  AN2D0 U5215 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [14]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ) );
  AN2D0 U5216 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [13]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N66 ) );
  AN2D0 U5217 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [12]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ) );
  AN2D0 U5218 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [11]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N64 ) );
  AN2D0 U5219 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [10]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ) );
  AN2D0 U5220 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [9]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N62 ) );
  AN2D0 U5221 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [8]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ) );
  AN2D0 U5222 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [7]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N60 ) );
  AN2D0 U5223 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [6]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ) );
  AN2D0 U5224 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [5]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N58 ) );
  AN2D0 U5225 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [4]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ) );
  AN2D0 U5226 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [3]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N56 ) );
  AN2D0 U5227 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [2]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ) );
  AN2D0 U5228 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [1]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N54 ) );
  AN2D0 U5229 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr [0]), .A2(
        n3580), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ) );
  OAI31D0 U5230 ( .A1(n5053), .A2(n5054), .A3(n5055), .B(n5056), .ZN(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 ) );
  OAI21D0 U5231 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ), .A2(n5057), .B(n5058), .ZN(n5056) );
  MUX2ND0 U5232 ( .I0(n5059), .I1(n5060), .S(n5057), .ZN(n5058) );
  MUX3ND0 U5233 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ), .I1(n5061), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N24 ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .S1(n5062), .ZN(n5060) );
  NR2D0 U5234 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .ZN(n5062) );
  MUX2D0 U5235 ( .I0(n5063), .I1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N26 ), .S(n5054), 
        .Z(n5061) );
  AN2D0 U5236 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ), .A2(n5055), .Z(n5063)
         );
  IND2D0 U5237 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .B1(n5055), .ZN(
        n5057) );
  CKND0 U5238 ( .CLK(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), .CN(n5055) );
  OAI21D0 U5239 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .B(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .ZN(n5054) );
  MUX2ND0 U5240 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N28 ), .S(n5059), .ZN(n5053) );
  CKND0 U5241 ( .CLK(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .CN(n5059) );
  CKND0 U5242 ( .CLK(ClockA), .CN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U5243 ( .A1(n4699), .A2(n4704), .A3(n1010), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ) );
  OAI21D0 U5244 ( .A1(n4723), .A2(n5064), .B(n5065), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ) );
  MUX2ND0 U5245 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .I1(n5066), 
        .S(n4704), .ZN(n5065) );
  NR2D0 U5246 ( .A1(n1010), .A2(n4768), .ZN(n5066) );
  CKND0 U5247 ( .CLK(n4720), .CN(n4768) );
  OAI21D0 U5248 ( .A1(n4764), .A2(n4754), .B(n4747), .ZN(n4720) );
  CKND0 U5249 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .CN(n4754)
         );
  OAI21D0 U5250 ( .A1(n4745), .A2(n5064), .B(n5067), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ) );
  MUX2ND0 U5251 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .I1(n5068), 
        .S(n4704), .ZN(n5067) );
  NR2D0 U5252 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n5069), 
        .ZN(n5068) );
  OAI21D0 U5253 ( .A1(n4704), .A2(n4499), .B(n5064), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ) );
  CKND2D0 U5254 ( .A1(n5070), .A2(n4704), .ZN(n5064) );
  CKND2D0 U5255 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A2(
        n4707), .ZN(n4704) );
  NR2D0 U5256 ( .A1(n4716), .A2(n4719), .ZN(n4707) );
  NR2D0 U5257 ( .A1(n4742), .A2(n4728), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ) );
  XNR2D0 U5258 ( .A1(n4501), .A2(n5071), .ZN(n4742) );
  CKND2D0 U5259 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n5071) );
  CKND2D0 U5260 ( .A1(n1015), .A2(n4699), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ) );
  CKND0 U5261 ( .CLK(n4710), .CN(n4699) );
  MUX2ND0 U5262 ( .I0(n5072), .I1(n5073), .S(n4500), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ) );
  CKND2D0 U5263 ( .A1(n5074), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(n5073) );
  CKND0 U5264 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ), .CN(n5072) );
  NR2D0 U5265 ( .A1(n4728), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ) );
  CKND0 U5266 ( .CLK(n5074), .CN(n4728) );
  NR2D0 U5267 ( .A1(n4710), .A2(n1015), .ZN(n5074) );
  NR2D0 U5268 ( .A1(n4702), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .ZN(n4710) );
  CKND2D0 U5269 ( .A1(n4716), .A2(n4719), .ZN(n4702) );
  CKND0 U5270 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .CN(
        n4719) );
  CKND0 U5271 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .CN(
        n4716) );
  NR3D0 U5272 ( .A1(n5075), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ) );
  NR3D0 U5273 ( .A1(n5069), .A2(n4723), .A3(n4745), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ) );
  NR3D0 U5274 ( .A1(n5075), .A2(n4723), .A3(n4745), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ) );
  CKND2D0 U5275 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n4745), 
        .ZN(n4747) );
  CKND0 U5276 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .CN(n4745)
         );
  CKND0 U5277 ( .CLK(n5070), .CN(n5075) );
  NR2D0 U5278 ( .A1(n1010), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n5070) );
  CKND2D0 U5279 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n4723), 
        .ZN(n4764) );
  CKND0 U5280 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .CN(n4723)
         );
  NR3D0 U5281 ( .A1(n5069), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ) );
  IND2D0 U5282 ( .A1(n1010), .B1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n5069) );
  AO22D0 U5283 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ), .A2(
        n4793), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ), .B2(n4789), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ) );
  MUX2ND0 U5284 ( .I0(n5076), .I1(n5077), .S(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .ZN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ) );
  CKND2D0 U5285 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        n4790), .ZN(n5077) );
  ND3D0 U5286 ( .A1(n5078), .A2(n4792), .A3(n5079), .ZN(n4790) );
  ND4D0 U5287 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .ZN(n5079) );
  IND3D0 U5288 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .B1(
        n4792), .B2(n4791), .ZN(n5076) );
  CKND2D0 U5289 ( .A1(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n4791) );
  AO22D0 U5290 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ), .A2(
        n4793), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ), .B2(n4789), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ) );
  AO22D0 U5291 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ), .A2(
        n4793), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ), .B2(n4789), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ) );
  AN2D0 U5292 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .Z(n4789) );
  NR2D0 U5293 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .ZN(n4793) );
  AN2D0 U5294 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ), .A2(n4782), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ) );
  AN2D0 U5295 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ), .A2(n4782), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ) );
  AN2D0 U5296 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ), .A2(n4782), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ) );
  AN2D0 U5297 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ), .A2(n4782), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ) );
  AN2D0 U5298 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ), .A2(n4782), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ) );
  AN2D0 U5299 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ), .A2(n4782), 
        .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ) );
  OAI21D0 U5300 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), 
        .A2(n4792), .B(n5080), .ZN(n4782) );
  IOA22D0 U5301 ( .B1(n5081), .B2(n5082), .A1(n4792), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .ZN(n5080)
         );
  AOI221D0 U5302 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .A2(n5078), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .B2(n5083), .C(n5084), .ZN(n5082) );
  AOI221D0 U5303 ( .A1(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(n5085), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B2(n5086), 
        .C(n5087), .ZN(n5084) );
  IAO21D0 U5304 ( .A1(n5086), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .ZN(n5087)
         );
  OAI32D0 U5305 ( .A1(n5088), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .A3(n5089), 
        .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .B2(
        n5090), .ZN(n5086) );
  AN2D0 U5306 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), 
        .A2(n5090), .Z(n5089) );
  CKND0 U5307 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .CN(n5090) );
  CKND0 U5308 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .CN(n5088) );
  CKND0 U5309 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .CN(n5085) );
  CKND0 U5310 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .CN(n5083) );
  NR2D0 U5311 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), 
        .A2(n5078), .ZN(n5081) );
  CKND0 U5312 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .CN(n5078) );
  CKND0 U5313 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .CN(n4792) );
  AN2D0 U5314 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]), .A2(
        n4440), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ) );
  CKXOR2D0 U5315 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ) );
  XNR2D0 U5316 ( .A1(n5091), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ) );
  AO221D0 U5317 ( .A1(n5092), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .B1(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), .B2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .C(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ) );
  NR2D0 U5318 ( .A1(n5091), .A2(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .ZN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ) );
  CKND0 U5319 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ) );
  IOA21D0 U5320 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .B(n5091), 
        .ZN(n5092) );
  CKND0 U5321 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .CN(n5091) );
  CKND2D0 U5322 ( .A1(\SerDes_U1/Rx_ParClk ), .A2(ClockB), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U5323 ( .A1(n5093), .A2(n4858), .A3(n4850), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ) );
  OAI22D0 U5324 ( .A1(n4563), .A2(n4858), .B1(n4862), .B2(n4850), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ) );
  OA211D0 U5325 ( .A1(n5094), .A2(n4812), .B(n5095), .C(n4832), .Z(n4862) );
  OAI22D0 U5326 ( .A1(n4562), .A2(n4858), .B1(n4864), .B2(n4850), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ) );
  XNR2D0 U5327 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n5094), 
        .ZN(n4864) );
  OAI22D0 U5328 ( .A1(n4561), .A2(n4858), .B1(n4863), .B2(n4850), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ) );
  AN2D0 U5329 ( .A1(n5096), .A2(n5097), .Z(n4863) );
  OAI22D0 U5330 ( .A1(n4560), .A2(n4858), .B1(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .B2(n4850), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ) );
  CKND2D0 U5331 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .A2(n4858), 
        .ZN(n4850) );
  CKND2D0 U5332 ( .A1(n4827), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .ZN(n4858) );
  CKND0 U5333 ( .CLK(n4802), .CN(n4827) );
  CKND2D0 U5334 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .ZN(n4802) );
  NR2D0 U5335 ( .A1(n4844), .A2(n5098), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ) );
  XNR2D0 U5336 ( .A1(n5099), .A2(n4563), .ZN(n4844) );
  CKND2D0 U5337 ( .A1(n5093), .A2(n5098), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ) );
  CKND0 U5338 ( .CLK(n4799), .CN(n5093) );
  NR2D0 U5339 ( .A1(n4845), .A2(n5098), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ) );
  OAI21D0 U5340 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .A2(n5100), 
        .B(n5099), .ZN(n4845) );
  CKND2D0 U5341 ( .A1(n5100), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), 
        .ZN(n5099) );
  NR2D0 U5342 ( .A1(n4560), .A2(n4561), .ZN(n5100) );
  MUX2ND0 U5343 ( .I0(n5101), .I1(n5102), .S(n4561), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ) );
  CKND2D0 U5344 ( .A1(n5103), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), 
        .ZN(n5102) );
  CKND0 U5345 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .CN(n5101) );
  NR2D0 U5346 ( .A1(n5098), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), 
        .ZN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ) );
  CKND0 U5347 ( .CLK(n5103), .CN(n5098) );
  NR2D0 U5348 ( .A1(n869), .A2(n4799), .ZN(n5103) );
  NR3D0 U5349 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[2] ), .ZN(n4799) );
  ND3D0 U5350 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), .A3(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .ZN(n5105) );
  OR2D0 U5351 ( .A1(n4832), .A2(n863), .Z(n5107) );
  CKND2D0 U5352 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .A2(n4846), 
        .ZN(n4832) );
  ND3D0 U5353 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n4812), 
        .A3(n5094), .ZN(n5095) );
  ND3D0 U5354 ( .A1(n4812), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), 
        .A3(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .ZN(n5108) );
  CKND0 U5355 ( .CLK(n5094), .CN(n5104) );
  NR2D0 U5356 ( .A1(n4842), .A2(n4854), .ZN(n5094) );
  CKND2D0 U5357 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n4842), 
        .ZN(n5097) );
  CKND2D0 U5358 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .A2(n4854), 
        .ZN(n5096) );
  ND3D0 U5359 ( .A1(n4812), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_MemWriteCmd ), 
        .A3(n4846), .ZN(n5109) );
  CKND0 U5360 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .CN(n4846)
         );
  CKND0 U5361 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .CN(n4812)
         );
  CKND2D0 U5362 ( .A1(n4842), .A2(n4854), .ZN(n5106) );
  CKND0 U5363 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .CN(n4854)
         );
  CKND0 U5364 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .CN(n4842)
         );
  NR2D0 U5365 ( .A1(n5110), .A2(n5111), .ZN(\SerDes_U1/Des_U1/DesDec_Rx1/N47 )
         );
  CKND2D0 U5366 ( .A1(n5112), .A2(n5113), .ZN(n5111) );
  NR4D0 U5367 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ), .ZN(n5113) );
  NR4D0 U5368 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ), .ZN(n5112) );
  AN4D0 U5369 ( .A1(n5114), .A2(n5115), .A3(n5116), .A4(n5117), .Z(n5110) );
  NR4D0 U5370 ( .A1(n5118), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ), 
        .A3(n1003), .A4(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ), .ZN(n5117)
         );
  ND3D0 U5371 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ), .ZN(n5118) );
  NR4D0 U5372 ( .A1(n5119), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ), .ZN(n5116) );
  ND3D0 U5373 ( .A1(n989), .A2(n985), .A3(n990), .ZN(n5119) );
  NR4D0 U5374 ( .A1(n5120), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ), .ZN(n5115) );
  ND3D0 U5375 ( .A1(n4611), .A2(n997), .A3(n4612), .ZN(n5120) );
  NR4D0 U5376 ( .A1(n5121), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ), .ZN(n5114) );
  ND3D0 U5377 ( .A1(n4614), .A2(n4613), .A3(n4615), .ZN(n5121) );
  OA21D0 U5378 ( .A1(n5122), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .B(
        \SerDes_U1/SerLineValid ), .Z(\SerDes_U1/Des_U1/DesDec_Rx1/N43 ) );
  NR4D0 U5379 ( .A1(n5123), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ), .ZN(n5122) );
  OR2D0 U5380 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ), .Z(n5123) );
  INR2D0 U5381 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N34 ), .B1(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N42 ) );
  INR2D0 U5382 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N33 ), .B1(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N41 ) );
  INR2D0 U5383 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N32 ), .B1(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N40 ) );
  INR2D0 U5384 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N31 ), .B1(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N39 ) );
  INR2D0 U5385 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N30 ), .B1(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N38 ) );
  NR2D0 U5386 ( .A1(\SerDes_U1/Rx_ParClk ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/doParSync ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N37 ) );
endmodule


module FullDup_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_4 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_5 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_6 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_7 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_8 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_9 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_3 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_10 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_11 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_12 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_13 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_4 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_5 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

