library verilog;
use verilog.vl_types.all;
entity uart_byte_rx_tb is
end uart_byte_rx_tb;
