/* Copyright Cadence Design Systems (c) 2015  */

package clock_and_reset_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "clock_and_reset.svh"

endpackage
