// =============================================
// Level4.  Lab problem in parameter passing
// by `define.
//
// 2006-06-07 jmw:  v. 1.1 Fixed Wid4 typo.
// 2005-02-02 jmw:  v. 1.0 completed.
// =============================================
`define Wid    4
//
module Level4 (inout[`Wid-1:0] DataB, input[3:0] Ctl, input Clk) ;
  always@(negedge Clk)
    ...
endmodule

