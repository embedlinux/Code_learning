
`ifndef RKV_I2C_DEFINES_SVH
`define RKV_I2C_DEFINES_SVH

parameter IC_INTR_NUM          = 12; 
parameter IC_RX_OVER_INTR_ID   = 0 ;  
parameter IC_RX_UNDER_INTR_ID  = 1 ;    
parameter IC_TX_OVER_INTR_ID   = 2 ;  
parameter IC_TX_ABRT_INTR_ID   = 3 ;  
parameter IC_RX_DONE_INTR_ID   = 4 ;  
parameter IC_TX_EMPTY_INTR_ID  = 5 ;  
parameter IC_ACTIVITY_INTR_ID  = 6 ;  
parameter IC_STOP_DET_INTR_ID  = 7 ;  
parameter IC_START_DET_INTR_ID = 8 ;  
parameter IC_RD_REQ_INTR_ID    = 9 ;  
parameter IC_RX_FULL_INTR_ID   = 10;  
parameter IC_GEN_CALL_INTR_ID  = 11;  



`endif // RKV_I2C_DEFINES_SVH
