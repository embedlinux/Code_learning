
module rr16 ( clk, rst, aw, ar, d, wr_n, full, do_m );
input  [3:0] aw;
input  [3:0] ar;
input  [7:0] d;
output [7:0] do_m;
input  clk, rst, wr_n, full;
    wire \re0[7] , \re0[6] , \re0[5] , \re0[4] , \re0[3] , \re0[2] , \re0[1] , 
        \re0[0] , \re1[7] , \re1[6] , \re1[5] , \re1[4] , \re1[3] , \re1[2] , 
        \re1[1] , \re1[0] , \re2[7] , \re2[6] , \re2[5] , \re2[4] , \re2[3] , 
        \re2[2] , \re2[1] , \re2[0] , \re3[7] , \re3[6] , \re3[5] , \re3[4] , 
        \re3[3] , \re3[2] , \re3[1] , \re3[0] , \re4[7] , \re4[6] , \re4[5] , 
        \re4[4] , \re4[3] , \re4[2] , \re4[1] , \re4[0] , \re5[7] , \re5[6] , 
        \re5[5] , \re5[4] , \re5[3] , \re5[2] , \re5[1] , \re5[0] , \re6[7] , 
        \re6[6] , \re6[5] , \re6[4] , \re6[3] , \re6[2] , \re6[1] , \re6[0] , 
        \re7[7] , \re7[6] , \re7[5] , \re7[4] , \re7[3] , \re7[2] , \re7[1] , 
        \re7[0] , \re8[7] , \re8[6] , \re8[5] , \re8[4] , \re8[3] , \re8[2] , 
        \re8[1] , \re8[0] , \re9[7] , \re9[6] , \re9[5] , \re9[4] , \re9[3] , 
        \re9[2] , \re9[1] , \re9[0] , \re10[7] , \re10[6] , \re10[5] , 
        \re10[4] , \re10[3] , \re10[2] , \re10[1] , \re10[0] , \re11[7] , 
        \re11[6] , \re11[5] , \re11[4] , \re11[3] , \re11[2] , \re11[1] , 
        \re11[0] , \re12[7] , \re12[6] , \re12[5] , \re12[4] , \re12[3] , 
        \re12[2] , \re12[1] , \re12[0] , \re13[7] , \re13[6] , \re13[5] , 
        \re13[4] , \re13[3] , \re13[2] , \re13[1] , \re13[0] , \re14[7] , 
        \re14[6] , \re14[5] , \re14[4] , \re14[3] , \re14[2] , \re14[1] , 
        \re14[0] , \re15[7] , \re15[6] , \re15[5] , \re15[4] , \re15[3] , 
        \re15[2] , \re15[1] , \re15[0] , n34, n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
        n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
        n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
        n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
        n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
        n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
        n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
        n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
        n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
        n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
        n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
        n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
        n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
        n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
        n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
        n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
        n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
        n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
        n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
        n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
        n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
        n373, n374;
    OR3P U2 ( .O(n34), .I1(aw[3]), .I2(n342), .I3(n343) );
    AN2B1P U3 ( .O(n105), .I1(ar[0]), .B1(ar[1]) );
    ND4 U4 ( .O(do_m[7]), .I1(n354), .I2(n351), .I3(n313), .I4(n314) );
    ND4 U5 ( .O(do_m[3]), .I1(n368), .I2(n367), .I3(n321), .I4(n322) );
    ND4 U6 ( .O(do_m[2]), .I1(n370), .I2(n369), .I3(n323), .I4(n324) );
    ND4 U7 ( .O(do_m[4]), .I1(n366), .I2(n365), .I3(n319), .I4(n320) );
    ND4 U8 ( .O(do_m[1]), .I1(n372), .I2(n371), .I3(n325), .I4(n326) );
    ND4 U9 ( .O(do_m[5]), .I1(n364), .I2(n363), .I3(n317), .I4(n318) );
    ND4 U10 ( .O(do_m[0]), .I1(n374), .I2(n373), .I3(n327), .I4(n328) );
    ND4 U11 ( .O(do_m[6]), .I1(n362), .I2(n361), .I3(n315), .I4(n316) );
    AN2P U12 ( .O(n101), .I1(ar[2]), .I2(ar[3]) );
    AN2 U13 ( .O(n66), .I1(ar[3]), .I2(n85) );
    AN2 U14 ( .O(n103), .I1(ar[2]), .I2(ar[3]) );
    AN2 U15 ( .O(n65), .I1(ar[2]), .I2(n329) );
    AN2 U16 ( .O(n95), .I1(aw[1]), .I2(n346) );
    AN2 U17 ( .O(n89), .I1(n346), .I2(n341) );
    OR2P U18 ( .O(n333), .I1(n100), .I2(n35) );
    INV2 U19 ( .O(n35), .I(n101) );
    OR2P U20 ( .O(n336), .I1(n36), .I2(n100) );
    INV2 U21 ( .O(n36), .I(n96) );
    OR2P U22 ( .O(n332), .I1(ar[1]), .I2(ar[0]) );
    BUF2 U23 ( .O(n96), .I(n66) );
    INV2 U24 ( .O(n100), .I(n334) );
    INV1 U25 ( .O(n330), .I(ar[0]) );
    OR2P U26 ( .O(n337), .I1(n39), .I2(n37) );
    INV2 U27 ( .O(n37), .I(n98) );
    BUF3 U28 ( .O(n98), .I(n104) );
    BUF2 U29 ( .O(n97), .I(n65) );
    OR2P U30 ( .O(n340), .I1(n38), .I2(n332) );
    INV2 U31 ( .O(n38), .I(n84) );
    OR2P U32 ( .O(n338), .I1(n39), .I2(n332) );
    INV2 U33 ( .O(n39), .I(n97) );
    INV2 U34 ( .O(n334), .I(n332) );
    INV2 U35 ( .O(n345), .I(n343) );
    AN2 U36 ( .O(n40), .I1(aw[0]), .I2(n341) );
    INV2 U37 ( .O(n347), .I(n40) );
    AN2 U38 ( .O(n41), .I1(aw[0]), .I2(aw[1]) );
    INV2 U39 ( .O(n349), .I(n41) );
    OR2P U40 ( .O(n343), .I1(full), .I2(wr_n) );
    OR2 U41 ( .O(n183), .I1(n344), .I2(n90) );
    INV2 U42 ( .O(n179), .I(n90) );
    INV2 U43 ( .O(n90), .I(n89) );
    INV2 U44 ( .O(n178), .I(n344) );
    INV2 U45 ( .O(n184), .I(rst) );
    BUF2 U46 ( .O(n169), .I(n175) );
    AN2P U47 ( .O(n67), .I1(n329), .I2(n85) );
    INV2 U48 ( .O(n329), .I(ar[3]) );
    AN2P U49 ( .O(n102), .I1(ar[0]), .I2(ar[1]) );
    BUF3 U50 ( .O(n114), .I(n57) );
    INV2 U51 ( .O(n85), .I(ar[2]) );
    AN2P U52 ( .O(n109), .I1(ar[0]), .I2(ar[1]) );
    BUF3 U53 ( .O(n112), .I(n59) );
    BUF3 U54 ( .O(n111), .I(n60) );
    BUF3 U55 ( .O(n113), .I(n58) );
    BUF2 U56 ( .O(n99), .I(n105) );
    OR3B2P U57 ( .O(n348), .I1(aw[2]), .B1(aw[3]), .B2(n345) );
    OR3B2P U58 ( .O(n350), .I1(aw[3]), .B1(n342), .B2(n345) );
    INV2 U59 ( .O(n341), .I(aw[1]) );
    OR3B2P U60 ( .O(n344), .I1(n342), .B1(aw[3]), .B2(n345) );
    BUF3 U61 ( .O(n127), .I(n44) );
    BUF3 U62 ( .O(n128), .I(n43) );
    BUF3 U63 ( .O(n126), .I(n45) );
    BUF3 U64 ( .O(n120), .I(n51) );
    BUF3 U65 ( .O(n125), .I(n46) );
    BUF3 U66 ( .O(n117), .I(n54) );
    INV3 U67 ( .O(n180), .I(n348) );
    BUF3 U68 ( .O(n123), .I(n48) );
    BUF3 U69 ( .O(n119), .I(n52) );
    BUF3 U70 ( .O(n121), .I(n50) );
    BUF3 U71 ( .O(n115), .I(n56) );
    INV3 U72 ( .O(n181), .I(n34) );
    BUF3 U73 ( .O(n122), .I(n49) );
    BUF3 U74 ( .O(n118), .I(n53) );
    INV3 U75 ( .O(n94), .I(n93) );
    INV2 U76 ( .O(n93), .I(n95) );
    BUF3 U77 ( .O(n124), .I(n47) );
    INV3 U78 ( .O(n92), .I(n347) );
    BUF3 U79 ( .O(n116), .I(n55) );
    INV3 U80 ( .O(n182), .I(n350) );
    BUF3 U81 ( .O(n129), .I(n42) );
    INV3 U82 ( .O(n91), .I(n349) );
    AN2T U83 ( .O(n42), .I1(n178), .I2(n91) );
    AN2T U84 ( .O(n43), .I1(n178), .I2(n92) );
    AN2T U85 ( .O(n44), .I1(n178), .I2(n94) );
    AN2T U86 ( .O(n45), .I1(n91), .I2(n180) );
    AN2T U87 ( .O(n46), .I1(n92), .I2(n180) );
    AN2T U88 ( .O(n47), .I1(n92), .I2(n182) );
    AN2T U89 ( .O(n48), .I1(n91), .I2(n181) );
    AN2T U90 ( .O(n49), .I1(n91), .I2(n182) );
    AN2T U91 ( .O(n50), .I1(n92), .I2(n181) );
    AN2T U92 ( .O(n51), .I1(n94), .I2(n180) );
    AN2T U93 ( .O(n52), .I1(n94), .I2(n181) );
    AN2T U94 ( .O(n53), .I1(n94), .I2(n182) );
    AN2T U95 ( .O(n54), .I1(n179), .I2(n180) );
    AN2T U96 ( .O(n55), .I1(n179), .I2(n182) );
    AN2T U97 ( .O(n56), .I1(n179), .I2(n181) );
    AN2T U98 ( .O(n57), .I1(n103), .I2(n109) );
    AN2T U99 ( .O(n58), .I1(n97), .I2(n102) );
    AN2T U100 ( .O(n59), .I1(n96), .I2(n109) );
    AN2T U101 ( .O(n60), .I1(n67), .I2(n102) );
    AN2 U102 ( .O(n61), .I1(n99), .I2(n103) );
    AN2 U103 ( .O(n62), .I1(n65), .I2(n105) );
    AN2 U104 ( .O(n63), .I1(n66), .I2(n99) );
    AN2 U105 ( .O(n64), .I1(n67), .I2(n99) );
    AN2 U106 ( .O(n104), .I1(ar[1]), .I2(n330) );
    BUF2 U107 ( .O(n176), .I(n177) );
    BUF4 U108 ( .O(n172), .I(n174) );
    BUF4 U109 ( .O(n165), .I(n169) );
    BUF1 U110 ( .O(n177), .I(n184) );
    BUF2 U111 ( .O(n174), .I(n176) );
    BUF2 U112 ( .O(n175), .I(n176) );
    BUF2 U113 ( .O(n166), .I(n184) );
    BUF2 U114 ( .O(n167), .I(n175) );
    BUF2 U115 ( .O(n168), .I(n175) );
    BUF2 U116 ( .O(n170), .I(n166) );
    BUF2 U117 ( .O(n171), .I(n174) );
    BUF2 U118 ( .O(n173), .I(n177) );
    INV1 U119 ( .O(n346), .I(aw[0]) );
    BUF4 U120 ( .O(n68), .I(d[6]) );
    BUF4 U121 ( .O(n69), .I(d[6]) );
    BUF4 U122 ( .O(n70), .I(d[2]) );
    BUF4 U123 ( .O(n71), .I(d[2]) );
    BUF4 U124 ( .O(n72), .I(d[1]) );
    BUF4 U125 ( .O(n73), .I(d[1]) );
    BUF4 U126 ( .O(n74), .I(d[5]) );
    BUF4 U127 ( .O(n75), .I(d[5]) );
    BUF4 U128 ( .O(n76), .I(d[7]) );
    BUF4 U129 ( .O(n77), .I(d[7]) );
    BUF4 U130 ( .O(n78), .I(d[3]) );
    BUF4 U131 ( .O(n79), .I(d[3]) );
    BUF4 U132 ( .O(n80), .I(d[0]) );
    BUF4 U133 ( .O(n81), .I(d[0]) );
    BUF4 U134 ( .O(n82), .I(d[4]) );
    BUF4 U135 ( .O(n83), .I(d[4]) );
    BUF2 U136 ( .O(n84), .I(n67) );
    MUX2 U137 ( .O(n242), .S(n48), .A(\re7[1] ), .B(n72) );
    MUX2 U138 ( .O(n250), .S(n52), .A(\re6[1] ), .B(n72) );
    MUX2 U139 ( .O(n234), .S(n54), .A(\re8[1] ), .B(n72) );
    MUX2 U140 ( .O(n258), .S(n50), .A(\re5[1] ), .B(n73) );
    MUX2 U141 ( .O(n226), .S(n46), .A(\re9[1] ), .B(n72) );
    MUX2 U142 ( .O(n266), .S(n56), .A(\re4[1] ), .B(n73) );
    MUX2 U143 ( .O(n218), .S(n51), .A(\re10[1] ), .B(n72) );
    MUX2 U144 ( .O(n274), .S(n49), .A(\re3[1] ), .B(n73) );
    MUX2 U145 ( .O(n210), .S(n45), .A(\re11[1] ), .B(n73) );
    MUX2 U146 ( .O(n282), .S(n53), .A(\re2[1] ), .B(n72) );
    MUX2 U147 ( .O(n202), .S(n131), .A(\re12[1] ), .B(n72) );
    MUX2 U148 ( .O(n290), .S(n47), .A(\re1[1] ), .B(n73) );
    MUX2 U149 ( .O(n194), .S(n43), .A(\re13[1] ), .B(n73) );
    MUX2 U150 ( .O(n298), .S(n55), .A(\re0[1] ), .B(n73) );
    MUX2 U151 ( .O(n186), .S(n44), .A(\re14[1] ), .B(n72) );
    MUX2 U152 ( .O(n306), .S(n42), .A(\re15[1] ), .B(n73) );
    MUX2 U153 ( .O(n245), .S(n48), .A(\re7[4] ), .B(n82) );
    MUX2 U154 ( .O(n253), .S(n52), .A(\re6[4] ), .B(n82) );
    MUX2 U155 ( .O(n237), .S(n54), .A(\re8[4] ), .B(n82) );
    MUX2 U156 ( .O(n261), .S(n50), .A(\re5[4] ), .B(n83) );
    MUX2 U157 ( .O(n229), .S(n46), .A(\re9[4] ), .B(n82) );
    MUX2 U158 ( .O(n269), .S(n56), .A(\re4[4] ), .B(n83) );
    MUX2 U159 ( .O(n221), .S(n51), .A(\re10[4] ), .B(n82) );
    MUX2 U160 ( .O(n277), .S(n49), .A(\re3[4] ), .B(n83) );
    MUX2 U161 ( .O(n213), .S(n45), .A(\re11[4] ), .B(n83) );
    MUX2 U162 ( .O(n285), .S(n53), .A(\re2[4] ), .B(n82) );
    MUX2 U163 ( .O(n205), .S(n131), .A(\re12[4] ), .B(n82) );
    MUX2 U164 ( .O(n293), .S(n47), .A(\re1[4] ), .B(n83) );
    MUX2 U165 ( .O(n197), .S(n43), .A(\re13[4] ), .B(n83) );
    MUX2 U166 ( .O(n301), .S(n55), .A(\re0[4] ), .B(n83) );
    MUX2 U167 ( .O(n189), .S(n44), .A(\re14[4] ), .B(n82) );
    MUX2 U168 ( .O(n309), .S(n42), .A(\re15[4] ), .B(n83) );
    BUF2 U169 ( .O(n86), .I(n339) );
    ND2 U170 ( .O(n339), .I1(n84), .I2(n98) );
    BUF2 U171 ( .O(n87), .I(n335) );
    ND2 U172 ( .O(n335), .I1(n96), .I2(n98) );
    BUF2 U173 ( .O(n88), .I(n331) );
    ND2 U174 ( .O(n331), .I1(n98), .I2(n101) );
    INV4 U175 ( .O(n360), .I(n340) );
    INV4 U176 ( .O(n359), .I(n86) );
    INV4 U177 ( .O(n356), .I(n336) );
    INV4 U178 ( .O(n353), .I(n333) );
    INV4 U179 ( .O(n355), .I(n87) );
    INV4 U180 ( .O(n352), .I(n88) );
    INV4 U181 ( .O(n358), .I(n338) );
    INV4 U182 ( .O(n357), .I(n337) );
    BUF4 U183 ( .O(n106), .I(n64) );
    BUF4 U184 ( .O(n107), .I(n63) );
    BUF4 U185 ( .O(n108), .I(n62) );
    BUF4 U186 ( .O(n110), .I(n61) );
    MUX2 U187 ( .O(n271), .S(n115), .A(\re4[6] ), .B(n68) );
    MUX2 U188 ( .O(n267), .S(n115), .A(\re4[2] ), .B(n70) );
    MUX2 U189 ( .O(n272), .S(n115), .A(\re4[7] ), .B(n76) );
    MUX2 U190 ( .O(n270), .S(n115), .A(\re4[5] ), .B(n74) );
    MUX2 U191 ( .O(n265), .S(n115), .A(\re4[0] ), .B(n80) );
    MUX2 U192 ( .O(n268), .S(n56), .A(\re4[3] ), .B(n78) );
    MUX2 U193 ( .O(n303), .S(n116), .A(\re0[6] ), .B(n68) );
    MUX2 U194 ( .O(n299), .S(n116), .A(\re0[2] ), .B(n70) );
    MUX2 U195 ( .O(n304), .S(n116), .A(\re0[7] ), .B(n76) );
    MUX2 U196 ( .O(n302), .S(n116), .A(\re0[5] ), .B(n74) );
    MUX2 U197 ( .O(n297), .S(n116), .A(\re0[0] ), .B(n80) );
    MUX2 U198 ( .O(n300), .S(n55), .A(\re0[3] ), .B(n78) );
    MUX2 U199 ( .O(n239), .S(n117), .A(\re8[6] ), .B(n68) );
    MUX2 U200 ( .O(n235), .S(n117), .A(\re8[2] ), .B(n70) );
    MUX2 U201 ( .O(n240), .S(n117), .A(\re8[7] ), .B(n76) );
    MUX2 U202 ( .O(n238), .S(n117), .A(\re8[5] ), .B(n74) );
    MUX2 U203 ( .O(n233), .S(n117), .A(\re8[0] ), .B(n80) );
    MUX2 U204 ( .O(n236), .S(n54), .A(\re8[3] ), .B(n78) );
    MUX2 U205 ( .O(n287), .S(n118), .A(\re2[6] ), .B(n69) );
    MUX2 U206 ( .O(n283), .S(n118), .A(\re2[2] ), .B(n71) );
    MUX2 U207 ( .O(n288), .S(n118), .A(\re2[7] ), .B(n77) );
    MUX2 U208 ( .O(n286), .S(n118), .A(\re2[5] ), .B(n75) );
    MUX2 U209 ( .O(n281), .S(n118), .A(\re2[0] ), .B(n81) );
    MUX2 U210 ( .O(n284), .S(n53), .A(\re2[3] ), .B(n79) );
    MUX2 U211 ( .O(n255), .S(n119), .A(\re6[6] ), .B(n68) );
    MUX2 U212 ( .O(n251), .S(n119), .A(\re6[2] ), .B(n70) );
    MUX2 U213 ( .O(n256), .S(n119), .A(\re6[7] ), .B(n76) );
    MUX2 U214 ( .O(n254), .S(n119), .A(\re6[5] ), .B(n74) );
    MUX2 U215 ( .O(n249), .S(n119), .A(\re6[0] ), .B(n80) );
    MUX2 U216 ( .O(n252), .S(n52), .A(\re6[3] ), .B(n78) );
    MUX2 U217 ( .O(n223), .S(n120), .A(\re10[6] ), .B(n69) );
    MUX2 U218 ( .O(n219), .S(n120), .A(\re10[2] ), .B(n71) );
    MUX2 U219 ( .O(n224), .S(n120), .A(\re10[7] ), .B(n77) );
    MUX2 U220 ( .O(n222), .S(n120), .A(\re10[5] ), .B(n75) );
    MUX2 U221 ( .O(n217), .S(n120), .A(\re10[0] ), .B(n81) );
    MUX2 U222 ( .O(n220), .S(n51), .A(\re10[3] ), .B(n79) );
    MUX2 U223 ( .O(n263), .S(n121), .A(\re5[6] ), .B(n68) );
    MUX2 U224 ( .O(n259), .S(n121), .A(\re5[2] ), .B(n70) );
    MUX2 U225 ( .O(n264), .S(n121), .A(\re5[7] ), .B(n76) );
    MUX2 U226 ( .O(n262), .S(n121), .A(\re5[5] ), .B(n74) );
    MUX2 U227 ( .O(n257), .S(n121), .A(\re5[0] ), .B(n80) );
    MUX2 U228 ( .O(n260), .S(n50), .A(\re5[3] ), .B(n78) );
    MUX2 U229 ( .O(n279), .S(n122), .A(\re3[6] ), .B(n69) );
    MUX2 U230 ( .O(n275), .S(n122), .A(\re3[2] ), .B(n71) );
    MUX2 U231 ( .O(n280), .S(n122), .A(\re3[7] ), .B(n77) );
    MUX2 U232 ( .O(n278), .S(n122), .A(\re3[5] ), .B(n75) );
    MUX2 U233 ( .O(n273), .S(n122), .A(\re3[0] ), .B(n81) );
    MUX2 U234 ( .O(n276), .S(n49), .A(\re3[3] ), .B(n79) );
    MUX2 U235 ( .O(n247), .S(n123), .A(\re7[6] ), .B(n69) );
    MUX2 U236 ( .O(n243), .S(n123), .A(\re7[2] ), .B(n71) );
    MUX2 U237 ( .O(n248), .S(n123), .A(\re7[7] ), .B(n77) );
    MUX2 U238 ( .O(n246), .S(n123), .A(\re7[5] ), .B(n75) );
    MUX2 U239 ( .O(n241), .S(n123), .A(\re7[0] ), .B(n81) );
    MUX2 U240 ( .O(n244), .S(n48), .A(\re7[3] ), .B(n79) );
    MUX2 U241 ( .O(n295), .S(n124), .A(\re1[6] ), .B(n68) );
    MUX2 U242 ( .O(n291), .S(n124), .A(\re1[2] ), .B(n70) );
    MUX2 U243 ( .O(n296), .S(n124), .A(\re1[7] ), .B(n76) );
    MUX2 U244 ( .O(n294), .S(n124), .A(\re1[5] ), .B(n74) );
    MUX2 U245 ( .O(n289), .S(n124), .A(\re1[0] ), .B(n80) );
    MUX2 U246 ( .O(n292), .S(n47), .A(\re1[3] ), .B(n78) );
    MUX2 U247 ( .O(n231), .S(n125), .A(\re9[6] ), .B(n68) );
    MUX2 U248 ( .O(n227), .S(n125), .A(\re9[2] ), .B(n70) );
    MUX2 U249 ( .O(n232), .S(n125), .A(\re9[7] ), .B(n76) );
    MUX2 U250 ( .O(n230), .S(n125), .A(\re9[5] ), .B(n74) );
    MUX2 U251 ( .O(n225), .S(n125), .A(\re9[0] ), .B(n80) );
    MUX2 U252 ( .O(n228), .S(n46), .A(\re9[3] ), .B(n78) );
    MUX2 U253 ( .O(n215), .S(n126), .A(\re11[6] ), .B(n69) );
    MUX2 U254 ( .O(n211), .S(n126), .A(\re11[2] ), .B(n71) );
    MUX2 U255 ( .O(n216), .S(n126), .A(\re11[7] ), .B(n77) );
    MUX2 U256 ( .O(n214), .S(n126), .A(\re11[5] ), .B(n75) );
    MUX2 U257 ( .O(n209), .S(n126), .A(\re11[0] ), .B(n81) );
    MUX2 U258 ( .O(n212), .S(n45), .A(\re11[3] ), .B(n79) );
    MUX2 U259 ( .O(n191), .S(n127), .A(\re14[6] ), .B(n69) );
    MUX2 U260 ( .O(n187), .S(n127), .A(\re14[2] ), .B(n71) );
    MUX2 U261 ( .O(n192), .S(n127), .A(\re14[7] ), .B(n77) );
    MUX2 U262 ( .O(n190), .S(n127), .A(\re14[5] ), .B(n75) );
    MUX2 U263 ( .O(n185), .S(n127), .A(\re14[0] ), .B(n81) );
    MUX2 U264 ( .O(n188), .S(n44), .A(\re14[3] ), .B(n79) );
    MUX2 U265 ( .O(n199), .S(n128), .A(\re13[6] ), .B(n69) );
    MUX2 U266 ( .O(n195), .S(n128), .A(\re13[2] ), .B(n71) );
    MUX2 U267 ( .O(n200), .S(n128), .A(\re13[7] ), .B(n77) );
    MUX2 U268 ( .O(n198), .S(n128), .A(\re13[5] ), .B(n75) );
    MUX2 U269 ( .O(n193), .S(n128), .A(\re13[0] ), .B(n81) );
    MUX2 U270 ( .O(n196), .S(n43), .A(\re13[3] ), .B(n79) );
    MUX2 U271 ( .O(n311), .S(n129), .A(\re15[6] ), .B(n68) );
    MUX2 U272 ( .O(n307), .S(n129), .A(\re15[2] ), .B(n70) );
    MUX2 U273 ( .O(n312), .S(n129), .A(\re15[7] ), .B(n76) );
    MUX2 U274 ( .O(n310), .S(n129), .A(\re15[5] ), .B(n74) );
    MUX2 U275 ( .O(n305), .S(n129), .A(\re15[0] ), .B(n80) );
    MUX2 U276 ( .O(n308), .S(n42), .A(\re15[3] ), .B(n78) );
    BUF3 U277 ( .O(n130), .I(n183) );
    INV2 U278 ( .O(n131), .I(n130) );
    INV4 U279 ( .O(n132), .I(n130) );
    MUX2 U280 ( .O(n207), .S(n132), .A(\re12[6] ), .B(n69) );
    MUX2 U281 ( .O(n203), .S(n132), .A(\re12[2] ), .B(n71) );
    MUX2 U282 ( .O(n208), .S(n132), .A(\re12[7] ), .B(n77) );
    MUX2 U283 ( .O(n206), .S(n132), .A(\re12[5] ), .B(n75) );
    MUX2 U284 ( .O(n201), .S(n132), .A(\re12[0] ), .B(n81) );
    MUX2 U285 ( .O(n204), .S(n132), .A(\re12[3] ), .B(n79) );
    BUF4 U286 ( .O(n133), .I(n171) );
    BUF4 U287 ( .O(n134), .I(n168) );
    BUF4 U288 ( .O(n135), .I(n184) );
    BUF4 U289 ( .O(n136), .I(n173) );
    BUF4 U290 ( .O(n137), .I(n173) );
    BUF4 U291 ( .O(n138), .I(n174) );
    BUF4 U292 ( .O(n139), .I(n167) );
    BUF4 U293 ( .O(n140), .I(n172) );
    BUF4 U294 ( .O(n141), .I(n172) );
    BUF4 U295 ( .O(n142), .I(n171) );
    BUF4 U296 ( .O(n143), .I(n171) );
    BUF4 U297 ( .O(n144), .I(n165) );
    BUF4 U298 ( .O(n145), .I(n165) );
    BUF4 U299 ( .O(n146), .I(n176) );
    BUF4 U300 ( .O(n147), .I(n165) );
    BUF4 U301 ( .O(n148), .I(n170) );
    BUF4 U302 ( .O(n149), .I(n170) );
    BUF4 U303 ( .O(n150), .I(n169) );
    BUF4 U304 ( .O(n151), .I(n169) );
    BUF4 U305 ( .O(n152), .I(n168) );
    BUF4 U306 ( .O(n153), .I(n168) );
    BUF4 U307 ( .O(n154), .I(n167) );
    BUF4 U308 ( .O(n155), .I(n167) );
    BUF4 U309 ( .O(n156), .I(n172) );
    BUF4 U310 ( .O(n157), .I(n172) );
    BUF4 U311 ( .O(n158), .I(n170) );
    BUF4 U312 ( .O(n159), .I(n173) );
    BUF4 U313 ( .O(n160), .I(n166) );
    BUF4 U314 ( .O(n161), .I(n166) );
    BUF4 U315 ( .O(n162), .I(n165) );
    BUF4 U316 ( .O(n163), .I(n165) );
    BUF4 U317 ( .O(n164), .I(n172) );
    DFFRBN \re14_reg[0]  ( .Q(\re14[0] ), .D(n185), .CK(clk), .RB(n153) );
    DFFRBN \re14_reg[1]  ( .Q(\re14[1] ), .D(n186), .CK(clk), .RB(n163) );
    DFFRBN \re14_reg[2]  ( .Q(\re14[2] ), .D(n187), .CK(clk), .RB(n153) );
    DFFRBN \re14_reg[3]  ( .Q(\re14[3] ), .D(n188), .CK(clk), .RB(n163) );
    DFFRBN \re14_reg[4]  ( .Q(\re14[4] ), .D(n189), .CK(clk), .RB(n154) );
    DFFRBN \re14_reg[5]  ( .Q(\re14[5] ), .D(n190), .CK(clk), .RB(n164) );
    DFFRBN \re14_reg[6]  ( .Q(\re14[6] ), .D(n191), .CK(clk), .RB(n154) );
    DFFRBN \re14_reg[7]  ( .Q(\re14[7] ), .D(n192), .CK(clk), .RB(n156) );
    DFFRBN \re13_reg[0]  ( .Q(\re13[0] ), .D(n193), .CK(clk), .RB(n155) );
    DFFRBN \re13_reg[1]  ( .Q(\re13[1] ), .D(n194), .CK(clk), .RB(n162) );
    DFFRBN \re13_reg[2]  ( .Q(\re13[2] ), .D(n195), .CK(clk), .RB(n155) );
    DFFRBN \re13_reg[3]  ( .Q(\re13[3] ), .D(n196), .CK(clk), .RB(n164) );
    DFFRBN \re13_reg[4]  ( .Q(\re13[4] ), .D(n197), .CK(clk), .RB(n155) );
    DFFRBN \re13_reg[5]  ( .Q(\re13[5] ), .D(n198), .CK(clk), .RB(n164) );
    DFFRBN \re13_reg[6]  ( .Q(\re13[6] ), .D(n199), .CK(clk), .RB(n153) );
    DFFRBN \re13_reg[7]  ( .Q(\re13[7] ), .D(n200), .CK(clk), .RB(n164) );
    DFFRBN \re12_reg[0]  ( .Q(\re12[0] ), .D(n201), .CK(clk), .RB(n147) );
    DFFRBN \re12_reg[1]  ( .Q(\re12[1] ), .D(n202), .CK(clk), .RB(n163) );
    DFFRBN \re12_reg[2]  ( .Q(\re12[2] ), .D(n203), .CK(clk), .RB(n155) );
    DFFRBN \re12_reg[3]  ( .Q(\re12[3] ), .D(n204), .CK(clk), .RB(n163) );
    DFFRBN \re12_reg[4]  ( .Q(\re12[4] ), .D(n205), .CK(clk), .RB(n154) );
    DFFRBN \re12_reg[5]  ( .Q(\re12[5] ), .D(n206), .CK(clk), .RB(n162) );
    DFFRBN \re12_reg[6]  ( .Q(\re12[6] ), .D(n207), .CK(clk), .RB(n154) );
    DFFRBN \re12_reg[7]  ( .Q(\re12[7] ), .D(n208), .CK(clk), .RB(n162) );
    DFFRBN \re11_reg[0]  ( .Q(\re11[0] ), .D(n209), .CK(clk), .RB(n147) );
    DFFRBN \re11_reg[1]  ( .Q(\re11[1] ), .D(n210), .CK(clk), .RB(n160) );
    DFFRBN \re11_reg[2]  ( .Q(\re11[2] ), .D(n211), .CK(clk), .RB(n147) );
    DFFRBN \re11_reg[3]  ( .Q(\re11[3] ), .D(n212), .CK(clk), .RB(n160) );
    DFFRBN \re11_reg[4]  ( .Q(\re11[4] ), .D(n213), .CK(clk), .RB(n148) );
    DFFRBN \re11_reg[5]  ( .Q(\re11[5] ), .D(n214), .CK(clk), .RB(n161) );
    DFFRBN \re11_reg[6]  ( .Q(\re11[6] ), .D(n215), .CK(clk), .RB(n148) );
    DFFRBN \re11_reg[7]  ( .Q(\re11[7] ), .D(n216), .CK(clk), .RB(n162) );
    DFFRBN \re10_reg[0]  ( .Q(\re10[0] ), .D(n217), .CK(clk), .RB(n149) );
    DFFRBN \re10_reg[1]  ( .Q(\re10[1] ), .D(n218), .CK(clk), .RB(n150) );
    DFFRBN \re10_reg[2]  ( .Q(\re10[2] ), .D(n219), .CK(clk), .RB(n149) );
    DFFRBN \re10_reg[3]  ( .Q(\re10[3] ), .D(n220), .CK(clk), .RB(n161) );
    DFFRBN \re10_reg[4]  ( .Q(\re10[4] ), .D(n221), .CK(clk), .RB(n149) );
    DFFRBN \re10_reg[5]  ( .Q(\re10[5] ), .D(n222), .CK(clk), .RB(n161) );
    DFFRBN \re10_reg[6]  ( .Q(\re10[6] ), .D(n223), .CK(clk), .RB(n147) );
    DFFRBN \re10_reg[7]  ( .Q(\re10[7] ), .D(n224), .CK(clk), .RB(n161) );
    DFFRBN \re9_reg[0]  ( .Q(\re9[0] ), .D(n225), .CK(clk), .RB(n144) );
    DFFRBN \re9_reg[1]  ( .Q(\re9[1] ), .D(n226), .CK(clk), .RB(n133) );
    DFFRBN \re9_reg[2]  ( .Q(\re9[2] ), .D(n227), .CK(clk), .RB(n143) );
    DFFRBN \re9_reg[3]  ( .Q(\re9[3] ), .D(n228), .CK(clk), .RB(n134) );
    DFFRBN \re9_reg[4]  ( .Q(\re9[4] ), .D(n229), .CK(clk), .RB(n143) );
    DFFRBN \re9_reg[5]  ( .Q(\re9[5] ), .D(n230), .CK(clk), .RB(n133) );
    DFFRBN \re9_reg[6]  ( .Q(\re9[6] ), .D(n231), .CK(clk), .RB(n143) );
    DFFRBN \re9_reg[7]  ( .Q(\re9[7] ), .D(n232), .CK(clk), .RB(n133) );
    DFFRBN \re8_reg[0]  ( .Q(\re8[0] ), .D(n233), .CK(clk), .RB(n144) );
    DFFRBN \re8_reg[1]  ( .Q(\re8[1] ), .D(n234), .CK(clk), .RB(n137) );
    DFFRBN \re8_reg[2]  ( .Q(\re8[2] ), .D(n235), .CK(clk), .RB(n144) );
    DFFRBN \re8_reg[3]  ( .Q(\re8[3] ), .D(n236), .CK(clk), .RB(n137) );
    DFFRBN \re8_reg[4]  ( .Q(\re8[4] ), .D(n237), .CK(clk), .RB(n145) );
    DFFRBN \re8_reg[5]  ( .Q(\re8[5] ), .D(n238), .CK(clk), .RB(n137) );
    DFFRBN \re8_reg[6]  ( .Q(\re8[6] ), .D(n239), .CK(clk), .RB(n145) );
    DFFRBN \re8_reg[7]  ( .Q(\re8[7] ), .D(n240), .CK(clk), .RB(n133) );
    DFFRBN \re7_reg[0]  ( .Q(\re7[0] ), .D(n241), .CK(clk), .RB(n146) );
    DFFRBN \re7_reg[1]  ( .Q(\re7[1] ), .D(n242), .CK(clk), .RB(n136) );
    DFFRBN \re7_reg[2]  ( .Q(\re7[2] ), .D(n243), .CK(clk), .RB(n146) );
    DFFRBN \re7_reg[3]  ( .Q(\re7[3] ), .D(n244), .CK(clk), .RB(n138) );
    DFFRBN \re7_reg[4]  ( .Q(\re7[4] ), .D(n245), .CK(clk), .RB(n146) );
    DFFRBN \re7_reg[5]  ( .Q(\re7[5] ), .D(n246), .CK(clk), .RB(n138) );
    DFFRBN \re7_reg[6]  ( .Q(\re7[6] ), .D(n247), .CK(clk), .RB(n144) );
    DFFRBN \re7_reg[7]  ( .Q(\re7[7] ), .D(n248), .CK(clk), .RB(n138) );
    DFFRBN \re6_reg[0]  ( .Q(\re6[0] ), .D(n249), .CK(clk), .RB(n139) );
    DFFRBN \re6_reg[1]  ( .Q(\re6[1] ), .D(n250), .CK(clk), .RB(n136) );
    DFFRBN \re6_reg[2]  ( .Q(\re6[2] ), .D(n251), .CK(clk), .RB(n146) );
    DFFRBN \re6_reg[3]  ( .Q(\re6[3] ), .D(n252), .CK(clk), .RB(n137) );
    DFFRBN \re6_reg[4]  ( .Q(\re6[4] ), .D(n253), .CK(clk), .RB(n145) );
    DFFRBN \re6_reg[5]  ( .Q(\re6[5] ), .D(n254), .CK(clk), .RB(n135) );
    DFFRBN \re6_reg[6]  ( .Q(\re6[6] ), .D(n255), .CK(clk), .RB(n145) );
    DFFRBN \re6_reg[7]  ( .Q(\re6[7] ), .D(n256), .CK(clk), .RB(n136) );
    DFFRBN \re5_reg[0]  ( .Q(\re5[0] ), .D(n257), .CK(clk), .RB(n139) );
    DFFRBN \re5_reg[1]  ( .Q(\re5[1] ), .D(n258), .CK(clk), .RB(n134) );
    DFFRBN \re5_reg[2]  ( .Q(\re5[2] ), .D(n259), .CK(clk), .RB(n138) );
    DFFRBN \re5_reg[3]  ( .Q(\re5[3] ), .D(n260), .CK(clk), .RB(n134) );
    DFFRBN \re5_reg[4]  ( .Q(\re5[4] ), .D(n261), .CK(clk), .RB(n140) );
    DFFRBN \re5_reg[5]  ( .Q(\re5[5] ), .D(n262), .CK(clk), .RB(n134) );
    DFFRBN \re5_reg[6]  ( .Q(\re5[6] ), .D(n263), .CK(clk), .RB(n139) );
    DFFRBN \re5_reg[7]  ( .Q(\re5[7] ), .D(n264), .CK(clk), .RB(n136) );
    DFFRBN \re4_reg[0]  ( .Q(\re4[0] ), .D(n265), .CK(clk), .RB(n141) );
    DFFRBN \re4_reg[1]  ( .Q(\re4[1] ), .D(n266), .CK(clk), .RB(n159) );
    DFFRBN \re4_reg[2]  ( .Q(\re4[2] ), .D(n267), .CK(clk), .RB(n141) );
    DFFRBN \re4_reg[3]  ( .Q(\re4[3] ), .D(n268), .CK(clk), .RB(n135) );
    DFFRBN \re4_reg[4]  ( .Q(\re4[4] ), .D(n269), .CK(clk), .RB(n141) );
    DFFRBN \re4_reg[5]  ( .Q(\re4[5] ), .D(n270), .CK(clk), .RB(n135) );
    DFFRBN \re4_reg[6]  ( .Q(\re4[6] ), .D(n271), .CK(clk), .RB(n139) );
    DFFRBN \re4_reg[7]  ( .Q(\re4[7] ), .D(n272), .CK(clk), .RB(n135) );
    DFFRBN \re3_reg[0]  ( .Q(\re3[0] ), .D(n273), .CK(clk), .RB(n142) );
    DFFRBN \re3_reg[1]  ( .Q(\re3[1] ), .D(n274), .CK(clk), .RB(n160) );
    DFFRBN \re3_reg[2]  ( .Q(\re3[2] ), .D(n275), .CK(clk), .RB(n140) );
    DFFRBN \re3_reg[3]  ( .Q(\re3[3] ), .D(n276), .CK(clk), .RB(n160) );
    DFFRBN \re3_reg[4]  ( .Q(\re3[4] ), .D(n277), .CK(clk), .RB(n140) );
    DFFRBN \re3_reg[5]  ( .Q(\re3[5] ), .D(n278), .CK(clk), .RB(n159) );
    DFFRBN \re3_reg[6]  ( .Q(\re3[6] ), .D(n279), .CK(clk), .RB(n140) );
    DFFRBN \re3_reg[7]  ( .Q(\re3[7] ), .D(n280), .CK(clk), .RB(n159) );
    DFFRBN \re2_reg[0]  ( .Q(\re2[0] ), .D(n281), .CK(clk), .RB(n142) );
    DFFRBN \re2_reg[1]  ( .Q(\re2[1] ), .D(n282), .CK(clk), .RB(n157) );
    DFFRBN \re2_reg[2]  ( .Q(\re2[2] ), .D(n283), .CK(clk), .RB(n141) );
    DFFRBN \re2_reg[3]  ( .Q(\re2[3] ), .D(n284), .CK(clk), .RB(n157) );
    DFFRBN \re2_reg[4]  ( .Q(\re2[4] ), .D(n285), .CK(clk), .RB(n143) );
    DFFRBN \re2_reg[5]  ( .Q(\re2[5] ), .D(n286), .CK(clk), .RB(n158) );
    DFFRBN \re2_reg[6]  ( .Q(\re2[6] ), .D(n287), .CK(clk), .RB(n142) );
    DFFRBN \re2_reg[7]  ( .Q(\re2[7] ), .D(n288), .CK(clk), .RB(n159) );
    DFFRBN \re1_reg[0]  ( .Q(\re1[0] ), .D(n289), .CK(clk), .RB(n152) );
    DFFRBN \re1_reg[1]  ( .Q(\re1[1] ), .D(n290), .CK(clk), .RB(n156) );
    DFFRBN \re1_reg[2]  ( .Q(\re1[2] ), .D(n291), .CK(clk), .RB(n152) );
    DFFRBN \re1_reg[3]  ( .Q(\re1[3] ), .D(n292), .CK(clk), .RB(n158) );
    DFFRBN \re1_reg[4]  ( .Q(\re1[4] ), .D(n293), .CK(clk), .RB(n152) );
    DFFRBN \re1_reg[5]  ( .Q(\re1[5] ), .D(n294), .CK(clk), .RB(n158) );
    DFFRBN \re1_reg[6]  ( .Q(\re1[6] ), .D(n295), .CK(clk), .RB(n142) );
    DFFRBN \re1_reg[7]  ( .Q(\re1[7] ), .D(n296), .CK(clk), .RB(n158) );
    DFFRBN \re0_reg[0]  ( .Q(\re0[0] ), .D(n297), .CK(clk), .RB(n150) );
    DFFRBN \re0_reg[1]  ( .Q(\re0[1] ), .D(n298), .CK(clk), .RB(n151) );
    DFFRBN \re0_reg[2]  ( .Q(\re0[2] ), .D(n299), .CK(clk), .RB(n149) );
    DFFRBN \re0_reg[3]  ( .Q(\re0[3] ), .D(n300), .CK(clk), .RB(n151) );
    DFFRBN \re0_reg[4]  ( .Q(\re0[4] ), .D(n301), .CK(clk), .RB(n148) );
    DFFRBN \re0_reg[5]  ( .Q(\re0[5] ), .D(n302), .CK(clk), .RB(n150) );
    DFFRBN \re0_reg[6]  ( .Q(\re0[6] ), .D(n303), .CK(clk), .RB(n148) );
    DFFRBN \re0_reg[7]  ( .Q(\re0[7] ), .D(n304), .CK(clk), .RB(n150) );
    DFFRBN \re15_reg[0]  ( .Q(\re15[0] ), .D(n305), .CK(clk), .RB(n153) );
    DFFRBN \re15_reg[1]  ( .Q(\re15[1] ), .D(n306), .CK(clk), .RB(n157) );
    DFFRBN \re15_reg[2]  ( .Q(\re15[2] ), .D(n307), .CK(clk), .RB(n152) );
    DFFRBN \re15_reg[3]  ( .Q(\re15[3] ), .D(n308), .CK(clk), .RB(n157) );
    DFFRBN \re15_reg[4]  ( .Q(\re15[4] ), .D(n309), .CK(clk), .RB(n151) );
    DFFRBN \re15_reg[5]  ( .Q(\re15[5] ), .D(n310), .CK(clk), .RB(n156) );
    DFFRBN \re15_reg[6]  ( .Q(\re15[6] ), .D(n311), .CK(clk), .RB(n151) );
    DFFRBN \re15_reg[7]  ( .Q(\re15[7] ), .D(n312), .CK(clk), .RB(n156) );
    INV2 U318 ( .O(n342), .I(aw[2]) );
    AOI2222 U319 ( .O(n351), .A1(n114), .A2(\re15[7] ), .B1(n352), .B2(
        \re14[7] ), .C1(n110), .C2(\re13[7] ), .D1(n353), .D2(\re12[7] ) );
    AOI2222 U320 ( .O(n354), .A1(n112), .A2(\re11[7] ), .B1(n355), .B2(
        \re10[7] ), .C1(n107), .C2(\re9[7] ), .D1(n356), .D2(\re8[7] ) );
    AOI2222 U321 ( .O(n313), .A1(n113), .A2(\re7[7] ), .B1(n357), .B2(\re6[7] 
        ), .C1(n108), .C2(\re5[7] ), .D1(n358), .D2(\re4[7] ) );
    AOI2222 U322 ( .O(n314), .A1(n111), .A2(\re3[7] ), .B1(n359), .B2(\re2[7] 
        ), .C1(n106), .C2(\re1[7] ), .D1(n360), .D2(\re0[7] ) );
    AOI2222 U323 ( .O(n361), .A1(\re15[6] ), .A2(n57), .B1(\re14[6] ), .B2(
        n352), .C1(\re13[6] ), .C2(n110), .D1(\re12[6] ), .D2(n353) );
    AOI2222 U324 ( .O(n362), .A1(\re11[6] ), .A2(n59), .B1(\re10[6] ), .B2(
        n355), .C1(\re9[6] ), .C2(n107), .D1(\re8[6] ), .D2(n356) );
    AOI2222 U325 ( .O(n315), .A1(\re7[6] ), .A2(n58), .B1(\re6[6] ), .B2(n357), 
        .C1(\re5[6] ), .C2(n108), .D1(\re4[6] ), .D2(n358) );
    AOI2222 U326 ( .O(n316), .A1(\re3[6] ), .A2(n60), .B1(\re2[6] ), .B2(n359), 
        .C1(\re1[6] ), .C2(n106), .D1(\re0[6] ), .D2(n360) );
    AOI2222 U327 ( .O(n363), .A1(\re15[5] ), .A2(n114), .B1(\re14[5] ), .B2(
        n352), .C1(\re13[5] ), .C2(n110), .D1(\re12[5] ), .D2(n353) );
    AOI2222 U328 ( .O(n364), .A1(\re11[5] ), .A2(n112), .B1(\re10[5] ), .B2(
        n355), .C1(\re9[5] ), .C2(n107), .D1(\re8[5] ), .D2(n356) );
    AOI2222 U329 ( .O(n317), .A1(\re7[5] ), .A2(n113), .B1(\re6[5] ), .B2(n357
        ), .C1(\re5[5] ), .C2(n108), .D1(\re4[5] ), .D2(n358) );
    AOI2222 U330 ( .O(n318), .A1(\re3[5] ), .A2(n111), .B1(\re2[5] ), .B2(n359
        ), .C1(\re1[5] ), .C2(n106), .D1(\re0[5] ), .D2(n360) );
    AOI2222 U331 ( .O(n365), .A1(\re15[4] ), .A2(n114), .B1(\re14[4] ), .B2(
        n352), .C1(\re13[4] ), .C2(n110), .D1(\re12[4] ), .D2(n353) );
    AOI2222 U332 ( .O(n366), .A1(\re11[4] ), .A2(n112), .B1(\re10[4] ), .B2(
        n355), .C1(\re9[4] ), .C2(n107), .D1(\re8[4] ), .D2(n356) );
    AOI2222 U333 ( .O(n319), .A1(\re7[4] ), .A2(n113), .B1(\re6[4] ), .B2(n357
        ), .C1(\re5[4] ), .C2(n108), .D1(\re4[4] ), .D2(n358) );
    AOI2222 U334 ( .O(n320), .A1(\re3[4] ), .A2(n111), .B1(\re2[4] ), .B2(n359
        ), .C1(\re1[4] ), .C2(n106), .D1(\re0[4] ), .D2(n360) );
    AOI2222 U335 ( .O(n367), .A1(\re15[3] ), .A2(n57), .B1(\re14[3] ), .B2(
        n352), .C1(\re13[3] ), .C2(n110), .D1(\re12[3] ), .D2(n353) );
    AOI2222 U336 ( .O(n368), .A1(\re11[3] ), .A2(n59), .B1(\re10[3] ), .B2(
        n355), .C1(\re9[3] ), .C2(n107), .D1(\re8[3] ), .D2(n356) );
    AOI2222 U337 ( .O(n321), .A1(\re7[3] ), .A2(n58), .B1(\re6[3] ), .B2(n357), 
        .C1(\re5[3] ), .C2(n108), .D1(\re4[3] ), .D2(n358) );
    AOI2222 U338 ( .O(n322), .A1(\re3[3] ), .A2(n60), .B1(\re2[3] ), .B2(n359), 
        .C1(\re1[3] ), .C2(n106), .D1(\re0[3] ), .D2(n360) );
    AOI2222 U339 ( .O(n369), .A1(\re15[2] ), .A2(n114), .B1(\re14[2] ), .B2(
        n352), .C1(\re13[2] ), .C2(n110), .D1(\re12[2] ), .D2(n353) );
    AOI2222 U340 ( .O(n370), .A1(\re11[2] ), .A2(n112), .B1(\re10[2] ), .B2(
        n355), .C1(\re9[2] ), .C2(n107), .D1(\re8[2] ), .D2(n356) );
    AOI2222 U341 ( .O(n323), .A1(\re7[2] ), .A2(n113), .B1(\re6[2] ), .B2(n357
        ), .C1(\re5[2] ), .C2(n108), .D1(\re4[2] ), .D2(n358) );
    AOI2222 U342 ( .O(n324), .A1(\re3[2] ), .A2(n111), .B1(\re2[2] ), .B2(n359
        ), .C1(\re1[2] ), .C2(n106), .D1(\re0[2] ), .D2(n360) );
    AOI2222 U343 ( .O(n371), .A1(\re15[1] ), .A2(n114), .B1(\re14[1] ), .B2(
        n352), .C1(\re13[1] ), .C2(n110), .D1(\re12[1] ), .D2(n353) );
    AOI2222 U344 ( .O(n372), .A1(\re11[1] ), .A2(n112), .B1(\re10[1] ), .B2(
        n355), .C1(\re9[1] ), .C2(n107), .D1(\re8[1] ), .D2(n356) );
    AOI2222 U345 ( .O(n325), .A1(\re7[1] ), .A2(n113), .B1(\re6[1] ), .B2(n357
        ), .C1(\re5[1] ), .C2(n108), .D1(\re4[1] ), .D2(n358) );
    AOI2222 U346 ( .O(n326), .A1(\re3[1] ), .A2(n111), .B1(\re2[1] ), .B2(n359
        ), .C1(\re1[1] ), .C2(n106), .D1(\re0[1] ), .D2(n360) );
    AOI2222 U347 ( .O(n373), .A1(\re15[0] ), .A2(n114), .B1(\re14[0] ), .B2(
        n352), .C1(\re13[0] ), .C2(n110), .D1(\re12[0] ), .D2(n353) );
    AOI2222 U348 ( .O(n374), .A1(\re11[0] ), .A2(n112), .B1(\re10[0] ), .B2(
        n355), .C1(\re9[0] ), .C2(n107), .D1(\re8[0] ), .D2(n356) );
    AOI2222 U349 ( .O(n327), .A1(\re7[0] ), .A2(n113), .B1(\re6[0] ), .B2(n357
        ), .C1(\re5[0] ), .C2(n108), .D1(\re4[0] ), .D2(n358) );
    AOI2222 U350 ( .O(n328), .A1(\re3[0] ), .A2(n111), .B1(\re2[0] ), .B2(n359
        ), .C1(\re1[0] ), .C2(n106), .D1(\re0[0] ), .D2(n360) );
endmodule


module fifo16x8 ( rst, clk, clr, rd_n, wr_n, di, \do , full, empty );
input  [7:0] di;
output [7:0] \do ;
input  rst, clk, clr, rd_n, wr_n;
output full, empty;
    wire n114, n115, \p_wr[3] , \p_wr[2] , \p_wr[1] , \p_wr[0] , \p_rd[3] , 
        \p_rd[2] , \p_rd[1] , \p_rd[0] , \do_m[7] , \do_m[6] , \do_m[5] , 
        \do_m[4] , \do_m[3] , \do_m[2] , \do_m[1] , \do_m[0] , N169, N170, n10, 
        n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
        n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39, 
        n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
        n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
        n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
        n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
        n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
        n109, n110, n111, n112, n113;
    rr16 fifo_regs ( .clk(clk), .rst(n31), .aw({n52, \p_wr[2] , n40, n48}), 
        .ar({n42, n47, n49, n53}), .d(di), .wr_n(n65), .full(n114), .do_m({
        \do_m[7] , \do_m[6] , \do_m[5] , \do_m[4] , \do_m[3] , \do_m[2] , 
        \do_m[1] , \do_m[0] }) );
    OR2P U3 ( .O(n103), .I1(n24), .I2(n25) );
    OR3 U4 ( .O(n74), .I1(n103), .I2(n27), .I3(n12) );
    OR2 U5 ( .O(n92), .I1(n103), .I2(n12) );
    XNR2 U6 ( .O(n80), .I1(n47), .I2(n81) );
    INV2 U7 ( .O(n14), .I(n12) );
    OR2 U8 ( .O(n10), .I1(n30), .I2(n26) );
    INV2 U9 ( .O(n39), .I(n10) );
    BUF1 U10 ( .O(n55), .I(\p_rd[0] ) );
    XOR2 U11 ( .O(N169), .I1(n13), .I2(n106) );
    XOR2 U12 ( .O(n109), .I1(\p_wr[1] ), .I2(n11) );
    OA12 U13 ( .O(n11), .A1(n106), .B1(n26), .B2(n30) );
    OR2P U14 ( .O(n12), .I1(n65), .I2(full) );
    BUF2 U15 ( .O(n48), .I(\p_wr[0] ) );
    INV3 U16 ( .O(full), .I(n36) );
    INV1 U17 ( .O(n107), .I(n65) );
    DFFRBP \p_wr_reg[2]  ( .Q(\p_wr[2] ), .QB(n27), .D(n21), .CK(clk), .RB(n59
        ) );
    AN2P U18 ( .O(n104), .I1(n39), .I2(\p_rd[2] ) );
    XOR3 U19 ( .O(n70), .I1(n46), .I2(n13), .I3(n39) );
    BUF2 U20 ( .O(n34), .I(n66) );
    MUX2 U21 ( .O(n101), .S(n66), .A(\do [6]), .B(\do_m[6] ) );
    INV2 U22 ( .O(n67), .I(n66) );
    MUX2 U23 ( .O(n99), .S(n34), .A(\do [4]), .B(\do_m[4] ) );
    INV3 U24 ( .O(n41), .I(\p_rd[3] ) );
    INV2 U25 ( .O(n89), .I(clr) );
    NR2P U26 ( .O(n105), .I1(\p_rd[2] ), .I2(n106) );
    INV3 U27 ( .O(n42), .I(n41) );
    ND2 U28 ( .O(n76), .I1(n14), .I2(n48) );
    ND2 U29 ( .O(n81), .I1(n38), .I2(n39) );
    ND2 U30 ( .O(n83), .I1(n38), .I2(n55) );
    BUF2 U31 ( .O(n38), .I(n29) );
    XOR2 U32 ( .O(N170), .I1(n43), .I2(n105) );
    BUF2 U33 ( .O(n40), .I(\p_wr[1] ) );
    INV2 U34 ( .O(n46), .I(n45) );
    BUF1 U35 ( .O(n45), .I(\p_wr[2] ) );
    ND2 U36 ( .O(n88), .I1(n85), .I2(n24) );
    DFFRBP \p_wr_reg[3]  ( .Q(\p_wr[3] ), .QB(n51), .D(n23), .CK(clk), .RB(n61
        ) );
    BUF2 U37 ( .O(n57), .I(n89) );
    BUF2 U38 ( .O(n58), .I(n89) );
    BUF3 U39 ( .O(n31), .I(rst) );
    BUF3 U40 ( .O(n47), .I(\p_rd[2] ) );
    BUF2 U41 ( .O(n50), .I(\p_rd[1] ) );
    BUF3 U42 ( .O(n49), .I(\p_rd[1] ) );
    INV2 U43 ( .O(n113), .I(\p_wr[3] ) );
    DFFRBP \p_rd_reg[3]  ( .Q(\p_rd[3] ), .D(n18), .CK(clk), .RB(n35) );
    DFFRBP \p_rd_reg[0]  ( .Q(\p_rd[0] ), .QB(n26), .D(n15), .CK(clk), .RB(n61
        ) );
    BUF1 U44 ( .O(n54), .I(\p_rd[0] ) );
    INV2 U45 ( .O(n43), .I(n41) );
    AN2 U46 ( .O(n15), .I1(n84), .I2(n58) );
    AN2 U47 ( .O(n16), .I1(n82), .I2(n57) );
    AN2 U48 ( .O(n17), .I1(n80), .I2(n58) );
    AN2 U49 ( .O(n18), .I1(n78), .I2(n57) );
    AN2 U50 ( .O(n19), .I1(n77), .I2(n57) );
    AN2 U51 ( .O(n20), .I1(n75), .I2(n58) );
    AN2 U52 ( .O(n21), .I1(n90), .I2(n58) );
    AOI12 U53 ( .O(n22), .A1(n63), .B1(n108), .B2(n91) );
    AN2 U54 ( .O(n23), .I1(n73), .I2(n57) );
    DFFRBP \p_wr_reg[1]  ( .Q(\p_wr[1] ), .QB(n25), .D(n20), .CK(clk), .RB(n62
        ) );
    INV2 U55 ( .O(n64), .I(wr_n) );
    DFFRBP \p_wr_reg[0]  ( .Q(\p_wr[0] ), .QB(n24), .D(n19), .CK(clk), .RB(n59
        ) );
    DFFRBP \p_rd_reg[2]  ( .Q(\p_rd[2] ), .QB(n13), .D(n17), .CK(clk), .RB(n60
        ) );
    BUF2 U56 ( .O(empty), .I(n115) );
    INV3 U57 ( .O(n65), .I(n64) );
    AN2P U58 ( .O(n29), .I1(n66), .I2(n28) );
    DFFRBP \p_rd_reg[1]  ( .Q(\p_rd[1] ), .QB(n30), .D(n16), .CK(clk), .RB(n35
        ) );
    INV2 U59 ( .O(n63), .I(n56) );
    BUF3 U60 ( .O(n60), .I(n93) );
    BUF3 U61 ( .O(n61), .I(n93) );
    BUF1 U62 ( .O(n32), .I(n71) );
    BUF1 U63 ( .O(n33), .I(n70) );
    ND2 U64 ( .O(n79), .I1(n104), .I2(n38) );
    XOR2 U65 ( .O(n112), .I1(n24), .I2(n26) );
    XOR2 U66 ( .O(n110), .I1(n46), .I2(N169) );
    XOR2 U67 ( .O(n111), .I1(n113), .I2(N170) );
    XOR2 U68 ( .O(n82), .I1(n30), .I2(n83) );
    XOR2 U69 ( .O(n78), .I1(n41), .I2(n79) );
    XOR2 U70 ( .O(n73), .I1(n113), .I2(n74) );
    XOR2 U71 ( .O(n75), .I1(n25), .I2(n76) );
    XOR2 U72 ( .O(n90), .I1(n92), .I2(n27) );
    OR2P U73 ( .O(n106), .I1(n54), .I2(n50) );
    BUF4 U74 ( .O(n35), .I(n93) );
    DFFRBP full_reg ( .Q(n114), .QB(n36), .D(n22), .CK(clk), .RB(n59) );
    DFFRBT \do_reg[1]  ( .Q(\do [1]), .D(n96), .CK(clk), .RB(n35) );
    DFFRBT \do_reg[0]  ( .Q(\do [0]), .D(n95), .CK(clk), .RB(n62) );
    DFFRBT \do_reg[2]  ( .Q(\do [2]), .D(n97), .CK(clk), .RB(n60) );
    XOR2 U75 ( .O(n77), .I1(\p_wr[0] ), .I2(n14) );
    ND2 U76 ( .O(n86), .I1(n87), .I2(\p_wr[0] ) );
    XOR2 U77 ( .O(n87), .I1(n25), .I2(n50) );
    XOR2 U78 ( .O(n85), .I1(n50), .I2(\p_wr[1] ) );
    INV3 U79 ( .O(n52), .I(n51) );
    BUF3 U80 ( .O(n53), .I(\p_rd[0] ) );
    XOR2 U81 ( .O(n84), .I1(n54), .I2(n29) );
    BUF1 U82 ( .O(n56), .I(n89) );
    BUF4 U83 ( .O(n59), .I(n93) );
    BUF4 U84 ( .O(n62), .I(n93) );
    DFFRBT \do_reg[4]  ( .Q(\do [4]), .D(n99), .CK(clk), .RB(n62) );
    DFFRBT \do_reg[6]  ( .Q(\do [6]), .D(n101), .CK(clk), .RB(n35) );
    DFFRBT \do_reg[7]  ( .Q(\do [7]), .D(n102), .CK(clk), .RB(n59) );
    DFFRBT \do_reg[5]  ( .Q(\do [5]), .D(n100), .CK(clk), .RB(n60) );
    DFFRBT \do_reg[3]  ( .Q(\do [3]), .D(n98), .CK(clk), .RB(n61) );
    INV4 U85 ( .O(n93), .I(n31) );
    INV3 U86 ( .O(n66), .I(rd_n) );
    INV4 U87 ( .O(n68), .I(n34) );
    ND2 U88 ( .O(n91), .I1(n67), .I2(n114) );
    AO112 U89 ( .O(n94), .A1(n63), .B1(n69), .C1(empty), .C2(n65) );
    NR5 U90 ( .O(n69), .I1(n68), .I2(n33), .I3(n107), .I4(n32), .I5(n72) );
    XOR3 U91 ( .O(n71), .I1(n43), .I2(\p_wr[3] ), .I3(n104) );
    MUX2 U92 ( .O(n72), .S(n55), .A(n86), .B(n88) );
    MUX2 U93 ( .O(n102), .S(n68), .A(\do_m[7] ), .B(\do [7]) );
    MUX2 U94 ( .O(n100), .S(n68), .A(\do_m[5] ), .B(\do [5]) );
    MUX2 U95 ( .O(n98), .S(n67), .A(\do_m[3] ), .B(\do [3]) );
    MUX2 U96 ( .O(n97), .S(n68), .A(\do_m[2] ), .B(\do [2]) );
    MUX2 U97 ( .O(n96), .S(n68), .A(\do_m[1] ), .B(\do [1]) );
    MUX2 U98 ( .O(n95), .S(n67), .A(\do_m[0] ), .B(\do [0]) );
    DFFSBN empty_reg ( .Q(n115), .QB(n28), .D(n94), .CK(clk), .SB(n62) );
    ND6 U99 ( .O(n108), .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n107), 
        .I6(n68) );
endmodule

