library verilog;
use verilog.vl_types.all;
entity ROUTINES is
end ROUTINES;
