
`ifndef RKV_I2C_TESTS_SVH
`define RKV_I2C_TESTS_SVH

`include "rkv_i2c_base_test.sv"
`include "rkv_i2c_quick_reg_access_test.sv"
`include "rkv_i2c_directed_tx_test.sv"
`include "rkv_i2c_directed_rx_test.sv"

`endif // RKV_I2C_TESTS_SVH
