/************************************************************************\
|*                                                                      *|
|*    Copyright (c) 2005  Springer. All rights reserved.                *|
|*                                                                      *|
|*  This example code shouyld be used only for illustration purpose     *| 
|*  This material is not to reproduced,  copied,  or used  in any       *|
|*  manner without the authorization of the author's/publishers         *|
|*  written permission                                                  *|
|*                                                                      *|
\************************************************************************/

// Author: Srikanth Vijayaraghavan and Meyyappan Ramanathan


module xpose_b(

input logic signed [15:0] d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28, d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61,d62,d63,d64,

output logic signed [15:0] q1,q2,q3,q4,q5,q6,q7,q8,q9,q10, q11,q12,q13,q14,q15,q16,q17,q18,q19,q20,q21,q22,q23,q24,q25, q26,q27,q28, q29,q30,q31,q32,q33,q34,q35,q36,q37,q38,q39,q40,q41,q42,q43,q44,q45,q46,q47,q48,q49,q50,q51,q52,q53,q54,q55,q56,q57,q58,q59,q60,q61,q62,q63,q64);


always@(*)
begin
q1 <= d1;
q9 <= d2;
q17 <= d3;
q25 <= d4;
q33 <= d5;
q41 <= d6;
q49 <= d7;
q57 <= d8;
q2 <= d9;
q10 <= d10;
q18 <= d11;
q26 <= d12;
q34 <= d13;
q42 <= d14;
q50 <= d15;
q58 <= d16;
q3 <= d17;
q11 <= d18;
q19 <= d19;
q27 <= d20;
q35 <= d21;
q43 <= d22;
q51 <= d23;
q59 <= d24;
q4 <= d25;
q12 <= d26;
q20 <= d27;
q28 <= d28;
q36 <= d29;
q44 <= d30;
q52 <= d31;
q60 <= d32;
q5 <= d33;
q13 <= d34;
q21 <= d35;
q29 <= d36;
q37 <= d37;
q45 <= d38;
q53 <= d39;
q61 <= d40;
q6 <= d41;
q14 <= d42;
q22 <= d43;
q30 <= d44;
q38 <= d45;
q46 <= d46;
q54 <= d47;
q62 <= d48;
q7 <= d49;
q15 <= d50;
q23 <= d51;
q31 <= d52;
q39 <= d53;
q47 <= d54;
q55 <= d54;
q63 <= d56;
q8 <= d57;
q16 <= d58;
q24 <= d59;
q32 <= d60;
q40 <= d61;
q48 <= d62;
q56 <= d63;
q64 <= d64;
end

endmodule









