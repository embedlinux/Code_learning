library verilog;
use verilog.vl_types.all;
entity myscfifo_tb is
end myscfifo_tb;
