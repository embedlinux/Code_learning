//----------------------------------------------------------------------------------------------------------
// Design Unit : Byte input FF received CRC
// Version : v0.1 2007/05/20
//----------------------------------------------------------------------------------------------------------
module ff_rcv_fcs_1b(clk,rst,en,d,fok);
input clk;
input rst;
input en;
input d;
output fok;
//-----------------------------------------------------------------------------------------------------------
//-----------------------------------------------------------------------------------------------------------
reg[15:0] q;
wire[15:0] qi;
wire fok;
//-----------------------------------------------------------------------------------------------------------
//-----------------------------------------------------------------------------------------------------------
always @(posedge clk or posedge rst)
begin
    if(rst == 1'b1)
        q <= 16'hffff;
    else if(en == 1'b1)
        q <= qi;
end
//------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------
wire iw;
assign iw = d ^ q[15];
assign qi[0]  = iw; 
assign qi[1]  = iw ^ q[0]; 
assign qi[2]  = iw ^ q[1];
assign qi[3]  = iw ^ q[2];
assign qi[4]  = q[3];
assign qi[5]  = q[4];
assign qi[6]  = iw ^ q[5];
assign qi[7]  = iw ^ q[6];
assign qi[8]  = iw ^ q[7];
assign qi[9]  = q[8];
assign qi[10] = iw ^ q[9];
assign qi[11] = iw ^ q[10];
assign qi[12] = iw ^ q[11];
assign qi[13] = q[12];
assign qi[14] = q[13];
assign qi[15] = q[14];
//-----------------------------------------------------------------------------------------------------------
assign fok = !q[0] & !q[1] & q[2] & !q[3] & q[4] & !q[5] & !q[6] & q[7] 
             & q[8] & q[9] & !q[10] & !q[11] & !q[12] & q[13] & q[14] & q[15];
//------------------------------------------------------------------------------------------------------------
endmodule
 