/*-----------------------------------------------------------------
File name     : top.sv
Description   : lab02_uvc top level module template file
Notes         : From the Cadence "SystemVerilog Accelerated Verification with UVM" training
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2015
-----------------------------------------------------------------*/

module top ();

  // import the UVM library
  import uvm_pkg::*;

  // include the UVM macros
  `include "uvm_macros.svh"

  // import the yapp package

  // define an environment handle
  // create an environment instance
  // run the test


  // code required for second part of lab02
  //uvm_config_wrapper::set(null, "<path>.run_phase",
  //                        "default_sequence",
  //                        yapp_5_packets::type_id::get());


endmodule : top
