library verilog;
use verilog.vl_types.all;
entity UART_DPRAM_tb is
end UART_DPRAM_tb;
