
module Mem ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, ClkR, ClkW, 
        ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, n716, ClockR, ClockW, Dreadyr,
         \Storage[31][32] , \Storage[31][31] , \Storage[31][30] ,
         \Storage[31][29] , \Storage[31][28] , \Storage[31][27] ,
         \Storage[31][26] , \Storage[31][25] , \Storage[31][24] ,
         \Storage[31][23] , \Storage[31][22] , \Storage[31][21] ,
         \Storage[31][20] , \Storage[31][19] , \Storage[31][18] ,
         \Storage[31][17] , \Storage[31][16] , \Storage[31][15] ,
         \Storage[31][14] , \Storage[31][13] , \Storage[31][12] ,
         \Storage[31][11] , \Storage[31][10] , \Storage[31][9] ,
         \Storage[31][8] , \Storage[31][7] , \Storage[31][6] ,
         \Storage[31][5] , \Storage[31][4] , \Storage[31][3] ,
         \Storage[31][2] , \Storage[31][1] , \Storage[31][0] ,
         \Storage[30][32] , \Storage[30][31] , \Storage[30][30] ,
         \Storage[30][29] , \Storage[30][28] , \Storage[30][27] ,
         \Storage[30][26] , \Storage[30][25] , \Storage[30][24] ,
         \Storage[30][23] , \Storage[30][22] , \Storage[30][21] ,
         \Storage[30][20] , \Storage[30][19] , \Storage[30][18] ,
         \Storage[30][17] , \Storage[30][16] , \Storage[30][15] ,
         \Storage[30][14] , \Storage[30][13] , \Storage[30][12] ,
         \Storage[30][11] , \Storage[30][10] , \Storage[30][9] ,
         \Storage[30][8] , \Storage[30][7] , \Storage[30][6] ,
         \Storage[30][5] , \Storage[30][4] , \Storage[30][3] ,
         \Storage[30][2] , \Storage[30][1] , \Storage[30][0] ,
         \Storage[29][32] , \Storage[29][31] , \Storage[29][30] ,
         \Storage[29][29] , \Storage[29][28] , \Storage[29][27] ,
         \Storage[29][26] , \Storage[29][25] , \Storage[29][24] ,
         \Storage[29][23] , \Storage[29][22] , \Storage[29][21] ,
         \Storage[29][20] , \Storage[29][19] , \Storage[29][18] ,
         \Storage[29][17] , \Storage[29][16] , \Storage[29][15] ,
         \Storage[29][14] , \Storage[29][13] , \Storage[29][12] ,
         \Storage[29][11] , \Storage[29][10] , \Storage[29][9] ,
         \Storage[29][8] , \Storage[29][7] , \Storage[29][6] ,
         \Storage[29][5] , \Storage[29][4] , \Storage[29][3] ,
         \Storage[29][2] , \Storage[29][1] , \Storage[29][0] ,
         \Storage[28][32] , \Storage[28][31] , \Storage[28][30] ,
         \Storage[28][29] , \Storage[28][28] , \Storage[28][27] ,
         \Storage[28][26] , \Storage[28][25] , \Storage[28][24] ,
         \Storage[28][23] , \Storage[28][22] , \Storage[28][21] ,
         \Storage[28][20] , \Storage[28][19] , \Storage[28][18] ,
         \Storage[28][17] , \Storage[28][16] , \Storage[28][15] ,
         \Storage[28][14] , \Storage[28][13] , \Storage[28][12] ,
         \Storage[28][11] , \Storage[28][10] , \Storage[28][9] ,
         \Storage[28][8] , \Storage[28][7] , \Storage[28][6] ,
         \Storage[28][5] , \Storage[28][4] , \Storage[28][3] ,
         \Storage[28][2] , \Storage[28][1] , \Storage[28][0] ,
         \Storage[27][32] , \Storage[27][31] , \Storage[27][30] ,
         \Storage[27][29] , \Storage[27][28] , \Storage[27][27] ,
         \Storage[27][26] , \Storage[27][25] , \Storage[27][24] ,
         \Storage[27][23] , \Storage[27][22] , \Storage[27][21] ,
         \Storage[27][20] , \Storage[27][19] , \Storage[27][18] ,
         \Storage[27][17] , \Storage[27][16] , \Storage[27][15] ,
         \Storage[27][14] , \Storage[27][13] , \Storage[27][12] ,
         \Storage[27][11] , \Storage[27][10] , \Storage[27][9] ,
         \Storage[27][8] , \Storage[27][7] , \Storage[27][6] ,
         \Storage[27][5] , \Storage[27][4] , \Storage[27][3] ,
         \Storage[27][2] , \Storage[27][1] , \Storage[27][0] ,
         \Storage[26][32] , \Storage[26][31] , \Storage[26][30] ,
         \Storage[26][29] , \Storage[26][28] , \Storage[26][27] ,
         \Storage[26][26] , \Storage[26][25] , \Storage[26][24] ,
         \Storage[26][23] , \Storage[26][22] , \Storage[26][21] ,
         \Storage[26][20] , \Storage[26][19] , \Storage[26][18] ,
         \Storage[26][17] , \Storage[26][16] , \Storage[26][15] ,
         \Storage[26][14] , \Storage[26][13] , \Storage[26][12] ,
         \Storage[26][11] , \Storage[26][10] , \Storage[26][9] ,
         \Storage[26][8] , \Storage[26][7] , \Storage[26][6] ,
         \Storage[26][5] , \Storage[26][4] , \Storage[26][3] ,
         \Storage[26][2] , \Storage[26][1] , \Storage[26][0] ,
         \Storage[25][32] , \Storage[25][31] , \Storage[25][30] ,
         \Storage[25][29] , \Storage[25][28] , \Storage[25][27] ,
         \Storage[25][26] , \Storage[25][25] , \Storage[25][24] ,
         \Storage[25][23] , \Storage[25][22] , \Storage[25][21] ,
         \Storage[25][20] , \Storage[25][19] , \Storage[25][18] ,
         \Storage[25][17] , \Storage[25][16] , \Storage[25][15] ,
         \Storage[25][14] , \Storage[25][13] , \Storage[25][12] ,
         \Storage[25][11] , \Storage[25][10] , \Storage[25][9] ,
         \Storage[25][8] , \Storage[25][7] , \Storage[25][6] ,
         \Storage[25][5] , \Storage[25][4] , \Storage[25][3] ,
         \Storage[25][2] , \Storage[25][1] , \Storage[25][0] ,
         \Storage[24][32] , \Storage[24][31] , \Storage[24][30] ,
         \Storage[24][29] , \Storage[24][28] , \Storage[24][27] ,
         \Storage[24][26] , \Storage[24][25] , \Storage[24][24] ,
         \Storage[24][23] , \Storage[24][22] , \Storage[24][21] ,
         \Storage[24][20] , \Storage[24][19] , \Storage[24][18] ,
         \Storage[24][17] , \Storage[24][16] , \Storage[24][15] ,
         \Storage[24][14] , \Storage[24][13] , \Storage[24][12] ,
         \Storage[24][11] , \Storage[24][10] , \Storage[24][9] ,
         \Storage[24][8] , \Storage[24][7] , \Storage[24][6] ,
         \Storage[24][5] , \Storage[24][4] , \Storage[24][3] ,
         \Storage[24][2] , \Storage[24][1] , \Storage[24][0] ,
         \Storage[23][32] , \Storage[23][31] , \Storage[23][30] ,
         \Storage[23][29] , \Storage[23][28] , \Storage[23][27] ,
         \Storage[23][26] , \Storage[23][25] , \Storage[23][24] ,
         \Storage[23][23] , \Storage[23][22] , \Storage[23][21] ,
         \Storage[23][20] , \Storage[23][19] , \Storage[23][18] ,
         \Storage[23][17] , \Storage[23][16] , \Storage[23][15] ,
         \Storage[23][14] , \Storage[23][13] , \Storage[23][12] ,
         \Storage[23][11] , \Storage[23][10] , \Storage[23][9] ,
         \Storage[23][8] , \Storage[23][7] , \Storage[23][6] ,
         \Storage[23][5] , \Storage[23][4] , \Storage[23][3] ,
         \Storage[23][2] , \Storage[23][1] , \Storage[23][0] ,
         \Storage[22][32] , \Storage[22][31] , \Storage[22][30] ,
         \Storage[22][29] , \Storage[22][28] , \Storage[22][27] ,
         \Storage[22][26] , \Storage[22][25] , \Storage[22][24] ,
         \Storage[22][23] , \Storage[22][22] , \Storage[22][21] ,
         \Storage[22][20] , \Storage[22][19] , \Storage[22][18] ,
         \Storage[22][17] , \Storage[22][16] , \Storage[22][15] ,
         \Storage[22][14] , \Storage[22][13] , \Storage[22][12] ,
         \Storage[22][11] , \Storage[22][10] , \Storage[22][9] ,
         \Storage[22][8] , \Storage[22][7] , \Storage[22][6] ,
         \Storage[22][5] , \Storage[22][4] , \Storage[22][3] ,
         \Storage[22][2] , \Storage[22][1] , \Storage[22][0] ,
         \Storage[21][32] , \Storage[21][31] , \Storage[21][30] ,
         \Storage[21][29] , \Storage[21][28] , \Storage[21][27] ,
         \Storage[21][26] , \Storage[21][25] , \Storage[21][24] ,
         \Storage[21][23] , \Storage[21][22] , \Storage[21][21] ,
         \Storage[21][20] , \Storage[21][19] , \Storage[21][18] ,
         \Storage[21][17] , \Storage[21][16] , \Storage[21][15] ,
         \Storage[21][14] , \Storage[21][13] , \Storage[21][12] ,
         \Storage[21][11] , \Storage[21][10] , \Storage[21][9] ,
         \Storage[21][8] , \Storage[21][7] , \Storage[21][6] ,
         \Storage[21][5] , \Storage[21][4] , \Storage[21][3] ,
         \Storage[21][2] , \Storage[21][1] , \Storage[21][0] ,
         \Storage[20][32] , \Storage[20][31] , \Storage[20][30] ,
         \Storage[20][29] , \Storage[20][28] , \Storage[20][27] ,
         \Storage[20][26] , \Storage[20][25] , \Storage[20][24] ,
         \Storage[20][23] , \Storage[20][22] , \Storage[20][21] ,
         \Storage[20][20] , \Storage[20][19] , \Storage[20][18] ,
         \Storage[20][17] , \Storage[20][16] , \Storage[20][15] ,
         \Storage[20][14] , \Storage[20][13] , \Storage[20][12] ,
         \Storage[20][11] , \Storage[20][10] , \Storage[20][9] ,
         \Storage[20][8] , \Storage[20][7] , \Storage[20][6] ,
         \Storage[20][5] , \Storage[20][4] , \Storage[20][3] ,
         \Storage[20][2] , \Storage[20][1] , \Storage[20][0] ,
         \Storage[19][32] , \Storage[19][31] , \Storage[19][30] ,
         \Storage[19][29] , \Storage[19][28] , \Storage[19][27] ,
         \Storage[19][26] , \Storage[19][25] , \Storage[19][24] ,
         \Storage[19][23] , \Storage[19][22] , \Storage[19][21] ,
         \Storage[19][20] , \Storage[19][19] , \Storage[19][18] ,
         \Storage[19][17] , \Storage[19][16] , \Storage[19][15] ,
         \Storage[19][14] , \Storage[19][13] , \Storage[19][12] ,
         \Storage[19][11] , \Storage[19][10] , \Storage[19][9] ,
         \Storage[19][8] , \Storage[19][7] , \Storage[19][6] ,
         \Storage[19][5] , \Storage[19][4] , \Storage[19][3] ,
         \Storage[19][2] , \Storage[19][1] , \Storage[19][0] ,
         \Storage[18][32] , \Storage[18][31] , \Storage[18][30] ,
         \Storage[18][29] , \Storage[18][28] , \Storage[18][27] ,
         \Storage[18][26] , \Storage[18][25] , \Storage[18][24] ,
         \Storage[18][23] , \Storage[18][22] , \Storage[18][21] ,
         \Storage[18][20] , \Storage[18][19] , \Storage[18][18] ,
         \Storage[18][17] , \Storage[18][16] , \Storage[18][15] ,
         \Storage[18][14] , \Storage[18][13] , \Storage[18][12] ,
         \Storage[18][11] , \Storage[18][10] , \Storage[18][9] ,
         \Storage[18][8] , \Storage[18][7] , \Storage[18][6] ,
         \Storage[18][5] , \Storage[18][4] , \Storage[18][3] ,
         \Storage[18][2] , \Storage[18][1] , \Storage[18][0] ,
         \Storage[17][32] , \Storage[17][31] , \Storage[17][30] ,
         \Storage[17][29] , \Storage[17][28] , \Storage[17][27] ,
         \Storage[17][26] , \Storage[17][25] , \Storage[17][24] ,
         \Storage[17][23] , \Storage[17][22] , \Storage[17][21] ,
         \Storage[17][20] , \Storage[17][19] , \Storage[17][18] ,
         \Storage[17][17] , \Storage[17][16] , \Storage[17][15] ,
         \Storage[17][14] , \Storage[17][13] , \Storage[17][12] ,
         \Storage[17][11] , \Storage[17][10] , \Storage[17][9] ,
         \Storage[17][8] , \Storage[17][7] , \Storage[17][6] ,
         \Storage[17][5] , \Storage[17][4] , \Storage[17][3] ,
         \Storage[17][2] , \Storage[17][1] , \Storage[17][0] ,
         \Storage[16][32] , \Storage[16][31] , \Storage[16][30] ,
         \Storage[16][29] , \Storage[16][28] , \Storage[16][27] ,
         \Storage[16][26] , \Storage[16][25] , \Storage[16][24] ,
         \Storage[16][23] , \Storage[16][22] , \Storage[16][21] ,
         \Storage[16][20] , \Storage[16][19] , \Storage[16][18] ,
         \Storage[16][17] , \Storage[16][16] , \Storage[16][15] ,
         \Storage[16][14] , \Storage[16][13] , \Storage[16][12] ,
         \Storage[16][11] , \Storage[16][10] , \Storage[16][9] ,
         \Storage[16][8] , \Storage[16][7] , \Storage[16][6] ,
         \Storage[16][5] , \Storage[16][4] , \Storage[16][3] ,
         \Storage[16][2] , \Storage[16][1] , \Storage[16][0] ,
         \Storage[15][32] , \Storage[15][31] , \Storage[15][30] ,
         \Storage[15][29] , \Storage[15][28] , \Storage[15][27] ,
         \Storage[15][26] , \Storage[15][25] , \Storage[15][24] ,
         \Storage[15][23] , \Storage[15][22] , \Storage[15][21] ,
         \Storage[15][20] , \Storage[15][19] , \Storage[15][18] ,
         \Storage[15][17] , \Storage[15][16] , \Storage[15][15] ,
         \Storage[15][14] , \Storage[15][13] , \Storage[15][12] ,
         \Storage[15][11] , \Storage[15][10] , \Storage[15][9] ,
         \Storage[15][8] , \Storage[15][7] , \Storage[15][6] ,
         \Storage[15][5] , \Storage[15][4] , \Storage[15][3] ,
         \Storage[15][2] , \Storage[15][1] , \Storage[15][0] ,
         \Storage[14][32] , \Storage[14][31] , \Storage[14][30] ,
         \Storage[14][29] , \Storage[14][28] , \Storage[14][27] ,
         \Storage[14][26] , \Storage[14][25] , \Storage[14][24] ,
         \Storage[14][23] , \Storage[14][22] , \Storage[14][21] ,
         \Storage[14][20] , \Storage[14][19] , \Storage[14][18] ,
         \Storage[14][17] , \Storage[14][16] , \Storage[14][15] ,
         \Storage[14][14] , \Storage[14][13] , \Storage[14][12] ,
         \Storage[14][11] , \Storage[14][10] , \Storage[14][9] ,
         \Storage[14][8] , \Storage[14][7] , \Storage[14][6] ,
         \Storage[14][5] , \Storage[14][4] , \Storage[14][3] ,
         \Storage[14][2] , \Storage[14][1] , \Storage[14][0] ,
         \Storage[13][32] , \Storage[13][31] , \Storage[13][30] ,
         \Storage[13][29] , \Storage[13][28] , \Storage[13][27] ,
         \Storage[13][26] , \Storage[13][25] , \Storage[13][24] ,
         \Storage[13][23] , \Storage[13][22] , \Storage[13][21] ,
         \Storage[13][20] , \Storage[13][19] , \Storage[13][18] ,
         \Storage[13][17] , \Storage[13][16] , \Storage[13][15] ,
         \Storage[13][14] , \Storage[13][13] , \Storage[13][12] ,
         \Storage[13][11] , \Storage[13][10] , \Storage[13][9] ,
         \Storage[13][8] , \Storage[13][7] , \Storage[13][6] ,
         \Storage[13][5] , \Storage[13][4] , \Storage[13][3] ,
         \Storage[13][2] , \Storage[13][1] , \Storage[13][0] ,
         \Storage[12][32] , \Storage[12][31] , \Storage[12][30] ,
         \Storage[12][29] , \Storage[12][28] , \Storage[12][27] ,
         \Storage[12][26] , \Storage[12][25] , \Storage[12][24] ,
         \Storage[12][23] , \Storage[12][22] , \Storage[12][21] ,
         \Storage[12][20] , \Storage[12][19] , \Storage[12][18] ,
         \Storage[12][17] , \Storage[12][16] , \Storage[12][15] ,
         \Storage[12][14] , \Storage[12][13] , \Storage[12][12] ,
         \Storage[12][11] , \Storage[12][10] , \Storage[12][9] ,
         \Storage[12][8] , \Storage[12][7] , \Storage[12][6] ,
         \Storage[12][5] , \Storage[12][4] , \Storage[12][3] ,
         \Storage[12][2] , \Storage[12][1] , \Storage[12][0] ,
         \Storage[11][32] , \Storage[11][31] , \Storage[11][30] ,
         \Storage[11][29] , \Storage[11][28] , \Storage[11][27] ,
         \Storage[11][26] , \Storage[11][25] , \Storage[11][24] ,
         \Storage[11][23] , \Storage[11][22] , \Storage[11][21] ,
         \Storage[11][20] , \Storage[11][19] , \Storage[11][18] ,
         \Storage[11][17] , \Storage[11][16] , \Storage[11][15] ,
         \Storage[11][14] , \Storage[11][13] , \Storage[11][12] ,
         \Storage[11][11] , \Storage[11][10] , \Storage[11][9] ,
         \Storage[11][8] , \Storage[11][7] , \Storage[11][6] ,
         \Storage[11][5] , \Storage[11][4] , \Storage[11][3] ,
         \Storage[11][2] , \Storage[11][1] , \Storage[11][0] ,
         \Storage[10][32] , \Storage[10][31] , \Storage[10][30] ,
         \Storage[10][29] , \Storage[10][28] , \Storage[10][27] ,
         \Storage[10][26] , \Storage[10][25] , \Storage[10][24] ,
         \Storage[10][23] , \Storage[10][22] , \Storage[10][21] ,
         \Storage[10][20] , \Storage[10][19] , \Storage[10][18] ,
         \Storage[10][17] , \Storage[10][16] , \Storage[10][15] ,
         \Storage[10][14] , \Storage[10][13] , \Storage[10][12] ,
         \Storage[10][11] , \Storage[10][10] , \Storage[10][9] ,
         \Storage[10][8] , \Storage[10][7] , \Storage[10][6] ,
         \Storage[10][5] , \Storage[10][4] , \Storage[10][3] ,
         \Storage[10][2] , \Storage[10][1] , \Storage[10][0] ,
         \Storage[9][32] , \Storage[9][31] , \Storage[9][30] ,
         \Storage[9][29] , \Storage[9][28] , \Storage[9][27] ,
         \Storage[9][26] , \Storage[9][25] , \Storage[9][24] ,
         \Storage[9][23] , \Storage[9][22] , \Storage[9][21] ,
         \Storage[9][20] , \Storage[9][19] , \Storage[9][18] ,
         \Storage[9][17] , \Storage[9][16] , \Storage[9][15] ,
         \Storage[9][14] , \Storage[9][13] , \Storage[9][12] ,
         \Storage[9][11] , \Storage[9][10] , \Storage[9][9] , \Storage[9][8] ,
         \Storage[9][7] , \Storage[9][6] , \Storage[9][5] , \Storage[9][4] ,
         \Storage[9][3] , \Storage[9][2] , \Storage[9][1] , \Storage[9][0] ,
         \Storage[8][32] , \Storage[8][31] , \Storage[8][30] ,
         \Storage[8][29] , \Storage[8][28] , \Storage[8][27] ,
         \Storage[8][26] , \Storage[8][25] , \Storage[8][24] ,
         \Storage[8][23] , \Storage[8][22] , \Storage[8][21] ,
         \Storage[8][20] , \Storage[8][19] , \Storage[8][18] ,
         \Storage[8][17] , \Storage[8][16] , \Storage[8][15] ,
         \Storage[8][14] , \Storage[8][13] , \Storage[8][12] ,
         \Storage[8][11] , \Storage[8][10] , \Storage[8][9] , \Storage[8][8] ,
         \Storage[8][7] , \Storage[8][6] , \Storage[8][5] , \Storage[8][4] ,
         \Storage[8][3] , \Storage[8][2] , \Storage[8][1] , \Storage[8][0] ,
         \Storage[7][32] , \Storage[7][31] , \Storage[7][30] ,
         \Storage[7][29] , \Storage[7][28] , \Storage[7][27] ,
         \Storage[7][26] , \Storage[7][25] , \Storage[7][24] ,
         \Storage[7][23] , \Storage[7][22] , \Storage[7][21] ,
         \Storage[7][20] , \Storage[7][19] , \Storage[7][18] ,
         \Storage[7][17] , \Storage[7][16] , \Storage[7][15] ,
         \Storage[7][14] , \Storage[7][13] , \Storage[7][12] ,
         \Storage[7][11] , \Storage[7][10] , \Storage[7][9] , \Storage[7][8] ,
         \Storage[7][7] , \Storage[7][6] , \Storage[7][5] , \Storage[7][4] ,
         \Storage[7][3] , \Storage[7][2] , \Storage[7][1] , \Storage[7][0] ,
         \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N85, N150, N183, N216, N249, N282, N315,
         N348, N381, N414, N447, N480, N513, N546, N579, N612, N645, N678,
         N711, N744, N777, N810, N843, N876, N909, N942, N975, N999, N1041,
         N1074, N1107, N1140, N1173, n107, n108, n109, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  EDFCNQD1 \Storage_reg[26][32]  ( .D(N85), .E(N999), .CP(n204), .CDN(n168), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(n123), .E(N999), .CP(n204), .CDN(n168), 
        .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(n142), .E(N999), .CP(n204), .CDN(n168), 
        .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(n139), .E(N999), .CP(n204), .CDN(n168), 
        .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(n117), .E(N999), .CP(n204), .CDN(n168), 
        .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(n111), .E(N999), .CP(n205), .CDN(n168), 
        .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(n138), .E(N999), .CP(n205), .CDN(n168), 
        .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(n135), .E(N999), .CP(n205), .CDN(n168), 
        .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(n121), .E(N999), .CP(n205), .CDN(n168), 
        .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(n119), .E(N999), .CP(n205), .CDN(n168), 
        .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n134), .E(N999), .CP(n205), .CDN(n169), 
        .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(n133), .E(N999), .CP(n205), .CDN(n169), 
        .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(n115), .E(N999), .CP(n205), .CDN(n169), 
        .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(n113), .E(N999), .CP(n205), .CDN(n169), 
        .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(n130), .E(N999), .CP(n205), .CDN(n169), 
        .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(n127), .E(N999), .CP(n204), .CDN(n169), 
        .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(n112), .E(N999), .CP(n190), .CDN(n169), 
        .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n136), .E(N999), .CP(n217), .CDN(n169), 
        .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n137), .E(N999), .CP(n211), .CDN(n169), 
        .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(n114), .E(N999), .CP(n207), .CDN(n169), 
        .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n116), .E(N999), .CP(n209), .CDN(n169), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(n128), .E(N999), .CP(n216), .CDN(n170), 
        .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(n129), .E(N999), .CP(n200), .CDN(n170), 
        .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n120), .E(N999), .CP(n188), .CDN(n170), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(n140), .E(N999), .CP(n199), .CDN(n170), 
        .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n141), .E(N999), .CP(n195), .CDN(n170), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n124), .E(N999), .CP(n205), .CDN(n170), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n118), .E(N999), .CP(n206), .CDN(n170), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n126), .E(N999), .CP(n188), .CDN(n170), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(n132), .E(N999), .CP(n215), .CDN(n170), 
        .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n125), .E(N999), .CP(n214), .CDN(n170), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(n131), .E(N999), .CP(n216), .CDN(n170), 
        .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n122), .E(N999), .CP(n208), .CDN(n171), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(N85), .E(N942), .CP(n206), .CDN(n167), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(n123), .E(N942), .CP(n206), .CDN(n166), 
        .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(n142), .E(N942), .CP(n206), .CDN(n167), 
        .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(n139), .E(N942), .CP(n206), .CDN(n168), 
        .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(n117), .E(N942), .CP(n206), .CDN(n173), 
        .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(n111), .E(N942), .CP(n206), .CDN(n162), 
        .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(n138), .E(N942), .CP(n206), .CDN(n163), 
        .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(n135), .E(N942), .CP(n206), .CDN(n164), 
        .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(n121), .E(N942), .CP(n206), .CDN(n165), 
        .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(n119), .E(N942), .CP(n209), .CDN(n155), 
        .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n134), .E(N942), .CP(n208), .CDN(n184), 
        .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(n133), .E(N942), .CP(n201), .CDN(n178), 
        .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(n115), .E(N942), .CP(n215), .CDN(n168), 
        .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(n113), .E(N942), .CP(n215), .CDN(n173), 
        .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(n130), .E(N942), .CP(n189), .CDN(n169), 
        .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(n127), .E(N942), .CP(n206), .CDN(n172), 
        .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(n112), .E(N942), .CP(n201), .CDN(n171), 
        .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n136), .E(N942), .CP(n205), .CDN(n170), 
        .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n137), .E(N942), .CP(n202), .CDN(n174), 
        .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(n114), .E(N942), .CP(n212), .CDN(n162), 
        .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n116), .E(N942), .CP(n208), .CDN(n163), 
        .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(n128), .E(N942), .CP(n207), .CDN(n186), 
        .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(n129), .E(N942), .CP(n190), .CDN(n178), 
        .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n120), .E(N942), .CP(n210), .CDN(n183), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(n140), .E(N942), .CP(n208), .CDN(n150), 
        .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n141), .E(N942), .CP(n200), .CDN(n160), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n124), .E(N942), .CP(n217), .CDN(n187), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n118), .E(N942), .CP(n188), .CDN(n181), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n126), .E(N942), .CP(n189), .CDN(n168), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(n132), .E(N942), .CP(n212), .CDN(n173), 
        .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n125), .E(N942), .CP(n213), .CDN(n167), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(n131), .E(N942), .CP(n214), .CDN(n166), 
        .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n122), .E(N942), .CP(n217), .CDN(n178), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(N85), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(n123), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(n142), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(n139), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(n117), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(n111), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(n138), .E(N1140), .CP(n191), .CDN(n156), 
        .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(n135), .E(N1140), .CP(n192), .CDN(n156), 
        .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(n121), .E(N1140), .CP(n192), .CDN(n156), 
        .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(n119), .E(N1140), .CP(n192), .CDN(n156), 
        .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(n134), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(n133), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(n115), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(n113), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(n130), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(n127), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(n112), .E(N1140), .CP(n192), .CDN(n157), 
        .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(n136), .E(N1140), .CP(n193), .CDN(n157), 
        .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(n137), .E(N1140), .CP(n193), .CDN(n157), 
        .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(n114), .E(N1140), .CP(n193), .CDN(n157), 
        .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(n116), .E(N1140), .CP(n193), .CDN(n157), 
        .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(n128), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(n129), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(n120), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(n140), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(n141), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n124), .E(N1140), .CP(n193), .CDN(n158), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(n118), .E(N1140), .CP(n194), .CDN(n158), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(n126), .E(N1140), .CP(n194), .CDN(n158), 
        .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(n132), .E(N1140), .CP(n194), .CDN(n158), 
        .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(n125), .E(N1140), .CP(n194), .CDN(n158), 
        .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(n131), .E(N1140), .CP(n194), .CDN(n158), 
        .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(n122), .E(N1140), .CP(n194), .CDN(n159), 
        .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(N85), .E(N1107), .CP(n194), .CDN(n159), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(n123), .E(N1107), .CP(n194), .CDN(n159), 
        .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(n142), .E(N1107), .CP(n194), .CDN(n159), 
        .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(n139), .E(N1107), .CP(n194), .CDN(n159), 
        .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(n117), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(n111), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(n138), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(n135), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(n121), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(n119), .E(N1107), .CP(n195), .CDN(n159), 
        .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(n134), .E(N1107), .CP(n195), .CDN(n160), 
        .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(n133), .E(N1107), .CP(n195), .CDN(n160), 
        .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(n115), .E(N1107), .CP(n195), .CDN(n160), 
        .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(n113), .E(N1107), .CP(n195), .CDN(n160), 
        .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(n130), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(n127), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(n112), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(n136), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(n137), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(n114), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(n116), .E(N1107), .CP(n196), .CDN(n160), 
        .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(n128), .E(N1107), .CP(n196), .CDN(n161), 
        .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(n129), .E(N1107), .CP(n196), .CDN(n161), 
        .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(n120), .E(N1107), .CP(n196), .CDN(n161), 
        .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(n140), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(n141), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(n124), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(n118), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(n126), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(n132), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(n125), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(n131), .E(N1107), .CP(n197), .CDN(n161), 
        .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(n122), .E(N1107), .CP(n197), .CDN(n162), 
        .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(N85), .E(N1074), .CP(n197), .CDN(n162), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(n123), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(n142), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(n139), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(n117), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(n111), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(n138), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(n135), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(n121), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(n119), .E(N1074), .CP(n198), .CDN(n162), 
        .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n134), .E(N1074), .CP(n198), .CDN(n163), 
        .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(n133), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(n115), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(n113), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(n130), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(n127), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(n112), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(n136), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(n137), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(n114), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n116), .E(N1074), .CP(n199), .CDN(n163), 
        .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(n128), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(n129), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n120), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(n140), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(n141), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n124), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n118), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n126), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(n132), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n125), .E(N1074), .CP(n200), .CDN(n164), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(n131), .E(N1074), .CP(n201), .CDN(n164), 
        .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n122), .E(N1074), .CP(n201), .CDN(n165), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(N85), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(n123), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(n142), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(n139), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(n117), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(n111), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(n138), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(n135), .E(N1041), .CP(n201), .CDN(n165), 
        .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(n121), .E(N1041), .CP(n202), .CDN(n165), 
        .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(n119), .E(N1041), .CP(n202), .CDN(n165), 
        .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n134), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(n133), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(n115), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(n113), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(n130), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(n127), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(n112), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n136), .E(N1041), .CP(n202), .CDN(n166), 
        .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n137), .E(N1041), .CP(n203), .CDN(n166), 
        .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(n114), .E(N1041), .CP(n203), .CDN(n166), 
        .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n116), .E(N1041), .CP(n203), .CDN(n166), 
        .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(n128), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(n129), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n120), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(n140), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n141), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n124), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n118), .E(N1041), .CP(n203), .CDN(n167), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n126), .E(N1041), .CP(n204), .CDN(n167), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(n132), .E(N1041), .CP(n204), .CDN(n167), 
        .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n125), .E(N1041), .CP(n204), .CDN(n167), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(n131), .E(N1041), .CP(n204), .CDN(n167), 
        .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n122), .E(N1041), .CP(n204), .CDN(n168), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(N85), .E(N975), .CP(n214), .CDN(n171), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(n123), .E(N975), .CP(n217), .CDN(n171), 
        .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(n142), .E(N975), .CP(n203), .CDN(n171), 
        .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(n139), .E(N975), .CP(n199), .CDN(n171), 
        .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(n117), .E(N975), .CP(n201), .CDN(n171), 
        .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(n111), .E(N975), .CP(n198), .CDN(n171), 
        .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(n138), .E(N975), .CP(n199), .CDN(n171), 
        .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(n135), .E(N975), .CP(n196), .CDN(n171), 
        .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(n121), .E(N975), .CP(n197), .CDN(n171), 
        .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(n119), .E(N975), .CP(n195), .CDN(n171), 
        .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n134), .E(N975), .CP(n194), .CDN(n172), 
        .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(n133), .E(N975), .CP(n190), .CDN(n172), 
        .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(n115), .E(N975), .CP(n211), .CDN(n172), 
        .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(n113), .E(N975), .CP(n212), .CDN(n172), 
        .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(n130), .E(N975), .CP(n214), .CDN(n172), 
        .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(n127), .E(N975), .CP(n213), .CDN(n172), 
        .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(n112), .E(N975), .CP(n188), .CDN(n172), 
        .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(n136), .E(N975), .CP(n199), .CDN(n172), 
        .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(n137), .E(N975), .CP(n201), .CDN(n172), 
        .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(n114), .E(N975), .CP(n203), .CDN(n172), 
        .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n116), .E(N975), .CP(n203), .CDN(n172), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(n128), .E(N975), .CP(n198), .CDN(n173), 
        .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(n129), .E(N975), .CP(n208), .CDN(n173), 
        .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n120), .E(N975), .CP(n207), .CDN(n173), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(n140), .E(N975), .CP(n210), .CDN(n173), 
        .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(n141), .E(N975), .CP(n211), .CDN(n173), 
        .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n124), .E(N975), .CP(n209), .CDN(n173), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n118), .E(N975), .CP(n212), .CDN(n173), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n126), .E(N975), .CP(n188), .CDN(n173), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(n132), .E(N975), .CP(n217), .CDN(n173), 
        .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n125), .E(N975), .CP(n213), .CDN(n173), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(n131), .E(N975), .CP(ClockW), .CDN(n173), 
        .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n122), .E(N975), .CP(n206), .CDN(n179), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(N85), .E(N876), .CP(n206), .CDN(n176), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n123), .E(N876), .CP(n190), .CDN(n176), 
        .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n142), .E(N876), .CP(n188), .CDN(n176), 
        .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(n139), .E(N876), .CP(n209), .CDN(n176), 
        .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(n117), .E(N876), .CP(n194), .CDN(n176), 
        .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(n111), .E(N876), .CP(n214), .CDN(n176), 
        .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n138), .E(N876), .CP(n200), .CDN(n176), 
        .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(n135), .E(N876), .CP(n192), .CDN(n176), 
        .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(n121), .E(N876), .CP(n191), .CDN(n176), 
        .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(n119), .E(N876), .CP(n194), .CDN(n176), 
        .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(n134), .E(N876), .CP(n215), .CDN(n177), 
        .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(n133), .E(N876), .CP(n216), .CDN(n177), 
        .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(n115), .E(N876), .CP(n213), .CDN(n177), 
        .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(n113), .E(N876), .CP(n191), .CDN(n177), 
        .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(n130), .E(N876), .CP(n190), .CDN(n177), 
        .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n127), .E(N876), .CP(n189), .CDN(n177), 
        .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(n112), .E(N876), .CP(n188), .CDN(n177), 
        .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(n136), .E(N876), .CP(n212), .CDN(n177), 
        .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(n137), .E(N876), .CP(n206), .CDN(n177), 
        .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n114), .E(N876), .CP(n189), .CDN(n177), 
        .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(n116), .E(N876), .CP(n202), .CDN(n177), 
        .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(n128), .E(N876), .CP(n192), .CDN(n162), 
        .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(n129), .E(N876), .CP(n214), .CDN(n178), 
        .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(n120), .E(N876), .CP(n196), .CDN(n177), 
        .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(n140), .E(N876), .CP(n201), .CDN(n175), 
        .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(n141), .E(N876), .CP(n210), .CDN(n174), 
        .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n124), .E(N876), .CP(n209), .CDN(n162), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n118), .E(N876), .CP(n208), .CDN(n163), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(n126), .E(N876), .CP(n207), .CDN(n164), 
        .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(n132), .E(N876), .CP(n212), .CDN(n165), 
        .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(n125), .E(N876), .CP(n190), .CDN(n166), 
        .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(n131), .E(N876), .CP(n206), .CDN(n167), 
        .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n122), .E(N876), .CP(n193), .CDN(n175), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(N85), .E(N843), .CP(n206), .CDN(n177), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n123), .E(N843), .CP(n212), .CDN(n150), 
        .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n142), .E(N843), .CP(n197), .CDN(n183), 
        .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n139), .E(N843), .CP(n199), .CDN(n181), 
        .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n117), .E(N843), .CP(n198), .CDN(n159), 
        .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(n111), .E(N843), .CP(n204), .CDN(n187), 
        .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n138), .E(N843), .CP(n205), .CDN(n154), 
        .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n135), .E(N843), .CP(n202), .CDN(n150), 
        .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n121), .E(N843), .CP(n203), .CDN(n186), 
        .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(n119), .E(N843), .CP(n201), .CDN(n161), 
        .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n134), .E(N843), .CP(n191), .CDN(n166), 
        .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n133), .E(N843), .CP(n192), .CDN(n162), 
        .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n115), .E(N843), .CP(n193), .CDN(n163), 
        .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n113), .E(N843), .CP(n199), .CDN(n164), 
        .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(n130), .E(N843), .CP(n198), .CDN(n165), 
        .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n127), .E(N843), .CP(n197), .CDN(n153), 
        .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n112), .E(N843), .CP(n196), .CDN(n180), 
        .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n136), .E(N843), .CP(n195), .CDN(n174), 
        .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n137), .E(N843), .CP(n194), .CDN(n167), 
        .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n114), .E(N843), .CP(n208), .CDN(n178), 
        .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n116), .E(N843), .CP(n189), .CDN(n152), 
        .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n128), .E(N843), .CP(n204), .CDN(n160), 
        .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n129), .E(N843), .CP(n216), .CDN(n159), 
        .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n120), .E(N843), .CP(n217), .CDN(n187), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n140), .E(N843), .CP(ClockW), .CDN(n154), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n141), .E(N843), .CP(n215), .CDN(n186), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n124), .E(N843), .CP(n195), .CDN(n185), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n118), .E(N843), .CP(n198), .CDN(n108), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n126), .E(N843), .CP(n193), .CDN(n184), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(n132), .E(N843), .CP(n196), .CDN(n179), 
        .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n125), .E(N843), .CP(n188), .CDN(n184), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n131), .E(N843), .CP(n211), .CDN(n180), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n122), .E(N843), .CP(n211), .CDN(n173), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N85), .E(N744), .CP(n194), .CDN(n170), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(n123), .E(N744), .CP(n211), .CDN(n168), 
        .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(n142), .E(N744), .CP(n203), .CDN(n175), 
        .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(n139), .E(N744), .CP(n197), .CDN(n176), 
        .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(n117), .E(N744), .CP(n205), .CDN(n177), 
        .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(n111), .E(N744), .CP(n201), .CDN(n178), 
        .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(n138), .E(N744), .CP(n200), .CDN(n152), 
        .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(n135), .E(N744), .CP(n211), .CDN(n154), 
        .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(n121), .E(N744), .CP(n202), .CDN(n155), 
        .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(n119), .E(N744), .CP(n206), .CDN(n154), 
        .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n134), .E(N744), .CP(n191), .CDN(n184), 
        .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(n133), .E(N744), .CP(n188), .CDN(n155), 
        .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(n115), .E(N744), .CP(n204), .CDN(n171), 
        .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(n113), .E(N744), .CP(n217), .CDN(n172), 
        .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(n130), .E(N744), .CP(n214), .CDN(n162), 
        .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(n127), .E(N744), .CP(n213), .CDN(n180), 
        .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(n112), .E(N744), .CP(n212), .CDN(n170), 
        .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(n136), .E(N744), .CP(n211), .CDN(n161), 
        .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(n137), .E(N744), .CP(n210), .CDN(n183), 
        .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n114), .E(N744), .CP(n209), .CDN(n179), 
        .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n116), .E(N744), .CP(n215), .CDN(n178), 
        .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(n128), .E(N744), .CP(n210), .CDN(n157), 
        .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(n129), .E(N744), .CP(n208), .CDN(n177), 
        .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n120), .E(N744), .CP(n203), .CDN(n167), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(n140), .E(N744), .CP(n211), .CDN(n182), 
        .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(n141), .E(N744), .CP(n195), .CDN(n182), 
        .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n124), .E(N744), .CP(n217), .CDN(n178), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n118), .E(N744), .CP(n193), .CDN(n160), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n126), .E(N744), .CP(n196), .CDN(n179), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(n132), .E(N744), .CP(n212), .CDN(n183), 
        .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n125), .E(N744), .CP(n201), .CDN(n181), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(n131), .E(N744), .CP(n190), .CDN(n180), 
        .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n122), .E(N744), .CP(n217), .CDN(n150), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(N85), .E(N711), .CP(n207), .CDN(n159), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n123), .E(N711), .CP(n210), .CDN(n158), 
        .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n142), .E(N711), .CP(n205), .CDN(n159), 
        .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(n139), .E(N711), .CP(n210), .CDN(n160), 
        .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(n117), .E(N711), .CP(n214), .CDN(n161), 
        .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n111), .E(N711), .CP(n194), .CDN(n162), 
        .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n138), .E(N711), .CP(n211), .CDN(n163), 
        .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(n135), .E(N711), .CP(n195), .CDN(n166), 
        .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(n121), .E(N711), .CP(n210), .CDN(n167), 
        .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n119), .E(N711), .CP(n214), .CDN(n170), 
        .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n134), .E(N711), .CP(n192), .CDN(n161), 
        .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(n133), .E(N711), .CP(ClockW), .CDN(n176), 
        .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(n115), .E(N711), .CP(n215), .CDN(n176), 
        .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(n113), .E(N711), .CP(n216), .CDN(n151), 
        .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n130), .E(N711), .CP(n204), .CDN(n152), 
        .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n127), .E(N711), .CP(n190), .CDN(n168), 
        .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(n112), .E(N711), .CP(n207), .CDN(n183), 
        .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(n136), .E(N711), .CP(n194), .CDN(n181), 
        .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(n137), .E(N711), .CP(n204), .CDN(n180), 
        .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n114), .E(N711), .CP(n216), .CDN(n164), 
        .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n116), .E(N711), .CP(n199), .CDN(n179), 
        .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(n128), .E(N711), .CP(n198), .CDN(n158), 
        .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(n129), .E(N711), .CP(n197), .CDN(n160), 
        .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n120), .E(N711), .CP(n196), .CDN(n172), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(n140), .E(N711), .CP(n195), .CDN(n150), 
        .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(n141), .E(N711), .CP(n194), .CDN(n154), 
        .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n124), .E(N711), .CP(n192), .CDN(n169), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n118), .E(N711), .CP(n193), .CDN(n184), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n126), .E(N711), .CP(n205), .CDN(n185), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n132), .E(N711), .CP(n206), .CDN(n186), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n125), .E(N711), .CP(n194), .CDN(n152), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(n131), .E(N711), .CP(n212), .CDN(n156), 
        .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n122), .E(N711), .CP(n189), .CDN(n166), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N85), .E(N612), .CP(n214), .CDN(n156), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n123), .E(N612), .CP(n194), .CDN(n156), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n142), .E(N612), .CP(n195), .CDN(n164), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n139), .E(N612), .CP(n196), .CDN(n165), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n117), .E(N612), .CP(n197), .CDN(n169), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n111), .E(N612), .CP(n198), .CDN(n168), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n138), .E(N612), .CP(n199), .CDN(n167), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n135), .E(N612), .CP(n192), .CDN(n166), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n121), .E(N612), .CP(n193), .CDN(n173), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n119), .E(N612), .CP(n196), .CDN(n171), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n134), .E(N612), .CP(n210), .CDN(n187), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n133), .E(N612), .CP(n188), .CDN(n167), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n115), .E(N612), .CP(n189), .CDN(n160), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n113), .E(N612), .CP(n190), .CDN(n153), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n130), .E(N612), .CP(n191), .CDN(n181), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n127), .E(N612), .CP(n192), .CDN(n160), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n112), .E(N612), .CP(n193), .CDN(n169), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n136), .E(N612), .CP(n194), .CDN(n153), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n137), .E(N612), .CP(n195), .CDN(n181), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n114), .E(N612), .CP(n194), .CDN(n186), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n116), .E(N612), .CP(n216), .CDN(n161), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n128), .E(N612), .CP(n191), .CDN(n185), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n129), .E(N612), .CP(n204), .CDN(n177), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n120), .E(N612), .CP(n201), .CDN(n179), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n140), .E(N612), .CP(n204), .CDN(n162), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n141), .E(N612), .CP(n205), .CDN(n178), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n124), .E(N612), .CP(n213), .CDN(n150), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n118), .E(N612), .CP(n203), .CDN(n156), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n126), .E(N612), .CP(n189), .CDN(n108), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n132), .E(N612), .CP(n214), .CDN(n169), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n125), .E(N612), .CP(n200), .CDN(n150), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n131), .E(N612), .CP(n197), .CDN(n184), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n122), .E(N612), .CP(n215), .CDN(n180), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N85), .E(N579), .CP(n190), .CDN(n165), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n123), .E(N579), .CP(n200), .CDN(n172), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n142), .E(N579), .CP(n189), .CDN(n175), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n139), .E(N579), .CP(n190), .CDN(n182), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n117), .E(N579), .CP(n198), .CDN(n183), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n111), .E(N579), .CP(n215), .CDN(n182), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n138), .E(N579), .CP(n206), .CDN(n175), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n135), .E(N579), .CP(n190), .CDN(n151), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n121), .E(N579), .CP(n204), .CDN(n181), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n119), .E(N579), .CP(n212), .CDN(n174), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n134), .E(N579), .CP(n215), .CDN(n178), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n133), .E(N579), .CP(n196), .CDN(n180), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n115), .E(N579), .CP(n198), .CDN(n172), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n113), .E(N579), .CP(n209), .CDN(n184), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n130), .E(N579), .CP(n211), .CDN(n156), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n127), .E(N579), .CP(n198), .CDN(n153), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n112), .E(N579), .CP(ClockW), .CDN(n176), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n136), .E(N579), .CP(n214), .CDN(n150), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n137), .E(N579), .CP(n213), .CDN(n171), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n114), .E(N579), .CP(n209), .CDN(n168), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n116), .E(N579), .CP(n204), .CDN(n169), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n128), .E(N579), .CP(n206), .CDN(n169), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n129), .E(N579), .CP(n191), .CDN(n171), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n120), .E(N579), .CP(n212), .CDN(n158), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n140), .E(N579), .CP(ClockW), .CDN(n159), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n141), .E(N579), .CP(n206), .CDN(n160), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n124), .E(N579), .CP(ClockW), .CDN(n161), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n118), .E(N579), .CP(n203), .CDN(n162), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n126), .E(N579), .CP(n200), .CDN(n163), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n132), .E(N579), .CP(n189), .CDN(n164), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n125), .E(N579), .CP(n214), .CDN(n165), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n131), .E(N579), .CP(n213), .CDN(n166), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n122), .E(N579), .CP(n207), .CDN(n168), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N85), .E(N480), .CP(ClockW), .CDN(n156), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n123), .E(N480), .CP(n210), .CDN(n171), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n142), .E(N480), .CP(n214), .CDN(n154), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n139), .E(N480), .CP(n197), .CDN(n155), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n117), .E(N480), .CP(n203), .CDN(n156), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n111), .E(N480), .CP(n194), .CDN(n177), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n138), .E(N480), .CP(n195), .CDN(n182), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n135), .E(N480), .CP(n208), .CDN(n169), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n121), .E(N480), .CP(n208), .CDN(n161), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n119), .E(N480), .CP(n195), .CDN(n184), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n134), .E(N480), .CP(n208), .CDN(n151), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n133), .E(N480), .CP(n207), .CDN(n160), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n115), .E(N480), .CP(n212), .CDN(n182), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n113), .E(N480), .CP(n209), .CDN(n175), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n130), .E(N480), .CP(n193), .CDN(n171), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n127), .E(N480), .CP(n191), .CDN(n178), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n112), .E(N480), .CP(n209), .CDN(n153), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n136), .E(N480), .CP(n196), .CDN(n183), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n137), .E(N480), .CP(n213), .CDN(n155), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n114), .E(N480), .CP(n214), .CDN(n154), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n116), .E(N480), .CP(n215), .CDN(n164), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n128), .E(N480), .CP(n190), .CDN(n176), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n129), .E(N480), .CP(n206), .CDN(n181), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n120), .E(N480), .CP(n216), .CDN(n187), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n140), .E(N480), .CP(n203), .CDN(n151), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n141), .E(N480), .CP(n205), .CDN(n180), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n124), .E(N480), .CP(ClockW), .CDN(n180), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n118), .E(N480), .CP(n211), .CDN(n164), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n126), .E(N480), .CP(n201), .CDN(n169), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n132), .E(N480), .CP(ClockW), .CDN(n185), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n125), .E(N480), .CP(n214), .CDN(n174), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n131), .E(N480), .CP(n217), .CDN(n175), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n122), .E(N480), .CP(n212), .CDN(n180), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N85), .E(N447), .CP(n213), .CDN(n169), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n123), .E(N447), .CP(n214), .CDN(n177), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n142), .E(N447), .CP(n209), .CDN(n162), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n139), .E(N447), .CP(n210), .CDN(n163), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n117), .E(N447), .CP(n216), .CDN(n164), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n111), .E(N447), .CP(n202), .CDN(n165), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n138), .E(N447), .CP(ClockW), .CDN(n158), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n135), .E(N447), .CP(n217), .CDN(n159), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n121), .E(N447), .CP(n214), .CDN(n160), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n119), .E(N447), .CP(n213), .CDN(n161), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n134), .E(N447), .CP(n212), .CDN(n174), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n133), .E(N447), .CP(n211), .CDN(n184), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n115), .E(N447), .CP(n210), .CDN(n182), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n113), .E(N447), .CP(n209), .CDN(n177), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n130), .E(N447), .CP(n206), .CDN(n178), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n127), .E(N447), .CP(n206), .CDN(n180), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n112), .E(N447), .CP(n195), .CDN(n183), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n136), .E(N447), .CP(n188), .CDN(n152), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n137), .E(N447), .CP(n191), .CDN(n168), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n114), .E(N447), .CP(n212), .CDN(n157), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n116), .E(N447), .CP(n205), .CDN(n176), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n128), .E(N447), .CP(n208), .CDN(n185), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n129), .E(N447), .CP(n217), .CDN(n157), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n120), .E(N447), .CP(n202), .CDN(n108), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n140), .E(N447), .CP(ClockW), .CDN(n174), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n141), .E(N447), .CP(n193), .CDN(n186), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n124), .E(N447), .CP(ClockW), .CDN(n150), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n118), .E(N447), .CP(n216), .CDN(n170), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n126), .E(N447), .CP(n199), .CDN(n178), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n132), .E(N447), .CP(n196), .CDN(n161), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n125), .E(N447), .CP(n202), .CDN(n179), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n131), .E(N447), .CP(n193), .CDN(n151), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n122), .E(N447), .CP(n216), .CDN(n168), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N85), .E(N348), .CP(n208), .CDN(n156), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n123), .E(N348), .CP(n197), .CDN(n177), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n142), .E(N348), .CP(n200), .CDN(n155), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n139), .E(N348), .CP(n197), .CDN(n180), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n117), .E(N348), .CP(n205), .CDN(n171), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n111), .E(N348), .CP(n200), .CDN(n181), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n138), .E(N348), .CP(n193), .CDN(n160), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n135), .E(N348), .CP(n193), .CDN(n175), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n121), .E(N348), .CP(n217), .CDN(n170), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n119), .E(N348), .CP(n192), .CDN(n167), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n134), .E(N348), .CP(n192), .CDN(n151), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n133), .E(N348), .CP(n205), .CDN(n157), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n115), .E(N348), .CP(n204), .CDN(n183), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n113), .E(N348), .CP(n209), .CDN(n183), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n130), .E(N348), .CP(n209), .CDN(n182), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n127), .E(N348), .CP(n208), .CDN(n176), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n112), .E(N348), .CP(n188), .CDN(n179), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n136), .E(N348), .CP(n217), .CDN(n178), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n137), .E(N348), .CP(n214), .CDN(n186), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n114), .E(N348), .CP(n213), .CDN(n157), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n116), .E(N348), .CP(n212), .CDN(n152), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n128), .E(N348), .CP(n211), .CDN(n173), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n129), .E(N348), .CP(n210), .CDN(n174), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n120), .E(N348), .CP(n209), .CDN(n187), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n140), .E(N348), .CP(n213), .CDN(n152), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n141), .E(N348), .CP(n208), .CDN(n184), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n124), .E(N348), .CP(n205), .CDN(n178), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n118), .E(N348), .CP(n200), .CDN(n181), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n126), .E(N348), .CP(n202), .CDN(n154), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n132), .E(N348), .CP(n203), .CDN(n186), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n125), .E(N348), .CP(n194), .CDN(n185), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n131), .E(N348), .CP(n203), .CDN(n163), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n122), .E(N348), .CP(n213), .CDN(n178), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N85), .E(N315), .CP(n210), .CDN(n168), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n123), .E(N315), .CP(n207), .CDN(n157), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n142), .E(N315), .CP(n217), .CDN(n184), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n139), .E(N315), .CP(n201), .CDN(n179), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n117), .E(N315), .CP(n193), .CDN(n108), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n111), .E(N315), .CP(n205), .CDN(n181), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n138), .E(N315), .CP(n195), .CDN(n180), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n135), .E(N315), .CP(n211), .CDN(n183), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n121), .E(N315), .CP(n196), .CDN(n153), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n119), .E(N315), .CP(n209), .CDN(n179), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n134), .E(N315), .CP(n195), .CDN(n160), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n133), .E(N315), .CP(n207), .CDN(n174), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n115), .E(N315), .CP(n202), .CDN(n187), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n113), .E(N315), .CP(n205), .CDN(n169), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n130), .E(N315), .CP(n203), .CDN(n156), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n127), .E(N315), .CP(ClockW), .CDN(n172), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n112), .E(N315), .CP(n208), .CDN(n152), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n136), .E(N315), .CP(n209), .CDN(n108), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n137), .E(N315), .CP(n192), .CDN(n174), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n114), .E(N315), .CP(n214), .CDN(n163), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n116), .E(N315), .CP(n192), .CDN(n181), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n128), .E(N315), .CP(n208), .CDN(n157), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n129), .E(N315), .CP(n191), .CDN(n187), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n120), .E(N315), .CP(n214), .CDN(n156), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n140), .E(N315), .CP(n207), .CDN(n151), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n141), .E(N315), .CP(ClockW), .CDN(n170), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n124), .E(N315), .CP(n216), .CDN(n171), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n118), .E(N315), .CP(n188), .CDN(n163), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n126), .E(N315), .CP(n198), .CDN(n187), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n132), .E(N315), .CP(n216), .CDN(n177), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n125), .E(N315), .CP(n213), .CDN(n159), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n131), .E(N315), .CP(n210), .CDN(n164), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n122), .E(N315), .CP(n208), .CDN(n153), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(N216), .CP(n193), .CDN(n165), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n123), .E(N216), .CP(n199), .CDN(n185), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n142), .E(N216), .CP(n215), .CDN(n178), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n139), .E(N216), .CP(n217), .CDN(n187), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n117), .E(N216), .CP(n189), .CDN(n184), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n111), .E(N216), .CP(n190), .CDN(n166), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n138), .E(N216), .CP(n188), .CDN(n168), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n135), .E(N216), .CP(n206), .CDN(n185), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n121), .E(N216), .CP(n199), .CDN(n186), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n119), .E(N216), .CP(n202), .CDN(n187), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n134), .E(N216), .CP(n189), .CDN(n153), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n133), .E(N216), .CP(n209), .CDN(n187), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n115), .E(N216), .CP(n201), .CDN(n108), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n113), .E(N216), .CP(n208), .CDN(n184), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n130), .E(N216), .CP(n212), .CDN(n185), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n127), .E(N216), .CP(n204), .CDN(n186), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n112), .E(N216), .CP(n192), .CDN(n175), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n136), .E(N216), .CP(n204), .CDN(n171), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n137), .E(N216), .CP(n196), .CDN(n157), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n114), .E(N216), .CP(n204), .CDN(n150), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n116), .E(N216), .CP(n192), .CDN(n186), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n128), .E(N216), .CP(n210), .CDN(n187), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n129), .E(N216), .CP(n207), .CDN(n150), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n120), .E(N216), .CP(n208), .CDN(n165), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n140), .E(N216), .CP(n207), .CDN(n153), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n141), .E(N216), .CP(n193), .CDN(n182), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n124), .E(N216), .CP(n209), .CDN(n164), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n118), .E(N216), .CP(n216), .CDN(n108), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n126), .E(N216), .CP(n197), .CDN(n182), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n132), .E(N216), .CP(n205), .CDN(n182), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n125), .E(N216), .CP(n200), .CDN(n186), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n131), .E(N216), .CP(n193), .CDN(n184), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n122), .E(N216), .CP(n210), .CDN(n182), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N85), .E(N183), .CP(n191), .CDN(n184), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n123), .E(N183), .CP(n202), .CDN(n156), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n142), .E(N183), .CP(n211), .CDN(n154), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n139), .E(N183), .CP(n210), .CDN(n172), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n117), .E(N183), .CP(n209), .CDN(n156), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n111), .E(N183), .CP(n214), .CDN(n155), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n138), .E(N183), .CP(n213), .CDN(n185), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n135), .E(N183), .CP(n212), .CDN(n186), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n121), .E(N183), .CP(n207), .CDN(n174), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n119), .E(N183), .CP(n211), .CDN(n158), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n134), .E(N183), .CP(n197), .CDN(n179), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n133), .E(N183), .CP(n197), .CDN(n108), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n115), .E(N183), .CP(n197), .CDN(n171), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n113), .E(N183), .CP(n213), .CDN(n183), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n130), .E(N183), .CP(n207), .CDN(n182), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n127), .E(N183), .CP(n207), .CDN(n170), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n112), .E(N183), .CP(n202), .CDN(n184), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n136), .E(N183), .CP(n212), .CDN(n172), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n137), .E(N183), .CP(n188), .CDN(n162), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n114), .E(N183), .CP(n198), .CDN(n152), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n116), .E(N183), .CP(n208), .CDN(n167), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n128), .E(N183), .CP(n208), .CDN(n178), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n129), .E(N183), .CP(n207), .CDN(n179), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n120), .E(N183), .CP(n194), .CDN(n180), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n140), .E(N183), .CP(n200), .CDN(n152), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n141), .E(N183), .CP(n212), .CDN(n161), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n124), .E(N183), .CP(n188), .CDN(n152), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n118), .E(N183), .CP(n202), .CDN(n164), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n126), .E(N183), .CP(n189), .CDN(n180), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n132), .E(N183), .CP(n200), .CDN(n181), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n125), .E(N183), .CP(n216), .CDN(n157), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n131), .E(N183), .CP(n214), .CDN(n179), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n122), .E(N183), .CP(n209), .CDN(n155), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n118), .E(N150), .CP(n202), .CDN(n185), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n126), .E(N150), .CP(n213), .CDN(n181), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n132), .E(N150), .CP(n203), .CDN(n164), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n125), .E(N150), .CP(n200), .CDN(n184), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n131), .E(N150), .CP(n215), .CDN(n187), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n122), .E(N150), .CP(n193), .CDN(n179), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(N85), .E(N909), .CP(n199), .CDN(n165), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(n123), .E(N909), .CP(n216), .CDN(n177), 
        .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(n142), .E(N909), .CP(n215), .CDN(n161), 
        .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(n139), .E(N909), .CP(n211), .CDN(n159), 
        .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(n117), .E(N909), .CP(n208), .CDN(n158), 
        .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(n111), .E(N909), .CP(n194), .CDN(n176), 
        .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(n138), .E(N909), .CP(n195), .CDN(n182), 
        .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(n135), .E(N909), .CP(n197), .CDN(n179), 
        .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(n121), .E(N909), .CP(n196), .CDN(n156), 
        .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(n119), .E(N909), .CP(n195), .CDN(n180), 
        .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n134), .E(N909), .CP(n198), .CDN(n174), 
        .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(n133), .E(N909), .CP(n192), .CDN(n174), 
        .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(n115), .E(N909), .CP(n193), .CDN(n174), 
        .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(n113), .E(N909), .CP(n190), .CDN(n174), 
        .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(n130), .E(N909), .CP(n191), .CDN(n174), 
        .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(n127), .E(N909), .CP(n188), .CDN(n174), 
        .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(n112), .E(N909), .CP(n213), .CDN(n174), 
        .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(n136), .E(N909), .CP(n209), .CDN(n174), 
        .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(n137), .E(N909), .CP(n210), .CDN(n174), 
        .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n114), .E(N909), .CP(n214), .CDN(n174), 
        .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n116), .E(N909), .CP(n216), .CDN(n174), 
        .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(n128), .E(N909), .CP(n215), .CDN(n175), 
        .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(n129), .E(N909), .CP(n210), .CDN(n175), 
        .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n120), .E(N909), .CP(n217), .CDN(n175), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(n140), .E(N909), .CP(n202), .CDN(n175), 
        .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(n141), .E(N909), .CP(n204), .CDN(n175), 
        .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n124), .E(N909), .CP(n189), .CDN(n175), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n118), .E(N909), .CP(n216), .CDN(n175), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n126), .E(N909), .CP(n216), .CDN(n175), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(n132), .E(N909), .CP(n190), .CDN(n175), 
        .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n125), .E(N909), .CP(n215), .CDN(n175), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(n131), .E(N909), .CP(n217), .CDN(n175), 
        .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n122), .E(N909), .CP(n189), .CDN(n176), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N85), .E(N810), .CP(n196), .CDN(n158), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(n123), .E(N810), .CP(n215), .CDN(n187), 
        .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(n142), .E(N810), .CP(n217), .CDN(n159), 
        .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(n139), .E(N810), .CP(n190), .CDN(n151), 
        .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(n117), .E(N810), .CP(n208), .CDN(n152), 
        .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(n111), .E(N810), .CP(n207), .CDN(n153), 
        .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(n138), .E(N810), .CP(n197), .CDN(n176), 
        .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(n135), .E(N810), .CP(n214), .CDN(n159), 
        .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(n121), .E(N810), .CP(n206), .CDN(n167), 
        .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(n119), .E(N810), .CP(n197), .CDN(n181), 
        .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n134), .E(N810), .CP(n211), .CDN(n161), 
        .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(n133), .E(N810), .CP(n196), .CDN(n166), 
        .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(n115), .E(N810), .CP(n212), .CDN(n185), 
        .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(n113), .E(N810), .CP(n213), .CDN(n163), 
        .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(n130), .E(N810), .CP(n214), .CDN(n169), 
        .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(n127), .E(N810), .CP(n209), .CDN(n176), 
        .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(n112), .E(N810), .CP(n210), .CDN(n158), 
        .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(n136), .E(N810), .CP(n188), .CDN(n172), 
        .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(n137), .E(N810), .CP(n189), .CDN(n171), 
        .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(n114), .E(N810), .CP(n190), .CDN(n170), 
        .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n116), .E(N810), .CP(n191), .CDN(n169), 
        .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(n128), .E(N810), .CP(n193), .CDN(n158), 
        .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(n129), .E(N810), .CP(n192), .CDN(n163), 
        .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n120), .E(N810), .CP(n213), .CDN(n164), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(n140), .E(N810), .CP(n198), .CDN(n165), 
        .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(n141), .E(N810), .CP(n199), .CDN(n169), 
        .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n124), .E(N810), .CP(n196), .CDN(n168), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n118), .E(N810), .CP(n197), .CDN(n170), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n126), .E(N810), .CP(n198), .CDN(n166), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(n132), .E(N810), .CP(n207), .CDN(n170), 
        .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n125), .E(N810), .CP(n207), .CDN(n171), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(n131), .E(N810), .CP(n192), .CDN(n172), 
        .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n122), .E(N810), .CP(n216), .CDN(n185), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(N85), .E(N777), .CP(n215), .CDN(n157), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(n123), .E(N777), .CP(n191), .CDN(n153), 
        .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(n142), .E(N777), .CP(n211), .CDN(n151), 
        .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(n139), .E(N777), .CP(n203), .CDN(n182), 
        .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(n117), .E(N777), .CP(n197), .CDN(n172), 
        .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(n111), .E(N777), .CP(n216), .CDN(n173), 
        .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(n138), .E(N777), .CP(n191), .CDN(n183), 
        .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(n135), .E(N777), .CP(n205), .CDN(n171), 
        .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(n121), .E(N777), .CP(n208), .CDN(n179), 
        .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(n119), .E(N777), .CP(n190), .CDN(n178), 
        .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n134), .E(N777), .CP(n206), .CDN(n167), 
        .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(n133), .E(N777), .CP(n213), .CDN(n185), 
        .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(n115), .E(N777), .CP(n195), .CDN(n181), 
        .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(n113), .E(N777), .CP(n194), .CDN(n180), 
        .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(n130), .E(N777), .CP(n212), .CDN(n175), 
        .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(n127), .E(N777), .CP(n198), .CDN(n178), 
        .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(n112), .E(N777), .CP(n199), .CDN(n182), 
        .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(n136), .E(N777), .CP(n189), .CDN(n150), 
        .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(n137), .E(N777), .CP(n188), .CDN(n182), 
        .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(n114), .E(N777), .CP(n191), .CDN(n161), 
        .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n116), .E(N777), .CP(n190), .CDN(n170), 
        .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(n128), .E(N777), .CP(n193), .CDN(n174), 
        .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(n129), .E(N777), .CP(n192), .CDN(n186), 
        .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n120), .E(N777), .CP(n213), .CDN(n161), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(n140), .E(N777), .CP(n192), .CDN(n160), 
        .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(n141), .E(N777), .CP(n210), .CDN(n159), 
        .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n124), .E(N777), .CP(n209), .CDN(n158), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n118), .E(N777), .CP(n212), .CDN(n165), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n126), .E(N777), .CP(n213), .CDN(n164), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(n132), .E(N777), .CP(n195), .CDN(n163), 
        .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n125), .E(N777), .CP(n210), .CDN(n162), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(n131), .E(N777), .CP(n199), .CDN(n170), 
        .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n122), .E(N777), .CP(n211), .CDN(n155), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(N678), .CP(n195), .CDN(n157), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(n123), .E(N678), .CP(n200), .CDN(n153), 
        .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(n142), .E(N678), .CP(n201), .CDN(n169), 
        .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(n139), .E(N678), .CP(n202), .CDN(n179), 
        .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(n117), .E(N678), .CP(n195), .CDN(n154), 
        .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(n111), .E(N678), .CP(n205), .CDN(n150), 
        .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(n138), .E(N678), .CP(n215), .CDN(n184), 
        .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(n135), .E(N678), .CP(n211), .CDN(n185), 
        .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(n121), .E(N678), .CP(n214), .CDN(n179), 
        .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(n119), .E(N678), .CP(n192), .CDN(n152), 
        .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n134), .E(N678), .CP(n194), .CDN(n156), 
        .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(n133), .E(N678), .CP(n195), .CDN(n183), 
        .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(n115), .E(N678), .CP(n217), .CDN(n160), 
        .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(n113), .E(N678), .CP(n206), .CDN(n178), 
        .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(n130), .E(N678), .CP(n192), .CDN(n180), 
        .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(n127), .E(N678), .CP(n188), .CDN(n181), 
        .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(n112), .E(N678), .CP(n216), .CDN(n180), 
        .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(n136), .E(N678), .CP(n210), .CDN(n182), 
        .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(n137), .E(N678), .CP(n198), .CDN(n150), 
        .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(n114), .E(N678), .CP(n199), .CDN(n153), 
        .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n116), .E(N678), .CP(n216), .CDN(n155), 
        .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(n128), .E(N678), .CP(n191), .CDN(n155), 
        .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(n129), .E(N678), .CP(n206), .CDN(n151), 
        .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n120), .E(N678), .CP(n217), .CDN(n158), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(n140), .E(N678), .CP(n210), .CDN(n170), 
        .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(n141), .E(N678), .CP(n214), .CDN(n169), 
        .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n124), .E(N678), .CP(n211), .CDN(n168), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n118), .E(N678), .CP(n199), .CDN(n185), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n126), .E(N678), .CP(n205), .CDN(n161), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(n132), .E(N678), .CP(n204), .CDN(n160), 
        .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n125), .E(N678), .CP(n195), .CDN(n159), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(n131), .E(N678), .CP(n189), .CDN(n176), 
        .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n122), .E(N678), .CP(n194), .CDN(n164), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N85), .E(N645), .CP(n192), .CDN(n163), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n123), .E(N645), .CP(n194), .CDN(n162), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n142), .E(N645), .CP(n191), .CDN(n171), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n139), .E(N645), .CP(n216), .CDN(n172), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n117), .E(N645), .CP(ClockW), .CDN(n173), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n111), .E(N645), .CP(ClockW), .CDN(n166), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n138), .E(N645), .CP(n210), .CDN(n174), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n135), .E(N645), .CP(n201), .CDN(n175), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n121), .E(N645), .CP(n210), .CDN(n177), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n119), .E(N645), .CP(n193), .CDN(n154), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n134), .E(N645), .CP(n196), .CDN(n158), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n133), .E(N645), .CP(n201), .CDN(n186), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n115), .E(N645), .CP(n197), .CDN(n186), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n113), .E(N645), .CP(n193), .CDN(n187), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n130), .E(N645), .CP(n213), .CDN(n176), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n127), .E(N645), .CP(n197), .CDN(n172), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n112), .E(N645), .CP(n203), .CDN(n179), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n136), .E(N645), .CP(n199), .CDN(n154), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n137), .E(N645), .CP(n207), .CDN(n155), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n114), .E(N645), .CP(n208), .CDN(n156), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n116), .E(N645), .CP(n198), .CDN(n157), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n128), .E(N645), .CP(n195), .CDN(n163), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n129), .E(N645), .CP(n209), .CDN(n166), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n120), .E(N645), .CP(n200), .CDN(n174), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n140), .E(N645), .CP(ClockW), .CDN(n175), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n141), .E(N645), .CP(n211), .CDN(n177), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n124), .E(N645), .CP(n200), .CDN(n166), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n118), .E(N645), .CP(n198), .CDN(n183), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n126), .E(N645), .CP(n201), .CDN(n155), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n132), .E(N645), .CP(n209), .CDN(n159), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n125), .E(N645), .CP(ClockW), .CDN(n186), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n131), .E(N645), .CP(n212), .CDN(n159), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n122), .E(N645), .CP(n190), .CDN(n170), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(N546), .CP(n202), .CDN(n151), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n123), .E(N546), .CP(n211), .CDN(n161), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n142), .E(N546), .CP(n197), .CDN(n179), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n139), .E(N546), .CP(n191), .CDN(n157), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n117), .E(N546), .CP(n191), .CDN(n181), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n111), .E(N546), .CP(ClockW), .CDN(n179), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n138), .E(N546), .CP(n202), .CDN(n177), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n135), .E(N546), .CP(n208), .CDN(n183), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n121), .E(N546), .CP(n207), .CDN(n182), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n119), .E(N546), .CP(n212), .CDN(n180), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n134), .E(N546), .CP(n200), .CDN(n186), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n133), .E(N546), .CP(n203), .CDN(n182), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n115), .E(N546), .CP(n189), .CDN(n162), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n113), .E(N546), .CP(n198), .CDN(n175), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n130), .E(N546), .CP(n215), .CDN(n153), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n127), .E(N546), .CP(n192), .CDN(n153), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n112), .E(N546), .CP(n216), .CDN(n150), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n136), .E(N546), .CP(n213), .CDN(n108), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n137), .E(N546), .CP(n215), .CDN(n108), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n114), .E(N546), .CP(n216), .CDN(n157), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n116), .E(N546), .CP(n207), .CDN(n185), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n128), .E(N546), .CP(n207), .CDN(n161), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n129), .E(N546), .CP(n212), .CDN(n162), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n120), .E(N546), .CP(n213), .CDN(n170), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n140), .E(N546), .CP(n215), .CDN(n183), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n141), .E(N546), .CP(n212), .CDN(n172), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n124), .E(N546), .CP(n202), .CDN(n162), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n118), .E(N546), .CP(n199), .CDN(n187), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n126), .E(N546), .CP(ClockW), .CDN(n172), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n132), .E(N546), .CP(n211), .CDN(n175), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n125), .E(N546), .CP(n210), .CDN(n176), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n131), .E(N546), .CP(n209), .CDN(n177), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n122), .E(N546), .CP(n212), .CDN(n176), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N85), .E(N513), .CP(n192), .CDN(n167), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n123), .E(N513), .CP(n189), .CDN(n170), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n142), .E(N513), .CP(n205), .CDN(n171), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n139), .E(N513), .CP(n191), .CDN(n173), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n117), .E(N513), .CP(n193), .CDN(n160), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n111), .E(N513), .CP(n209), .CDN(n159), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n138), .E(N513), .CP(n201), .CDN(n158), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n135), .E(N513), .CP(n190), .CDN(n186), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n121), .E(N513), .CP(n217), .CDN(n173), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n119), .E(N513), .CP(n205), .CDN(n151), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n134), .E(N513), .CP(n205), .CDN(n152), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n133), .E(N513), .CP(n201), .CDN(n185), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n115), .E(N513), .CP(ClockW), .CDN(n172), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n113), .E(N513), .CP(n196), .CDN(n157), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n130), .E(N513), .CP(n210), .CDN(n186), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n127), .E(N513), .CP(n200), .CDN(n150), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n112), .E(N513), .CP(n188), .CDN(n173), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n136), .E(N513), .CP(n205), .CDN(n187), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n137), .E(N513), .CP(n213), .CDN(n153), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n114), .E(N513), .CP(n217), .CDN(n184), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n116), .E(N513), .CP(n208), .CDN(n185), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n128), .E(N513), .CP(n200), .CDN(n155), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n129), .E(N513), .CP(n205), .CDN(n158), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n120), .E(N513), .CP(n214), .CDN(n179), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n140), .E(N513), .CP(n188), .CDN(n170), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n141), .E(N513), .CP(ClockW), .CDN(n180), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n124), .E(N513), .CP(ClockW), .CDN(n176), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n118), .E(N513), .CP(n215), .CDN(n181), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n126), .E(N513), .CP(n216), .CDN(n157), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n132), .E(N513), .CP(n189), .CDN(n160), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n125), .E(N513), .CP(n201), .CDN(n157), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n131), .E(N513), .CP(n204), .CDN(n153), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n122), .E(N513), .CP(n217), .CDN(n171), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(N414), .CP(n217), .CDN(n174), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n123), .E(N414), .CP(n215), .CDN(n178), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n142), .E(N414), .CP(n204), .CDN(n173), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n139), .E(N414), .CP(n217), .CDN(n178), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n117), .E(N414), .CP(ClockW), .CDN(n184), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n111), .E(N414), .CP(n209), .CDN(n158), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n138), .E(N414), .CP(n210), .CDN(n184), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n135), .E(N414), .CP(n211), .CDN(n169), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n121), .E(N414), .CP(n213), .CDN(n184), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n119), .E(N414), .CP(n214), .CDN(n186), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n134), .E(N414), .CP(n212), .CDN(n175), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n133), .E(N414), .CP(n207), .CDN(n183), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n115), .E(N414), .CP(n207), .CDN(n182), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n113), .E(N414), .CP(n203), .CDN(n184), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n130), .E(N414), .CP(n206), .CDN(n175), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n127), .E(N414), .CP(n204), .CDN(n108), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n112), .E(N414), .CP(n191), .CDN(n154), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n136), .E(N414), .CP(n210), .CDN(n162), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n137), .E(N414), .CP(n217), .CDN(n173), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n114), .E(N414), .CP(n201), .CDN(n185), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n116), .E(N414), .CP(n209), .CDN(n184), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n128), .E(N414), .CP(n215), .CDN(n181), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n129), .E(N414), .CP(n194), .CDN(n174), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n120), .E(N414), .CP(n216), .CDN(n173), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n140), .E(N414), .CP(n204), .CDN(n168), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n141), .E(N414), .CP(n211), .CDN(n159), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n124), .E(N414), .CP(n199), .CDN(n186), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n118), .E(N414), .CP(n191), .CDN(n156), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n126), .E(N414), .CP(n198), .CDN(n176), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n132), .E(N414), .CP(n205), .CDN(n187), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n125), .E(N414), .CP(n190), .CDN(n180), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n131), .E(N414), .CP(n200), .CDN(n172), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n122), .E(N414), .CP(n212), .CDN(n159), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N85), .E(N381), .CP(n213), .CDN(n165), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n123), .E(N381), .CP(n212), .CDN(n174), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n142), .E(N381), .CP(n211), .CDN(n183), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n139), .E(N381), .CP(n210), .CDN(n182), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n117), .E(N381), .CP(n209), .CDN(n166), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n111), .E(N381), .CP(n208), .CDN(n165), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n138), .E(N381), .CP(n207), .CDN(n157), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n135), .E(N381), .CP(n207), .CDN(n158), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n121), .E(N381), .CP(n196), .CDN(n182), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n119), .E(N381), .CP(n212), .CDN(n166), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n134), .E(N381), .CP(n194), .CDN(n172), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n133), .E(N381), .CP(n202), .CDN(n180), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n115), .E(N381), .CP(n197), .CDN(n179), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n113), .E(N381), .CP(n189), .CDN(n151), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n130), .E(N381), .CP(n214), .CDN(n178), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n127), .E(N381), .CP(n203), .CDN(n171), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n112), .E(N381), .CP(n213), .CDN(n163), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n136), .E(N381), .CP(n201), .CDN(n108), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n137), .E(N381), .CP(n215), .CDN(n155), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n114), .E(N381), .CP(n207), .CDN(n187), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n116), .E(N381), .CP(n200), .CDN(n152), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n128), .E(N381), .CP(n211), .CDN(n187), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n129), .E(N381), .CP(n189), .CDN(n187), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n120), .E(N381), .CP(n190), .CDN(n165), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n140), .E(N381), .CP(n215), .CDN(n159), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n141), .E(N381), .CP(n191), .CDN(n185), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n124), .E(N381), .CP(ClockW), .CDN(n177), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n118), .E(N381), .CP(n215), .CDN(n164), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n126), .E(N381), .CP(n204), .CDN(n184), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n132), .E(N381), .CP(n216), .CDN(n186), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n125), .E(N381), .CP(n204), .CDN(n156), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n131), .E(N381), .CP(n207), .CDN(n168), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n122), .E(N381), .CP(n213), .CDN(n169), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(N282), .CP(n194), .CDN(n151), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n123), .E(N282), .CP(n208), .CDN(n158), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n142), .E(N282), .CP(n203), .CDN(n155), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n139), .E(N282), .CP(n188), .CDN(n185), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n117), .E(N282), .CP(n216), .CDN(n155), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n111), .E(N282), .CP(ClockW), .CDN(n177), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n138), .E(N282), .CP(n191), .CDN(n151), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n135), .E(N282), .CP(n215), .CDN(n181), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n121), .E(N282), .CP(n205), .CDN(n108), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n119), .E(N282), .CP(n198), .CDN(n173), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n134), .E(N282), .CP(n195), .CDN(n187), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n133), .E(N282), .CP(n204), .CDN(n154), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n115), .E(N282), .CP(n217), .CDN(n176), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n113), .E(N282), .CP(n202), .CDN(n181), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n130), .E(N282), .CP(n207), .CDN(n173), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n127), .E(N282), .CP(n215), .CDN(n166), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n112), .E(N282), .CP(n199), .CDN(n187), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n136), .E(N282), .CP(n197), .CDN(n165), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n137), .E(N282), .CP(n194), .CDN(n179), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n114), .E(N282), .CP(n193), .CDN(n179), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n116), .E(N282), .CP(n206), .CDN(n151), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n128), .E(N282), .CP(n196), .CDN(n186), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n129), .E(N282), .CP(n193), .CDN(n185), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n120), .E(N282), .CP(n196), .CDN(n182), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n140), .E(N282), .CP(n209), .CDN(n183), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n141), .E(N282), .CP(n217), .CDN(n181), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n124), .E(N282), .CP(n206), .CDN(n180), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n118), .E(N282), .CP(n217), .CDN(n178), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n126), .E(N282), .CP(n189), .CDN(n178), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n132), .E(N282), .CP(n206), .CDN(n166), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n125), .E(N282), .CP(n199), .CDN(n152), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n131), .E(N282), .CP(n217), .CDN(n179), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n122), .E(N282), .CP(n198), .CDN(n154), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N85), .E(N249), .CP(n196), .CDN(n180), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n123), .E(N249), .CP(n188), .CDN(n184), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n142), .E(N249), .CP(ClockW), .CDN(n158), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n139), .E(N249), .CP(n207), .CDN(n151), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n117), .E(N249), .CP(n192), .CDN(n174), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n111), .E(N249), .CP(n200), .CDN(n173), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n138), .E(N249), .CP(n203), .CDN(n187), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n135), .E(N249), .CP(n196), .CDN(n184), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n121), .E(N249), .CP(n203), .CDN(n185), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n119), .E(N249), .CP(n196), .CDN(n185), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n134), .E(N249), .CP(n214), .CDN(n152), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n133), .E(N249), .CP(n211), .CDN(n187), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n115), .E(N249), .CP(n189), .CDN(n164), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n113), .E(N249), .CP(n200), .CDN(n108), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n130), .E(N249), .CP(n202), .CDN(n187), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n127), .E(N249), .CP(ClockW), .CDN(n167), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n112), .E(N249), .CP(n199), .CDN(n154), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n136), .E(N249), .CP(n211), .CDN(n178), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n137), .E(N249), .CP(n213), .CDN(n167), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n114), .E(N249), .CP(n208), .CDN(n185), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n116), .E(N249), .CP(n209), .CDN(n167), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n128), .E(N249), .CP(n206), .CDN(n181), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n129), .E(N249), .CP(n194), .CDN(n155), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n120), .E(N249), .CP(n214), .CDN(n167), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n140), .E(N249), .CP(ClockW), .CDN(n185), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n141), .E(N249), .CP(n198), .CDN(n176), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n124), .E(N249), .CP(n201), .CDN(n187), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n118), .E(N249), .CP(n216), .CDN(n182), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n126), .E(N249), .CP(n215), .CDN(n183), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n132), .E(N249), .CP(n203), .CDN(n162), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n125), .E(N249), .CP(n216), .CDN(n178), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n131), .E(N249), .CP(n217), .CDN(n180), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n122), .E(N249), .CP(n192), .CDN(n186), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(N150), .CP(n211), .CDN(n151), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n123), .E(N150), .CP(n217), .CDN(n152), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n142), .E(N150), .CP(n214), .CDN(n161), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n139), .E(N150), .CP(n190), .CDN(n165), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n117), .E(N150), .CP(ClockW), .CDN(n183), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n111), .E(N150), .CP(ClockW), .CDN(n163), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n138), .E(N150), .CP(n215), .CDN(n183), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n135), .E(N150), .CP(n199), .CDN(n182), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n121), .E(N150), .CP(n216), .CDN(n154), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n119), .E(N150), .CP(ClockW), .CDN(n153), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n134), .E(N150), .CP(n201), .CDN(n184), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n133), .E(N150), .CP(ClockW), .CDN(n173), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n115), .E(N150), .CP(ClockW), .CDN(n165), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n113), .E(N150), .CP(n197), .CDN(n181), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n130), .E(N150), .CP(n209), .CDN(n168), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n127), .E(N150), .CP(n188), .CDN(n163), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n112), .E(N150), .CP(n211), .CDN(n185), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n136), .E(N150), .CP(n195), .CDN(n183), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n137), .E(N150), .CP(n210), .CDN(n175), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n114), .E(N150), .CP(n198), .CDN(n154), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n116), .E(N150), .CP(n199), .CDN(n168), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n128), .E(N150), .CP(n210), .CDN(n175), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n129), .E(N150), .CP(n212), .CDN(n186), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n120), .E(N150), .CP(n204), .CDN(n156), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n140), .E(N150), .CP(n208), .CDN(n186), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n141), .E(N150), .CP(n203), .CDN(n186), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n124), .E(N150), .CP(n202), .CDN(n177), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(N85), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(n123), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(n142), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(n139), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(n117), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(n111), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(n138), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(n135), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(n121), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(n119), .E(N1173), .CP(n188), .CDN(n153), 
        .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(n134), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(n133), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(n115), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(n113), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(n130), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(n127), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(n112), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(n136), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(n137), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(n114), .E(N1173), .CP(n189), .CDN(n154), 
        .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(n116), .E(N1173), .CP(n190), .CDN(n154), 
        .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(n128), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(n129), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(n120), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(n140), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(n141), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n124), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(n118), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(n126), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(n132), .E(N1173), .CP(n190), .CDN(n155), 
        .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(n125), .E(N1173), .CP(n191), .CDN(n155), 
        .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(n131), .E(N1173), .CP(n191), .CDN(n155), 
        .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(n122), .E(N1173), .CP(n191), .CDN(n156), 
        .Q(\Storage[31][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n107), .CP(ClockR), .CDN(n150), .Q(Dreadyr) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N51), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N52), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N53), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N54), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N55), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N56), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N57), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N58), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N59), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N60), .E(Read), .CP(ClockR), .CDN(n150), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N61), .E(Read), .CP(ClockR), .CDN(n151), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N62), .E(Read), .CP(ClockR), .CDN(n151), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N63), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N64), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N65), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N66), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N67), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N68), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N69), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N70), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N71), .E(n143), .CP(ClockR), .CDN(n151), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N72), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N73), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N74), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N75), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N76), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N77), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N78), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N79), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N80), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N81), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N82), .E(n143), .CP(ClockR), .CDN(n152), .Q(
        DataOr[0]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOr[29]), .OE(n146), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOr[2]), .OE(n146), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOr[28]), .OE(n146), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOr[3]), .OE(n146), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOr[27]), .OE(n146), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOr[4]), .OE(n146), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOr[26]), .OE(n146), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOr[5]), .OE(n146), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOr[25]), .OE(n146), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOr[6]), .OE(n146), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOr[24]), .OE(n146), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOr[7]), .OE(n146), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOr[23]), .OE(n146), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOr[8]), .OE(n146), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOr[22]), .OE(n146), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOr[9]), .OE(n146), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOr[21]), .OE(n146), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOr[10]), .OE(n146), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOr[20]), .OE(n146), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOr[11]), .OE(n146), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOr[19]), .OE(n146), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOr[12]), .OE(n146), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOr[18]), .OE(n146), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOr[13]), .OE(n146), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOr[17]), .OE(n146), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOr[14]), .OE(n146), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  EDFCNQD1 Parityr_reg ( .D(N83), .E(Read), .CP(ClockR), .CDN(n153), .Q(n716)
         );
  CKND2D0 U83 ( .A1(n146), .A2(Dreadyr), .ZN(n109) );
  CKNXD16 U84 ( .I(n109), .ZN(Dready) );
  AN2D1 U85 ( .A1(ClkW), .A2(n146), .Z(ClockW) );
  XOR3D1 U86 ( .A1(n125), .A2(n131), .A3(n682), .Z(N85) );
  BUFFD1 U87 ( .I(DataI[27]), .Z(n111) );
  BUFFD1 U88 ( .I(DataI[16]), .Z(n112) );
  BUFFD1 U89 ( .I(DataI[19]), .Z(n113) );
  BUFFD1 U90 ( .I(DataI[13]), .Z(n114) );
  BUFFD1 U91 ( .I(DataI[20]), .Z(n115) );
  BUFFD1 U92 ( .I(DataI[12]), .Z(n116) );
  BUFFD1 U93 ( .I(DataI[28]), .Z(n117) );
  BUFFD1 U94 ( .I(DataI[5]), .Z(n118) );
  BUFFD1 U95 ( .I(DataI[23]), .Z(n119) );
  BUFFD1 U96 ( .I(DataI[9]), .Z(n120) );
  BUFFD1 U97 ( .I(DataI[24]), .Z(n121) );
  BUFFD1 U98 ( .I(DataI[0]), .Z(n122) );
  BUFFD1 U99 ( .I(DataI[31]), .Z(n123) );
  BUFFD1 U100 ( .I(DataI[6]), .Z(n124) );
  BUFFD1 U101 ( .I(DataI[2]), .Z(n125) );
  BUFFD1 U102 ( .I(DataI[4]), .Z(n126) );
  BUFFD1 U103 ( .I(DataI[17]), .Z(n127) );
  BUFFD1 U104 ( .I(DataI[11]), .Z(n128) );
  BUFFD1 U105 ( .I(DataI[10]), .Z(n129) );
  BUFFD1 U106 ( .I(DataI[18]), .Z(n130) );
  BUFFD1 U107 ( .I(DataI[1]), .Z(n131) );
  BUFFD1 U108 ( .I(DataI[3]), .Z(n132) );
  BUFFD1 U109 ( .I(DataI[21]), .Z(n133) );
  BUFFD1 U110 ( .I(DataI[22]), .Z(n134) );
  BUFFD1 U111 ( .I(DataI[25]), .Z(n135) );
  BUFFD1 U112 ( .I(DataI[15]), .Z(n136) );
  BUFFD1 U113 ( .I(DataI[14]), .Z(n137) );
  BUFFD1 U114 ( .I(DataI[26]), .Z(n138) );
  BUFFD1 U115 ( .I(DataI[29]), .Z(n139) );
  BUFFD1 U116 ( .I(DataI[8]), .Z(n140) );
  BUFFD1 U117 ( .I(DataI[7]), .Z(n141) );
  BUFFD1 U118 ( .I(DataI[30]), .Z(n142) );
  BUFFD1 U119 ( .I(Read), .Z(n143) );
  BUFFD1 U120 ( .I(N48), .Z(n144) );
  BUFFD3 U121 ( .I(N47), .Z(n145) );
  BUFFD2 U122 ( .I(ChipEna), .Z(n146) );
  CKBD0 U123 ( .CLK(n149), .C(n147) );
  CKNXD16 U124 ( .I(n147), .ZN(ParityErr) );
  CKND0 U125 ( .CLK(n716), .CN(n149) );
  NR2D2P5 U126 ( .A1(n677), .A2(n710), .ZN(N447) );
  NR2D2P5 U127 ( .A1(n676), .A2(n707), .ZN(N1074) );
  NR2D2P5 U128 ( .A1(n681), .A2(n710), .ZN(N612) );
  ND3D1 U129 ( .A1(AddrW[3]), .A2(n711), .A3(Write), .ZN(n710) );
  NR2D2P5 U130 ( .A1(n694), .A2(n712), .ZN(N315) );
  NR2D2P5 U131 ( .A1(n676), .A2(n708), .ZN(N1041) );
  NR2D2P5 U132 ( .A1(n679), .A2(n680), .ZN(N909) );
  NR2D2P5 U133 ( .A1(n677), .A2(n712), .ZN(N183) );
  ND3D1 U134 ( .A1(n709), .A2(n711), .A3(Write), .ZN(n712) );
  NR2D2P5 U135 ( .A1(n676), .A2(n680), .ZN(N1173) );
  ND3D1 U136 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n676) );
  NR2D2P5 U137 ( .A1(n679), .A2(n681), .ZN(N876) );
  NR2D2P5 U138 ( .A1(n679), .A2(n694), .ZN(N843) );
  ND3D1 U139 ( .A1(AddrW[4]), .A2(n709), .A3(Write), .ZN(n679) );
  NR2D2P5 U140 ( .A1(n707), .A2(n710), .ZN(N546) );
  NR2D2P5 U141 ( .A1(n708), .A2(n712), .ZN(N249) );
  NR2D2P5 U142 ( .A1(n676), .A2(n681), .ZN(N1140) );
  NR2D2P5 U143 ( .A1(n679), .A2(n707), .ZN(N810) );
  NR2D2P5 U144 ( .A1(n680), .A2(n712), .ZN(N381) );
  NR2D2P5 U145 ( .A1(n675), .A2(n710), .ZN(N480) );
  NR2D2P5 U146 ( .A1(n676), .A2(n677), .ZN(N975) );
  NR2D2P5 U147 ( .A1(n679), .A2(n708), .ZN(N777) );
  NR2D2P5 U148 ( .A1(n694), .A2(n710), .ZN(N579) );
  NR2D2P5 U149 ( .A1(n675), .A2(n712), .ZN(N216) );
  NR2D2P5 U150 ( .A1(n676), .A2(n678), .ZN(N942) );
  NR2D2P5 U151 ( .A1(n675), .A2(n679), .ZN(N744) );
  NR2D2P5 U152 ( .A1(n680), .A2(n710), .ZN(N645) );
  NR2D2P5 U153 ( .A1(n681), .A2(n712), .ZN(N348) );
  NR2D2P5 U154 ( .A1(n676), .A2(n694), .ZN(N1107) );
  NR2D2P5 U155 ( .A1(n678), .A2(n679), .ZN(N678) );
  NR2D2P5 U156 ( .A1(n708), .A2(n710), .ZN(N513) );
  NR2D2P5 U157 ( .A1(n707), .A2(n712), .ZN(N282) );
  AN2D1 U158 ( .A1(ClkR), .A2(n146), .Z(ClockR) );
  NR2D2P5 U159 ( .A1(n675), .A2(n676), .ZN(N999) );
  ND3D1 U160 ( .A1(n713), .A2(n714), .A3(AddrW[1]), .ZN(n675) );
  NR2D2P5 U161 ( .A1(n677), .A2(n679), .ZN(N711) );
  NR2D2P5 U162 ( .A1(n678), .A2(n710), .ZN(N414) );
  NR2D2P5 U163 ( .A1(n678), .A2(n712), .ZN(N150) );
  ND3D1 U164 ( .A1(n715), .A2(n714), .A3(n713), .ZN(n678) );
  BUFFD1 U165 ( .I(n201), .Z(n206) );
  BUFFD1 U166 ( .I(n215), .Z(n205) );
  BUFFD1 U167 ( .I(n202), .Z(n204) );
  BUFFD1 U168 ( .I(n207), .Z(n203) );
  BUFFD1 U169 ( .I(n207), .Z(n202) );
  BUFFD1 U170 ( .I(n208), .Z(n201) );
  BUFFD1 U171 ( .I(n208), .Z(n200) );
  BUFFD1 U172 ( .I(n209), .Z(n199) );
  BUFFD1 U173 ( .I(n209), .Z(n198) );
  BUFFD1 U174 ( .I(n210), .Z(n197) );
  BUFFD1 U175 ( .I(n210), .Z(n196) );
  BUFFD1 U176 ( .I(n211), .Z(n195) );
  BUFFD1 U177 ( .I(n211), .Z(n194) );
  BUFFD1 U178 ( .I(n212), .Z(n193) );
  BUFFD1 U179 ( .I(n212), .Z(n192) );
  BUFFD1 U180 ( .I(n213), .Z(n191) );
  BUFFD1 U181 ( .I(n213), .Z(n190) );
  BUFFD1 U182 ( .I(n214), .Z(n189) );
  BUFFD1 U183 ( .I(n214), .Z(n188) );
  BUFFD1 U184 ( .I(n181), .Z(n177) );
  BUFFD1 U185 ( .I(n178), .Z(n176) );
  BUFFD1 U186 ( .I(n183), .Z(n175) );
  BUFFD1 U187 ( .I(n150), .Z(n174) );
  BUFFD1 U188 ( .I(n179), .Z(n173) );
  BUFFD1 U189 ( .I(n179), .Z(n172) );
  BUFFD1 U190 ( .I(n179), .Z(n171) );
  BUFFD1 U191 ( .I(n179), .Z(n170) );
  BUFFD1 U192 ( .I(n160), .Z(n169) );
  BUFFD1 U193 ( .I(n187), .Z(n168) );
  BUFFD1 U194 ( .I(n183), .Z(n167) );
  BUFFD1 U195 ( .I(n150), .Z(n166) );
  BUFFD1 U196 ( .I(n180), .Z(n165) );
  BUFFD1 U197 ( .I(n180), .Z(n164) );
  BUFFD1 U198 ( .I(n180), .Z(n163) );
  BUFFD1 U199 ( .I(n180), .Z(n162) );
  BUFFD1 U200 ( .I(n181), .Z(n161) );
  BUFFD1 U201 ( .I(n181), .Z(n160) );
  BUFFD1 U202 ( .I(n181), .Z(n159) );
  BUFFD1 U203 ( .I(n181), .Z(n158) );
  BUFFD1 U204 ( .I(n217), .Z(n207) );
  BUFFD1 U205 ( .I(n213), .Z(n208) );
  BUFFD1 U206 ( .I(n216), .Z(n209) );
  BUFFD1 U207 ( .I(n216), .Z(n210) );
  BUFFD1 U208 ( .I(n216), .Z(n211) );
  BUFFD1 U209 ( .I(n215), .Z(n212) );
  BUFFD1 U210 ( .I(n215), .Z(n213) );
  BUFFD1 U211 ( .I(n215), .Z(n214) );
  BUFFD1 U212 ( .I(n183), .Z(n150) );
  BUFFD1 U213 ( .I(n182), .Z(n157) );
  BUFFD1 U214 ( .I(n182), .Z(n156) );
  BUFFD1 U215 ( .I(n182), .Z(n155) );
  BUFFD1 U216 ( .I(n182), .Z(n154) );
  BUFFD1 U217 ( .I(n183), .Z(n153) );
  BUFFD1 U218 ( .I(n183), .Z(n152) );
  BUFFD1 U219 ( .I(n183), .Z(n151) );
  BUFFD1 U220 ( .I(n217), .Z(n216) );
  BUFFD1 U221 ( .I(n217), .Z(n215) );
  BUFFD1 U222 ( .I(n160), .Z(n178) );
  BUFFD1 U223 ( .I(n186), .Z(n179) );
  BUFFD1 U224 ( .I(n185), .Z(n180) );
  BUFFD1 U225 ( .I(n185), .Z(n181) );
  BUFFD1 U226 ( .I(n240), .Z(n236) );
  BUFFD1 U227 ( .I(n240), .Z(n235) );
  BUFFD1 U228 ( .I(n241), .Z(n234) );
  BUFFD1 U229 ( .I(n241), .Z(n233) );
  BUFFD1 U230 ( .I(n230), .Z(n223) );
  BUFFD1 U231 ( .I(n229), .Z(n224) );
  BUFFD1 U232 ( .I(n229), .Z(n225) );
  BUFFD1 U233 ( .I(n228), .Z(n226) );
  BUFFD1 U234 ( .I(n228), .Z(n227) );
  BUFFD1 U235 ( .I(ClockW), .Z(n217) );
  BUFFD1 U236 ( .I(n183), .Z(n186) );
  BUFFD1 U237 ( .I(n150), .Z(n185) );
  BUFFD1 U238 ( .I(n184), .Z(n182) );
  BUFFD1 U239 ( .I(n184), .Z(n183) );
  BUFFD1 U240 ( .I(n239), .Z(n237) );
  BUFFD1 U241 ( .I(n242), .Z(n232) );
  BUFFD1 U242 ( .I(n243), .Z(n242) );
  BUFFD1 U243 ( .I(n222), .Z(n219) );
  BUFFD1 U244 ( .I(n221), .Z(n218) );
  BUFFD1 U245 ( .I(n221), .Z(n220) );
  BUFFD1 U246 ( .I(n239), .Z(n238) );
  BUFFD1 U247 ( .I(n243), .Z(n240) );
  BUFFD1 U248 ( .I(n243), .Z(n241) );
  BUFFD1 U249 ( .I(n231), .Z(n228) );
  BUFFD1 U250 ( .I(n231), .Z(n229) );
  BUFFD1 U251 ( .I(n231), .Z(n230) );
  BUFFD1 U252 ( .I(n187), .Z(n184) );
  BUFFD1 U253 ( .I(n108), .Z(n187) );
  MUX4ND0 U254 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n240), .S1(N45), .ZN(
        n665) );
  MUX4ND0 U255 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n238), .S1(N45), .ZN(
        n262) );
  MUX4ND0 U256 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n234), .S1(n228), .ZN(
        n275) );
  MUX4ND0 U257 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n241), .S1(n226), .ZN(
        n288) );
  MUX4ND0 U258 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n239), .S1(n231), .ZN(
        n301) );
  MUX4ND0 U259 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n243), .S1(n229), .ZN(
        n314) );
  MUX4ND0 U260 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n241), .S1(n224), .ZN(
        n327) );
  MUX4ND0 U261 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n240), .S1(n229), .ZN(
        n340) );
  MUX4ND0 U262 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n242), .S1(n231), .ZN(
        n353) );
  MUX4ND0 U263 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n245), .S1(n231), .ZN(
        n366) );
  MUX4ND0 U264 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n242), .S1(n230), .ZN(
        n379) );
  MUX4ND0 U265 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n240), .S1(n231), .ZN(
        n392) );
  MUX4ND0 U266 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n245), .S1(n231), .ZN(
        n405) );
  MUX4ND0 U267 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n245), .S1(N45), .ZN(
        n418) );
  MUX4ND0 U268 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n240), .S1(n229), .ZN(
        n431) );
  MUX4ND0 U269 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n241), .S1(n227), .ZN(
        n444) );
  MUX4ND0 U270 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(N44), .S1(N45), .ZN(
        n457) );
  MUX4ND0 U271 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n236), .S1(n226), .ZN(
        n470) );
  MUX4ND0 U272 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n244), .S1(n231), .ZN(
        n483) );
  MUX4ND0 U273 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n243), .S1(n223), .ZN(
        n496) );
  MUX4ND0 U274 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n244), .S1(n225), .ZN(
        n509) );
  MUX4ND0 U275 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n243), .S1(n228), .ZN(
        n522) );
  MUX4ND0 U276 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n238), .S1(n229), .ZN(
        n535) );
  MUX4ND0 U277 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n234), .S1(n228), .ZN(
        n548) );
  MUX4ND0 U278 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n234), .S1(n230), .ZN(
        n561) );
  MUX4ND0 U279 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n241), .S1(n225), .ZN(
        n574) );
  MUX4ND0 U280 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n240), .S1(n231), .ZN(
        n587) );
  MUX4ND0 U281 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n241), .S1(N45), .ZN(
        n600) );
  MUX4ND0 U282 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n239), .S1(n231), .ZN(
        n613) );
  MUX4ND0 U283 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n243), .S1(n230), .ZN(
        n249) );
  MUX4ND0 U284 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n242), .S1(n227), .ZN(
        n626) );
  MUX4ND0 U285 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n245), .S1(n230), .ZN(
        n639) );
  MUX4ND0 U286 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n232), .S1(n228), .ZN(
        n652) );
  MUX4D0 U287 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n232), .S1(n223), .Z(
        n666) );
  MUX4D0 U288 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n241), .S1(n225), .Z(
        n250) );
  MUX4D0 U289 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n239), .S1(n223), .Z(
        n263) );
  MUX4D0 U290 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n240), .S1(n229), .Z(
        n276) );
  MUX4D0 U291 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n237), .S1(n230), .Z(
        n289) );
  MUX4D0 U292 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(N44), .S1(n228), .Z(n302) );
  MUX4D0 U293 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n245), .S1(n230), .Z(
        n315) );
  MUX4D0 U294 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n245), .S1(n230), .Z(
        n328) );
  MUX4D0 U295 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n242), .S1(n227), .Z(
        n341) );
  MUX4D0 U296 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n232), .S1(n223), .Z(
        n354) );
  MUX4D0 U297 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n244), .S1(n224), .Z(
        n367) );
  MUX4D0 U298 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n233), .S1(n225), .Z(
        n380) );
  MUX4D0 U299 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n245), .S1(n229), .Z(
        n393) );
  MUX4D0 U300 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n242), .S1(n230), .Z(
        n406) );
  MUX4D0 U301 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n237), .S1(n230), .Z(
        n419) );
  MUX4D0 U302 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n244), .S1(n226), .Z(
        n432) );
  MUX4D0 U303 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n244), .S1(n224), .Z(
        n445) );
  MUX4D0 U304 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n243), .S1(n228), .Z(
        n458) );
  MUX4D0 U305 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n244), .S1(n231), .Z(
        n471) );
  MUX4D0 U306 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n244), .S1(n225), .Z(
        n484) );
  MUX4D0 U307 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n241), .S1(n225), .Z(
        n497) );
  MUX4D0 U308 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n239), .S1(n226), .Z(
        n510) );
  MUX4D0 U309 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n242), .S1(n225), .Z(
        n523) );
  MUX4D0 U310 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n239), .S1(n226), .Z(
        n536) );
  MUX4D0 U311 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n244), .S1(n227), .Z(
        n549) );
  MUX4D0 U312 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n236), .S1(n230), .Z(
        n562) );
  MUX4D0 U313 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n236), .S1(N45), .Z(
        n575) );
  MUX4D0 U314 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n235), .S1(n226), .Z(
        n588) );
  MUX4D0 U315 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n235), .S1(n228), .Z(
        n601) );
  MUX4D0 U316 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n234), .S1(n231), .Z(
        n614) );
  MUX4D0 U317 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n234), .S1(n231), .Z(
        n627) );
  MUX4D0 U318 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n233), .S1(n228), .Z(
        n640) );
  MUX4D0 U319 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n233), .S1(n230), .Z(
        n653) );
  BUFFD1 U320 ( .I(N44), .Z(n244) );
  BUFFD1 U321 ( .I(N44), .Z(n243) );
  MUX4D0 U322 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n232), .S1(n230), .Z(
        n668) );
  MUX4D0 U323 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n232), .S1(n225), .Z(
        n670) );
  MUX4D0 U324 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n236), .S1(N45), .Z(n252) );
  MUX4D0 U325 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n233), .S1(n231), .Z(n254)
         );
  MUX4D0 U326 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n240), .S1(n228), .Z(
        n265) );
  MUX4D0 U327 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n237), .S1(n228), .Z(n267)
         );
  MUX4D0 U328 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n245), .S1(n224), .Z(
        n278) );
  MUX4D0 U329 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n235), .S1(n223), .Z(n280)
         );
  MUX4D0 U330 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n233), .S1(n229), .Z(
        n291) );
  MUX4D0 U331 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n236), .S1(n223), .Z(n293)
         );
  MUX4D0 U332 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n239), .S1(n223), .Z(
        n304) );
  MUX4D0 U333 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n241), .S1(n225), .Z(n306)
         );
  MUX4D0 U334 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n244), .S1(n224), .Z(
        n317) );
  MUX4D0 U335 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n232), .S1(n226), .Z(n319)
         );
  MUX4D0 U336 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n240), .S1(n223), .Z(
        n330) );
  MUX4D0 U337 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n236), .S1(n228), .Z(n332)
         );
  MUX4D0 U338 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n233), .S1(n224), .Z(
        n343) );
  MUX4D0 U339 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n243), .S1(n223), .Z(n345)
         );
  MUX4D0 U340 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n238), .S1(n227), .Z(
        n356) );
  MUX4D0 U341 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n238), .S1(n225), .Z(n358)
         );
  MUX4D0 U342 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(N44), .S1(n227), .Z(n369) );
  MUX4D0 U343 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n239), .S1(n227), .Z(n371)
         );
  MUX4D0 U344 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n235), .S1(n226), .Z(
        n382) );
  MUX4D0 U345 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n239), .S1(N45), .Z(n384) );
  MUX4D0 U346 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n240), .S1(n231), .Z(
        n395) );
  MUX4D0 U347 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n245), .S1(n230), .Z(
        n397) );
  MUX4D0 U348 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n237), .S1(n231), .Z(
        n408) );
  MUX4D0 U349 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(N44), .S1(n226), .Z(n410) );
  MUX4D0 U350 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n233), .S1(n228), .Z(
        n421) );
  MUX4D0 U351 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n243), .S1(n229), .Z(
        n423) );
  MUX4D0 U352 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n243), .S1(N45), .Z(
        n434) );
  MUX4D0 U353 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n244), .S1(n228), .Z(
        n436) );
  MUX4D0 U354 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n234), .S1(n229), .Z(
        n447) );
  MUX4D0 U355 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(N44), .S1(n227), .Z(n449) );
  MUX4D0 U356 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n245), .S1(n231), .Z(
        n460) );
  MUX4D0 U357 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n244), .S1(n227), .Z(
        n462) );
  MUX4D0 U358 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n239), .S1(n224), .Z(
        n473) );
  MUX4D0 U359 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n232), .S1(n231), .Z(
        n475) );
  MUX4D0 U360 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n244), .S1(n225), .Z(
        n486) );
  MUX4D0 U361 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n243), .S1(n227), .Z(
        n488) );
  MUX4D0 U362 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n241), .S1(n225), .Z(
        n499) );
  MUX4D0 U363 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n239), .S1(n226), .Z(
        n501) );
  MUX4D0 U364 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n238), .S1(n225), .Z(
        n512) );
  MUX4D0 U365 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n234), .S1(n225), .Z(
        n514) );
  MUX4D0 U366 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n236), .S1(n229), .Z(
        n525) );
  MUX4D0 U367 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n233), .S1(n226), .Z(
        n527) );
  MUX4D0 U368 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n243), .S1(n227), .Z(
        n538) );
  MUX4D0 U369 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n245), .S1(n227), .Z(
        n540) );
  MUX4D0 U370 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n242), .S1(n227), .Z(
        n551) );
  MUX4D0 U371 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n241), .S1(n228), .Z(
        n553) );
  MUX4D0 U372 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n236), .S1(n226), .Z(
        n564) );
  MUX4D0 U373 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n236), .S1(n226), .Z(
        n566) );
  MUX4D0 U374 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n236), .S1(n229), .Z(
        n577) );
  MUX4D0 U375 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n235), .S1(n228), .Z(
        n579) );
  MUX4D0 U376 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n235), .S1(n230), .Z(
        n590) );
  MUX4D0 U377 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n235), .S1(n227), .Z(
        n592) );
  MUX4D0 U378 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n235), .S1(n229), .Z(
        n603) );
  MUX4D0 U379 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n234), .S1(n230), .Z(
        n605) );
  MUX4D0 U380 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n234), .S1(n231), .Z(
        n616) );
  MUX4D0 U381 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n234), .S1(n228), .Z(
        n618) );
  MUX4D0 U382 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n233), .S1(n229), .Z(
        n629) );
  MUX4D0 U383 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n233), .S1(n227), .Z(
        n631) );
  MUX4D0 U384 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n233), .S1(n228), .Z(
        n642) );
  MUX4D0 U385 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n233), .S1(n228), .Z(
        n644) );
  MUX4D0 U386 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n232), .S1(n229), .Z(
        n655) );
  MUX4D0 U387 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n232), .S1(n230), .Z(
        n657) );
  BUFFD1 U388 ( .I(N46), .Z(n221) );
  BUFFD1 U389 ( .I(N46), .Z(n222) );
  MUX4D0 U390 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n232), .S1(n225), .Z(
        n667) );
  MUX4D0 U391 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n245), .S1(n227), .Z(
        n251) );
  MUX4D0 U392 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n233), .S1(n230), .Z(
        n264) );
  MUX4D0 U393 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n234), .S1(n223), .Z(
        n277) );
  MUX4D0 U394 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n238), .S1(n227), .Z(
        n290) );
  MUX4D0 U395 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n239), .S1(n224), .Z(
        n303) );
  MUX4D0 U396 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n242), .S1(n229), .Z(
        n316) );
  MUX4D0 U397 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(N44), .S1(n230), .Z(n329) );
  MUX4D0 U398 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n240), .S1(n226), .Z(
        n342) );
  MUX4D0 U399 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n242), .S1(n228), .Z(
        n355) );
  MUX4D0 U400 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n241), .S1(n225), .Z(
        n368) );
  MUX4D0 U401 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n235), .S1(n224), .Z(
        n381) );
  MUX4D0 U402 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n240), .S1(n231), .Z(
        n394) );
  MUX4D0 U403 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n243), .S1(n230), .Z(
        n407) );
  MUX4D0 U404 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n242), .S1(n226), .Z(
        n420) );
  MUX4D0 U405 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n245), .S1(n225), .Z(
        n433) );
  MUX4D0 U406 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n242), .S1(n228), .Z(
        n446) );
  MUX4D0 U407 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n239), .S1(n229), .Z(
        n459) );
  MUX4D0 U408 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n242), .S1(n230), .Z(
        n472) );
  MUX4D0 U409 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n238), .S1(n226), .Z(
        n485) );
  MUX4D0 U410 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n238), .S1(n227), .Z(
        n498) );
  MUX4D0 U411 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n235), .S1(n225), .Z(
        n511) );
  MUX4D0 U412 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n245), .S1(n226), .Z(
        n524) );
  MUX4D0 U413 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n241), .S1(n227), .Z(
        n537) );
  MUX4D0 U414 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n243), .S1(n227), .Z(
        n550) );
  MUX4D0 U415 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n236), .S1(n226), .Z(
        n563) );
  MUX4D0 U416 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n236), .S1(n228), .Z(
        n576) );
  MUX4D0 U417 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n235), .S1(n230), .Z(
        n589) );
  MUX4D0 U418 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n235), .S1(n231), .Z(
        n602) );
  MUX4D0 U419 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n234), .S1(n223), .Z(
        n615) );
  MUX4D0 U420 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n234), .S1(n228), .Z(
        n628) );
  MUX4D0 U421 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n233), .S1(n228), .Z(
        n641) );
  MUX4D0 U422 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n232), .S1(n225), .Z(
        n654) );
  MUX4D0 U423 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n232), .S1(n229), .Z(
        n669) );
  MUX4D0 U424 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n232), .S1(n226), .Z(
        n671) );
  MUX4D0 U425 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n235), .S1(n229), .Z(
        n253) );
  MUX4D0 U426 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n234), .S1(n225), .Z(n255)
         );
  MUX4D0 U427 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n236), .S1(n226), .Z(
        n266) );
  MUX4D0 U428 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n238), .S1(n224), .Z(n268)
         );
  MUX4D0 U429 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n242), .S1(n228), .Z(
        n279) );
  MUX4D0 U430 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n232), .S1(n229), .Z(n281)
         );
  MUX4D0 U431 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n232), .S1(n226), .Z(
        n292) );
  MUX4D0 U432 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n243), .S1(n227), .Z(n294)
         );
  MUX4D0 U433 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n244), .S1(n225), .Z(
        n305) );
  MUX4D0 U434 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n235), .S1(n228), .Z(n307)
         );
  MUX4D0 U435 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n239), .S1(n224), .Z(
        n318) );
  MUX4D0 U436 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n241), .S1(n231), .Z(n320)
         );
  MUX4D0 U437 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n241), .S1(n225), .Z(
        n331) );
  MUX4D0 U438 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n238), .S1(n225), .Z(n333)
         );
  MUX4D0 U439 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n245), .S1(n229), .Z(
        n344) );
  MUX4D0 U440 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n240), .S1(n230), .Z(n346)
         );
  MUX4D0 U441 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n245), .S1(n229), .Z(
        n357) );
  MUX4D0 U442 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n239), .S1(n223), .Z(n359)
         );
  MUX4D0 U443 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n244), .S1(n223), .Z(
        n370) );
  MUX4D0 U444 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n235), .S1(N45), .Z(n372)
         );
  MUX4D0 U445 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n240), .S1(n226), .Z(
        n383) );
  MUX4D0 U446 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n240), .S1(n227), .Z(
        n385) );
  MUX4D0 U447 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n242), .S1(n225), .Z(
        n396) );
  MUX4D0 U448 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n241), .S1(n231), .Z(
        n398) );
  MUX4D0 U449 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n243), .S1(n224), .Z(
        n409) );
  MUX4D0 U450 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n237), .S1(n231), .Z(
        n411) );
  MUX4D0 U451 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n240), .S1(n226), .Z(
        n422) );
  MUX4D0 U452 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n244), .S1(n224), .Z(
        n424) );
  MUX4D0 U453 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n239), .S1(n229), .Z(
        n435) );
  MUX4D0 U454 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n236), .S1(n229), .Z(
        n437) );
  MUX4D0 U455 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n244), .S1(N45), .Z(
        n448) );
  MUX4D0 U456 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n242), .S1(n228), .Z(
        n450) );
  MUX4D0 U457 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n234), .S1(n231), .Z(
        n461) );
  MUX4D0 U458 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n236), .S1(n227), .Z(
        n463) );
  MUX4D0 U459 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n233), .S1(n229), .Z(
        n474) );
  MUX4D0 U460 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n235), .S1(n224), .Z(
        n476) );
  MUX4D0 U461 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n243), .S1(n226), .Z(
        n487) );
  MUX4D0 U462 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n240), .S1(n225), .Z(
        n489) );
  MUX4D0 U463 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n244), .S1(n225), .Z(
        n500) );
  MUX4D0 U464 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n237), .S1(n227), .Z(
        n502) );
  MUX4D0 U465 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n232), .S1(n226), .Z(
        n513) );
  MUX4D0 U466 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n240), .S1(n226), .Z(
        n515) );
  MUX4D0 U467 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n239), .S1(n226), .Z(
        n526) );
  MUX4D0 U468 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n241), .S1(n226), .Z(
        n528) );
  MUX4D0 U469 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n232), .S1(n227), .Z(
        n539) );
  MUX4D0 U470 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n242), .S1(n227), .Z(
        n541) );
  MUX4D0 U471 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n239), .S1(n231), .Z(
        n552) );
  MUX4D0 U472 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n236), .S1(n223), .Z(
        n554) );
  MUX4D0 U473 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n236), .S1(N45), .Z(
        n565) );
  MUX4D0 U474 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n236), .S1(n231), .Z(
        n567) );
  MUX4D0 U475 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n236), .S1(n227), .Z(
        n578) );
  MUX4D0 U476 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n235), .S1(n230), .Z(
        n580) );
  MUX4D0 U477 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n235), .S1(n231), .Z(
        n591) );
  MUX4D0 U478 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n235), .S1(N45), .Z(n593) );
  MUX4D0 U479 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n234), .S1(n229), .Z(
        n604) );
  MUX4D0 U480 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n234), .S1(n230), .Z(
        n606) );
  MUX4D0 U481 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n234), .S1(n225), .Z(
        n617) );
  MUX4D0 U482 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n234), .S1(n229), .Z(
        n619) );
  MUX4D0 U483 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n233), .S1(n230), .Z(
        n630) );
  MUX4D0 U484 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n233), .S1(N45), .Z(n632) );
  MUX4D0 U485 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n233), .S1(n223), .Z(
        n643) );
  MUX4D0 U486 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n233), .S1(n225), .Z(
        n645) );
  MUX4D0 U487 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n232), .S1(n230), .Z(
        n656) );
  MUX4D0 U488 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n232), .S1(n227), .Z(
        n658) );
  BUFFD1 U489 ( .I(N45), .Z(n231) );
  BUFFD1 U490 ( .I(n245), .Z(n239) );
  BUFFD1 U491 ( .I(N44), .Z(n245) );
  MUX3ND0 U492 ( .I0(n247), .I1(n248), .I2(n249), .S0(n223), .S1(n221), .ZN(
        n246) );
  MUX3ND0 U493 ( .I0(n256), .I1(n257), .I2(n258), .S0(n145), .S1(n144), .ZN(
        N82) );
  MUX3ND0 U494 ( .I0(n260), .I1(n261), .I2(n262), .S0(n223), .S1(N46), .ZN(
        n259) );
  MUX3ND0 U495 ( .I0(n269), .I1(n270), .I2(n271), .S0(n145), .S1(n144), .ZN(
        N81) );
  MUX3ND0 U496 ( .I0(n273), .I1(n274), .I2(n275), .S0(n223), .S1(n222), .ZN(
        n272) );
  MUX3ND0 U497 ( .I0(n282), .I1(n283), .I2(n284), .S0(n145), .S1(n144), .ZN(
        N80) );
  MUX3ND0 U498 ( .I0(n286), .I1(n287), .I2(n288), .S0(n229), .S1(n221), .ZN(
        n285) );
  MUX3ND0 U499 ( .I0(n295), .I1(n296), .I2(n297), .S0(n145), .S1(n144), .ZN(
        N79) );
  MUX3ND0 U500 ( .I0(n299), .I1(n300), .I2(n301), .S0(n223), .S1(n220), .ZN(
        n298) );
  MUX3ND0 U501 ( .I0(n308), .I1(n309), .I2(n310), .S0(n145), .S1(n144), .ZN(
        N78) );
  MUX3ND0 U502 ( .I0(n312), .I1(n313), .I2(n314), .S0(n224), .S1(n221), .ZN(
        n311) );
  MUX3ND0 U503 ( .I0(n321), .I1(n322), .I2(n323), .S0(n145), .S1(n144), .ZN(
        N77) );
  MUX3ND0 U504 ( .I0(n325), .I1(n326), .I2(n327), .S0(n230), .S1(n218), .ZN(
        n324) );
  MUX3ND0 U505 ( .I0(n334), .I1(n335), .I2(n336), .S0(n145), .S1(n144), .ZN(
        N76) );
  MUX3ND0 U506 ( .I0(n338), .I1(n339), .I2(n340), .S0(n224), .S1(n219), .ZN(
        n337) );
  MUX3ND0 U507 ( .I0(n347), .I1(n348), .I2(n349), .S0(n145), .S1(n144), .ZN(
        N75) );
  MUX3ND0 U508 ( .I0(n351), .I1(n352), .I2(n353), .S0(n224), .S1(n220), .ZN(
        n350) );
  MUX3ND0 U509 ( .I0(n360), .I1(n361), .I2(n362), .S0(n145), .S1(n144), .ZN(
        N74) );
  MUX3ND0 U510 ( .I0(n364), .I1(n365), .I2(n366), .S0(n224), .S1(n221), .ZN(
        n363) );
  MUX3ND0 U511 ( .I0(n373), .I1(n374), .I2(n375), .S0(n145), .S1(n144), .ZN(
        N73) );
  MUX3ND0 U512 ( .I0(n377), .I1(n378), .I2(n379), .S0(n223), .S1(n222), .ZN(
        n376) );
  MUX3ND0 U513 ( .I0(n386), .I1(n387), .I2(n388), .S0(n145), .S1(n144), .ZN(
        N72) );
  MUX3ND0 U514 ( .I0(n390), .I1(n391), .I2(n392), .S0(n224), .S1(n222), .ZN(
        n389) );
  MUX3ND0 U515 ( .I0(n399), .I1(n400), .I2(n401), .S0(n145), .S1(n144), .ZN(
        N71) );
  MUX3ND0 U516 ( .I0(n403), .I1(n404), .I2(n405), .S0(n224), .S1(N46), .ZN(
        n402) );
  MUX3ND0 U517 ( .I0(n412), .I1(n413), .I2(n414), .S0(n145), .S1(n144), .ZN(
        N70) );
  MUX3ND0 U518 ( .I0(n416), .I1(n417), .I2(n418), .S0(n223), .S1(n219), .ZN(
        n415) );
  MUX3ND0 U519 ( .I0(n425), .I1(n426), .I2(n427), .S0(n145), .S1(n144), .ZN(
        N69) );
  MUX3ND0 U520 ( .I0(n429), .I1(n430), .I2(n431), .S0(n223), .S1(n219), .ZN(
        n428) );
  MUX3ND0 U521 ( .I0(n438), .I1(n439), .I2(n440), .S0(n145), .S1(n144), .ZN(
        N68) );
  MUX3ND0 U522 ( .I0(n442), .I1(n443), .I2(n444), .S0(n224), .S1(n218), .ZN(
        n441) );
  MUX3ND0 U523 ( .I0(n451), .I1(n452), .I2(n453), .S0(n145), .S1(n144), .ZN(
        N67) );
  MUX3ND0 U524 ( .I0(n455), .I1(n456), .I2(n457), .S0(n225), .S1(n219), .ZN(
        n454) );
  MUX3ND0 U525 ( .I0(n464), .I1(n465), .I2(n466), .S0(n145), .S1(n144), .ZN(
        N66) );
  MUX3ND0 U526 ( .I0(n468), .I1(n469), .I2(n470), .S0(n223), .S1(n222), .ZN(
        n467) );
  MUX3ND0 U527 ( .I0(n477), .I1(n478), .I2(n479), .S0(n145), .S1(n144), .ZN(
        N65) );
  MUX3ND0 U528 ( .I0(n481), .I1(n482), .I2(n483), .S0(n223), .S1(n220), .ZN(
        n480) );
  MUX3ND0 U529 ( .I0(n490), .I1(n491), .I2(n492), .S0(n145), .S1(n144), .ZN(
        N64) );
  MUX3ND0 U530 ( .I0(n494), .I1(n495), .I2(n496), .S0(n223), .S1(n218), .ZN(
        n493) );
  MUX3ND0 U531 ( .I0(n503), .I1(n504), .I2(n505), .S0(n145), .S1(n144), .ZN(
        N63) );
  MUX3ND0 U532 ( .I0(n507), .I1(n508), .I2(n509), .S0(n227), .S1(n221), .ZN(
        n506) );
  MUX3ND0 U533 ( .I0(n516), .I1(n517), .I2(n518), .S0(n145), .S1(N48), .ZN(N62) );
  MUX3ND0 U534 ( .I0(n520), .I1(n521), .I2(n522), .S0(n226), .S1(N46), .ZN(
        n519) );
  MUX3ND0 U535 ( .I0(n529), .I1(n530), .I2(n531), .S0(n145), .S1(N48), .ZN(N61) );
  MUX3ND0 U536 ( .I0(n533), .I1(n534), .I2(n535), .S0(n231), .S1(n220), .ZN(
        n532) );
  MUX3ND0 U537 ( .I0(n542), .I1(n543), .I2(n544), .S0(n145), .S1(N48), .ZN(N60) );
  MUX3ND0 U538 ( .I0(n546), .I1(n547), .I2(n548), .S0(n228), .S1(n220), .ZN(
        n545) );
  MUX3ND0 U539 ( .I0(n555), .I1(n556), .I2(n557), .S0(n145), .S1(N48), .ZN(N59) );
  MUX3ND0 U540 ( .I0(n559), .I1(n560), .I2(n561), .S0(n224), .S1(n221), .ZN(
        n558) );
  MUX3ND0 U541 ( .I0(n568), .I1(n569), .I2(n570), .S0(n145), .S1(N48), .ZN(N58) );
  MUX3ND0 U542 ( .I0(n572), .I1(n573), .I2(n574), .S0(n224), .S1(n222), .ZN(
        n571) );
  MUX3ND0 U543 ( .I0(n581), .I1(n582), .I2(n583), .S0(n145), .S1(N48), .ZN(N57) );
  MUX3ND0 U544 ( .I0(n585), .I1(n586), .I2(n587), .S0(n224), .S1(N46), .ZN(
        n584) );
  MUX3ND0 U545 ( .I0(n594), .I1(n595), .I2(n596), .S0(n145), .S1(N48), .ZN(N56) );
  MUX3ND0 U546 ( .I0(n598), .I1(n599), .I2(n600), .S0(n224), .S1(n222), .ZN(
        n597) );
  MUX3ND0 U547 ( .I0(n607), .I1(n608), .I2(n609), .S0(n145), .S1(N48), .ZN(N55) );
  MUX3ND0 U548 ( .I0(n611), .I1(n612), .I2(n613), .S0(n223), .S1(n220), .ZN(
        n610) );
  MUX3ND0 U549 ( .I0(n620), .I1(n621), .I2(n622), .S0(n145), .S1(N48), .ZN(N54) );
  MUX3ND0 U550 ( .I0(n624), .I1(n625), .I2(n626), .S0(n224), .S1(n221), .ZN(
        n623) );
  MUX3ND0 U551 ( .I0(n633), .I1(n634), .I2(n635), .S0(n145), .S1(N48), .ZN(N53) );
  MUX3ND0 U552 ( .I0(n637), .I1(n638), .I2(n639), .S0(n230), .S1(n222), .ZN(
        n636) );
  MUX3ND0 U553 ( .I0(n646), .I1(n647), .I2(n648), .S0(n145), .S1(N48), .ZN(N52) );
  MUX3ND0 U554 ( .I0(n650), .I1(n651), .I2(n652), .S0(n224), .S1(n221), .ZN(
        n649) );
  MUX3ND0 U555 ( .I0(n659), .I1(n660), .I2(n661), .S0(n145), .S1(N48), .ZN(N51) );
  MUX3ND0 U556 ( .I0(n663), .I1(n664), .I2(n665), .S0(n223), .S1(N46), .ZN(
        n662) );
  MUX3ND0 U557 ( .I0(n672), .I1(n673), .I2(n674), .S0(n145), .S1(n144), .ZN(
        N50) );
  MUX2ND0 U558 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n238), .ZN(
        n248) );
  MUX2ND0 U559 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n238), .ZN(
        n247) );
  MUX3ND0 U560 ( .I0(n251), .I1(n250), .I2(n246), .S0(n219), .S1(n145), .ZN(
        n258) );
  MUX2ND0 U561 ( .I0(n253), .I1(n252), .S(N46), .ZN(n257) );
  MUX2ND0 U562 ( .I0(n255), .I1(n254), .S(n220), .ZN(n256) );
  MUX2ND0 U563 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n238), .ZN(
        n261) );
  MUX2ND0 U564 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n237), .ZN(
        n260) );
  MUX3ND0 U565 ( .I0(n264), .I1(n263), .I2(n259), .S0(n219), .S1(n145), .ZN(
        n271) );
  MUX2ND0 U566 ( .I0(n266), .I1(n265), .S(n221), .ZN(n270) );
  MUX2ND0 U567 ( .I0(n268), .I1(n267), .S(n222), .ZN(n269) );
  MUX2ND0 U568 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n237), .ZN(
        n274) );
  MUX2ND0 U569 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n237), .ZN(
        n273) );
  MUX3ND0 U570 ( .I0(n277), .I1(n276), .I2(n272), .S0(n219), .S1(n145), .ZN(
        n284) );
  MUX2ND0 U571 ( .I0(n279), .I1(n278), .S(N46), .ZN(n283) );
  MUX2ND0 U572 ( .I0(n281), .I1(n280), .S(N46), .ZN(n282) );
  MUX2ND0 U573 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n237), .ZN(
        n287) );
  MUX2ND0 U574 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n244), .ZN(
        n286) );
  MUX3ND0 U575 ( .I0(n290), .I1(n289), .I2(n285), .S0(n222), .S1(n145), .ZN(
        n297) );
  MUX2ND0 U576 ( .I0(n292), .I1(n291), .S(n218), .ZN(n296) );
  MUX2ND0 U577 ( .I0(n294), .I1(n293), .S(n221), .ZN(n295) );
  MUX2ND0 U578 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(N44), .ZN(
        n300) );
  MUX2ND0 U579 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n242), .ZN(
        n299) );
  MUX3ND0 U580 ( .I0(n303), .I1(n302), .I2(n298), .S0(n219), .S1(n145), .ZN(
        n310) );
  MUX2ND0 U581 ( .I0(n305), .I1(n304), .S(n222), .ZN(n309) );
  MUX2ND0 U582 ( .I0(n307), .I1(n306), .S(n221), .ZN(n308) );
  MUX2ND0 U583 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n233), .ZN(
        n313) );
  MUX2ND0 U584 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n245), .ZN(
        n312) );
  MUX3ND0 U585 ( .I0(n316), .I1(n315), .I2(n311), .S0(n218), .S1(n145), .ZN(
        n323) );
  MUX2ND0 U586 ( .I0(n318), .I1(n317), .S(n220), .ZN(n322) );
  MUX2ND0 U587 ( .I0(n320), .I1(n319), .S(N46), .ZN(n321) );
  MUX2ND0 U588 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n239), .ZN(
        n326) );
  MUX2ND0 U589 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n235), .ZN(
        n325) );
  MUX3ND0 U590 ( .I0(n329), .I1(n328), .I2(n324), .S0(n219), .S1(n145), .ZN(
        n336) );
  MUX2ND0 U591 ( .I0(n331), .I1(n330), .S(n219), .ZN(n335) );
  MUX2ND0 U592 ( .I0(n333), .I1(n332), .S(n218), .ZN(n334) );
  MUX2ND0 U593 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n238), .ZN(
        n339) );
  MUX2ND0 U594 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(N44), .ZN(
        n338) );
  MUX3ND0 U595 ( .I0(n342), .I1(n341), .I2(n337), .S0(n220), .S1(n145), .ZN(
        n349) );
  MUX2ND0 U596 ( .I0(n344), .I1(n343), .S(n221), .ZN(n348) );
  MUX2ND0 U597 ( .I0(n346), .I1(n345), .S(n222), .ZN(n347) );
  MUX2ND0 U598 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n239), .ZN(
        n352) );
  MUX2ND0 U599 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n243), .ZN(
        n351) );
  MUX3ND0 U600 ( .I0(n355), .I1(n354), .I2(n350), .S0(n218), .S1(n145), .ZN(
        n362) );
  MUX2ND0 U601 ( .I0(n357), .I1(n356), .S(N46), .ZN(n361) );
  MUX2ND0 U602 ( .I0(n359), .I1(n358), .S(N46), .ZN(n360) );
  MUX2ND0 U603 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n233), .ZN(
        n365) );
  MUX2ND0 U604 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(N44), .ZN(
        n364) );
  MUX3ND0 U605 ( .I0(n368), .I1(n367), .I2(n363), .S0(n219), .S1(n145), .ZN(
        n375) );
  MUX2ND0 U606 ( .I0(n370), .I1(n369), .S(n220), .ZN(n374) );
  MUX2ND0 U607 ( .I0(n372), .I1(n371), .S(n219), .ZN(n373) );
  MUX2ND0 U608 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n244), 
        .ZN(n378) );
  MUX2ND0 U609 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n240), 
        .ZN(n377) );
  MUX3ND0 U610 ( .I0(n381), .I1(n380), .I2(n376), .S0(n219), .S1(n145), .ZN(
        n388) );
  MUX2ND0 U611 ( .I0(n383), .I1(n382), .S(n222), .ZN(n387) );
  MUX2ND0 U612 ( .I0(n385), .I1(n384), .S(n221), .ZN(n386) );
  MUX2ND0 U613 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n240), 
        .ZN(n391) );
  MUX2ND0 U614 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n241), 
        .ZN(n390) );
  MUX3ND0 U615 ( .I0(n394), .I1(n393), .I2(n389), .S0(n221), .S1(n145), .ZN(
        n401) );
  MUX2ND0 U616 ( .I0(n396), .I1(n395), .S(n222), .ZN(n400) );
  MUX2ND0 U617 ( .I0(n398), .I1(n397), .S(n221), .ZN(n399) );
  MUX2ND0 U618 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n241), 
        .ZN(n404) );
  MUX2ND0 U619 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n243), 
        .ZN(n403) );
  MUX3ND0 U620 ( .I0(n407), .I1(n406), .I2(n402), .S0(n222), .S1(n145), .ZN(
        n414) );
  MUX2ND0 U621 ( .I0(n409), .I1(n408), .S(n222), .ZN(n413) );
  MUX2ND0 U622 ( .I0(n411), .I1(n410), .S(n222), .ZN(n412) );
  MUX2ND0 U623 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n243), 
        .ZN(n417) );
  MUX2ND0 U624 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n242), 
        .ZN(n416) );
  MUX3ND0 U625 ( .I0(n420), .I1(n419), .I2(n415), .S0(n218), .S1(n145), .ZN(
        n427) );
  MUX2ND0 U626 ( .I0(n422), .I1(n421), .S(n221), .ZN(n426) );
  MUX2ND0 U627 ( .I0(n424), .I1(n423), .S(n219), .ZN(n425) );
  MUX2ND0 U628 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n236), 
        .ZN(n430) );
  MUX2ND0 U629 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n245), 
        .ZN(n429) );
  MUX3ND0 U630 ( .I0(n433), .I1(n432), .I2(n428), .S0(n219), .S1(n145), .ZN(
        n440) );
  MUX2ND0 U631 ( .I0(n435), .I1(n434), .S(n219), .ZN(n439) );
  MUX2ND0 U632 ( .I0(n437), .I1(n436), .S(n220), .ZN(n438) );
  MUX2ND0 U633 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n245), 
        .ZN(n443) );
  MUX2ND0 U634 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n244), 
        .ZN(n442) );
  MUX3ND0 U635 ( .I0(n446), .I1(n445), .I2(n441), .S0(n218), .S1(n145), .ZN(
        n453) );
  MUX2ND0 U636 ( .I0(n448), .I1(n447), .S(n218), .ZN(n452) );
  MUX2ND0 U637 ( .I0(n450), .I1(n449), .S(n221), .ZN(n451) );
  MUX2ND0 U638 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n242), 
        .ZN(n456) );
  MUX2ND0 U639 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n241), 
        .ZN(n455) );
  MUX3ND0 U640 ( .I0(n459), .I1(n458), .I2(n454), .S0(n222), .S1(n145), .ZN(
        n466) );
  MUX2ND0 U641 ( .I0(n461), .I1(n460), .S(n220), .ZN(n465) );
  MUX2ND0 U642 ( .I0(n463), .I1(n462), .S(n220), .ZN(n464) );
  MUX2ND0 U643 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n232), 
        .ZN(n469) );
  MUX2ND0 U644 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n241), 
        .ZN(n468) );
  MUX3ND0 U645 ( .I0(n472), .I1(n471), .I2(n467), .S0(n218), .S1(n145), .ZN(
        n479) );
  MUX2ND0 U646 ( .I0(n474), .I1(n473), .S(n220), .ZN(n478) );
  MUX2ND0 U647 ( .I0(n476), .I1(n475), .S(n220), .ZN(n477) );
  MUX2ND0 U648 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n240), 
        .ZN(n482) );
  MUX2ND0 U649 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n234), 
        .ZN(n481) );
  MUX3ND0 U650 ( .I0(n485), .I1(n484), .I2(n480), .S0(n219), .S1(n145), .ZN(
        n492) );
  MUX2ND0 U651 ( .I0(n487), .I1(n486), .S(n220), .ZN(n491) );
  MUX2ND0 U652 ( .I0(n489), .I1(n488), .S(n222), .ZN(n490) );
  MUX2ND0 U653 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n239), 
        .ZN(n495) );
  MUX2ND0 U654 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n238), 
        .ZN(n494) );
  MUX3ND0 U655 ( .I0(n498), .I1(n497), .I2(n493), .S0(n221), .S1(n145), .ZN(
        n505) );
  MUX2ND0 U656 ( .I0(n500), .I1(n499), .S(n222), .ZN(n504) );
  MUX2ND0 U657 ( .I0(n502), .I1(n501), .S(n220), .ZN(n503) );
  MUX2ND0 U658 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n238), 
        .ZN(n508) );
  MUX2ND0 U659 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n245), 
        .ZN(n507) );
  MUX3ND0 U660 ( .I0(n511), .I1(n510), .I2(n506), .S0(n220), .S1(n145), .ZN(
        n518) );
  MUX2ND0 U661 ( .I0(n513), .I1(n512), .S(n222), .ZN(n517) );
  MUX2ND0 U662 ( .I0(n515), .I1(n514), .S(n220), .ZN(n516) );
  MUX2ND0 U663 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n243), 
        .ZN(n521) );
  MUX2ND0 U664 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n242), 
        .ZN(n520) );
  MUX3ND0 U665 ( .I0(n524), .I1(n523), .I2(n519), .S0(n218), .S1(n145), .ZN(
        n531) );
  MUX2ND0 U666 ( .I0(n526), .I1(n525), .S(n219), .ZN(n530) );
  MUX2ND0 U667 ( .I0(n528), .I1(n527), .S(n220), .ZN(n529) );
  MUX2ND0 U668 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n244), 
        .ZN(n534) );
  MUX2ND0 U669 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n237), 
        .ZN(n533) );
  MUX3ND0 U670 ( .I0(n537), .I1(n536), .I2(n532), .S0(n219), .S1(n145), .ZN(
        n544) );
  MUX2ND0 U671 ( .I0(n539), .I1(n538), .S(n218), .ZN(n543) );
  MUX2ND0 U672 ( .I0(n541), .I1(n540), .S(n220), .ZN(n542) );
  MUX2ND0 U673 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n237), 
        .ZN(n547) );
  MUX2ND0 U674 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n237), 
        .ZN(n546) );
  MUX3ND0 U675 ( .I0(n550), .I1(n549), .I2(n545), .S0(n219), .S1(n145), .ZN(
        n557) );
  MUX2ND0 U676 ( .I0(n552), .I1(n551), .S(n222), .ZN(n556) );
  MUX2ND0 U677 ( .I0(n554), .I1(n553), .S(n218), .ZN(n555) );
  MUX2ND0 U678 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n237), 
        .ZN(n560) );
  MUX2ND0 U679 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n237), 
        .ZN(n559) );
  MUX3ND0 U680 ( .I0(n563), .I1(n562), .I2(n558), .S0(n219), .S1(n145), .ZN(
        n570) );
  MUX2ND0 U681 ( .I0(n565), .I1(n564), .S(n221), .ZN(n569) );
  MUX2ND0 U682 ( .I0(n567), .I1(n566), .S(n220), .ZN(n568) );
  MUX2ND0 U683 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n237), 
        .ZN(n573) );
  MUX2ND0 U684 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n237), 
        .ZN(n572) );
  MUX3ND0 U685 ( .I0(n576), .I1(n575), .I2(n571), .S0(n219), .S1(n145), .ZN(
        n583) );
  MUX2ND0 U686 ( .I0(n578), .I1(n577), .S(n218), .ZN(n582) );
  MUX2ND0 U687 ( .I0(n580), .I1(n579), .S(n222), .ZN(n581) );
  MUX2ND0 U688 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n237), 
        .ZN(n586) );
  MUX2ND0 U689 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n237), 
        .ZN(n585) );
  MUX3ND0 U690 ( .I0(n589), .I1(n588), .I2(n584), .S0(n218), .S1(n145), .ZN(
        n596) );
  MUX2ND0 U691 ( .I0(n591), .I1(n590), .S(n221), .ZN(n595) );
  MUX2ND0 U692 ( .I0(n593), .I1(n592), .S(n218), .ZN(n594) );
  MUX2ND0 U693 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n237), 
        .ZN(n599) );
  MUX2ND0 U694 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n237), 
        .ZN(n598) );
  MUX3ND0 U695 ( .I0(n602), .I1(n601), .I2(n597), .S0(n218), .S1(n145), .ZN(
        n609) );
  MUX2ND0 U696 ( .I0(n604), .I1(n603), .S(n220), .ZN(n608) );
  MUX2ND0 U697 ( .I0(n606), .I1(n605), .S(n222), .ZN(n607) );
  MUX2ND0 U698 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n237), 
        .ZN(n612) );
  MUX2ND0 U699 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n237), 
        .ZN(n611) );
  MUX3ND0 U700 ( .I0(n615), .I1(n614), .I2(n610), .S0(n218), .S1(n145), .ZN(
        n622) );
  MUX2ND0 U701 ( .I0(n617), .I1(n616), .S(n219), .ZN(n621) );
  MUX2ND0 U702 ( .I0(n619), .I1(n618), .S(n221), .ZN(n620) );
  MUX2ND0 U703 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n238), 
        .ZN(n625) );
  MUX2ND0 U704 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n238), 
        .ZN(n624) );
  MUX3ND0 U705 ( .I0(n628), .I1(n627), .I2(n623), .S0(n218), .S1(n145), .ZN(
        n635) );
  MUX2ND0 U706 ( .I0(n630), .I1(n629), .S(n221), .ZN(n634) );
  MUX2ND0 U707 ( .I0(n632), .I1(n631), .S(n221), .ZN(n633) );
  MUX2ND0 U708 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n238), 
        .ZN(n638) );
  MUX2ND0 U709 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n238), 
        .ZN(n637) );
  MUX3ND0 U710 ( .I0(n641), .I1(n640), .I2(n636), .S0(n218), .S1(n145), .ZN(
        n648) );
  MUX2ND0 U711 ( .I0(n643), .I1(n642), .S(n222), .ZN(n647) );
  MUX2ND0 U712 ( .I0(n645), .I1(n644), .S(n219), .ZN(n646) );
  MUX2ND0 U713 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n238), 
        .ZN(n651) );
  MUX2ND0 U714 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n238), 
        .ZN(n650) );
  MUX3ND0 U715 ( .I0(n654), .I1(n653), .I2(n649), .S0(n218), .S1(n145), .ZN(
        n661) );
  MUX2ND0 U716 ( .I0(n656), .I1(n655), .S(n220), .ZN(n660) );
  MUX2ND0 U717 ( .I0(n658), .I1(n657), .S(n218), .ZN(n659) );
  MUX2ND0 U718 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n238), 
        .ZN(n664) );
  MUX2ND0 U719 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(N44), .ZN(
        n663) );
  MUX3ND0 U720 ( .I0(n667), .I1(n666), .I2(n662), .S0(n218), .S1(n145), .ZN(
        n674) );
  MUX2ND0 U721 ( .I0(n669), .I1(n668), .S(n220), .ZN(n673) );
  MUX2ND0 U722 ( .I0(n671), .I1(n670), .S(N46), .ZN(n672) );
  CKND0 U723 ( .CLK(Reset), .CN(n108) );
  OR2D0 U724 ( .A1(n143), .A2(Dreadyr), .Z(n107) );
  XOR3D0 U725 ( .A1(n122), .A2(n683), .A3(n684), .Z(n682) );
  XOR3D0 U726 ( .A1(n118), .A2(n126), .A3(n685), .Z(n684) );
  XOR3D0 U727 ( .A1(n686), .A2(n132), .A3(n687), .Z(n685) );
  XOR3D0 U728 ( .A1(n116), .A2(n128), .A3(n688), .Z(n687) );
  XOR3D0 U729 ( .A1(n689), .A2(n129), .A3(n690), .Z(n688) );
  XOR3D0 U730 ( .A1(n113), .A2(n130), .A3(n691), .Z(n690) );
  XOR3D0 U731 ( .A1(n692), .A2(n127), .A3(n693), .Z(n691) );
  XNR4D0 U732 ( .A1(n135), .A2(n121), .A3(n111), .A4(n138), .ZN(n693) );
  XOR4D0 U733 ( .A1(n139), .A2(n117), .A3(n123), .A4(n142), .Z(n692) );
  XOR4D0 U734 ( .A1(n133), .A2(n115), .A3(n119), .A4(n134), .Z(n689) );
  XOR4D0 U735 ( .A1(n137), .A2(n114), .A3(n112), .A4(n136), .Z(n686) );
  XNR4D0 U736 ( .A1(n141), .A2(n124), .A3(n120), .A4(n140), .ZN(n683) );
  XOR4D0 U737 ( .A1(n695), .A2(N79), .A3(n696), .A4(n697), .Z(N83) );
  XNR4D0 U738 ( .A1(N76), .A2(N75), .A3(N78), .A4(N77), .ZN(n697) );
  XNR3D0 U739 ( .A1(N82), .A2(N81), .A3(N80), .ZN(n696) );
  XOR3D0 U740 ( .A1(N74), .A2(N73), .A3(n698), .Z(n695) );
  XOR3D0 U741 ( .A1(N72), .A2(n699), .A3(n700), .Z(n698) );
  XOR3D0 U742 ( .A1(N67), .A2(N66), .A3(n701), .Z(n700) );
  XOR3D0 U743 ( .A1(n702), .A2(N65), .A3(n703), .Z(n701) );
  XOR3D0 U744 ( .A1(N60), .A2(N59), .A3(n704), .Z(n703) );
  XOR3D0 U745 ( .A1(n705), .A2(N58), .A3(n706), .Z(n704) );
  XNR4D0 U746 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n706) );
  XOR4D0 U747 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n705) );
  XOR4D0 U748 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .Z(n702) );
  XNR4D0 U749 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n699) );
  ND3D0 U750 ( .A1(n715), .A2(n714), .A3(AddrW[0]), .ZN(n677) );
  CKND0 U751 ( .CLK(AddrW[4]), .CN(n711) );
  CKND0 U752 ( .CLK(AddrW[3]), .CN(n709) );
  ND3D0 U753 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n680) );
  ND3D0 U754 ( .A1(AddrW[1]), .A2(n713), .A3(AddrW[2]), .ZN(n681) );
  ND3D0 U755 ( .A1(AddrW[0]), .A2(n715), .A3(AddrW[2]), .ZN(n694) );
  ND3D0 U756 ( .A1(n713), .A2(n715), .A3(AddrW[2]), .ZN(n707) );
  CKND0 U757 ( .CLK(AddrW[1]), .CN(n715) );
  CKND0 U758 ( .CLK(AddrW[0]), .CN(n713) );
  ND3D0 U759 ( .A1(AddrW[1]), .A2(n714), .A3(AddrW[0]), .ZN(n708) );
  CKND0 U760 ( .CLK(AddrW[2]), .CN(n714) );
endmodule

