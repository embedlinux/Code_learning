
module SerFrameEnc ( FrameOut, BusIn, DoFrame );
  output [63:0] FrameOut;
  input [31:0] BusIn;
  input DoFrame;
  wire   n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n1, n2, n4, n6,
         n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34,
         n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62,
         n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97;

  DFQD1 \FrameReg_reg[63]  ( .D(BusIn[31]), .CP(n1), .Q(n98) );
  DFQD1 \FrameReg_reg[9]  ( .D(BusIn[1]), .CP(n1), .Q(n128) );
  DFQD1 \FrameReg_reg[8]  ( .D(BusIn[0]), .CP(n1), .Q(n129) );
  DFQD1 \FrameReg_reg[62]  ( .D(BusIn[30]), .CP(n1), .Q(n99) );
  DFQD1 \FrameReg_reg[61]  ( .D(BusIn[29]), .CP(n1), .Q(n100) );
  DFQD1 \FrameReg_reg[10]  ( .D(BusIn[2]), .CP(n1), .Q(n127) );
  DFQD1 \FrameReg_reg[11]  ( .D(BusIn[3]), .CP(n1), .Q(n126) );
  DFQD1 \FrameReg_reg[60]  ( .D(BusIn[28]), .CP(n1), .Q(n101) );
  DFQD1 \FrameReg_reg[59]  ( .D(BusIn[27]), .CP(n1), .Q(n102) );
  DFQD1 \FrameReg_reg[12]  ( .D(BusIn[4]), .CP(n1), .Q(n125) );
  DFQD1 \FrameReg_reg[13]  ( .D(BusIn[5]), .CP(n1), .Q(n124) );
  DFQD1 \FrameReg_reg[58]  ( .D(BusIn[26]), .CP(n1), .Q(n103) );
  DFQD1 \FrameReg_reg[57]  ( .D(BusIn[25]), .CP(n1), .Q(n104) );
  DFQD1 \FrameReg_reg[14]  ( .D(BusIn[6]), .CP(n1), .Q(n123) );
  DFQD1 \FrameReg_reg[15]  ( .D(BusIn[7]), .CP(n1), .Q(n122) );
  DFQD1 \FrameReg_reg[56]  ( .D(BusIn[24]), .CP(n1), .Q(n105) );
  DFQD1 \FrameReg_reg[47]  ( .D(BusIn[23]), .CP(n1), .Q(n106) );
  DFQD1 \FrameReg_reg[24]  ( .D(BusIn[8]), .CP(n1), .Q(n121) );
  DFQD1 \FrameReg_reg[25]  ( .D(BusIn[9]), .CP(n1), .Q(n120) );
  DFQD1 \FrameReg_reg[46]  ( .D(BusIn[22]), .CP(n1), .Q(n107) );
  DFQD1 \FrameReg_reg[45]  ( .D(BusIn[21]), .CP(n1), .Q(n108) );
  DFQD1 \FrameReg_reg[26]  ( .D(BusIn[10]), .CP(n1), .Q(n119) );
  DFQD1 \FrameReg_reg[27]  ( .D(BusIn[11]), .CP(n1), .Q(n118) );
  DFQD1 \FrameReg_reg[44]  ( .D(BusIn[20]), .CP(n1), .Q(n109) );
  DFQD1 \FrameReg_reg[43]  ( .D(BusIn[19]), .CP(n1), .Q(n110) );
  DFQD1 \FrameReg_reg[28]  ( .D(BusIn[12]), .CP(n1), .Q(n117) );
  DFQD1 \FrameReg_reg[29]  ( .D(BusIn[13]), .CP(n1), .Q(n116) );
  DFQD1 \FrameReg_reg[42]  ( .D(BusIn[18]), .CP(n1), .Q(n111) );
  DFQD1 \FrameReg_reg[41]  ( .D(BusIn[17]), .CP(n1), .Q(n112) );
  DFQD1 \FrameReg_reg[30]  ( .D(BusIn[14]), .CP(n1), .Q(n115) );
  DFQD1 \FrameReg_reg[31]  ( .D(BusIn[15]), .CP(n1), .Q(n114) );
  DFQD1 \FrameReg_reg[40]  ( .D(BusIn[16]), .CP(n1), .Q(n113) );
  BUFFD1 U35 ( .I(DoFrame), .Z(n1) );
  CKBD0 U36 ( .CLK(n68), .C(n2) );
  CKNXD16 U37 ( .I(n2), .ZN(FrameOut[30]) );
  CKND0 U38 ( .CLK(n115), .CN(n68) );
  CKBD0 U39 ( .CLK(n72), .C(n4) );
  CKNXD16 U40 ( .I(n4), .ZN(FrameOut[28]) );
  CKND0 U41 ( .CLK(n117), .CN(n72) );
  CKBD0 U42 ( .CLK(n70), .C(n6) );
  CKNXD16 U43 ( .I(n6), .ZN(FrameOut[42]) );
  CKND0 U44 ( .CLK(n111), .CN(n70) );
  CKBD0 U45 ( .CLK(n76), .C(n8) );
  CKNXD16 U46 ( .I(n8), .ZN(FrameOut[26]) );
  CKND0 U47 ( .CLK(n119), .CN(n76) );
  CKBD0 U48 ( .CLK(n74), .C(n10) );
  CKNXD16 U49 ( .I(n10), .ZN(FrameOut[44]) );
  CKND0 U50 ( .CLK(n109), .CN(n74) );
  CKBD0 U51 ( .CLK(n80), .C(n12) );
  CKNXD16 U52 ( .I(n12), .ZN(FrameOut[24]) );
  CKND0 U53 ( .CLK(n121), .CN(n80) );
  CKBD0 U54 ( .CLK(n78), .C(n14) );
  CKNXD16 U55 ( .I(n14), .ZN(FrameOut[46]) );
  CKND0 U56 ( .CLK(n107), .CN(n78) );
  CKBD0 U57 ( .CLK(n84), .C(n16) );
  CKNXD16 U58 ( .I(n16), .ZN(FrameOut[14]) );
  CKND0 U59 ( .CLK(n123), .CN(n84) );
  CKBD0 U60 ( .CLK(n82), .C(n18) );
  CKNXD16 U61 ( .I(n18), .ZN(FrameOut[56]) );
  CKND0 U62 ( .CLK(n105), .CN(n82) );
  CKBD0 U63 ( .CLK(n88), .C(n20) );
  CKNXD16 U64 ( .I(n20), .ZN(FrameOut[12]) );
  CKND0 U65 ( .CLK(n125), .CN(n88) );
  CKBD0 U66 ( .CLK(n86), .C(n22) );
  CKNXD16 U67 ( .I(n22), .ZN(FrameOut[58]) );
  CKND0 U68 ( .CLK(n103), .CN(n86) );
  CKBD0 U69 ( .CLK(n92), .C(n24) );
  CKNXD16 U70 ( .I(n24), .ZN(FrameOut[10]) );
  CKND0 U71 ( .CLK(n127), .CN(n92) );
  CKBD0 U72 ( .CLK(n90), .C(n26) );
  CKNXD16 U73 ( .I(n26), .ZN(FrameOut[60]) );
  CKND0 U74 ( .CLK(n101), .CN(n90) );
  CKBD0 U75 ( .CLK(n96), .C(n28) );
  CKNXD16 U76 ( .I(n28), .ZN(FrameOut[9]) );
  CKND0 U77 ( .CLK(n128), .CN(n96) );
  CKBD0 U78 ( .CLK(n94), .C(n30) );
  CKNXD16 U79 ( .I(n30), .ZN(FrameOut[62]) );
  CKND0 U80 ( .CLK(n99), .CN(n94) );
  CKBD0 U81 ( .CLK(n97), .C(n32) );
  CKNXD16 U82 ( .I(n32), .ZN(FrameOut[63]) );
  CKND0 U83 ( .CLK(n98), .CN(n97) );
  CKBD0 U84 ( .CLK(n95), .C(n34) );
  CKNXD16 U85 ( .I(n34), .ZN(FrameOut[8]) );
  CKND0 U86 ( .CLK(n129), .CN(n95) );
  CKBD0 U87 ( .CLK(n93), .C(n36) );
  CKNXD16 U88 ( .I(n36), .ZN(FrameOut[61]) );
  CKND0 U89 ( .CLK(n100), .CN(n93) );
  CKBD0 U90 ( .CLK(n91), .C(n38) );
  CKNXD16 U91 ( .I(n38), .ZN(FrameOut[11]) );
  CKND0 U92 ( .CLK(n126), .CN(n91) );
  CKBD0 U93 ( .CLK(n89), .C(n40) );
  CKNXD16 U94 ( .I(n40), .ZN(FrameOut[59]) );
  CKND0 U95 ( .CLK(n102), .CN(n89) );
  CKBD0 U96 ( .CLK(n87), .C(n42) );
  CKNXD16 U97 ( .I(n42), .ZN(FrameOut[13]) );
  CKND0 U98 ( .CLK(n124), .CN(n87) );
  CKBD0 U99 ( .CLK(n85), .C(n44) );
  CKNXD16 U100 ( .I(n44), .ZN(FrameOut[57]) );
  CKND0 U101 ( .CLK(n104), .CN(n85) );
  CKBD0 U102 ( .CLK(n83), .C(n46) );
  CKNXD16 U103 ( .I(n46), .ZN(FrameOut[15]) );
  CKND0 U104 ( .CLK(n122), .CN(n83) );
  CKBD0 U105 ( .CLK(n81), .C(n48) );
  CKNXD16 U106 ( .I(n48), .ZN(FrameOut[47]) );
  CKND0 U107 ( .CLK(n106), .CN(n81) );
  CKBD0 U108 ( .CLK(n79), .C(n50) );
  CKNXD16 U109 ( .I(n50), .ZN(FrameOut[25]) );
  CKND0 U110 ( .CLK(n120), .CN(n79) );
  CKBD0 U111 ( .CLK(n77), .C(n52) );
  CKNXD16 U112 ( .I(n52), .ZN(FrameOut[45]) );
  CKND0 U113 ( .CLK(n108), .CN(n77) );
  CKBD0 U114 ( .CLK(n75), .C(n54) );
  CKNXD16 U115 ( .I(n54), .ZN(FrameOut[27]) );
  CKND0 U116 ( .CLK(n118), .CN(n75) );
  CKBD0 U117 ( .CLK(n73), .C(n56) );
  CKNXD16 U118 ( .I(n56), .ZN(FrameOut[43]) );
  CKND0 U119 ( .CLK(n110), .CN(n73) );
  CKBD0 U120 ( .CLK(n71), .C(n58) );
  CKNXD16 U121 ( .I(n58), .ZN(FrameOut[29]) );
  CKND0 U122 ( .CLK(n116), .CN(n71) );
  CKBD0 U123 ( .CLK(n67), .C(n60) );
  CKNXD16 U124 ( .I(n60), .ZN(FrameOut[31]) );
  CKND0 U125 ( .CLK(n114), .CN(n67) );
  CKBD0 U126 ( .CLK(n66), .C(n62) );
  CKNXD16 U127 ( .I(n62), .ZN(FrameOut[40]) );
  CKBD0 U128 ( .CLK(n69), .C(n64) );
  CKNXD16 U129 ( .I(n64), .ZN(FrameOut[41]) );
  CKND0 U130 ( .CLK(n113), .CN(n66) );
  CKND0 U131 ( .CLK(n112), .CN(n69) );
  TIEL U132 ( .ZN(FrameOut[0]) );
  TIEL U133 ( .ZN(FrameOut[1]) );
  TIEL U134 ( .ZN(FrameOut[2]) );
  TIEL U135 ( .ZN(FrameOut[3]) );
  TIEL U136 ( .ZN(FrameOut[4]) );
  TIEL U137 ( .ZN(FrameOut[5]) );
  TIEL U138 ( .ZN(FrameOut[6]) );
  TIEL U139 ( .ZN(FrameOut[7]) );
  TIEL U140 ( .ZN(FrameOut[16]) );
  TIEL U141 ( .ZN(FrameOut[17]) );
  TIEL U142 ( .ZN(FrameOut[18]) );
  TIEH U143 ( .Z(FrameOut[19]) );
  TIEL U144 ( .ZN(FrameOut[20]) );
  TIEL U145 ( .ZN(FrameOut[21]) );
  TIEL U146 ( .ZN(FrameOut[22]) );
  TIEL U147 ( .ZN(FrameOut[23]) );
  TIEL U148 ( .ZN(FrameOut[32]) );
  TIEL U149 ( .ZN(FrameOut[33]) );
  TIEL U150 ( .ZN(FrameOut[34]) );
  TIEL U151 ( .ZN(FrameOut[35]) );
  TIEH U152 ( .Z(FrameOut[36]) );
  TIEL U153 ( .ZN(FrameOut[37]) );
  TIEL U154 ( .ZN(FrameOut[38]) );
  TIEL U155 ( .ZN(FrameOut[39]) );
  TIEL U156 ( .ZN(FrameOut[48]) );
  TIEL U157 ( .ZN(FrameOut[49]) );
  TIEL U158 ( .ZN(FrameOut[50]) );
  TIEH U159 ( .Z(FrameOut[51]) );
  TIEH U160 ( .Z(FrameOut[52]) );
  TIEL U161 ( .ZN(FrameOut[53]) );
  TIEL U162 ( .ZN(FrameOut[54]) );
  TIEL U163 ( .ZN(FrameOut[55]) );
endmodule

