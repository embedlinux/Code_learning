
module Decoder1024 ( AdrEna, Address );
  output [1023:0] AdrEna;
  input [9:0] Address;
  wire   \*Logic0* , \DL2[0].tempL2[15] , \DL2[0].tempL2[14] ,
         \DL2[0].tempL2[13] , \DL2[0].tempL2[12] , \DL2[0].tempL2[11] ,
         \DL2[0].tempL2[10] , \DL2[0].tempL2[9] , \DL2[0].tempL2[8] ,
         \DL2[0].tempL2[7] , \DL2[0].tempL2[6] , \DL2[0].tempL2[5] ,
         \DL2[0].tempL2[4] , \DL2[0].tempL2[3] , \DL2[0].tempL2[2] ,
         \DL2[0].tempL2[1] , \DL2[0].tempL2[0] , \DL2[1].tempL2[15] ,
         \DL2[1].tempL2[14] , \DL2[1].tempL2[13] , \DL2[1].tempL2[12] ,
         \DL2[1].tempL2[11] , \DL2[1].tempL2[10] , \DL2[1].tempL2[9] ,
         \DL2[1].tempL2[8] , \DL2[1].tempL2[7] , \DL2[1].tempL2[6] ,
         \DL2[1].tempL2[5] , \DL2[1].tempL2[4] , \DL2[1].tempL2[3] ,
         \DL2[1].tempL2[2] , \DL2[1].tempL2[1] , \DL2[1].tempL2[0] ,
         \DL2[2].tempL2[15] , \DL2[2].tempL2[14] , \DL2[2].tempL2[13] ,
         \DL2[2].tempL2[12] , \DL2[2].tempL2[11] , \DL2[2].tempL2[10] ,
         \DL2[2].tempL2[9] , \DL2[2].tempL2[8] , \DL2[2].tempL2[7] ,
         \DL2[2].tempL2[6] , \DL2[2].tempL2[5] , \DL2[2].tempL2[4] ,
         \DL2[2].tempL2[3] , \DL2[2].tempL2[2] , \DL2[2].tempL2[1] ,
         \DL2[2].tempL2[0] , \DL2[3].tempL2[15] , \DL2[3].tempL2[14] ,
         \DL2[3].tempL2[13] , \DL2[3].tempL2[12] , \DL2[3].tempL2[11] ,
         \DL2[3].tempL2[10] , \DL2[3].tempL2[9] , \DL2[3].tempL2[8] ,
         \DL2[3].tempL2[7] , \DL2[3].tempL2[6] , \DL2[3].tempL2[5] ,
         \DL2[3].tempL2[4] , \DL2[3].tempL2[3] , \DL2[3].tempL2[2] ,
         \DL2[3].tempL2[1] , \DL2[3].tempL2[0] , \DL3[0].tempL3[15] ,
         \DL3[0].tempL3[14] , \DL3[0].tempL3[13] , \DL3[0].tempL3[12] ,
         \DL3[0].tempL3[11] , \DL3[0].tempL3[10] , \DL3[0].tempL3[9] ,
         \DL3[0].tempL3[8] , \DL3[0].tempL3[7] , \DL3[0].tempL3[6] ,
         \DL3[0].tempL3[5] , \DL3[0].tempL3[4] , \DL3[0].tempL3[3] ,
         \DL3[0].tempL3[2] , \DL3[0].tempL3[1] , \DL3[0].tempL3[0] ,
         \DL3[1].tempL3[15] , \DL3[1].tempL3[14] , \DL3[1].tempL3[13] ,
         \DL3[1].tempL3[12] , \DL3[1].tempL3[11] , \DL3[1].tempL3[10] ,
         \DL3[1].tempL3[9] , \DL3[1].tempL3[8] , \DL3[1].tempL3[7] ,
         \DL3[1].tempL3[6] , \DL3[1].tempL3[5] , \DL3[1].tempL3[4] ,
         \DL3[1].tempL3[3] , \DL3[1].tempL3[2] , \DL3[1].tempL3[1] ,
         \DL3[1].tempL3[0] , \DL3[2].tempL3[15] , \DL3[2].tempL3[14] ,
         \DL3[2].tempL3[13] , \DL3[2].tempL3[12] , \DL3[2].tempL3[11] ,
         \DL3[2].tempL3[10] , \DL3[2].tempL3[9] , \DL3[2].tempL3[8] ,
         \DL3[2].tempL3[7] , \DL3[2].tempL3[6] , \DL3[2].tempL3[5] ,
         \DL3[2].tempL3[4] , \DL3[2].tempL3[3] , \DL3[2].tempL3[2] ,
         \DL3[2].tempL3[1] , \DL3[2].tempL3[0] , \DL3[3].tempL3[15] ,
         \DL3[3].tempL3[14] , \DL3[3].tempL3[13] , \DL3[3].tempL3[12] ,
         \DL3[3].tempL3[11] , \DL3[3].tempL3[10] , \DL3[3].tempL3[9] ,
         \DL3[3].tempL3[8] , \DL3[3].tempL3[7] , \DL3[3].tempL3[6] ,
         \DL3[3].tempL3[5] , \DL3[3].tempL3[4] , \DL3[3].tempL3[3] ,
         \DL3[3].tempL3[2] , \DL3[3].tempL3[1] , \DL3[3].tempL3[0] ,
         \DL3[4].tempL3[15] , \DL3[4].tempL3[14] , \DL3[4].tempL3[13] ,
         \DL3[4].tempL3[12] , \DL3[4].tempL3[11] , \DL3[4].tempL3[10] ,
         \DL3[4].tempL3[9] , \DL3[4].tempL3[8] , \DL3[4].tempL3[7] ,
         \DL3[4].tempL3[6] , \DL3[4].tempL3[5] , \DL3[4].tempL3[4] ,
         \DL3[4].tempL3[3] , \DL3[4].tempL3[2] , \DL3[4].tempL3[1] ,
         \DL3[4].tempL3[0] , \DL3[5].tempL3[15] , \DL3[5].tempL3[14] ,
         \DL3[5].tempL3[13] , \DL3[5].tempL3[12] , \DL3[5].tempL3[11] ,
         \DL3[5].tempL3[10] , \DL3[5].tempL3[9] , \DL3[5].tempL3[8] ,
         \DL3[5].tempL3[7] , \DL3[5].tempL3[6] , \DL3[5].tempL3[5] ,
         \DL3[5].tempL3[4] , \DL3[5].tempL3[3] , \DL3[5].tempL3[2] ,
         \DL3[5].tempL3[1] , \DL3[5].tempL3[0] , \DL3[6].tempL3[15] ,
         \DL3[6].tempL3[14] , \DL3[6].tempL3[13] , \DL3[6].tempL3[12] ,
         \DL3[6].tempL3[11] , \DL3[6].tempL3[10] , \DL3[6].tempL3[9] ,
         \DL3[6].tempL3[8] , \DL3[6].tempL3[7] , \DL3[6].tempL3[6] ,
         \DL3[6].tempL3[5] , \DL3[6].tempL3[4] , \DL3[6].tempL3[3] ,
         \DL3[6].tempL3[2] , \DL3[6].tempL3[1] , \DL3[6].tempL3[0] ,
         \DL3[7].tempL3[15] , \DL3[7].tempL3[14] , \DL3[7].tempL3[13] ,
         \DL3[7].tempL3[12] , \DL3[7].tempL3[11] , \DL3[7].tempL3[10] ,
         \DL3[7].tempL3[9] , \DL3[7].tempL3[8] , \DL3[7].tempL3[7] ,
         \DL3[7].tempL3[6] , \DL3[7].tempL3[5] , \DL3[7].tempL3[4] ,
         \DL3[7].tempL3[3] , \DL3[7].tempL3[2] , \DL3[7].tempL3[1] ,
         \DL3[7].tempL3[0] , \DL3[8].tempL3[15] , \DL3[8].tempL3[14] ,
         \DL3[8].tempL3[13] , \DL3[8].tempL3[12] , \DL3[8].tempL3[11] ,
         \DL3[8].tempL3[10] , \DL3[8].tempL3[9] , \DL3[8].tempL3[8] ,
         \DL3[8].tempL3[7] , \DL3[8].tempL3[6] , \DL3[8].tempL3[5] ,
         \DL3[8].tempL3[4] , \DL3[8].tempL3[3] , \DL3[8].tempL3[2] ,
         \DL3[8].tempL3[1] , \DL3[8].tempL3[0] , \DL3[9].tempL3[15] ,
         \DL3[9].tempL3[14] , \DL3[9].tempL3[13] , \DL3[9].tempL3[12] ,
         \DL3[9].tempL3[11] , \DL3[9].tempL3[10] , \DL3[9].tempL3[9] ,
         \DL3[9].tempL3[8] , \DL3[9].tempL3[7] , \DL3[9].tempL3[6] ,
         \DL3[9].tempL3[5] , \DL3[9].tempL3[4] , \DL3[9].tempL3[3] ,
         \DL3[9].tempL3[2] , \DL3[9].tempL3[1] , \DL3[9].tempL3[0] ,
         \DL3[10].tempL3[15] , \DL3[10].tempL3[14] , \DL3[10].tempL3[13] ,
         \DL3[10].tempL3[12] , \DL3[10].tempL3[11] , \DL3[10].tempL3[10] ,
         \DL3[10].tempL3[9] , \DL3[10].tempL3[8] , \DL3[10].tempL3[7] ,
         \DL3[10].tempL3[6] , \DL3[10].tempL3[5] , \DL3[10].tempL3[4] ,
         \DL3[10].tempL3[3] , \DL3[10].tempL3[2] , \DL3[10].tempL3[1] ,
         \DL3[10].tempL3[0] , \DL3[11].tempL3[15] , \DL3[11].tempL3[14] ,
         \DL3[11].tempL3[13] , \DL3[11].tempL3[12] , \DL3[11].tempL3[11] ,
         \DL3[11].tempL3[10] , \DL3[11].tempL3[9] , \DL3[11].tempL3[8] ,
         \DL3[11].tempL3[7] , \DL3[11].tempL3[6] , \DL3[11].tempL3[5] ,
         \DL3[11].tempL3[4] , \DL3[11].tempL3[3] , \DL3[11].tempL3[2] ,
         \DL3[11].tempL3[1] , \DL3[11].tempL3[0] , \DL3[12].tempL3[15] ,
         \DL3[12].tempL3[14] , \DL3[12].tempL3[13] , \DL3[12].tempL3[12] ,
         \DL3[12].tempL3[11] , \DL3[12].tempL3[10] , \DL3[12].tempL3[9] ,
         \DL3[12].tempL3[8] , \DL3[12].tempL3[7] , \DL3[12].tempL3[6] ,
         \DL3[12].tempL3[5] , \DL3[12].tempL3[4] , \DL3[12].tempL3[3] ,
         \DL3[12].tempL3[2] , \DL3[12].tempL3[1] , \DL3[12].tempL3[0] ,
         \DL3[13].tempL3[15] , \DL3[13].tempL3[14] , \DL3[13].tempL3[13] ,
         \DL3[13].tempL3[12] , \DL3[13].tempL3[11] , \DL3[13].tempL3[10] ,
         \DL3[13].tempL3[9] , \DL3[13].tempL3[8] , \DL3[13].tempL3[7] ,
         \DL3[13].tempL3[6] , \DL3[13].tempL3[5] , \DL3[13].tempL3[4] ,
         \DL3[13].tempL3[3] , \DL3[13].tempL3[2] , \DL3[13].tempL3[1] ,
         \DL3[13].tempL3[0] , \DL3[14].tempL3[15] , \DL3[14].tempL3[14] ,
         \DL3[14].tempL3[13] , \DL3[14].tempL3[12] , \DL3[14].tempL3[11] ,
         \DL3[14].tempL3[10] , \DL3[14].tempL3[9] , \DL3[14].tempL3[8] ,
         \DL3[14].tempL3[7] , \DL3[14].tempL3[6] , \DL3[14].tempL3[5] ,
         \DL3[14].tempL3[4] , \DL3[14].tempL3[3] , \DL3[14].tempL3[2] ,
         \DL3[14].tempL3[1] , \DL3[14].tempL3[0] , \DL3[15].tempL3[15] ,
         \DL3[15].tempL3[14] , \DL3[15].tempL3[13] , \DL3[15].tempL3[12] ,
         \DL3[15].tempL3[11] , \DL3[15].tempL3[10] , \DL3[15].tempL3[9] ,
         \DL3[15].tempL3[8] , \DL3[15].tempL3[7] , \DL3[15].tempL3[6] ,
         \DL3[15].tempL3[5] , \DL3[15].tempL3[4] , \DL3[15].tempL3[3] ,
         \DL3[15].tempL3[2] , \DL3[15].tempL3[1] , \DL3[15].tempL3[0] ,
         \DL3[16].tempL3[15] , \DL3[16].tempL3[14] , \DL3[16].tempL3[13] ,
         \DL3[16].tempL3[12] , \DL3[16].tempL3[11] , \DL3[16].tempL3[10] ,
         \DL3[16].tempL3[9] , \DL3[16].tempL3[8] , \DL3[16].tempL3[7] ,
         \DL3[16].tempL3[6] , \DL3[16].tempL3[5] , \DL3[16].tempL3[4] ,
         \DL3[16].tempL3[3] , \DL3[16].tempL3[2] , \DL3[16].tempL3[1] ,
         \DL3[16].tempL3[0] , \DL3[17].tempL3[15] , \DL3[17].tempL3[14] ,
         \DL3[17].tempL3[13] , \DL3[17].tempL3[12] , \DL3[17].tempL3[11] ,
         \DL3[17].tempL3[10] , \DL3[17].tempL3[9] , \DL3[17].tempL3[8] ,
         \DL3[17].tempL3[7] , \DL3[17].tempL3[6] , \DL3[17].tempL3[5] ,
         \DL3[17].tempL3[4] , \DL3[17].tempL3[3] , \DL3[17].tempL3[2] ,
         \DL3[17].tempL3[1] , \DL3[17].tempL3[0] , \DL3[18].tempL3[15] ,
         \DL3[18].tempL3[14] , \DL3[18].tempL3[13] , \DL3[18].tempL3[12] ,
         \DL3[18].tempL3[11] , \DL3[18].tempL3[10] , \DL3[18].tempL3[9] ,
         \DL3[18].tempL3[8] , \DL3[18].tempL3[7] , \DL3[18].tempL3[6] ,
         \DL3[18].tempL3[5] , \DL3[18].tempL3[4] , \DL3[18].tempL3[3] ,
         \DL3[18].tempL3[2] , \DL3[18].tempL3[1] , \DL3[18].tempL3[0] ,
         \DL3[19].tempL3[15] , \DL3[19].tempL3[14] , \DL3[19].tempL3[13] ,
         \DL3[19].tempL3[12] , \DL3[19].tempL3[11] , \DL3[19].tempL3[10] ,
         \DL3[19].tempL3[9] , \DL3[19].tempL3[8] , \DL3[19].tempL3[7] ,
         \DL3[19].tempL3[6] , \DL3[19].tempL3[5] , \DL3[19].tempL3[4] ,
         \DL3[19].tempL3[3] , \DL3[19].tempL3[2] , \DL3[19].tempL3[1] ,
         \DL3[19].tempL3[0] , \DL3[20].tempL3[15] , \DL3[20].tempL3[14] ,
         \DL3[20].tempL3[13] , \DL3[20].tempL3[12] , \DL3[20].tempL3[11] ,
         \DL3[20].tempL3[10] , \DL3[20].tempL3[9] , \DL3[20].tempL3[8] ,
         \DL3[20].tempL3[7] , \DL3[20].tempL3[6] , \DL3[20].tempL3[5] ,
         \DL3[20].tempL3[4] , \DL3[20].tempL3[3] , \DL3[20].tempL3[2] ,
         \DL3[20].tempL3[1] , \DL3[20].tempL3[0] , \DL3[21].tempL3[15] ,
         \DL3[21].tempL3[14] , \DL3[21].tempL3[13] , \DL3[21].tempL3[12] ,
         \DL3[21].tempL3[11] , \DL3[21].tempL3[10] , \DL3[21].tempL3[9] ,
         \DL3[21].tempL3[8] , \DL3[21].tempL3[7] , \DL3[21].tempL3[6] ,
         \DL3[21].tempL3[5] , \DL3[21].tempL3[4] , \DL3[21].tempL3[3] ,
         \DL3[21].tempL3[2] , \DL3[21].tempL3[1] , \DL3[21].tempL3[0] ,
         \DL3[22].tempL3[15] , \DL3[22].tempL3[14] , \DL3[22].tempL3[13] ,
         \DL3[22].tempL3[12] , \DL3[22].tempL3[11] , \DL3[22].tempL3[10] ,
         \DL3[22].tempL3[9] , \DL3[22].tempL3[8] , \DL3[22].tempL3[7] ,
         \DL3[22].tempL3[6] , \DL3[22].tempL3[5] , \DL3[22].tempL3[4] ,
         \DL3[22].tempL3[3] , \DL3[22].tempL3[2] , \DL3[22].tempL3[1] ,
         \DL3[22].tempL3[0] , \DL3[23].tempL3[15] , \DL3[23].tempL3[14] ,
         \DL3[23].tempL3[13] , \DL3[23].tempL3[12] , \DL3[23].tempL3[11] ,
         \DL3[23].tempL3[10] , \DL3[23].tempL3[9] , \DL3[23].tempL3[8] ,
         \DL3[23].tempL3[7] , \DL3[23].tempL3[6] , \DL3[23].tempL3[5] ,
         \DL3[23].tempL3[4] , \DL3[23].tempL3[3] , \DL3[23].tempL3[2] ,
         \DL3[23].tempL3[1] , \DL3[23].tempL3[0] , \DL3[24].tempL3[15] ,
         \DL3[24].tempL3[14] , \DL3[24].tempL3[13] , \DL3[24].tempL3[12] ,
         \DL3[24].tempL3[11] , \DL3[24].tempL3[10] , \DL3[24].tempL3[9] ,
         \DL3[24].tempL3[8] , \DL3[24].tempL3[7] , \DL3[24].tempL3[6] ,
         \DL3[24].tempL3[5] , \DL3[24].tempL3[4] , \DL3[24].tempL3[3] ,
         \DL3[24].tempL3[2] , \DL3[24].tempL3[1] , \DL3[24].tempL3[0] ,
         \DL3[25].tempL3[15] , \DL3[25].tempL3[14] , \DL3[25].tempL3[13] ,
         \DL3[25].tempL3[12] , \DL3[25].tempL3[11] , \DL3[25].tempL3[10] ,
         \DL3[25].tempL3[9] , \DL3[25].tempL3[8] , \DL3[25].tempL3[7] ,
         \DL3[25].tempL3[6] , \DL3[25].tempL3[5] , \DL3[25].tempL3[4] ,
         \DL3[25].tempL3[3] , \DL3[25].tempL3[2] , \DL3[25].tempL3[1] ,
         \DL3[25].tempL3[0] , \DL3[26].tempL3[15] , \DL3[26].tempL3[14] ,
         \DL3[26].tempL3[13] , \DL3[26].tempL3[12] , \DL3[26].tempL3[11] ,
         \DL3[26].tempL3[10] , \DL3[26].tempL3[9] , \DL3[26].tempL3[8] ,
         \DL3[26].tempL3[7] , \DL3[26].tempL3[6] , \DL3[26].tempL3[5] ,
         \DL3[26].tempL3[4] , \DL3[26].tempL3[3] , \DL3[26].tempL3[2] ,
         \DL3[26].tempL3[1] , \DL3[26].tempL3[0] , \DL3[27].tempL3[15] ,
         \DL3[27].tempL3[14] , \DL3[27].tempL3[13] , \DL3[27].tempL3[12] ,
         \DL3[27].tempL3[11] , \DL3[27].tempL3[10] , \DL3[27].tempL3[9] ,
         \DL3[27].tempL3[8] , \DL3[27].tempL3[7] , \DL3[27].tempL3[6] ,
         \DL3[27].tempL3[5] , \DL3[27].tempL3[4] , \DL3[27].tempL3[3] ,
         \DL3[27].tempL3[2] , \DL3[27].tempL3[1] , \DL3[27].tempL3[0] ,
         \DL3[28].tempL3[15] , \DL3[28].tempL3[14] , \DL3[28].tempL3[13] ,
         \DL3[28].tempL3[12] , \DL3[28].tempL3[11] , \DL3[28].tempL3[10] ,
         \DL3[28].tempL3[9] , \DL3[28].tempL3[8] , \DL3[28].tempL3[7] ,
         \DL3[28].tempL3[6] , \DL3[28].tempL3[5] , \DL3[28].tempL3[4] ,
         \DL3[28].tempL3[3] , \DL3[28].tempL3[2] , \DL3[28].tempL3[1] ,
         \DL3[28].tempL3[0] , \DL3[29].tempL3[15] , \DL3[29].tempL3[14] ,
         \DL3[29].tempL3[13] , \DL3[29].tempL3[12] , \DL3[29].tempL3[11] ,
         \DL3[29].tempL3[10] , \DL3[29].tempL3[9] , \DL3[29].tempL3[8] ,
         \DL3[29].tempL3[7] , \DL3[29].tempL3[6] , \DL3[29].tempL3[5] ,
         \DL3[29].tempL3[4] , \DL3[29].tempL3[3] , \DL3[29].tempL3[2] ,
         \DL3[29].tempL3[1] , \DL3[29].tempL3[0] , \DL3[30].tempL3[15] ,
         \DL3[30].tempL3[14] , \DL3[30].tempL3[13] , \DL3[30].tempL3[12] ,
         \DL3[30].tempL3[11] , \DL3[30].tempL3[10] , \DL3[30].tempL3[9] ,
         \DL3[30].tempL3[8] , \DL3[30].tempL3[7] , \DL3[30].tempL3[6] ,
         \DL3[30].tempL3[5] , \DL3[30].tempL3[4] , \DL3[30].tempL3[3] ,
         \DL3[30].tempL3[2] , \DL3[30].tempL3[1] , \DL3[30].tempL3[0] ,
         \DL3[31].tempL3[15] , \DL3[31].tempL3[14] , \DL3[31].tempL3[13] ,
         \DL3[31].tempL3[12] , \DL3[31].tempL3[11] , \DL3[31].tempL3[10] ,
         \DL3[31].tempL3[9] , \DL3[31].tempL3[8] , \DL3[31].tempL3[7] ,
         \DL3[31].tempL3[6] , \DL3[31].tempL3[5] , \DL3[31].tempL3[4] ,
         \DL3[31].tempL3[3] , \DL3[31].tempL3[2] , \DL3[31].tempL3[1] ,
         \DL3[31].tempL3[0] , \DL3[32].tempL3[15] , \DL3[32].tempL3[14] ,
         \DL3[32].tempL3[13] , \DL3[32].tempL3[12] , \DL3[32].tempL3[11] ,
         \DL3[32].tempL3[10] , \DL3[32].tempL3[9] , \DL3[32].tempL3[8] ,
         \DL3[32].tempL3[7] , \DL3[32].tempL3[6] , \DL3[32].tempL3[5] ,
         \DL3[32].tempL3[4] , \DL3[32].tempL3[3] , \DL3[32].tempL3[2] ,
         \DL3[32].tempL3[1] , \DL3[32].tempL3[0] , \DL3[33].tempL3[15] ,
         \DL3[33].tempL3[14] , \DL3[33].tempL3[13] , \DL3[33].tempL3[12] ,
         \DL3[33].tempL3[11] , \DL3[33].tempL3[10] , \DL3[33].tempL3[9] ,
         \DL3[33].tempL3[8] , \DL3[33].tempL3[7] , \DL3[33].tempL3[6] ,
         \DL3[33].tempL3[5] , \DL3[33].tempL3[4] , \DL3[33].tempL3[3] ,
         \DL3[33].tempL3[2] , \DL3[33].tempL3[1] , \DL3[33].tempL3[0] ,
         \DL3[34].tempL3[15] , \DL3[34].tempL3[14] , \DL3[34].tempL3[13] ,
         \DL3[34].tempL3[12] , \DL3[34].tempL3[11] , \DL3[34].tempL3[10] ,
         \DL3[34].tempL3[9] , \DL3[34].tempL3[8] , \DL3[34].tempL3[7] ,
         \DL3[34].tempL3[6] , \DL3[34].tempL3[5] , \DL3[34].tempL3[4] ,
         \DL3[34].tempL3[3] , \DL3[34].tempL3[2] , \DL3[34].tempL3[1] ,
         \DL3[34].tempL3[0] , \DL3[35].tempL3[15] , \DL3[35].tempL3[14] ,
         \DL3[35].tempL3[13] , \DL3[35].tempL3[12] , \DL3[35].tempL3[11] ,
         \DL3[35].tempL3[10] , \DL3[35].tempL3[9] , \DL3[35].tempL3[8] ,
         \DL3[35].tempL3[7] , \DL3[35].tempL3[6] , \DL3[35].tempL3[5] ,
         \DL3[35].tempL3[4] , \DL3[35].tempL3[3] , \DL3[35].tempL3[2] ,
         \DL3[35].tempL3[1] , \DL3[35].tempL3[0] , \DL3[36].tempL3[15] ,
         \DL3[36].tempL3[14] , \DL3[36].tempL3[13] , \DL3[36].tempL3[12] ,
         \DL3[36].tempL3[11] , \DL3[36].tempL3[10] , \DL3[36].tempL3[9] ,
         \DL3[36].tempL3[8] , \DL3[36].tempL3[7] , \DL3[36].tempL3[6] ,
         \DL3[36].tempL3[5] , \DL3[36].tempL3[4] , \DL3[36].tempL3[3] ,
         \DL3[36].tempL3[2] , \DL3[36].tempL3[1] , \DL3[36].tempL3[0] ,
         \DL3[37].tempL3[15] , \DL3[37].tempL3[14] , \DL3[37].tempL3[13] ,
         \DL3[37].tempL3[12] , \DL3[37].tempL3[11] , \DL3[37].tempL3[10] ,
         \DL3[37].tempL3[9] , \DL3[37].tempL3[8] , \DL3[37].tempL3[7] ,
         \DL3[37].tempL3[6] , \DL3[37].tempL3[5] , \DL3[37].tempL3[4] ,
         \DL3[37].tempL3[3] , \DL3[37].tempL3[2] , \DL3[37].tempL3[1] ,
         \DL3[37].tempL3[0] , \DL3[38].tempL3[15] , \DL3[38].tempL3[14] ,
         \DL3[38].tempL3[13] , \DL3[38].tempL3[12] , \DL3[38].tempL3[11] ,
         \DL3[38].tempL3[10] , \DL3[38].tempL3[9] , \DL3[38].tempL3[8] ,
         \DL3[38].tempL3[7] , \DL3[38].tempL3[6] , \DL3[38].tempL3[5] ,
         \DL3[38].tempL3[4] , \DL3[38].tempL3[3] , \DL3[38].tempL3[2] ,
         \DL3[38].tempL3[1] , \DL3[38].tempL3[0] , \DL3[39].tempL3[15] ,
         \DL3[39].tempL3[14] , \DL3[39].tempL3[13] , \DL3[39].tempL3[12] ,
         \DL3[39].tempL3[11] , \DL3[39].tempL3[10] , \DL3[39].tempL3[9] ,
         \DL3[39].tempL3[8] , \DL3[39].tempL3[7] , \DL3[39].tempL3[6] ,
         \DL3[39].tempL3[5] , \DL3[39].tempL3[4] , \DL3[39].tempL3[3] ,
         \DL3[39].tempL3[2] , \DL3[39].tempL3[1] , \DL3[39].tempL3[0] ,
         \DL3[40].tempL3[15] , \DL3[40].tempL3[14] , \DL3[40].tempL3[13] ,
         \DL3[40].tempL3[12] , \DL3[40].tempL3[11] , \DL3[40].tempL3[10] ,
         \DL3[40].tempL3[9] , \DL3[40].tempL3[8] , \DL3[40].tempL3[7] ,
         \DL3[40].tempL3[6] , \DL3[40].tempL3[5] , \DL3[40].tempL3[4] ,
         \DL3[40].tempL3[3] , \DL3[40].tempL3[2] , \DL3[40].tempL3[1] ,
         \DL3[40].tempL3[0] , \DL3[41].tempL3[15] , \DL3[41].tempL3[14] ,
         \DL3[41].tempL3[13] , \DL3[41].tempL3[12] , \DL3[41].tempL3[11] ,
         \DL3[41].tempL3[10] , \DL3[41].tempL3[9] , \DL3[41].tempL3[8] ,
         \DL3[41].tempL3[7] , \DL3[41].tempL3[6] , \DL3[41].tempL3[5] ,
         \DL3[41].tempL3[4] , \DL3[41].tempL3[3] , \DL3[41].tempL3[2] ,
         \DL3[41].tempL3[1] , \DL3[41].tempL3[0] , \DL3[42].tempL3[15] ,
         \DL3[42].tempL3[14] , \DL3[42].tempL3[13] , \DL3[42].tempL3[12] ,
         \DL3[42].tempL3[11] , \DL3[42].tempL3[10] , \DL3[42].tempL3[9] ,
         \DL3[42].tempL3[8] , \DL3[42].tempL3[7] , \DL3[42].tempL3[6] ,
         \DL3[42].tempL3[5] , \DL3[42].tempL3[4] , \DL3[42].tempL3[3] ,
         \DL3[42].tempL3[2] , \DL3[42].tempL3[1] , \DL3[42].tempL3[0] ,
         \DL3[43].tempL3[15] , \DL3[43].tempL3[14] , \DL3[43].tempL3[13] ,
         \DL3[43].tempL3[12] , \DL3[43].tempL3[11] , \DL3[43].tempL3[10] ,
         \DL3[43].tempL3[9] , \DL3[43].tempL3[8] , \DL3[43].tempL3[7] ,
         \DL3[43].tempL3[6] , \DL3[43].tempL3[5] , \DL3[43].tempL3[4] ,
         \DL3[43].tempL3[3] , \DL3[43].tempL3[2] , \DL3[43].tempL3[1] ,
         \DL3[43].tempL3[0] , \DL3[44].tempL3[15] , \DL3[44].tempL3[14] ,
         \DL3[44].tempL3[13] , \DL3[44].tempL3[12] , \DL3[44].tempL3[11] ,
         \DL3[44].tempL3[10] , \DL3[44].tempL3[9] , \DL3[44].tempL3[8] ,
         \DL3[44].tempL3[7] , \DL3[44].tempL3[6] , \DL3[44].tempL3[5] ,
         \DL3[44].tempL3[4] , \DL3[44].tempL3[3] , \DL3[44].tempL3[2] ,
         \DL3[44].tempL3[1] , \DL3[44].tempL3[0] , \DL3[45].tempL3[15] ,
         \DL3[45].tempL3[14] , \DL3[45].tempL3[13] , \DL3[45].tempL3[12] ,
         \DL3[45].tempL3[11] , \DL3[45].tempL3[10] , \DL3[45].tempL3[9] ,
         \DL3[45].tempL3[8] , \DL3[45].tempL3[7] , \DL3[45].tempL3[6] ,
         \DL3[45].tempL3[5] , \DL3[45].tempL3[4] , \DL3[45].tempL3[3] ,
         \DL3[45].tempL3[2] , \DL3[45].tempL3[1] , \DL3[45].tempL3[0] ,
         \DL3[46].tempL3[15] , \DL3[46].tempL3[14] , \DL3[46].tempL3[13] ,
         \DL3[46].tempL3[12] , \DL3[46].tempL3[11] , \DL3[46].tempL3[10] ,
         \DL3[46].tempL3[9] , \DL3[46].tempL3[8] , \DL3[46].tempL3[7] ,
         \DL3[46].tempL3[6] , \DL3[46].tempL3[5] , \DL3[46].tempL3[4] ,
         \DL3[46].tempL3[3] , \DL3[46].tempL3[2] , \DL3[46].tempL3[1] ,
         \DL3[46].tempL3[0] , \DL3[47].tempL3[15] , \DL3[47].tempL3[14] ,
         \DL3[47].tempL3[13] , \DL3[47].tempL3[12] , \DL3[47].tempL3[11] ,
         \DL3[47].tempL3[10] , \DL3[47].tempL3[9] , \DL3[47].tempL3[8] ,
         \DL3[47].tempL3[7] , \DL3[47].tempL3[6] , \DL3[47].tempL3[5] ,
         \DL3[47].tempL3[4] , \DL3[47].tempL3[3] , \DL3[47].tempL3[2] ,
         \DL3[47].tempL3[1] , \DL3[47].tempL3[0] , \DL3[48].tempL3[15] ,
         \DL3[48].tempL3[14] , \DL3[48].tempL3[13] , \DL3[48].tempL3[12] ,
         \DL3[48].tempL3[11] , \DL3[48].tempL3[10] , \DL3[48].tempL3[9] ,
         \DL3[48].tempL3[8] , \DL3[48].tempL3[7] , \DL3[48].tempL3[6] ,
         \DL3[48].tempL3[5] , \DL3[48].tempL3[4] , \DL3[48].tempL3[3] ,
         \DL3[48].tempL3[2] , \DL3[48].tempL3[1] , \DL3[48].tempL3[0] ,
         \DL3[49].tempL3[15] , \DL3[49].tempL3[14] , \DL3[49].tempL3[13] ,
         \DL3[49].tempL3[12] , \DL3[49].tempL3[11] , \DL3[49].tempL3[10] ,
         \DL3[49].tempL3[9] , \DL3[49].tempL3[8] , \DL3[49].tempL3[7] ,
         \DL3[49].tempL3[6] , \DL3[49].tempL3[5] , \DL3[49].tempL3[4] ,
         \DL3[49].tempL3[3] , \DL3[49].tempL3[2] , \DL3[49].tempL3[1] ,
         \DL3[49].tempL3[0] , \DL3[50].tempL3[15] , \DL3[50].tempL3[14] ,
         \DL3[50].tempL3[13] , \DL3[50].tempL3[12] , \DL3[50].tempL3[11] ,
         \DL3[50].tempL3[10] , \DL3[50].tempL3[9] , \DL3[50].tempL3[8] ,
         \DL3[50].tempL3[7] , \DL3[50].tempL3[6] , \DL3[50].tempL3[5] ,
         \DL3[50].tempL3[4] , \DL3[50].tempL3[3] , \DL3[50].tempL3[2] ,
         \DL3[50].tempL3[1] , \DL3[50].tempL3[0] , \DL3[51].tempL3[15] ,
         \DL3[51].tempL3[14] , \DL3[51].tempL3[13] , \DL3[51].tempL3[12] ,
         \DL3[51].tempL3[11] , \DL3[51].tempL3[10] , \DL3[51].tempL3[9] ,
         \DL3[51].tempL3[8] , \DL3[51].tempL3[7] , \DL3[51].tempL3[6] ,
         \DL3[51].tempL3[5] , \DL3[51].tempL3[4] , \DL3[51].tempL3[3] ,
         \DL3[51].tempL3[2] , \DL3[51].tempL3[1] , \DL3[51].tempL3[0] ,
         \DL3[52].tempL3[15] , \DL3[52].tempL3[14] , \DL3[52].tempL3[13] ,
         \DL3[52].tempL3[12] , \DL3[52].tempL3[11] , \DL3[52].tempL3[10] ,
         \DL3[52].tempL3[9] , \DL3[52].tempL3[8] , \DL3[52].tempL3[7] ,
         \DL3[52].tempL3[6] , \DL3[52].tempL3[5] , \DL3[52].tempL3[4] ,
         \DL3[52].tempL3[3] , \DL3[52].tempL3[2] , \DL3[52].tempL3[1] ,
         \DL3[52].tempL3[0] , \DL3[53].tempL3[15] , \DL3[53].tempL3[14] ,
         \DL3[53].tempL3[13] , \DL3[53].tempL3[12] , \DL3[53].tempL3[11] ,
         \DL3[53].tempL3[10] , \DL3[53].tempL3[9] , \DL3[53].tempL3[8] ,
         \DL3[53].tempL3[7] , \DL3[53].tempL3[6] , \DL3[53].tempL3[5] ,
         \DL3[53].tempL3[4] , \DL3[53].tempL3[3] , \DL3[53].tempL3[2] ,
         \DL3[53].tempL3[1] , \DL3[53].tempL3[0] , \DL3[54].tempL3[15] ,
         \DL3[54].tempL3[14] , \DL3[54].tempL3[13] , \DL3[54].tempL3[12] ,
         \DL3[54].tempL3[11] , \DL3[54].tempL3[10] , \DL3[54].tempL3[9] ,
         \DL3[54].tempL3[8] , \DL3[54].tempL3[7] , \DL3[54].tempL3[6] ,
         \DL3[54].tempL3[5] , \DL3[54].tempL3[4] , \DL3[54].tempL3[3] ,
         \DL3[54].tempL3[2] , \DL3[54].tempL3[1] , \DL3[54].tempL3[0] ,
         \DL3[55].tempL3[15] , \DL3[55].tempL3[14] , \DL3[55].tempL3[13] ,
         \DL3[55].tempL3[12] , \DL3[55].tempL3[11] , \DL3[55].tempL3[10] ,
         \DL3[55].tempL3[9] , \DL3[55].tempL3[8] , \DL3[55].tempL3[7] ,
         \DL3[55].tempL3[6] , \DL3[55].tempL3[5] , \DL3[55].tempL3[4] ,
         \DL3[55].tempL3[3] , \DL3[55].tempL3[2] , \DL3[55].tempL3[1] ,
         \DL3[55].tempL3[0] , \DL3[56].tempL3[15] , \DL3[56].tempL3[14] ,
         \DL3[56].tempL3[13] , \DL3[56].tempL3[12] , \DL3[56].tempL3[11] ,
         \DL3[56].tempL3[10] , \DL3[56].tempL3[9] , \DL3[56].tempL3[8] ,
         \DL3[56].tempL3[7] , \DL3[56].tempL3[6] , \DL3[56].tempL3[5] ,
         \DL3[56].tempL3[4] , \DL3[56].tempL3[3] , \DL3[56].tempL3[2] ,
         \DL3[56].tempL3[1] , \DL3[56].tempL3[0] , \DL3[57].tempL3[15] ,
         \DL3[57].tempL3[14] , \DL3[57].tempL3[13] , \DL3[57].tempL3[12] ,
         \DL3[57].tempL3[11] , \DL3[57].tempL3[10] , \DL3[57].tempL3[9] ,
         \DL3[57].tempL3[8] , \DL3[57].tempL3[7] , \DL3[57].tempL3[6] ,
         \DL3[57].tempL3[5] , \DL3[57].tempL3[4] , \DL3[57].tempL3[3] ,
         \DL3[57].tempL3[2] , \DL3[57].tempL3[1] , \DL3[57].tempL3[0] ,
         \DL3[58].tempL3[15] , \DL3[58].tempL3[14] , \DL3[58].tempL3[13] ,
         \DL3[58].tempL3[12] , \DL3[58].tempL3[11] , \DL3[58].tempL3[10] ,
         \DL3[58].tempL3[9] , \DL3[58].tempL3[8] , \DL3[58].tempL3[7] ,
         \DL3[58].tempL3[6] , \DL3[58].tempL3[5] , \DL3[58].tempL3[4] ,
         \DL3[58].tempL3[3] , \DL3[58].tempL3[2] , \DL3[58].tempL3[1] ,
         \DL3[58].tempL3[0] , \DL3[59].tempL3[15] , \DL3[59].tempL3[14] ,
         \DL3[59].tempL3[13] , \DL3[59].tempL3[12] , \DL3[59].tempL3[11] ,
         \DL3[59].tempL3[10] , \DL3[59].tempL3[9] , \DL3[59].tempL3[8] ,
         \DL3[59].tempL3[7] , \DL3[59].tempL3[6] , \DL3[59].tempL3[5] ,
         \DL3[59].tempL3[4] , \DL3[59].tempL3[3] , \DL3[59].tempL3[2] ,
         \DL3[59].tempL3[1] , \DL3[59].tempL3[0] , \DL3[60].tempL3[15] ,
         \DL3[60].tempL3[14] , \DL3[60].tempL3[13] , \DL3[60].tempL3[12] ,
         \DL3[60].tempL3[11] , \DL3[60].tempL3[10] , \DL3[60].tempL3[9] ,
         \DL3[60].tempL3[8] , \DL3[60].tempL3[7] , \DL3[60].tempL3[6] ,
         \DL3[60].tempL3[5] , \DL3[60].tempL3[4] , \DL3[60].tempL3[3] ,
         \DL3[60].tempL3[2] , \DL3[60].tempL3[1] , \DL3[60].tempL3[0] ,
         \DL3[61].tempL3[15] , \DL3[61].tempL3[14] , \DL3[61].tempL3[13] ,
         \DL3[61].tempL3[12] , \DL3[61].tempL3[11] , \DL3[61].tempL3[10] ,
         \DL3[61].tempL3[9] , \DL3[61].tempL3[8] , \DL3[61].tempL3[7] ,
         \DL3[61].tempL3[6] , \DL3[61].tempL3[5] , \DL3[61].tempL3[4] ,
         \DL3[61].tempL3[3] , \DL3[61].tempL3[2] , \DL3[61].tempL3[1] ,
         \DL3[61].tempL3[0] , \DL3[62].tempL3[15] , \DL3[62].tempL3[14] ,
         \DL3[62].tempL3[13] , \DL3[62].tempL3[12] , \DL3[62].tempL3[11] ,
         \DL3[62].tempL3[10] , \DL3[62].tempL3[9] , \DL3[62].tempL3[8] ,
         \DL3[62].tempL3[7] , \DL3[62].tempL3[6] , \DL3[62].tempL3[5] ,
         \DL3[62].tempL3[4] , \DL3[62].tempL3[3] , \DL3[62].tempL3[2] ,
         \DL3[62].tempL3[1] , \DL3[62].tempL3[0] , \DL3[63].tempL3[15] ,
         \DL3[63].tempL3[14] , \DL3[63].tempL3[13] , \DL3[63].tempL3[12] ,
         \DL3[63].tempL3[11] , \DL3[63].tempL3[10] , \DL3[63].tempL3[9] ,
         \DL3[63].tempL3[8] , \DL3[63].tempL3[7] , \DL3[63].tempL3[6] ,
         \DL3[63].tempL3[5] , \DL3[63].tempL3[4] , \DL3[63].tempL3[3] ,
         \DL3[63].tempL3[2] , \DL3[63].tempL3[1] , \DL3[63].tempL3[0] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n225, n227, n229, n231, n233, n235, n237, n239, n241, n243,
         n245, n247, n249, n251, n253, n255, n257, n259, n261, n263, n265,
         n267, n269, n271, n273, n275, n277, n279, n281, n283, n285, n287,
         n289, n291, n293, n295, n297, n299, n301, n303, n305, n307, n309,
         n311, n313, n315, n317, n319, n321, n323, n325, n327, n329, n331,
         n333, n335, n337, n339, n341, n343, n345, n347, n349, n351, n353,
         n355, n357, n359, n361, n363, n365, n367, n369, n371, n373, n375,
         n377, n379, n381, n383, n385, n387, n389, n391, n393, n395, n397,
         n399, n401, n403, n405, n407, n409, n411, n413, n415, n417, n419,
         n421, n423, n425, n427, n429, n431, n433, n435, n437, n439, n441,
         n443, n445, n447, n449, n451, n453, n455, n457, n459, n461, n463,
         n465, n467, n469, n471, n473, n475, n477, n479, n481, n483, n485,
         n487, n489, n491, n493, n495, n497, n499, n501, n503, n505, n507,
         n509, n511, n513, n515, n517, n519, n521, n523, n525, n527, n529,
         n531, n533, n535, n537, n539, n541, n543, n545, n547, n549, n551,
         n553, n555, n557, n559, n561, n563, n565, n567, n569, n571, n573,
         n575, n577, n579, n581, n583, n585, n587, n589, n591, n593, n595,
         n597, n599, n601, n603, n605, n607, n609, n611, n613, n615, n617,
         n619, n621, n623, n625, n627, n629, n631, n633, n635, n637, n639,
         n641, n643, n645, n647, n649, n651, n653, n655, n657, n659, n661,
         n663, n665, n667, n669, n671, n673, n675, n677, n679, n681, n683,
         n685, n687, n689, n691, n693, n695, n697, n699, n701, n703, n705,
         n707, n709, n711, n713, n715, n717, n719, n721, n723, n725, n727,
         n729, n731, n733, n735, n737, n739, n741, n743, n745, n747, n749,
         n751, n753, n755, n757, n759, n761, n763, n765, n767, n769, n771,
         n773, n775, n777, n779, n781, n783, n785, n787, n789, n791, n793,
         n795, n797, n799, n801, n803, n805, n807, n809, n811, n813, n815,
         n817, n819, n821, n823, n825, n827, n829, n831, n833, n835, n837,
         n839, n841, n843, n845, n847, n849, n851, n853, n855, n857, n859,
         n861, n863, n865, n867, n869, n871, n873, n875, n877, n879, n881,
         n883, n885, n887, n889, n891, n893, n895, n897, n899, n901, n903,
         n905, n907, n909, n911, n913, n915, n917, n919, n921, n923, n925,
         n927, n929, n931, n933, n935, n937, n939, n941, n943, n945, n947,
         n949, n951, n953, n955, n957, n959, n961, n963, n965, n967, n969,
         n971, n973, n975, n977, n979, n981, n983, n985, n987, n989, n991,
         n993, n995, n997, n999, n1001, n1003, n1005, n1007, n1009, n1011,
         n1013, n1015, n1017, n1019, n1021, n1023, n1025, n1027, n1029, n1031,
         n1033, n1035, n1037, n1039, n1041, n1043, n1045, n1047, n1049, n1051,
         n1053, n1055, n1057, n1059, n1061, n1063, n1065, n1067, n1069, n1071,
         n1073, n1075, n1077, n1079, n1081, n1083, n1085, n1087, n1089, n1091,
         n1093, n1095, n1097, n1099, n1101, n1103, n1105, n1107, n1109, n1111,
         n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127, n1129, n1131,
         n1133, n1135, n1137, n1139, n1141, n1143, n1145, n1147, n1149, n1151,
         n1153, n1155, n1157, n1159, n1161, n1163, n1165, n1167, n1169, n1171,
         n1173, n1175, n1177, n1179, n1181, n1183, n1185, n1187, n1189, n1191,
         n1193, n1195, n1197, n1199, n1201, n1203, n1205, n1207, n1209, n1211,
         n1213, n1215, n1217, n1219, n1221, n1223, n1225, n1227, n1229, n1231,
         n1233, n1235, n1237, n1239, n1241, n1243, n1245, n1247, n1249, n1251,
         n1253, n1255, n1257, n1259, n1261, n1263, n1265, n1267, n1269, n1271,
         n1273, n1275, n1277, n1279, n1281, n1283, n1285, n1287, n1289, n1291,
         n1293, n1295, n1297, n1299, n1301, n1303, n1305, n1307, n1309, n1311,
         n1313, n1315, n1317, n1319, n1321, n1323, n1325, n1327, n1329, n1331,
         n1333, n1335, n1337, n1339, n1341, n1343, n1345, n1347, n1349, n1351,
         n1353, n1355, n1357, n1359, n1361, n1363, n1365, n1367, n1369, n1371,
         n1373, n1375, n1377, n1379, n1381, n1383, n1385, n1387, n1389, n1391,
         n1393, n1395, n1397, n1399, n1401, n1403, n1405, n1407, n1409, n1411,
         n1413, n1415, n1417, n1419, n1421, n1423, n1425, n1427, n1429, n1431,
         n1433, n1435, n1437, n1439, n1441, n1443, n1445, n1447, n1449, n1451,
         n1453, n1455, n1457, n1459, n1461, n1463, n1465, n1467, n1469, n1471,
         n1473, n1475, n1477, n1479, n1481, n1483, n1485, n1487, n1489, n1491,
         n1493, n1495, n1497, n1499, n1501, n1503, n1505, n1507, n1509, n1511,
         n1513, n1515, n1517, n1519, n1521, n1523, n1525, n1527, n1529, n1531,
         n1533, n1535, n1537, n1539, n1541, n1543, n1545, n1547, n1549, n1551,
         n1553, n1555, n1557, n1559, n1561, n1563, n1565, n1567, n1569, n1571,
         n1573, n1575, n1577, n1579, n1581, n1583, n1585, n1587, n1589, n1591,
         n1593, n1595, n1597, n1599, n1601, n1603, n1605, n1607, n1609, n1611,
         n1613, n1615, n1617, n1619, n1621, n1623, n1625, n1627, n1629, n1631,
         n1633, n1635, n1637, n1639, n1641, n1643, n1645, n1647, n1649, n1651,
         n1653, n1655, n1657, n1659, n1661, n1663, n1665, n1667, n1669, n1671,
         n1673, n1675, n1677, n1679, n1681, n1683, n1685, n1687, n1689, n1691,
         n1693, n1695, n1697, n1699, n1701, n1703, n1705, n1707, n1709, n1711,
         n1713, n1715, n1717, n1719, n1721, n1723, n1725, n1727, n1729, n1731,
         n1733, n1735, n1737, n1739, n1741, n1743, n1745, n1747, n1749, n1751,
         n1753, n1755, n1757, n1759, n1761, n1763, n1765, n1767, n1769, n1771,
         n1773, n1775, n1777, n1779, n1781, n1783, n1785, n1787, n1789, n1791,
         n1793, n1795, n1797, n1799, n1801, n1803, n1805, n1807, n1809, n1811,
         n1813, n1815, n1817, n1819, n1821, n1823, n1825, n1827, n1829, n1831,
         n1833, n1835, n1837, n1839, n1841, n1843, n1845, n1847, n1849, n1851,
         n1853, n1855, n1857, n1859, n1861, n1863, n1865, n1867, n1869, n1871,
         n1873, n1875, n1877, n1879, n1881, n1883, n1885, n1887, n1889, n1891,
         n1893, n1895, n1897, n1899, n1901, n1903, n1905, n1907, n1909, n1911,
         n1913, n1915, n1917, n1919, n1921, n1923, n1925, n1927, n1929, n1931,
         n1933, n1935, n1937, n1939, n1941, n1943, n1945, n1947, n1949, n1951,
         n1953, n1955, n1957, n1959, n1961, n1963, n1965, n1967, n1969, n1971,
         n1973, n1975, n1977, n1979, n1981, n1983, n1985, n1987, n1989, n1991,
         n1993, n1995, n1997, n1999, n2001, n2003, n2005, n2007, n2009, n2011,
         n2013, n2015, n2017, n2019, n2021, n2023, n2025, n2027, n2029, n2031,
         n2033, n2035, n2037, n2039, n2041, n2043, n2045, n2047, n2049, n2051,
         n2053, n2055, n2057, n2059, n2061, n2063, n2065, n2067, n2069, n2071,
         n2073, n2075, n2077, n2079, n2081, n2083, n2085, n2087, n2089, n2091,
         n2093, n2095, n2097, n2099, n2101, n2103, n2105, n2107, n2109, n2111,
         n2113, n2115, n2117, n2119, n2121, n2123, n2125, n2127, n2129, n2131,
         n2133, n2135, n2137, n2139, n2141, n2143, n2145, n2147, n2149, n2151,
         n2153, n2155, n2157, n2159, n2161, n2163, n2165, n2167, n2169, n2171,
         n2173, n2175, n2177, n2179, n2181, n2183, n2185, n2187, n2189, n2191,
         n2193, n2195, n2197, n2199, n2201, n2203, n2205, n2207, n2209, n2211,
         n2213, n2215, n2217, n2219, n2221, n2223, n2225, n2227, n2229, n2231,
         n2233, n2235, n2237, n2239, n2241, n2243, n2245, n2247, n2249, n2251,
         n2253, n2255, n2257, n2259, n2261, n2263, n2265, n2267, n2269, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296;
  wire   [3:0] DecodedL1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  Dec4_16_0 U1 ( .Hot({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, DecodedL1}), .Sel(
        {\*Logic0* , \*Logic0* , Address[1], n2274}) );
  Dec4_16_68 \DL2[0].U2  ( .Hot({\DL2[0].tempL2[15] , \DL2[0].tempL2[14] , 
        \DL2[0].tempL2[13] , \DL2[0].tempL2[12] , \DL2[0].tempL2[11] , 
        \DL2[0].tempL2[10] , \DL2[0].tempL2[9] , \DL2[0].tempL2[8] , 
        \DL2[0].tempL2[7] , \DL2[0].tempL2[6] , \DL2[0].tempL2[5] , 
        \DL2[0].tempL2[4] , \DL2[0].tempL2[3] , \DL2[0].tempL2[2] , 
        \DL2[0].tempL2[1] , \DL2[0].tempL2[0] }), .Sel({n2278, n2277, n2276, 
        n2275}) );
  Dec4_16_67 \DL2[1].U2  ( .Hot({\DL2[1].tempL2[15] , \DL2[1].tempL2[14] , 
        \DL2[1].tempL2[13] , \DL2[1].tempL2[12] , \DL2[1].tempL2[11] , 
        \DL2[1].tempL2[10] , \DL2[1].tempL2[9] , \DL2[1].tempL2[8] , 
        \DL2[1].tempL2[7] , \DL2[1].tempL2[6] , \DL2[1].tempL2[5] , 
        \DL2[1].tempL2[4] , \DL2[1].tempL2[3] , \DL2[1].tempL2[2] , 
        \DL2[1].tempL2[1] , \DL2[1].tempL2[0] }), .Sel({n2278, n2277, n2276, 
        n2275}) );
  Dec4_16_66 \DL2[2].U2  ( .Hot({\DL2[2].tempL2[15] , \DL2[2].tempL2[14] , 
        \DL2[2].tempL2[13] , \DL2[2].tempL2[12] , \DL2[2].tempL2[11] , 
        \DL2[2].tempL2[10] , \DL2[2].tempL2[9] , \DL2[2].tempL2[8] , 
        \DL2[2].tempL2[7] , \DL2[2].tempL2[6] , \DL2[2].tempL2[5] , 
        \DL2[2].tempL2[4] , \DL2[2].tempL2[3] , \DL2[2].tempL2[2] , 
        \DL2[2].tempL2[1] , \DL2[2].tempL2[0] }), .Sel({n2278, n2277, n2276, 
        n2275}) );
  Dec4_16_65 \DL2[3].U2  ( .Hot({\DL2[3].tempL2[15] , \DL2[3].tempL2[14] , 
        \DL2[3].tempL2[13] , \DL2[3].tempL2[12] , \DL2[3].tempL2[11] , 
        \DL2[3].tempL2[10] , \DL2[3].tempL2[9] , \DL2[3].tempL2[8] , 
        \DL2[3].tempL2[7] , \DL2[3].tempL2[6] , \DL2[3].tempL2[5] , 
        \DL2[3].tempL2[4] , \DL2[3].tempL2[3] , \DL2[3].tempL2[2] , 
        \DL2[3].tempL2[1] , \DL2[3].tempL2[0] }), .Sel({n2278, n2277, n2276, 
        n2275}) );
  Dec4_16_64 \DL3[0].U3  ( .Hot({\DL3[0].tempL3[15] , \DL3[0].tempL3[14] , 
        \DL3[0].tempL3[13] , \DL3[0].tempL3[12] , \DL3[0].tempL3[11] , 
        \DL3[0].tempL3[10] , \DL3[0].tempL3[9] , \DL3[0].tempL3[8] , 
        \DL3[0].tempL3[7] , \DL3[0].tempL3[6] , \DL3[0].tempL3[5] , 
        \DL3[0].tempL3[4] , \DL3[0].tempL3[3] , \DL3[0].tempL3[2] , 
        \DL3[0].tempL3[1] , \DL3[0].tempL3[0] }), .Sel({n2294, n2289, n2273, 
        n2281}) );
  Dec4_16_63 \DL3[1].U3  ( .Hot({\DL3[1].tempL3[15] , \DL3[1].tempL3[14] , 
        \DL3[1].tempL3[13] , \DL3[1].tempL3[12] , \DL3[1].tempL3[11] , 
        \DL3[1].tempL3[10] , \DL3[1].tempL3[9] , \DL3[1].tempL3[8] , 
        \DL3[1].tempL3[7] , \DL3[1].tempL3[6] , \DL3[1].tempL3[5] , 
        \DL3[1].tempL3[4] , \DL3[1].tempL3[3] , \DL3[1].tempL3[2] , 
        \DL3[1].tempL3[1] , \DL3[1].tempL3[0] }), .Sel({n2295, n2287, n2285, 
        n2272}) );
  Dec4_16_62 \DL3[2].U3  ( .Hot({\DL3[2].tempL3[15] , \DL3[2].tempL3[14] , 
        \DL3[2].tempL3[13] , \DL3[2].tempL3[12] , \DL3[2].tempL3[11] , 
        \DL3[2].tempL3[10] , \DL3[2].tempL3[9] , \DL3[2].tempL3[8] , 
        \DL3[2].tempL3[7] , \DL3[2].tempL3[6] , \DL3[2].tempL3[5] , 
        \DL3[2].tempL3[4] , \DL3[2].tempL3[3] , \DL3[2].tempL3[2] , 
        \DL3[2].tempL3[1] , \DL3[2].tempL3[0] }), .Sel({n2295, n2290, 
        Address[7], n2280}) );
  Dec4_16_61 \DL3[3].U3  ( .Hot({\DL3[3].tempL3[15] , \DL3[3].tempL3[14] , 
        \DL3[3].tempL3[13] , \DL3[3].tempL3[12] , \DL3[3].tempL3[11] , 
        \DL3[3].tempL3[10] , \DL3[3].tempL3[9] , \DL3[3].tempL3[8] , 
        \DL3[3].tempL3[7] , \DL3[3].tempL3[6] , \DL3[3].tempL3[5] , 
        \DL3[3].tempL3[4] , \DL3[3].tempL3[3] , \DL3[3].tempL3[2] , 
        \DL3[3].tempL3[1] , \DL3[3].tempL3[0] }), .Sel({n2293, n2287, n2285, 
        n2280}) );
  Dec4_16_60 \DL3[4].U3  ( .Hot({\DL3[4].tempL3[15] , \DL3[4].tempL3[14] , 
        \DL3[4].tempL3[13] , \DL3[4].tempL3[12] , \DL3[4].tempL3[11] , 
        \DL3[4].tempL3[10] , \DL3[4].tempL3[9] , \DL3[4].tempL3[8] , 
        \DL3[4].tempL3[7] , \DL3[4].tempL3[6] , \DL3[4].tempL3[5] , 
        \DL3[4].tempL3[4] , \DL3[4].tempL3[3] , \DL3[4].tempL3[2] , 
        \DL3[4].tempL3[1] , \DL3[4].tempL3[0] }), .Sel({n2294, n2287, n2273, 
        n2272}) );
  Dec4_16_59 \DL3[5].U3  ( .Hot({\DL3[5].tempL3[15] , \DL3[5].tempL3[14] , 
        \DL3[5].tempL3[13] , \DL3[5].tempL3[12] , \DL3[5].tempL3[11] , 
        \DL3[5].tempL3[10] , \DL3[5].tempL3[9] , \DL3[5].tempL3[8] , 
        \DL3[5].tempL3[7] , \DL3[5].tempL3[6] , \DL3[5].tempL3[5] , 
        \DL3[5].tempL3[4] , \DL3[5].tempL3[3] , \DL3[5].tempL3[2] , 
        \DL3[5].tempL3[1] , \DL3[5].tempL3[0] }), .Sel({n2295, n2287, n2273, 
        n2282}) );
  Dec4_16_58 \DL3[6].U3  ( .Hot({\DL3[6].tempL3[15] , \DL3[6].tempL3[14] , 
        \DL3[6].tempL3[13] , \DL3[6].tempL3[12] , \DL3[6].tempL3[11] , 
        \DL3[6].tempL3[10] , \DL3[6].tempL3[9] , \DL3[6].tempL3[8] , 
        \DL3[6].tempL3[7] , \DL3[6].tempL3[6] , \DL3[6].tempL3[5] , 
        \DL3[6].tempL3[4] , \DL3[6].tempL3[3] , \DL3[6].tempL3[2] , 
        \DL3[6].tempL3[1] , \DL3[6].tempL3[0] }), .Sel({n2293, n2287, n2273, 
        n2272}) );
  Dec4_16_57 \DL3[7].U3  ( .Hot({\DL3[7].tempL3[15] , \DL3[7].tempL3[14] , 
        \DL3[7].tempL3[13] , \DL3[7].tempL3[12] , \DL3[7].tempL3[11] , 
        \DL3[7].tempL3[10] , \DL3[7].tempL3[9] , \DL3[7].tempL3[8] , 
        \DL3[7].tempL3[7] , \DL3[7].tempL3[6] , \DL3[7].tempL3[5] , 
        \DL3[7].tempL3[4] , \DL3[7].tempL3[3] , \DL3[7].tempL3[2] , 
        \DL3[7].tempL3[1] , \DL3[7].tempL3[0] }), .Sel({n2295, n2287, n2285, 
        n2271}) );
  Dec4_16_56 \DL3[8].U3  ( .Hot({\DL3[8].tempL3[15] , \DL3[8].tempL3[14] , 
        \DL3[8].tempL3[13] , \DL3[8].tempL3[12] , \DL3[8].tempL3[11] , 
        \DL3[8].tempL3[10] , \DL3[8].tempL3[9] , \DL3[8].tempL3[8] , 
        \DL3[8].tempL3[7] , \DL3[8].tempL3[6] , \DL3[8].tempL3[5] , 
        \DL3[8].tempL3[4] , \DL3[8].tempL3[3] , \DL3[8].tempL3[2] , 
        \DL3[8].tempL3[1] , \DL3[8].tempL3[0] }), .Sel({n2292, n2290, n2285, 
        n2272}) );
  Dec4_16_55 \DL3[9].U3  ( .Hot({\DL3[9].tempL3[15] , \DL3[9].tempL3[14] , 
        \DL3[9].tempL3[13] , \DL3[9].tempL3[12] , \DL3[9].tempL3[11] , 
        \DL3[9].tempL3[10] , \DL3[9].tempL3[9] , \DL3[9].tempL3[8] , 
        \DL3[9].tempL3[7] , \DL3[9].tempL3[6] , \DL3[9].tempL3[5] , 
        \DL3[9].tempL3[4] , \DL3[9].tempL3[3] , \DL3[9].tempL3[2] , 
        \DL3[9].tempL3[1] , \DL3[9].tempL3[0] }), .Sel({n2293, n2290, n2285, 
        n2281}) );
  Dec4_16_54 \DL3[10].U3  ( .Hot({\DL3[10].tempL3[15] , \DL3[10].tempL3[14] , 
        \DL3[10].tempL3[13] , \DL3[10].tempL3[12] , \DL3[10].tempL3[11] , 
        \DL3[10].tempL3[10] , \DL3[10].tempL3[9] , \DL3[10].tempL3[8] , 
        \DL3[10].tempL3[7] , \DL3[10].tempL3[6] , \DL3[10].tempL3[5] , 
        \DL3[10].tempL3[4] , \DL3[10].tempL3[3] , \DL3[10].tempL3[2] , 
        \DL3[10].tempL3[1] , \DL3[10].tempL3[0] }), .Sel({n2294, n2289, n2273, 
        n2281}) );
  Dec4_16_53 \DL3[11].U3  ( .Hot({\DL3[11].tempL3[15] , \DL3[11].tempL3[14] , 
        \DL3[11].tempL3[13] , \DL3[11].tempL3[12] , \DL3[11].tempL3[11] , 
        \DL3[11].tempL3[10] , \DL3[11].tempL3[9] , \DL3[11].tempL3[8] , 
        \DL3[11].tempL3[7] , \DL3[11].tempL3[6] , \DL3[11].tempL3[5] , 
        \DL3[11].tempL3[4] , \DL3[11].tempL3[3] , \DL3[11].tempL3[2] , 
        \DL3[11].tempL3[1] , \DL3[11].tempL3[0] }), .Sel({n2295, n2288, n2285, 
        n2272}) );
  Dec4_16_52 \DL3[12].U3  ( .Hot({\DL3[12].tempL3[15] , \DL3[12].tempL3[14] , 
        \DL3[12].tempL3[13] , \DL3[12].tempL3[12] , \DL3[12].tempL3[11] , 
        \DL3[12].tempL3[10] , \DL3[12].tempL3[9] , \DL3[12].tempL3[8] , 
        \DL3[12].tempL3[7] , \DL3[12].tempL3[6] , \DL3[12].tempL3[5] , 
        \DL3[12].tempL3[4] , \DL3[12].tempL3[3] , \DL3[12].tempL3[2] , 
        \DL3[12].tempL3[1] , \DL3[12].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2271}) );
  Dec4_16_51 \DL3[13].U3  ( .Hot({\DL3[13].tempL3[15] , \DL3[13].tempL3[14] , 
        \DL3[13].tempL3[13] , \DL3[13].tempL3[12] , \DL3[13].tempL3[11] , 
        \DL3[13].tempL3[10] , \DL3[13].tempL3[9] , \DL3[13].tempL3[8] , 
        \DL3[13].tempL3[7] , \DL3[13].tempL3[6] , \DL3[13].tempL3[5] , 
        \DL3[13].tempL3[4] , \DL3[13].tempL3[3] , \DL3[13].tempL3[2] , 
        \DL3[13].tempL3[1] , \DL3[13].tempL3[0] }), .Sel({n2292, n2287, n2284, 
        n2282}) );
  Dec4_16_50 \DL3[14].U3  ( .Hot({\DL3[14].tempL3[15] , \DL3[14].tempL3[14] , 
        \DL3[14].tempL3[13] , \DL3[14].tempL3[12] , \DL3[14].tempL3[11] , 
        \DL3[14].tempL3[10] , \DL3[14].tempL3[9] , \DL3[14].tempL3[8] , 
        \DL3[14].tempL3[7] , \DL3[14].tempL3[6] , \DL3[14].tempL3[5] , 
        \DL3[14].tempL3[4] , \DL3[14].tempL3[3] , \DL3[14].tempL3[2] , 
        \DL3[14].tempL3[1] , \DL3[14].tempL3[0] }), .Sel({n2292, n2287, n2284, 
        n2280}) );
  Dec4_16_49 \DL3[15].U3  ( .Hot({\DL3[15].tempL3[15] , \DL3[15].tempL3[14] , 
        \DL3[15].tempL3[13] , \DL3[15].tempL3[12] , \DL3[15].tempL3[11] , 
        \DL3[15].tempL3[10] , \DL3[15].tempL3[9] , \DL3[15].tempL3[8] , 
        \DL3[15].tempL3[7] , \DL3[15].tempL3[6] , \DL3[15].tempL3[5] , 
        \DL3[15].tempL3[4] , \DL3[15].tempL3[3] , \DL3[15].tempL3[2] , 
        \DL3[15].tempL3[1] , \DL3[15].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2282}) );
  Dec4_16_48 \DL3[16].U3  ( .Hot({\DL3[16].tempL3[15] , \DL3[16].tempL3[14] , 
        \DL3[16].tempL3[13] , \DL3[16].tempL3[12] , \DL3[16].tempL3[11] , 
        \DL3[16].tempL3[10] , \DL3[16].tempL3[9] , \DL3[16].tempL3[8] , 
        \DL3[16].tempL3[7] , \DL3[16].tempL3[6] , \DL3[16].tempL3[5] , 
        \DL3[16].tempL3[4] , \DL3[16].tempL3[3] , \DL3[16].tempL3[2] , 
        \DL3[16].tempL3[1] , \DL3[16].tempL3[0] }), .Sel({n2292, n2287, 
        Address[7], n2272}) );
  Dec4_16_47 \DL3[17].U3  ( .Hot({\DL3[17].tempL3[15] , \DL3[17].tempL3[14] , 
        \DL3[17].tempL3[13] , \DL3[17].tempL3[12] , \DL3[17].tempL3[11] , 
        \DL3[17].tempL3[10] , \DL3[17].tempL3[9] , \DL3[17].tempL3[8] , 
        \DL3[17].tempL3[7] , \DL3[17].tempL3[6] , \DL3[17].tempL3[5] , 
        \DL3[17].tempL3[4] , \DL3[17].tempL3[3] , \DL3[17].tempL3[2] , 
        \DL3[17].tempL3[1] , \DL3[17].tempL3[0] }), .Sel({n2292, n2287, n2273, 
        n2282}) );
  Dec4_16_46 \DL3[18].U3  ( .Hot({\DL3[18].tempL3[15] , \DL3[18].tempL3[14] , 
        \DL3[18].tempL3[13] , \DL3[18].tempL3[12] , \DL3[18].tempL3[11] , 
        \DL3[18].tempL3[10] , \DL3[18].tempL3[9] , \DL3[18].tempL3[8] , 
        \DL3[18].tempL3[7] , \DL3[18].tempL3[6] , \DL3[18].tempL3[5] , 
        \DL3[18].tempL3[4] , \DL3[18].tempL3[3] , \DL3[18].tempL3[2] , 
        \DL3[18].tempL3[1] , \DL3[18].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2280}) );
  Dec4_16_45 \DL3[19].U3  ( .Hot({\DL3[19].tempL3[15] , \DL3[19].tempL3[14] , 
        \DL3[19].tempL3[13] , \DL3[19].tempL3[12] , \DL3[19].tempL3[11] , 
        \DL3[19].tempL3[10] , \DL3[19].tempL3[9] , \DL3[19].tempL3[8] , 
        \DL3[19].tempL3[7] , \DL3[19].tempL3[6] , \DL3[19].tempL3[5] , 
        \DL3[19].tempL3[4] , \DL3[19].tempL3[3] , \DL3[19].tempL3[2] , 
        \DL3[19].tempL3[1] , \DL3[19].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2271}) );
  Dec4_16_44 \DL3[20].U3  ( .Hot({\DL3[20].tempL3[15] , \DL3[20].tempL3[14] , 
        \DL3[20].tempL3[13] , \DL3[20].tempL3[12] , \DL3[20].tempL3[11] , 
        \DL3[20].tempL3[10] , \DL3[20].tempL3[9] , \DL3[20].tempL3[8] , 
        \DL3[20].tempL3[7] , \DL3[20].tempL3[6] , \DL3[20].tempL3[5] , 
        \DL3[20].tempL3[4] , \DL3[20].tempL3[3] , \DL3[20].tempL3[2] , 
        \DL3[20].tempL3[1] , \DL3[20].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2271}) );
  Dec4_16_43 \DL3[21].U3  ( .Hot({\DL3[21].tempL3[15] , \DL3[21].tempL3[14] , 
        \DL3[21].tempL3[13] , \DL3[21].tempL3[12] , \DL3[21].tempL3[11] , 
        \DL3[21].tempL3[10] , \DL3[21].tempL3[9] , \DL3[21].tempL3[8] , 
        \DL3[21].tempL3[7] , \DL3[21].tempL3[6] , \DL3[21].tempL3[5] , 
        \DL3[21].tempL3[4] , \DL3[21].tempL3[3] , \DL3[21].tempL3[2] , 
        \DL3[21].tempL3[1] , \DL3[21].tempL3[0] }), .Sel({n2292, n2287, n2285, 
        n2282}) );
  Dec4_16_42 \DL3[22].U3  ( .Hot({\DL3[22].tempL3[15] , \DL3[22].tempL3[14] , 
        \DL3[22].tempL3[13] , \DL3[22].tempL3[12] , \DL3[22].tempL3[11] , 
        \DL3[22].tempL3[10] , \DL3[22].tempL3[9] , \DL3[22].tempL3[8] , 
        \DL3[22].tempL3[7] , \DL3[22].tempL3[6] , \DL3[22].tempL3[5] , 
        \DL3[22].tempL3[4] , \DL3[22].tempL3[3] , \DL3[22].tempL3[2] , 
        \DL3[22].tempL3[1] , \DL3[22].tempL3[0] }), .Sel({n2292, n2287, 
        Address[7], n2281}) );
  Dec4_16_41 \DL3[23].U3  ( .Hot({\DL3[23].tempL3[15] , \DL3[23].tempL3[14] , 
        \DL3[23].tempL3[13] , \DL3[23].tempL3[12] , \DL3[23].tempL3[11] , 
        \DL3[23].tempL3[10] , \DL3[23].tempL3[9] , \DL3[23].tempL3[8] , 
        \DL3[23].tempL3[7] , \DL3[23].tempL3[6] , \DL3[23].tempL3[5] , 
        \DL3[23].tempL3[4] , \DL3[23].tempL3[3] , \DL3[23].tempL3[2] , 
        \DL3[23].tempL3[1] , \DL3[23].tempL3[0] }), .Sel({n2292, n2287, n2284, 
        n2280}) );
  Dec4_16_40 \DL3[24].U3  ( .Hot({\DL3[24].tempL3[15] , \DL3[24].tempL3[14] , 
        \DL3[24].tempL3[13] , \DL3[24].tempL3[12] , \DL3[24].tempL3[11] , 
        \DL3[24].tempL3[10] , \DL3[24].tempL3[9] , \DL3[24].tempL3[8] , 
        \DL3[24].tempL3[7] , \DL3[24].tempL3[6] , \DL3[24].tempL3[5] , 
        \DL3[24].tempL3[4] , \DL3[24].tempL3[3] , \DL3[24].tempL3[2] , 
        \DL3[24].tempL3[1] , \DL3[24].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2280}) );
  Dec4_16_39 \DL3[25].U3  ( .Hot({\DL3[25].tempL3[15] , \DL3[25].tempL3[14] , 
        \DL3[25].tempL3[13] , \DL3[25].tempL3[12] , \DL3[25].tempL3[11] , 
        \DL3[25].tempL3[10] , \DL3[25].tempL3[9] , \DL3[25].tempL3[8] , 
        \DL3[25].tempL3[7] , \DL3[25].tempL3[6] , \DL3[25].tempL3[5] , 
        \DL3[25].tempL3[4] , \DL3[25].tempL3[3] , \DL3[25].tempL3[2] , 
        \DL3[25].tempL3[1] , \DL3[25].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2271}) );
  Dec4_16_38 \DL3[26].U3  ( .Hot({\DL3[26].tempL3[15] , \DL3[26].tempL3[14] , 
        \DL3[26].tempL3[13] , \DL3[26].tempL3[12] , \DL3[26].tempL3[11] , 
        \DL3[26].tempL3[10] , \DL3[26].tempL3[9] , \DL3[26].tempL3[8] , 
        \DL3[26].tempL3[7] , \DL3[26].tempL3[6] , \DL3[26].tempL3[5] , 
        \DL3[26].tempL3[4] , \DL3[26].tempL3[3] , \DL3[26].tempL3[2] , 
        \DL3[26].tempL3[1] , \DL3[26].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2281}) );
  Dec4_16_37 \DL3[27].U3  ( .Hot({\DL3[27].tempL3[15] , \DL3[27].tempL3[14] , 
        \DL3[27].tempL3[13] , \DL3[27].tempL3[12] , \DL3[27].tempL3[11] , 
        \DL3[27].tempL3[10] , \DL3[27].tempL3[9] , \DL3[27].tempL3[8] , 
        \DL3[27].tempL3[7] , \DL3[27].tempL3[6] , \DL3[27].tempL3[5] , 
        \DL3[27].tempL3[4] , \DL3[27].tempL3[3] , \DL3[27].tempL3[2] , 
        \DL3[27].tempL3[1] , \DL3[27].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2272}) );
  Dec4_16_36 \DL3[28].U3  ( .Hot({\DL3[28].tempL3[15] , \DL3[28].tempL3[14] , 
        \DL3[28].tempL3[13] , \DL3[28].tempL3[12] , \DL3[28].tempL3[11] , 
        \DL3[28].tempL3[10] , \DL3[28].tempL3[9] , \DL3[28].tempL3[8] , 
        \DL3[28].tempL3[7] , \DL3[28].tempL3[6] , \DL3[28].tempL3[5] , 
        \DL3[28].tempL3[4] , \DL3[28].tempL3[3] , \DL3[28].tempL3[2] , 
        \DL3[28].tempL3[1] , \DL3[28].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2271}) );
  Dec4_16_35 \DL3[29].U3  ( .Hot({\DL3[29].tempL3[15] , \DL3[29].tempL3[14] , 
        \DL3[29].tempL3[13] , \DL3[29].tempL3[12] , \DL3[29].tempL3[11] , 
        \DL3[29].tempL3[10] , \DL3[29].tempL3[9] , \DL3[29].tempL3[8] , 
        \DL3[29].tempL3[7] , \DL3[29].tempL3[6] , \DL3[29].tempL3[5] , 
        \DL3[29].tempL3[4] , \DL3[29].tempL3[3] , \DL3[29].tempL3[2] , 
        \DL3[29].tempL3[1] , \DL3[29].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2281}) );
  Dec4_16_34 \DL3[30].U3  ( .Hot({\DL3[30].tempL3[15] , \DL3[30].tempL3[14] , 
        \DL3[30].tempL3[13] , \DL3[30].tempL3[12] , \DL3[30].tempL3[11] , 
        \DL3[30].tempL3[10] , \DL3[30].tempL3[9] , \DL3[30].tempL3[8] , 
        \DL3[30].tempL3[7] , \DL3[30].tempL3[6] , \DL3[30].tempL3[5] , 
        \DL3[30].tempL3[4] , \DL3[30].tempL3[3] , \DL3[30].tempL3[2] , 
        \DL3[30].tempL3[1] , \DL3[30].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2280}) );
  Dec4_16_33 \DL3[31].U3  ( .Hot({\DL3[31].tempL3[15] , \DL3[31].tempL3[14] , 
        \DL3[31].tempL3[13] , \DL3[31].tempL3[12] , \DL3[31].tempL3[11] , 
        \DL3[31].tempL3[10] , \DL3[31].tempL3[9] , \DL3[31].tempL3[8] , 
        \DL3[31].tempL3[7] , \DL3[31].tempL3[6] , \DL3[31].tempL3[5] , 
        \DL3[31].tempL3[4] , \DL3[31].tempL3[3] , \DL3[31].tempL3[2] , 
        \DL3[31].tempL3[1] , \DL3[31].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2272}) );
  Dec4_16_32 \DL3[32].U3  ( .Hot({\DL3[32].tempL3[15] , \DL3[32].tempL3[14] , 
        \DL3[32].tempL3[13] , \DL3[32].tempL3[12] , \DL3[32].tempL3[11] , 
        \DL3[32].tempL3[10] , \DL3[32].tempL3[9] , \DL3[32].tempL3[8] , 
        \DL3[32].tempL3[7] , \DL3[32].tempL3[6] , \DL3[32].tempL3[5] , 
        \DL3[32].tempL3[4] , \DL3[32].tempL3[3] , \DL3[32].tempL3[2] , 
        \DL3[32].tempL3[1] , \DL3[32].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2280}) );
  Dec4_16_31 \DL3[33].U3  ( .Hot({\DL3[33].tempL3[15] , \DL3[33].tempL3[14] , 
        \DL3[33].tempL3[13] , \DL3[33].tempL3[12] , \DL3[33].tempL3[11] , 
        \DL3[33].tempL3[10] , \DL3[33].tempL3[9] , \DL3[33].tempL3[8] , 
        \DL3[33].tempL3[7] , \DL3[33].tempL3[6] , \DL3[33].tempL3[5] , 
        \DL3[33].tempL3[4] , \DL3[33].tempL3[3] , \DL3[33].tempL3[2] , 
        \DL3[33].tempL3[1] , \DL3[33].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2280}) );
  Dec4_16_30 \DL3[34].U3  ( .Hot({\DL3[34].tempL3[15] , \DL3[34].tempL3[14] , 
        \DL3[34].tempL3[13] , \DL3[34].tempL3[12] , \DL3[34].tempL3[11] , 
        \DL3[34].tempL3[10] , \DL3[34].tempL3[9] , \DL3[34].tempL3[8] , 
        \DL3[34].tempL3[7] , \DL3[34].tempL3[6] , \DL3[34].tempL3[5] , 
        \DL3[34].tempL3[4] , \DL3[34].tempL3[3] , \DL3[34].tempL3[2] , 
        \DL3[34].tempL3[1] , \DL3[34].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2280}) );
  Dec4_16_29 \DL3[35].U3  ( .Hot({\DL3[35].tempL3[15] , \DL3[35].tempL3[14] , 
        \DL3[35].tempL3[13] , \DL3[35].tempL3[12] , \DL3[35].tempL3[11] , 
        \DL3[35].tempL3[10] , \DL3[35].tempL3[9] , \DL3[35].tempL3[8] , 
        \DL3[35].tempL3[7] , \DL3[35].tempL3[6] , \DL3[35].tempL3[5] , 
        \DL3[35].tempL3[4] , \DL3[35].tempL3[3] , \DL3[35].tempL3[2] , 
        \DL3[35].tempL3[1] , \DL3[35].tempL3[0] }), .Sel({n2293, n2288, n2284, 
        n2271}) );
  Dec4_16_28 \DL3[36].U3  ( .Hot({\DL3[36].tempL3[15] , \DL3[36].tempL3[14] , 
        \DL3[36].tempL3[13] , \DL3[36].tempL3[12] , \DL3[36].tempL3[11] , 
        \DL3[36].tempL3[10] , \DL3[36].tempL3[9] , \DL3[36].tempL3[8] , 
        \DL3[36].tempL3[7] , \DL3[36].tempL3[6] , \DL3[36].tempL3[5] , 
        \DL3[36].tempL3[4] , \DL3[36].tempL3[3] , \DL3[36].tempL3[2] , 
        \DL3[36].tempL3[1] , \DL3[36].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2281}) );
  Dec4_16_27 \DL3[37].U3  ( .Hot({\DL3[37].tempL3[15] , \DL3[37].tempL3[14] , 
        \DL3[37].tempL3[13] , \DL3[37].tempL3[12] , \DL3[37].tempL3[11] , 
        \DL3[37].tempL3[10] , \DL3[37].tempL3[9] , \DL3[37].tempL3[8] , 
        \DL3[37].tempL3[7] , \DL3[37].tempL3[6] , \DL3[37].tempL3[5] , 
        \DL3[37].tempL3[4] , \DL3[37].tempL3[3] , \DL3[37].tempL3[2] , 
        \DL3[37].tempL3[1] , \DL3[37].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2271}) );
  Dec4_16_26 \DL3[38].U3  ( .Hot({\DL3[38].tempL3[15] , \DL3[38].tempL3[14] , 
        \DL3[38].tempL3[13] , \DL3[38].tempL3[12] , \DL3[38].tempL3[11] , 
        \DL3[38].tempL3[10] , \DL3[38].tempL3[9] , \DL3[38].tempL3[8] , 
        \DL3[38].tempL3[7] , \DL3[38].tempL3[6] , \DL3[38].tempL3[5] , 
        \DL3[38].tempL3[4] , \DL3[38].tempL3[3] , \DL3[38].tempL3[2] , 
        \DL3[38].tempL3[1] , \DL3[38].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2272}) );
  Dec4_16_25 \DL3[39].U3  ( .Hot({\DL3[39].tempL3[15] , \DL3[39].tempL3[14] , 
        \DL3[39].tempL3[13] , \DL3[39].tempL3[12] , \DL3[39].tempL3[11] , 
        \DL3[39].tempL3[10] , \DL3[39].tempL3[9] , \DL3[39].tempL3[8] , 
        \DL3[39].tempL3[7] , \DL3[39].tempL3[6] , \DL3[39].tempL3[5] , 
        \DL3[39].tempL3[4] , \DL3[39].tempL3[3] , \DL3[39].tempL3[2] , 
        \DL3[39].tempL3[1] , \DL3[39].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2281}) );
  Dec4_16_24 \DL3[40].U3  ( .Hot({\DL3[40].tempL3[15] , \DL3[40].tempL3[14] , 
        \DL3[40].tempL3[13] , \DL3[40].tempL3[12] , \DL3[40].tempL3[11] , 
        \DL3[40].tempL3[10] , \DL3[40].tempL3[9] , \DL3[40].tempL3[8] , 
        \DL3[40].tempL3[7] , \DL3[40].tempL3[6] , \DL3[40].tempL3[5] , 
        \DL3[40].tempL3[4] , \DL3[40].tempL3[3] , \DL3[40].tempL3[2] , 
        \DL3[40].tempL3[1] , \DL3[40].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2271}) );
  Dec4_16_23 \DL3[41].U3  ( .Hot({\DL3[41].tempL3[15] , \DL3[41].tempL3[14] , 
        \DL3[41].tempL3[13] , \DL3[41].tempL3[12] , \DL3[41].tempL3[11] , 
        \DL3[41].tempL3[10] , \DL3[41].tempL3[9] , \DL3[41].tempL3[8] , 
        \DL3[41].tempL3[7] , \DL3[41].tempL3[6] , \DL3[41].tempL3[5] , 
        \DL3[41].tempL3[4] , \DL3[41].tempL3[3] , \DL3[41].tempL3[2] , 
        \DL3[41].tempL3[1] , \DL3[41].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2271}) );
  Dec4_16_22 \DL3[42].U3  ( .Hot({\DL3[42].tempL3[15] , \DL3[42].tempL3[14] , 
        \DL3[42].tempL3[13] , \DL3[42].tempL3[12] , \DL3[42].tempL3[11] , 
        \DL3[42].tempL3[10] , \DL3[42].tempL3[9] , \DL3[42].tempL3[8] , 
        \DL3[42].tempL3[7] , \DL3[42].tempL3[6] , \DL3[42].tempL3[5] , 
        \DL3[42].tempL3[4] , \DL3[42].tempL3[3] , \DL3[42].tempL3[2] , 
        \DL3[42].tempL3[1] , \DL3[42].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2271}) );
  Dec4_16_21 \DL3[43].U3  ( .Hot({\DL3[43].tempL3[15] , \DL3[43].tempL3[14] , 
        \DL3[43].tempL3[13] , \DL3[43].tempL3[12] , \DL3[43].tempL3[11] , 
        \DL3[43].tempL3[10] , \DL3[43].tempL3[9] , \DL3[43].tempL3[8] , 
        \DL3[43].tempL3[7] , \DL3[43].tempL3[6] , \DL3[43].tempL3[5] , 
        \DL3[43].tempL3[4] , \DL3[43].tempL3[3] , \DL3[43].tempL3[2] , 
        \DL3[43].tempL3[1] , \DL3[43].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2281}) );
  Dec4_16_20 \DL3[44].U3  ( .Hot({\DL3[44].tempL3[15] , \DL3[44].tempL3[14] , 
        \DL3[44].tempL3[13] , \DL3[44].tempL3[12] , \DL3[44].tempL3[11] , 
        \DL3[44].tempL3[10] , \DL3[44].tempL3[9] , \DL3[44].tempL3[8] , 
        \DL3[44].tempL3[7] , \DL3[44].tempL3[6] , \DL3[44].tempL3[5] , 
        \DL3[44].tempL3[4] , \DL3[44].tempL3[3] , \DL3[44].tempL3[2] , 
        \DL3[44].tempL3[1] , \DL3[44].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2281}) );
  Dec4_16_19 \DL3[45].U3  ( .Hot({\DL3[45].tempL3[15] , \DL3[45].tempL3[14] , 
        \DL3[45].tempL3[13] , \DL3[45].tempL3[12] , \DL3[45].tempL3[11] , 
        \DL3[45].tempL3[10] , \DL3[45].tempL3[9] , \DL3[45].tempL3[8] , 
        \DL3[45].tempL3[7] , \DL3[45].tempL3[6] , \DL3[45].tempL3[5] , 
        \DL3[45].tempL3[4] , \DL3[45].tempL3[3] , \DL3[45].tempL3[2] , 
        \DL3[45].tempL3[1] , \DL3[45].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2281}) );
  Dec4_16_18 \DL3[46].U3  ( .Hot({\DL3[46].tempL3[15] , \DL3[46].tempL3[14] , 
        \DL3[46].tempL3[13] , \DL3[46].tempL3[12] , \DL3[46].tempL3[11] , 
        \DL3[46].tempL3[10] , \DL3[46].tempL3[9] , \DL3[46].tempL3[8] , 
        \DL3[46].tempL3[7] , \DL3[46].tempL3[6] , \DL3[46].tempL3[5] , 
        \DL3[46].tempL3[4] , \DL3[46].tempL3[3] , \DL3[46].tempL3[2] , 
        \DL3[46].tempL3[1] , \DL3[46].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2272}) );
  Dec4_16_17 \DL3[47].U3  ( .Hot({\DL3[47].tempL3[15] , \DL3[47].tempL3[14] , 
        \DL3[47].tempL3[13] , \DL3[47].tempL3[12] , \DL3[47].tempL3[11] , 
        \DL3[47].tempL3[10] , \DL3[47].tempL3[9] , \DL3[47].tempL3[8] , 
        \DL3[47].tempL3[7] , \DL3[47].tempL3[6] , \DL3[47].tempL3[5] , 
        \DL3[47].tempL3[4] , \DL3[47].tempL3[3] , \DL3[47].tempL3[2] , 
        \DL3[47].tempL3[1] , \DL3[47].tempL3[0] }), .Sel({n2294, n2289, n2279, 
        n2280}) );
  Dec4_16_16 \DL3[48].U3  ( .Hot({\DL3[48].tempL3[15] , \DL3[48].tempL3[14] , 
        \DL3[48].tempL3[13] , \DL3[48].tempL3[12] , \DL3[48].tempL3[11] , 
        \DL3[48].tempL3[10] , \DL3[48].tempL3[9] , \DL3[48].tempL3[8] , 
        \DL3[48].tempL3[7] , \DL3[48].tempL3[6] , \DL3[48].tempL3[5] , 
        \DL3[48].tempL3[4] , \DL3[48].tempL3[3] , \DL3[48].tempL3[2] , 
        \DL3[48].tempL3[1] , \DL3[48].tempL3[0] }), .Sel({n2292, n2290, n2284, 
        n2280}) );
  Dec4_16_15 \DL3[49].U3  ( .Hot({\DL3[49].tempL3[15] , \DL3[49].tempL3[14] , 
        \DL3[49].tempL3[13] , \DL3[49].tempL3[12] , \DL3[49].tempL3[11] , 
        \DL3[49].tempL3[10] , \DL3[49].tempL3[9] , \DL3[49].tempL3[8] , 
        \DL3[49].tempL3[7] , \DL3[49].tempL3[6] , \DL3[49].tempL3[5] , 
        \DL3[49].tempL3[4] , \DL3[49].tempL3[3] , \DL3[49].tempL3[2] , 
        \DL3[49].tempL3[1] , \DL3[49].tempL3[0] }), .Sel({n2292, n2288, n2284, 
        n2282}) );
  Dec4_16_14 \DL3[50].U3  ( .Hot({\DL3[50].tempL3[15] , \DL3[50].tempL3[14] , 
        \DL3[50].tempL3[13] , \DL3[50].tempL3[12] , \DL3[50].tempL3[11] , 
        \DL3[50].tempL3[10] , \DL3[50].tempL3[9] , \DL3[50].tempL3[8] , 
        \DL3[50].tempL3[7] , \DL3[50].tempL3[6] , \DL3[50].tempL3[5] , 
        \DL3[50].tempL3[4] , \DL3[50].tempL3[3] , \DL3[50].tempL3[2] , 
        \DL3[50].tempL3[1] , \DL3[50].tempL3[0] }), .Sel({n2295, n2288, n2279, 
        n2271}) );
  Dec4_16_13 \DL3[51].U3  ( .Hot({\DL3[51].tempL3[15] , \DL3[51].tempL3[14] , 
        \DL3[51].tempL3[13] , \DL3[51].tempL3[12] , \DL3[51].tempL3[11] , 
        \DL3[51].tempL3[10] , \DL3[51].tempL3[9] , \DL3[51].tempL3[8] , 
        \DL3[51].tempL3[7] , \DL3[51].tempL3[6] , \DL3[51].tempL3[5] , 
        \DL3[51].tempL3[4] , \DL3[51].tempL3[3] , \DL3[51].tempL3[2] , 
        \DL3[51].tempL3[1] , \DL3[51].tempL3[0] }), .Sel({n2292, n2288, n2284, 
        n2282}) );
  Dec4_16_12 \DL3[52].U3  ( .Hot({\DL3[52].tempL3[15] , \DL3[52].tempL3[14] , 
        \DL3[52].tempL3[13] , \DL3[52].tempL3[12] , \DL3[52].tempL3[11] , 
        \DL3[52].tempL3[10] , \DL3[52].tempL3[9] , \DL3[52].tempL3[8] , 
        \DL3[52].tempL3[7] , \DL3[52].tempL3[6] , \DL3[52].tempL3[5] , 
        \DL3[52].tempL3[4] , \DL3[52].tempL3[3] , \DL3[52].tempL3[2] , 
        \DL3[52].tempL3[1] , \DL3[52].tempL3[0] }), .Sel({n2295, n2288, n2284, 
        n2282}) );
  Dec4_16_11 \DL3[53].U3  ( .Hot({\DL3[53].tempL3[15] , \DL3[53].tempL3[14] , 
        \DL3[53].tempL3[13] , \DL3[53].tempL3[12] , \DL3[53].tempL3[11] , 
        \DL3[53].tempL3[10] , \DL3[53].tempL3[9] , \DL3[53].tempL3[8] , 
        \DL3[53].tempL3[7] , \DL3[53].tempL3[6] , \DL3[53].tempL3[5] , 
        \DL3[53].tempL3[4] , \DL3[53].tempL3[3] , \DL3[53].tempL3[2] , 
        \DL3[53].tempL3[1] , \DL3[53].tempL3[0] }), .Sel({n2292, n2290, n2284, 
        n2282}) );
  Dec4_16_10 \DL3[54].U3  ( .Hot({\DL3[54].tempL3[15] , \DL3[54].tempL3[14] , 
        \DL3[54].tempL3[13] , \DL3[54].tempL3[12] , \DL3[54].tempL3[11] , 
        \DL3[54].tempL3[10] , \DL3[54].tempL3[9] , \DL3[54].tempL3[8] , 
        \DL3[54].tempL3[7] , \DL3[54].tempL3[6] , \DL3[54].tempL3[5] , 
        \DL3[54].tempL3[4] , \DL3[54].tempL3[3] , \DL3[54].tempL3[2] , 
        \DL3[54].tempL3[1] , \DL3[54].tempL3[0] }), .Sel({n2295, n2290, n2284, 
        n2271}) );
  Dec4_16_9 \DL3[55].U3  ( .Hot({\DL3[55].tempL3[15] , \DL3[55].tempL3[14] , 
        \DL3[55].tempL3[13] , \DL3[55].tempL3[12] , \DL3[55].tempL3[11] , 
        \DL3[55].tempL3[10] , \DL3[55].tempL3[9] , \DL3[55].tempL3[8] , 
        \DL3[55].tempL3[7] , \DL3[55].tempL3[6] , \DL3[55].tempL3[5] , 
        \DL3[55].tempL3[4] , \DL3[55].tempL3[3] , \DL3[55].tempL3[2] , 
        \DL3[55].tempL3[1] , \DL3[55].tempL3[0] }), .Sel({n2295, n2290, n2284, 
        n2282}) );
  Dec4_16_8 \DL3[56].U3  ( .Hot({\DL3[56].tempL3[15] , \DL3[56].tempL3[14] , 
        \DL3[56].tempL3[13] , \DL3[56].tempL3[12] , \DL3[56].tempL3[11] , 
        \DL3[56].tempL3[10] , \DL3[56].tempL3[9] , \DL3[56].tempL3[8] , 
        \DL3[56].tempL3[7] , \DL3[56].tempL3[6] , \DL3[56].tempL3[5] , 
        \DL3[56].tempL3[4] , \DL3[56].tempL3[3] , \DL3[56].tempL3[2] , 
        \DL3[56].tempL3[1] , \DL3[56].tempL3[0] }), .Sel({n2292, n2290, n2284, 
        n2282}) );
  Dec4_16_7 \DL3[57].U3  ( .Hot({\DL3[57].tempL3[15] , \DL3[57].tempL3[14] , 
        \DL3[57].tempL3[13] , \DL3[57].tempL3[12] , \DL3[57].tempL3[11] , 
        \DL3[57].tempL3[10] , \DL3[57].tempL3[9] , \DL3[57].tempL3[8] , 
        \DL3[57].tempL3[7] , \DL3[57].tempL3[6] , \DL3[57].tempL3[5] , 
        \DL3[57].tempL3[4] , \DL3[57].tempL3[3] , \DL3[57].tempL3[2] , 
        \DL3[57].tempL3[1] , \DL3[57].tempL3[0] }), .Sel({n2292, n2288, n2284, 
        n2282}) );
  Dec4_16_6 \DL3[58].U3  ( .Hot({\DL3[58].tempL3[15] , \DL3[58].tempL3[14] , 
        \DL3[58].tempL3[13] , \DL3[58].tempL3[12] , \DL3[58].tempL3[11] , 
        \DL3[58].tempL3[10] , \DL3[58].tempL3[9] , \DL3[58].tempL3[8] , 
        \DL3[58].tempL3[7] , \DL3[58].tempL3[6] , \DL3[58].tempL3[5] , 
        \DL3[58].tempL3[4] , \DL3[58].tempL3[3] , \DL3[58].tempL3[2] , 
        \DL3[58].tempL3[1] , \DL3[58].tempL3[0] }), .Sel({n2295, n2288, n2284, 
        n2271}) );
  Dec4_16_5 \DL3[59].U3  ( .Hot({\DL3[59].tempL3[15] , \DL3[59].tempL3[14] , 
        \DL3[59].tempL3[13] , \DL3[59].tempL3[12] , \DL3[59].tempL3[11] , 
        \DL3[59].tempL3[10] , \DL3[59].tempL3[9] , \DL3[59].tempL3[8] , 
        \DL3[59].tempL3[7] , \DL3[59].tempL3[6] , \DL3[59].tempL3[5] , 
        \DL3[59].tempL3[4] , \DL3[59].tempL3[3] , \DL3[59].tempL3[2] , 
        \DL3[59].tempL3[1] , \DL3[59].tempL3[0] }), .Sel({n2295, n2290, n2284, 
        n2282}) );
  Dec4_16_4 \DL3[60].U3  ( .Hot({\DL3[60].tempL3[15] , \DL3[60].tempL3[14] , 
        \DL3[60].tempL3[13] , \DL3[60].tempL3[12] , \DL3[60].tempL3[11] , 
        \DL3[60].tempL3[10] , \DL3[60].tempL3[9] , \DL3[60].tempL3[8] , 
        \DL3[60].tempL3[7] , \DL3[60].tempL3[6] , \DL3[60].tempL3[5] , 
        \DL3[60].tempL3[4] , \DL3[60].tempL3[3] , \DL3[60].tempL3[2] , 
        \DL3[60].tempL3[1] , \DL3[60].tempL3[0] }), .Sel({n2295, n2290, n2285, 
        n2282}) );
  Dec4_16_3 \DL3[61].U3  ( .Hot({\DL3[61].tempL3[15] , \DL3[61].tempL3[14] , 
        \DL3[61].tempL3[13] , \DL3[61].tempL3[12] , \DL3[61].tempL3[11] , 
        \DL3[61].tempL3[10] , \DL3[61].tempL3[9] , \DL3[61].tempL3[8] , 
        \DL3[61].tempL3[7] , \DL3[61].tempL3[6] , \DL3[61].tempL3[5] , 
        \DL3[61].tempL3[4] , \DL3[61].tempL3[3] , \DL3[61].tempL3[2] , 
        \DL3[61].tempL3[1] , \DL3[61].tempL3[0] }), .Sel({n2295, n2290, n2285, 
        n2282}) );
  Dec4_16_2 \DL3[62].U3  ( .Hot({\DL3[62].tempL3[15] , \DL3[62].tempL3[14] , 
        \DL3[62].tempL3[13] , \DL3[62].tempL3[12] , \DL3[62].tempL3[11] , 
        \DL3[62].tempL3[10] , \DL3[62].tempL3[9] , \DL3[62].tempL3[8] , 
        \DL3[62].tempL3[7] , \DL3[62].tempL3[6] , \DL3[62].tempL3[5] , 
        \DL3[62].tempL3[4] , \DL3[62].tempL3[3] , \DL3[62].tempL3[2] , 
        \DL3[62].tempL3[1] , \DL3[62].tempL3[0] }), .Sel({n2295, n2290, n2273, 
        n2282}) );
  Dec4_16_1 \DL3[63].U3  ( .Hot({\DL3[63].tempL3[15] , \DL3[63].tempL3[14] , 
        \DL3[63].tempL3[13] , \DL3[63].tempL3[12] , \DL3[63].tempL3[11] , 
        \DL3[63].tempL3[10] , \DL3[63].tempL3[9] , \DL3[63].tempL3[8] , 
        \DL3[63].tempL3[7] , \DL3[63].tempL3[6] , \DL3[63].tempL3[5] , 
        \DL3[63].tempL3[4] , \DL3[63].tempL3[3] , \DL3[63].tempL3[2] , 
        \DL3[63].tempL3[1] , \DL3[63].tempL3[0] }), .Sel({n2295, n2290, n2285, 
        n2282}) );
  ND2D1 U1091 ( .A1(\DL3[0].tempL3[11] ), .A2(n2), .ZN(n66) );
  ND2D1 U1092 ( .A1(\DL3[0].tempL3[14] ), .A2(n2), .ZN(n67) );
  ND2D1 U1093 ( .A1(\DL3[0].tempL3[15] ), .A2(n2), .ZN(n68) );
  ND2D1 U1094 ( .A1(\DL3[1].tempL3[11] ), .A2(n51), .ZN(n69) );
  ND2D1 U1095 ( .A1(\DL3[1].tempL3[13] ), .A2(n51), .ZN(n70) );
  ND2D1 U1096 ( .A1(\DL3[1].tempL3[14] ), .A2(n51), .ZN(n71) );
  ND2D1 U1097 ( .A1(\DL3[1].tempL3[15] ), .A2(n51), .ZN(n72) );
  ND2D1 U1098 ( .A1(\DL3[2].tempL3[11] ), .A2(n40), .ZN(n73) );
  ND2D1 U1099 ( .A1(\DL3[2].tempL3[13] ), .A2(n40), .ZN(n74) );
  ND2D1 U1100 ( .A1(\DL3[2].tempL3[14] ), .A2(n40), .ZN(n75) );
  ND2D1 U1101 ( .A1(\DL3[2].tempL3[15] ), .A2(n40), .ZN(n76) );
  ND2D1 U1102 ( .A1(\DL3[3].tempL3[11] ), .A2(n29), .ZN(n77) );
  ND2D1 U1103 ( .A1(\DL3[3].tempL3[13] ), .A2(n29), .ZN(n78) );
  ND2D1 U1104 ( .A1(\DL3[3].tempL3[14] ), .A2(n29), .ZN(n79) );
  ND2D1 U1105 ( .A1(\DL3[3].tempL3[15] ), .A2(n29), .ZN(n80) );
  ND2D1 U1106 ( .A1(\DL3[4].tempL3[11] ), .A2(n18), .ZN(n81) );
  ND2D1 U1107 ( .A1(\DL3[4].tempL3[13] ), .A2(n18), .ZN(n82) );
  ND2D1 U1108 ( .A1(\DL3[4].tempL3[14] ), .A2(n18), .ZN(n83) );
  ND2D1 U1109 ( .A1(\DL3[4].tempL3[15] ), .A2(n18), .ZN(n84) );
  ND2D1 U1110 ( .A1(\DL3[5].tempL3[11] ), .A2(n7), .ZN(n85) );
  ND2D1 U1111 ( .A1(\DL3[5].tempL3[13] ), .A2(n7), .ZN(n86) );
  ND2D1 U1112 ( .A1(\DL3[5].tempL3[14] ), .A2(n7), .ZN(n87) );
  ND2D1 U1113 ( .A1(\DL3[5].tempL3[15] ), .A2(n7), .ZN(n88) );
  ND2D1 U1114 ( .A1(\DL3[6].tempL3[11] ), .A2(n3), .ZN(n89) );
  ND2D1 U1115 ( .A1(\DL3[6].tempL3[13] ), .A2(n3), .ZN(n90) );
  ND2D1 U1116 ( .A1(\DL3[6].tempL3[14] ), .A2(n3), .ZN(n91) );
  ND2D1 U1117 ( .A1(\DL3[6].tempL3[15] ), .A2(n3), .ZN(n92) );
  ND2D1 U1118 ( .A1(\DL3[7].tempL3[11] ), .A2(n64), .ZN(n93) );
  ND2D1 U1119 ( .A1(\DL3[7].tempL3[13] ), .A2(n64), .ZN(n94) );
  ND2D1 U1120 ( .A1(\DL3[7].tempL3[14] ), .A2(n64), .ZN(n95) );
  ND2D1 U1121 ( .A1(\DL3[7].tempL3[15] ), .A2(n64), .ZN(n96) );
  ND2D1 U1122 ( .A1(\DL3[8].tempL3[11] ), .A2(n63), .ZN(n97) );
  ND2D1 U1123 ( .A1(\DL3[8].tempL3[13] ), .A2(n63), .ZN(n98) );
  ND2D1 U1124 ( .A1(\DL3[8].tempL3[14] ), .A2(n63), .ZN(n99) );
  ND2D1 U1125 ( .A1(\DL3[8].tempL3[15] ), .A2(n63), .ZN(n100) );
  ND2D1 U1126 ( .A1(\DL3[9].tempL3[11] ), .A2(n62), .ZN(n101) );
  ND2D1 U1127 ( .A1(\DL3[9].tempL3[13] ), .A2(n62), .ZN(n102) );
  ND2D1 U1128 ( .A1(\DL3[9].tempL3[14] ), .A2(n62), .ZN(n103) );
  ND2D1 U1129 ( .A1(\DL3[9].tempL3[15] ), .A2(n62), .ZN(n104) );
  ND2D1 U1130 ( .A1(\DL3[10].tempL3[11] ), .A2(n61), .ZN(n105) );
  ND2D1 U1131 ( .A1(\DL3[10].tempL3[13] ), .A2(n61), .ZN(n106) );
  ND2D1 U1132 ( .A1(\DL3[10].tempL3[14] ), .A2(n61), .ZN(n107) );
  ND2D1 U1133 ( .A1(\DL3[10].tempL3[15] ), .A2(n61), .ZN(n108) );
  ND2D1 U1134 ( .A1(\DL3[11].tempL3[13] ), .A2(n60), .ZN(n109) );
  ND2D1 U1135 ( .A1(\DL3[11].tempL3[14] ), .A2(n60), .ZN(n110) );
  ND2D1 U1136 ( .A1(\DL3[11].tempL3[15] ), .A2(n60), .ZN(n111) );
  ND2D1 U1137 ( .A1(\DL3[12].tempL3[13] ), .A2(n59), .ZN(n112) );
  ND2D1 U1138 ( .A1(\DL3[12].tempL3[14] ), .A2(n59), .ZN(n113) );
  ND2D1 U1139 ( .A1(\DL3[12].tempL3[15] ), .A2(n59), .ZN(n114) );
  ND2D1 U1140 ( .A1(\DL3[13].tempL3[13] ), .A2(n58), .ZN(n115) );
  ND2D1 U1141 ( .A1(\DL3[13].tempL3[14] ), .A2(n58), .ZN(n116) );
  ND2D1 U1142 ( .A1(\DL3[13].tempL3[15] ), .A2(n58), .ZN(n117) );
  ND2D1 U1143 ( .A1(\DL3[14].tempL3[13] ), .A2(n57), .ZN(n118) );
  ND2D1 U1144 ( .A1(\DL3[14].tempL3[14] ), .A2(n57), .ZN(n119) );
  ND2D1 U1145 ( .A1(\DL3[14].tempL3[15] ), .A2(n57), .ZN(n120) );
  ND2D1 U1146 ( .A1(\DL3[15].tempL3[13] ), .A2(n56), .ZN(n121) );
  ND2D1 U1147 ( .A1(\DL3[15].tempL3[14] ), .A2(n56), .ZN(n122) );
  ND2D1 U1148 ( .A1(\DL3[15].tempL3[15] ), .A2(n56), .ZN(n123) );
  ND2D1 U1149 ( .A1(\DL3[32].tempL3[10] ), .A2(n37), .ZN(n124) );
  ND2D1 U1150 ( .A1(\DL3[32].tempL3[11] ), .A2(n37), .ZN(n125) );
  ND2D1 U1151 ( .A1(\DL3[32].tempL3[12] ), .A2(n37), .ZN(n126) );
  ND2D1 U1152 ( .A1(\DL3[32].tempL3[13] ), .A2(n37), .ZN(n127) );
  ND2D1 U1153 ( .A1(\DL3[32].tempL3[14] ), .A2(n37), .ZN(n128) );
  ND2D1 U1154 ( .A1(\DL3[32].tempL3[15] ), .A2(n37), .ZN(n129) );
  ND2D1 U1155 ( .A1(\DL3[33].tempL3[10] ), .A2(n36), .ZN(n130) );
  ND2D1 U1156 ( .A1(\DL3[33].tempL3[11] ), .A2(n36), .ZN(n131) );
  ND2D1 U1157 ( .A1(\DL3[33].tempL3[12] ), .A2(n36), .ZN(n132) );
  ND2D1 U1158 ( .A1(\DL3[33].tempL3[13] ), .A2(n36), .ZN(n133) );
  ND2D1 U1159 ( .A1(\DL3[33].tempL3[14] ), .A2(n36), .ZN(n134) );
  ND2D1 U1160 ( .A1(\DL3[33].tempL3[15] ), .A2(n36), .ZN(n135) );
  ND2D1 U1161 ( .A1(\DL3[34].tempL3[10] ), .A2(n35), .ZN(n136) );
  ND2D1 U1162 ( .A1(\DL3[34].tempL3[11] ), .A2(n35), .ZN(n137) );
  ND2D1 U1163 ( .A1(\DL3[34].tempL3[12] ), .A2(n35), .ZN(n138) );
  ND2D1 U1164 ( .A1(\DL3[34].tempL3[13] ), .A2(n35), .ZN(n139) );
  ND2D1 U1165 ( .A1(\DL3[34].tempL3[14] ), .A2(n35), .ZN(n140) );
  ND2D1 U1166 ( .A1(\DL3[34].tempL3[15] ), .A2(n35), .ZN(n141) );
  ND2D1 U1167 ( .A1(\DL3[35].tempL3[10] ), .A2(n34), .ZN(n142) );
  ND2D1 U1168 ( .A1(\DL3[35].tempL3[11] ), .A2(n34), .ZN(n143) );
  ND2D1 U1169 ( .A1(\DL3[35].tempL3[12] ), .A2(n34), .ZN(n144) );
  ND2D1 U1170 ( .A1(\DL3[35].tempL3[13] ), .A2(n34), .ZN(n145) );
  ND2D1 U1171 ( .A1(\DL3[35].tempL3[14] ), .A2(n34), .ZN(n146) );
  ND2D1 U1172 ( .A1(\DL3[35].tempL3[15] ), .A2(n34), .ZN(n147) );
  ND2D1 U1173 ( .A1(\DL3[36].tempL3[10] ), .A2(n33), .ZN(n148) );
  ND2D1 U1174 ( .A1(\DL3[36].tempL3[11] ), .A2(n33), .ZN(n149) );
  ND2D1 U1175 ( .A1(\DL3[36].tempL3[12] ), .A2(n33), .ZN(n150) );
  ND2D1 U1176 ( .A1(\DL3[36].tempL3[13] ), .A2(n33), .ZN(n151) );
  ND2D1 U1177 ( .A1(\DL3[36].tempL3[14] ), .A2(n33), .ZN(n152) );
  ND2D1 U1178 ( .A1(\DL3[36].tempL3[15] ), .A2(n33), .ZN(n153) );
  ND2D1 U1179 ( .A1(\DL3[37].tempL3[10] ), .A2(n32), .ZN(n154) );
  ND2D1 U1180 ( .A1(\DL3[37].tempL3[11] ), .A2(n32), .ZN(n155) );
  ND2D1 U1181 ( .A1(\DL3[37].tempL3[12] ), .A2(n32), .ZN(n156) );
  ND2D1 U1182 ( .A1(\DL3[37].tempL3[13] ), .A2(n32), .ZN(n157) );
  ND2D1 U1183 ( .A1(\DL3[37].tempL3[14] ), .A2(n32), .ZN(n158) );
  ND2D1 U1184 ( .A1(\DL3[37].tempL3[15] ), .A2(n32), .ZN(n159) );
  ND2D1 U1185 ( .A1(\DL3[38].tempL3[10] ), .A2(n31), .ZN(n160) );
  ND2D1 U1186 ( .A1(\DL3[38].tempL3[11] ), .A2(n31), .ZN(n161) );
  ND2D1 U1187 ( .A1(\DL3[38].tempL3[12] ), .A2(n31), .ZN(n162) );
  ND2D1 U1188 ( .A1(\DL3[38].tempL3[13] ), .A2(n31), .ZN(n163) );
  ND2D1 U1189 ( .A1(\DL3[38].tempL3[14] ), .A2(n31), .ZN(n164) );
  ND2D1 U1190 ( .A1(\DL3[38].tempL3[15] ), .A2(n31), .ZN(n165) );
  ND2D1 U1191 ( .A1(\DL3[39].tempL3[10] ), .A2(n30), .ZN(n166) );
  ND2D1 U1192 ( .A1(\DL3[39].tempL3[11] ), .A2(n30), .ZN(n167) );
  ND2D1 U1193 ( .A1(\DL3[39].tempL3[12] ), .A2(n30), .ZN(n168) );
  ND2D1 U1194 ( .A1(\DL3[39].tempL3[13] ), .A2(n30), .ZN(n169) );
  ND2D1 U1195 ( .A1(\DL3[39].tempL3[14] ), .A2(n30), .ZN(n170) );
  ND2D1 U1196 ( .A1(\DL3[39].tempL3[15] ), .A2(n30), .ZN(n171) );
  ND2D1 U1197 ( .A1(\DL3[40].tempL3[10] ), .A2(n28), .ZN(n172) );
  ND2D1 U1198 ( .A1(\DL3[40].tempL3[11] ), .A2(n28), .ZN(n173) );
  ND2D1 U1199 ( .A1(\DL3[40].tempL3[12] ), .A2(n28), .ZN(n174) );
  ND2D1 U1200 ( .A1(\DL3[40].tempL3[13] ), .A2(n28), .ZN(n175) );
  ND2D1 U1201 ( .A1(\DL3[40].tempL3[14] ), .A2(n28), .ZN(n176) );
  ND2D1 U1202 ( .A1(\DL3[40].tempL3[15] ), .A2(n28), .ZN(n177) );
  ND2D1 U1203 ( .A1(\DL3[41].tempL3[10] ), .A2(n27), .ZN(n178) );
  ND2D1 U1204 ( .A1(\DL3[41].tempL3[11] ), .A2(n27), .ZN(n179) );
  ND2D1 U1205 ( .A1(\DL3[41].tempL3[12] ), .A2(n27), .ZN(n180) );
  ND2D1 U1206 ( .A1(\DL3[41].tempL3[13] ), .A2(n27), .ZN(n181) );
  ND2D1 U1207 ( .A1(\DL3[41].tempL3[14] ), .A2(n27), .ZN(n182) );
  ND2D1 U1208 ( .A1(\DL3[41].tempL3[15] ), .A2(n27), .ZN(n183) );
  ND2D1 U1209 ( .A1(\DL3[42].tempL3[10] ), .A2(n26), .ZN(n184) );
  ND2D1 U1210 ( .A1(\DL3[42].tempL3[11] ), .A2(n26), .ZN(n185) );
  ND2D1 U1211 ( .A1(\DL3[42].tempL3[12] ), .A2(n26), .ZN(n186) );
  ND2D1 U1212 ( .A1(\DL3[42].tempL3[13] ), .A2(n26), .ZN(n187) );
  ND2D1 U1213 ( .A1(\DL3[42].tempL3[14] ), .A2(n26), .ZN(n188) );
  ND2D1 U1214 ( .A1(\DL3[42].tempL3[15] ), .A2(n26), .ZN(n189) );
  ND2D1 U1215 ( .A1(\DL3[43].tempL3[10] ), .A2(n25), .ZN(n190) );
  ND2D1 U1216 ( .A1(\DL3[43].tempL3[11] ), .A2(n25), .ZN(n191) );
  ND2D1 U1217 ( .A1(\DL3[43].tempL3[12] ), .A2(n25), .ZN(n192) );
  ND2D1 U1218 ( .A1(\DL3[43].tempL3[13] ), .A2(n25), .ZN(n193) );
  ND2D1 U1219 ( .A1(\DL3[43].tempL3[14] ), .A2(n25), .ZN(n194) );
  ND2D1 U1220 ( .A1(\DL3[43].tempL3[15] ), .A2(n25), .ZN(n195) );
  ND2D1 U1221 ( .A1(\DL3[44].tempL3[10] ), .A2(n24), .ZN(n196) );
  ND2D1 U1222 ( .A1(\DL3[44].tempL3[11] ), .A2(n24), .ZN(n197) );
  ND2D1 U1223 ( .A1(\DL3[44].tempL3[12] ), .A2(n24), .ZN(n198) );
  ND2D1 U1224 ( .A1(\DL3[44].tempL3[13] ), .A2(n24), .ZN(n199) );
  ND2D1 U1225 ( .A1(\DL3[44].tempL3[14] ), .A2(n24), .ZN(n200) );
  ND2D1 U1226 ( .A1(\DL3[44].tempL3[15] ), .A2(n24), .ZN(n201) );
  ND2D1 U1227 ( .A1(\DL3[45].tempL3[10] ), .A2(n23), .ZN(n202) );
  ND2D1 U1228 ( .A1(\DL3[45].tempL3[11] ), .A2(n23), .ZN(n203) );
  ND2D1 U1229 ( .A1(\DL3[45].tempL3[12] ), .A2(n23), .ZN(n204) );
  ND2D1 U1230 ( .A1(\DL3[45].tempL3[13] ), .A2(n23), .ZN(n205) );
  ND2D1 U1231 ( .A1(\DL3[45].tempL3[14] ), .A2(n23), .ZN(n206) );
  ND2D1 U1232 ( .A1(\DL3[45].tempL3[15] ), .A2(n23), .ZN(n207) );
  ND2D1 U1233 ( .A1(\DL3[46].tempL3[10] ), .A2(n22), .ZN(n208) );
  ND2D1 U1234 ( .A1(\DL3[46].tempL3[11] ), .A2(n22), .ZN(n209) );
  ND2D1 U1235 ( .A1(\DL3[46].tempL3[12] ), .A2(n22), .ZN(n210) );
  ND2D1 U1236 ( .A1(\DL3[46].tempL3[13] ), .A2(n22), .ZN(n211) );
  ND2D1 U1237 ( .A1(\DL3[46].tempL3[14] ), .A2(n22), .ZN(n212) );
  ND2D1 U1238 ( .A1(\DL3[46].tempL3[15] ), .A2(n22), .ZN(n213) );
  ND2D1 U1239 ( .A1(\DL3[47].tempL3[11] ), .A2(n21), .ZN(n214) );
  ND2D1 U1240 ( .A1(\DL3[47].tempL3[12] ), .A2(n21), .ZN(n215) );
  ND2D1 U1241 ( .A1(\DL3[47].tempL3[13] ), .A2(n21), .ZN(n216) );
  ND2D1 U1242 ( .A1(\DL3[47].tempL3[14] ), .A2(n21), .ZN(n217) );
  ND2D1 U1243 ( .A1(\DL3[47].tempL3[15] ), .A2(n21), .ZN(n218) );
  ND2D1 U1244 ( .A1(\DL3[50].tempL3[15] ), .A2(n17), .ZN(n219) );
  ND2D1 U1245 ( .A1(\DL3[57].tempL3[15] ), .A2(n10), .ZN(n220) );
  ND2D1 U1246 ( .A1(\DL3[58].tempL3[15] ), .A2(n9), .ZN(n221) );
  ND2D1 U1247 ( .A1(\DL3[59].tempL3[15] ), .A2(n8), .ZN(n222) );
  BUFFD1 U1248 ( .I(Address[7]), .Z(n2279) );
  BUFFD1 U1249 ( .I(Address[3]), .Z(n2276) );
  BUFFD1 U1250 ( .I(Address[2]), .Z(n2275) );
  BUFFD1 U1251 ( .I(Address[5]), .Z(n2278) );
  BUFFD1 U1252 ( .I(Address[4]), .Z(n2277) );
  INVD1 U1253 ( .I(n2291), .ZN(n2287) );
  INVD1 U1254 ( .I(n2296), .ZN(n2293) );
  INVD1 U1255 ( .I(n2283), .ZN(n2281) );
  INVD1 U1256 ( .I(n2283), .ZN(n2272) );
  INVD1 U1257 ( .I(n2291), .ZN(n2289) );
  INVD1 U1258 ( .I(n2296), .ZN(n2294) );
  INVD1 U1259 ( .I(n2286), .ZN(n2285) );
  AN2D1 U1260 ( .A1(DecodedL1[0]), .A2(\DL2[0].tempL2[0] ), .Z(n2) );
  AN2D1 U1261 ( .A1(\DL2[0].tempL2[1] ), .A2(DecodedL1[0]), .Z(n51) );
  AN2D1 U1262 ( .A1(\DL2[0].tempL2[2] ), .A2(DecodedL1[0]), .Z(n40) );
  AN2D1 U1263 ( .A1(\DL2[0].tempL2[3] ), .A2(DecodedL1[0]), .Z(n29) );
  AN2D1 U1264 ( .A1(\DL2[0].tempL2[4] ), .A2(DecodedL1[0]), .Z(n18) );
  AN2D1 U1265 ( .A1(\DL2[0].tempL2[5] ), .A2(DecodedL1[0]), .Z(n7) );
  AN2D1 U1266 ( .A1(\DL2[0].tempL2[6] ), .A2(DecodedL1[0]), .Z(n3) );
  AN2D1 U1267 ( .A1(\DL2[0].tempL2[7] ), .A2(DecodedL1[0]), .Z(n64) );
  AN2D1 U1268 ( .A1(\DL2[0].tempL2[8] ), .A2(DecodedL1[0]), .Z(n63) );
  AN2D1 U1269 ( .A1(\DL2[0].tempL2[9] ), .A2(DecodedL1[0]), .Z(n62) );
  AN2D1 U1270 ( .A1(\DL2[0].tempL2[10] ), .A2(DecodedL1[0]), .Z(n61) );
  AN2D1 U1271 ( .A1(\DL2[0].tempL2[11] ), .A2(DecodedL1[0]), .Z(n60) );
  AN2D1 U1272 ( .A1(\DL2[0].tempL2[12] ), .A2(DecodedL1[0]), .Z(n59) );
  AN2D1 U1273 ( .A1(\DL2[0].tempL2[13] ), .A2(DecodedL1[0]), .Z(n58) );
  AN2D1 U1274 ( .A1(\DL2[0].tempL2[14] ), .A2(DecodedL1[0]), .Z(n57) );
  AN2D1 U1275 ( .A1(\DL2[0].tempL2[15] ), .A2(DecodedL1[0]), .Z(n56) );
  AN2D1 U1276 ( .A1(\DL2[1].tempL2[1] ), .A2(DecodedL1[1]), .Z(n54) );
  AN2D1 U1277 ( .A1(\DL2[1].tempL2[2] ), .A2(DecodedL1[1]), .Z(n53) );
  AN2D1 U1278 ( .A1(\DL2[1].tempL2[3] ), .A2(DecodedL1[1]), .Z(n52) );
  AN2D1 U1279 ( .A1(\DL2[1].tempL2[4] ), .A2(DecodedL1[1]), .Z(n50) );
  AN2D1 U1280 ( .A1(\DL2[1].tempL2[5] ), .A2(DecodedL1[1]), .Z(n49) );
  AN2D1 U1281 ( .A1(\DL2[1].tempL2[6] ), .A2(DecodedL1[1]), .Z(n48) );
  AN2D1 U1282 ( .A1(\DL2[1].tempL2[7] ), .A2(DecodedL1[1]), .Z(n47) );
  AN2D1 U1283 ( .A1(\DL2[1].tempL2[8] ), .A2(DecodedL1[1]), .Z(n46) );
  AN2D1 U1284 ( .A1(\DL2[1].tempL2[9] ), .A2(DecodedL1[1]), .Z(n45) );
  AN2D1 U1285 ( .A1(\DL2[1].tempL2[10] ), .A2(DecodedL1[1]), .Z(n44) );
  AN2D1 U1286 ( .A1(\DL2[1].tempL2[11] ), .A2(DecodedL1[1]), .Z(n43) );
  AN2D1 U1287 ( .A1(\DL2[1].tempL2[12] ), .A2(DecodedL1[1]), .Z(n42) );
  AN2D1 U1288 ( .A1(\DL2[1].tempL2[13] ), .A2(DecodedL1[1]), .Z(n41) );
  AN2D1 U1289 ( .A1(\DL2[1].tempL2[14] ), .A2(DecodedL1[1]), .Z(n39) );
  AN2D1 U1290 ( .A1(DecodedL1[1]), .A2(\DL2[1].tempL2[15] ), .Z(n38) );
  AN2D1 U1291 ( .A1(\DL2[2].tempL2[0] ), .A2(DecodedL1[2]), .Z(n37) );
  AN2D1 U1292 ( .A1(\DL2[2].tempL2[1] ), .A2(DecodedL1[2]), .Z(n36) );
  AN2D1 U1293 ( .A1(\DL2[2].tempL2[2] ), .A2(DecodedL1[2]), .Z(n35) );
  AN2D1 U1294 ( .A1(\DL2[2].tempL2[3] ), .A2(DecodedL1[2]), .Z(n34) );
  AN2D1 U1295 ( .A1(\DL2[2].tempL2[4] ), .A2(DecodedL1[2]), .Z(n33) );
  AN2D1 U1296 ( .A1(\DL2[2].tempL2[5] ), .A2(DecodedL1[2]), .Z(n32) );
  AN2D1 U1297 ( .A1(\DL2[2].tempL2[7] ), .A2(DecodedL1[2]), .Z(n30) );
  AN2D1 U1298 ( .A1(\DL2[2].tempL2[8] ), .A2(DecodedL1[2]), .Z(n28) );
  AN2D1 U1299 ( .A1(\DL2[2].tempL2[9] ), .A2(DecodedL1[2]), .Z(n27) );
  AN2D1 U1300 ( .A1(\DL2[2].tempL2[10] ), .A2(DecodedL1[2]), .Z(n26) );
  AN2D1 U1301 ( .A1(\DL2[2].tempL2[11] ), .A2(DecodedL1[2]), .Z(n25) );
  AN2D1 U1302 ( .A1(\DL2[2].tempL2[12] ), .A2(DecodedL1[2]), .Z(n24) );
  AN2D1 U1303 ( .A1(\DL2[2].tempL2[13] ), .A2(DecodedL1[2]), .Z(n23) );
  AN2D1 U1304 ( .A1(\DL2[2].tempL2[14] ), .A2(DecodedL1[2]), .Z(n22) );
  AN2D1 U1305 ( .A1(DecodedL1[2]), .A2(\DL2[2].tempL2[15] ), .Z(n21) );
  AN2D1 U1306 ( .A1(\DL2[3].tempL2[0] ), .A2(DecodedL1[3]), .Z(n20) );
  AN2D1 U1307 ( .A1(\DL2[3].tempL2[1] ), .A2(DecodedL1[3]), .Z(n19) );
  AN2D1 U1308 ( .A1(\DL2[3].tempL2[2] ), .A2(DecodedL1[3]), .Z(n17) );
  AN2D1 U1309 ( .A1(\DL2[3].tempL2[4] ), .A2(DecodedL1[3]), .Z(n15) );
  AN2D1 U1310 ( .A1(\DL2[3].tempL2[5] ), .A2(DecodedL1[3]), .Z(n14) );
  AN2D1 U1311 ( .A1(\DL2[3].tempL2[6] ), .A2(DecodedL1[3]), .Z(n13) );
  AN2D1 U1312 ( .A1(\DL2[3].tempL2[7] ), .A2(DecodedL1[3]), .Z(n12) );
  AN2D1 U1313 ( .A1(\DL2[3].tempL2[8] ), .A2(DecodedL1[3]), .Z(n11) );
  AN2D1 U1314 ( .A1(\DL2[3].tempL2[9] ), .A2(DecodedL1[3]), .Z(n10) );
  AN2D1 U1315 ( .A1(\DL2[3].tempL2[10] ), .A2(DecodedL1[3]), .Z(n9) );
  AN2D1 U1316 ( .A1(\DL2[3].tempL2[11] ), .A2(DecodedL1[3]), .Z(n8) );
  AN2D1 U1317 ( .A1(\DL2[3].tempL2[12] ), .A2(DecodedL1[3]), .Z(n6) );
  AN2D1 U1318 ( .A1(\DL2[3].tempL2[13] ), .A2(DecodedL1[3]), .Z(n5) );
  AN2D1 U1319 ( .A1(DecodedL1[3]), .A2(\DL2[3].tempL2[14] ), .Z(n4) );
  AN2D1 U1320 ( .A1(\DL2[3].tempL2[15] ), .A2(DecodedL1[3]), .Z(n65) );
  BUFFD1 U1321 ( .I(Address[0]), .Z(n2274) );
  INVD1 U1322 ( .I(Address[9]), .ZN(n2296) );
  INVD1 U1323 ( .I(n2296), .ZN(n2295) );
  INVD1 U1324 ( .I(n2296), .ZN(n2292) );
  INVD1 U1325 ( .I(n2279), .ZN(n2286) );
  INVD1 U1326 ( .I(n2286), .ZN(n2284) );
  INVD1 U1327 ( .I(Address[6]), .ZN(n2283) );
  INVD1 U1328 ( .I(n2283), .ZN(n2282) );
  INVD1 U1329 ( .I(n2283), .ZN(n2271) );
  INVD1 U1330 ( .I(n2283), .ZN(n2280) );
  INVD1 U1331 ( .I(Address[8]), .ZN(n2291) );
  INVD1 U1332 ( .I(n2291), .ZN(n2290) );
  INVD1 U1333 ( .I(n2291), .ZN(n2288) );
  CKND2D0 U1334 ( .A1(\DL3[62].tempL3[1] ), .A2(n4), .ZN(n223) );
  CKNXD16 U1335 ( .I(n223), .ZN(AdrEna[993]) );
  CKND2D0 U1336 ( .A1(\DL3[46].tempL3[2] ), .A2(n22), .ZN(n225) );
  CKNXD16 U1337 ( .I(n225), .ZN(AdrEna[738]) );
  CKND2D0 U1338 ( .A1(\DL3[62].tempL3[2] ), .A2(n4), .ZN(n227) );
  CKNXD16 U1339 ( .I(n227), .ZN(AdrEna[994]) );
  CKND2D0 U1340 ( .A1(\DL3[10].tempL3[10] ), .A2(n61), .ZN(n229) );
  CKNXD16 U1341 ( .I(n229), .ZN(AdrEna[170]) );
  CKND2D0 U1342 ( .A1(\DL3[33].tempL3[5] ), .A2(n36), .ZN(n231) );
  CKNXD16 U1343 ( .I(n231), .ZN(AdrEna[533]) );
  CKND2D0 U1344 ( .A1(\DL3[5].tempL3[2] ), .A2(n7), .ZN(n233) );
  CKNXD16 U1345 ( .I(n233), .ZN(AdrEna[82]) );
  CKND2D0 U1346 ( .A1(\DL3[62].tempL3[7] ), .A2(n4), .ZN(n235) );
  CKNXD16 U1347 ( .I(n235), .ZN(AdrEna[999]) );
  CKND2D0 U1348 ( .A1(\DL3[1].tempL3[12] ), .A2(n51), .ZN(n237) );
  CKNXD16 U1349 ( .I(n237), .ZN(AdrEna[28]) );
  CKND2D0 U1350 ( .A1(\DL3[62].tempL3[8] ), .A2(n4), .ZN(n239) );
  CKNXD16 U1351 ( .I(n239), .ZN(AdrEna[1000]) );
  CKND2D0 U1352 ( .A1(\DL3[63].tempL3[0] ), .A2(n65), .ZN(n241) );
  CKNXD16 U1353 ( .I(n241), .ZN(AdrEna[1008]) );
  CKND2D0 U1354 ( .A1(\DL3[62].tempL3[12] ), .A2(n4), .ZN(n243) );
  CKNXD16 U1355 ( .I(n243), .ZN(AdrEna[1004]) );
  CKND2D0 U1356 ( .A1(\DL3[1].tempL3[0] ), .A2(n51), .ZN(n245) );
  CKNXD16 U1357 ( .I(n245), .ZN(AdrEna[16]) );
  CKND2D0 U1358 ( .A1(\DL3[1].tempL3[6] ), .A2(n51), .ZN(n247) );
  CKNXD16 U1359 ( .I(n247), .ZN(AdrEna[22]) );
  CKND2D0 U1360 ( .A1(\DL3[0].tempL3[7] ), .A2(n2), .ZN(n249) );
  CKNXD16 U1361 ( .I(n249), .ZN(AdrEna[7]) );
  CKND2D0 U1362 ( .A1(\DL3[63].tempL3[1] ), .A2(n65), .ZN(n251) );
  CKNXD16 U1363 ( .I(n251), .ZN(AdrEna[1009]) );
  CKND2D0 U1364 ( .A1(\DL3[1].tempL3[5] ), .A2(n51), .ZN(n253) );
  CKNXD16 U1365 ( .I(n253), .ZN(AdrEna[21]) );
  CKND2D0 U1366 ( .A1(\DL3[0].tempL3[3] ), .A2(n2), .ZN(n255) );
  CKNXD16 U1367 ( .I(n255), .ZN(AdrEna[3]) );
  CKND2D0 U1368 ( .A1(\DL3[63].tempL3[5] ), .A2(n65), .ZN(n257) );
  CKNXD16 U1369 ( .I(n257), .ZN(AdrEna[1013]) );
  CKND2D0 U1370 ( .A1(\DL3[63].tempL3[3] ), .A2(n65), .ZN(n259) );
  CKNXD16 U1371 ( .I(n259), .ZN(AdrEna[1011]) );
  CKND2D0 U1372 ( .A1(\DL3[0].tempL3[13] ), .A2(n2), .ZN(n261) );
  CKNXD16 U1373 ( .I(n261), .ZN(AdrEna[13]) );
  CKND2D0 U1374 ( .A1(\DL3[0].tempL3[5] ), .A2(n2), .ZN(n263) );
  CKNXD16 U1375 ( .I(n263), .ZN(AdrEna[5]) );
  CKND2D0 U1376 ( .A1(\DL3[63].tempL3[13] ), .A2(n65), .ZN(n265) );
  CKNXD16 U1377 ( .I(n265), .ZN(AdrEna[1021]) );
  CKND2D0 U1378 ( .A1(\DL3[63].tempL3[9] ), .A2(n65), .ZN(n267) );
  CKNXD16 U1379 ( .I(n267), .ZN(AdrEna[1017]) );
  CKND2D0 U1380 ( .A1(\DL3[0].tempL3[6] ), .A2(n2), .ZN(n269) );
  CKNXD16 U1381 ( .I(n269), .ZN(AdrEna[6]) );
  CKND2D0 U1382 ( .A1(\DL3[0].tempL3[4] ), .A2(n2), .ZN(n271) );
  CKNXD16 U1383 ( .I(n271), .ZN(AdrEna[4]) );
  CKBD0 U1384 ( .CLK(n69), .C(n273) );
  CKNXD16 U1385 ( .I(n273), .ZN(AdrEna[27]) );
  CKBD0 U1386 ( .CLK(n213), .C(n275) );
  CKNXD16 U1387 ( .I(n275), .ZN(AdrEna[751]) );
  CKBD0 U1388 ( .CLK(n66), .C(n277) );
  CKNXD16 U1389 ( .I(n277), .ZN(AdrEna[11]) );
  CKBD0 U1390 ( .CLK(n73), .C(n279) );
  CKNXD16 U1391 ( .I(n279), .ZN(AdrEna[43]) );
  CKBD0 U1392 ( .CLK(n189), .C(n281) );
  CKNXD16 U1393 ( .I(n281), .ZN(AdrEna[687]) );
  CKBD0 U1394 ( .CLK(n195), .C(n283) );
  CKNXD16 U1395 ( .I(n283), .ZN(AdrEna[703]) );
  CKBD0 U1396 ( .CLK(n201), .C(n285) );
  CKNXD16 U1397 ( .I(n285), .ZN(AdrEna[719]) );
  CKBD0 U1398 ( .CLK(n207), .C(n287) );
  CKNXD16 U1399 ( .I(n287), .ZN(AdrEna[735]) );
  CKBD0 U1400 ( .CLK(n171), .C(n289) );
  CKNXD16 U1401 ( .I(n289), .ZN(AdrEna[639]) );
  CKBD0 U1402 ( .CLK(n177), .C(n291) );
  CKNXD16 U1403 ( .I(n291), .ZN(AdrEna[655]) );
  CKBD0 U1404 ( .CLK(n183), .C(n293) );
  CKNXD16 U1405 ( .I(n293), .ZN(AdrEna[671]) );
  CKBD0 U1406 ( .CLK(n147), .C(n295) );
  CKNXD16 U1407 ( .I(n295), .ZN(AdrEna[575]) );
  CKBD0 U1408 ( .CLK(n153), .C(n297) );
  CKNXD16 U1409 ( .I(n297), .ZN(AdrEna[591]) );
  CKBD0 U1410 ( .CLK(n159), .C(n299) );
  CKNXD16 U1411 ( .I(n299), .ZN(AdrEna[607]) );
  CKBD0 U1412 ( .CLK(n165), .C(n301) );
  CKNXD16 U1413 ( .I(n301), .ZN(AdrEna[623]) );
  CKBD0 U1414 ( .CLK(n129), .C(n303) );
  CKNXD16 U1415 ( .I(n303), .ZN(AdrEna[527]) );
  CKBD0 U1416 ( .CLK(n135), .C(n305) );
  CKNXD16 U1417 ( .I(n305), .ZN(AdrEna[543]) );
  CKBD0 U1418 ( .CLK(n141), .C(n307) );
  CKNXD16 U1419 ( .I(n307), .ZN(AdrEna[559]) );
  CKBD0 U1420 ( .CLK(n200), .C(n309) );
  CKNXD16 U1421 ( .I(n309), .ZN(AdrEna[718]) );
  CKBD0 U1422 ( .CLK(n206), .C(n311) );
  CKNXD16 U1423 ( .I(n311), .ZN(AdrEna[734]) );
  CKBD0 U1424 ( .CLK(n212), .C(n313) );
  CKNXD16 U1425 ( .I(n313), .ZN(AdrEna[750]) );
  CKBD0 U1426 ( .CLK(n218), .C(n315) );
  CKNXD16 U1427 ( .I(n315), .ZN(AdrEna[767]) );
  CKBD0 U1428 ( .CLK(n182), .C(n317) );
  CKNXD16 U1429 ( .I(n317), .ZN(AdrEna[670]) );
  CKBD0 U1430 ( .CLK(n188), .C(n319) );
  CKNXD16 U1431 ( .I(n319), .ZN(AdrEna[686]) );
  CKBD0 U1432 ( .CLK(n194), .C(n321) );
  CKNXD16 U1433 ( .I(n321), .ZN(AdrEna[702]) );
  CKBD0 U1434 ( .CLK(n158), .C(n323) );
  CKNXD16 U1435 ( .I(n323), .ZN(AdrEna[606]) );
  CKBD0 U1436 ( .CLK(n164), .C(n325) );
  CKNXD16 U1437 ( .I(n325), .ZN(AdrEna[622]) );
  CKBD0 U1438 ( .CLK(n170), .C(n327) );
  CKNXD16 U1439 ( .I(n327), .ZN(AdrEna[638]) );
  CKBD0 U1440 ( .CLK(n176), .C(n329) );
  CKNXD16 U1441 ( .I(n329), .ZN(AdrEna[654]) );
  CKBD0 U1442 ( .CLK(n140), .C(n331) );
  CKNXD16 U1443 ( .I(n331), .ZN(AdrEna[558]) );
  CKBD0 U1444 ( .CLK(n146), .C(n333) );
  CKNXD16 U1445 ( .I(n333), .ZN(AdrEna[574]) );
  CKBD0 U1446 ( .CLK(n152), .C(n335) );
  CKNXD16 U1447 ( .I(n335), .ZN(AdrEna[590]) );
  CKBD0 U1448 ( .CLK(n211), .C(n337) );
  CKNXD16 U1449 ( .I(n337), .ZN(AdrEna[749]) );
  CKBD0 U1450 ( .CLK(n217), .C(n339) );
  CKNXD16 U1451 ( .I(n339), .ZN(AdrEna[766]) );
  CKBD0 U1452 ( .CLK(n128), .C(n341) );
  CKNXD16 U1453 ( .I(n341), .ZN(AdrEna[526]) );
  CKBD0 U1454 ( .CLK(n134), .C(n343) );
  CKNXD16 U1455 ( .I(n343), .ZN(AdrEna[542]) );
  CKBD0 U1456 ( .CLK(n193), .C(n345) );
  CKNXD16 U1457 ( .I(n345), .ZN(AdrEna[701]) );
  CKBD0 U1458 ( .CLK(n199), .C(n347) );
  CKNXD16 U1459 ( .I(n347), .ZN(AdrEna[717]) );
  CKBD0 U1460 ( .CLK(n205), .C(n349) );
  CKNXD16 U1461 ( .I(n349), .ZN(AdrEna[733]) );
  CKBD0 U1462 ( .CLK(n169), .C(n351) );
  CKNXD16 U1463 ( .I(n351), .ZN(AdrEna[637]) );
  CKBD0 U1464 ( .CLK(n175), .C(n353) );
  CKNXD16 U1465 ( .I(n353), .ZN(AdrEna[653]) );
  CKBD0 U1466 ( .CLK(n181), .C(n355) );
  CKNXD16 U1467 ( .I(n355), .ZN(AdrEna[669]) );
  CKBD0 U1468 ( .CLK(n187), .C(n357) );
  CKNXD16 U1469 ( .I(n357), .ZN(AdrEna[685]) );
  CKBD0 U1470 ( .CLK(n151), .C(n359) );
  CKNXD16 U1471 ( .I(n359), .ZN(AdrEna[589]) );
  CKBD0 U1472 ( .CLK(n157), .C(n361) );
  CKNXD16 U1473 ( .I(n361), .ZN(AdrEna[605]) );
  CKBD0 U1474 ( .CLK(n163), .C(n363) );
  CKNXD16 U1475 ( .I(n363), .ZN(AdrEna[621]) );
  CKBD0 U1476 ( .CLK(n127), .C(n365) );
  CKNXD16 U1477 ( .I(n365), .ZN(AdrEna[525]) );
  CKBD0 U1478 ( .CLK(n133), .C(n367) );
  CKNXD16 U1479 ( .I(n367), .ZN(AdrEna[541]) );
  CKBD0 U1480 ( .CLK(n139), .C(n369) );
  CKNXD16 U1481 ( .I(n369), .ZN(AdrEna[557]) );
  CKBD0 U1482 ( .CLK(n145), .C(n371) );
  CKNXD16 U1483 ( .I(n371), .ZN(AdrEna[573]) );
  CKBD0 U1484 ( .CLK(n204), .C(n373) );
  CKNXD16 U1485 ( .I(n373), .ZN(AdrEna[732]) );
  CKBD0 U1486 ( .CLK(n210), .C(n375) );
  CKNXD16 U1487 ( .I(n375), .ZN(AdrEna[748]) );
  CKBD0 U1488 ( .CLK(n216), .C(n377) );
  CKNXD16 U1489 ( .I(n377), .ZN(AdrEna[765]) );
  CKBD0 U1490 ( .CLK(n180), .C(n379) );
  CKNXD16 U1491 ( .I(n379), .ZN(AdrEna[668]) );
  CKBD0 U1492 ( .CLK(n186), .C(n381) );
  CKNXD16 U1493 ( .I(n381), .ZN(AdrEna[684]) );
  CKBD0 U1494 ( .CLK(n192), .C(n383) );
  CKNXD16 U1495 ( .I(n383), .ZN(AdrEna[700]) );
  CKBD0 U1496 ( .CLK(n198), .C(n385) );
  CKNXD16 U1497 ( .I(n385), .ZN(AdrEna[716]) );
  CKBD0 U1498 ( .CLK(n162), .C(n387) );
  CKNXD16 U1499 ( .I(n387), .ZN(AdrEna[620]) );
  CKBD0 U1500 ( .CLK(n168), .C(n389) );
  CKNXD16 U1501 ( .I(n389), .ZN(AdrEna[636]) );
  CKBD0 U1502 ( .CLK(n174), .C(n391) );
  CKNXD16 U1503 ( .I(n391), .ZN(AdrEna[652]) );
  CKBD0 U1504 ( .CLK(n138), .C(n393) );
  CKNXD16 U1505 ( .I(n393), .ZN(AdrEna[556]) );
  CKBD0 U1506 ( .CLK(n144), .C(n395) );
  CKNXD16 U1507 ( .I(n395), .ZN(AdrEna[572]) );
  CKBD0 U1508 ( .CLK(n150), .C(n397) );
  CKNXD16 U1509 ( .I(n397), .ZN(AdrEna[588]) );
  CKBD0 U1510 ( .CLK(n156), .C(n399) );
  CKNXD16 U1511 ( .I(n399), .ZN(AdrEna[604]) );
  CKBD0 U1512 ( .CLK(n215), .C(n401) );
  CKNXD16 U1513 ( .I(n401), .ZN(AdrEna[764]) );
  CKBD0 U1514 ( .CLK(n126), .C(n403) );
  CKNXD16 U1515 ( .I(n403), .ZN(AdrEna[524]) );
  CKBD0 U1516 ( .CLK(n132), .C(n405) );
  CKNXD16 U1517 ( .I(n405), .ZN(AdrEna[540]) );
  CKBD0 U1518 ( .CLK(n191), .C(n407) );
  CKNXD16 U1519 ( .I(n407), .ZN(AdrEna[699]) );
  CKBD0 U1520 ( .CLK(n197), .C(n409) );
  CKNXD16 U1521 ( .I(n409), .ZN(AdrEna[715]) );
  CKBD0 U1522 ( .CLK(n203), .C(n411) );
  CKNXD16 U1523 ( .I(n411), .ZN(AdrEna[731]) );
  CKBD0 U1524 ( .CLK(n209), .C(n413) );
  CKNXD16 U1525 ( .I(n413), .ZN(AdrEna[747]) );
  CKBD0 U1526 ( .CLK(n173), .C(n415) );
  CKNXD16 U1527 ( .I(n415), .ZN(AdrEna[651]) );
  CKBD0 U1528 ( .CLK(n179), .C(n417) );
  CKNXD16 U1529 ( .I(n417), .ZN(AdrEna[667]) );
  CKBD0 U1530 ( .CLK(n185), .C(n419) );
  CKNXD16 U1531 ( .I(n419), .ZN(AdrEna[683]) );
  CKBD0 U1532 ( .CLK(n149), .C(n421) );
  CKNXD16 U1533 ( .I(n421), .ZN(AdrEna[587]) );
  CKBD0 U1534 ( .CLK(n155), .C(n423) );
  CKNXD16 U1535 ( .I(n423), .ZN(AdrEna[603]) );
  CKBD0 U1536 ( .CLK(n161), .C(n425) );
  CKNXD16 U1537 ( .I(n425), .ZN(AdrEna[619]) );
  CKBD0 U1538 ( .CLK(n167), .C(n427) );
  CKNXD16 U1539 ( .I(n427), .ZN(AdrEna[635]) );
  CKBD0 U1540 ( .CLK(n131), .C(n429) );
  CKNXD16 U1541 ( .I(n429), .ZN(AdrEna[539]) );
  CKBD0 U1542 ( .CLK(n137), .C(n431) );
  CKNXD16 U1543 ( .I(n431), .ZN(AdrEna[555]) );
  CKBD0 U1544 ( .CLK(n143), .C(n433) );
  CKNXD16 U1545 ( .I(n433), .ZN(AdrEna[571]) );
  CKBD0 U1546 ( .CLK(n202), .C(n435) );
  CKNXD16 U1547 ( .I(n435), .ZN(AdrEna[730]) );
  CKBD0 U1548 ( .CLK(n208), .C(n437) );
  CKNXD16 U1549 ( .I(n437), .ZN(AdrEna[746]) );
  CKBD0 U1550 ( .CLK(n214), .C(n439) );
  CKNXD16 U1551 ( .I(n439), .ZN(AdrEna[763]) );
  CKBD0 U1552 ( .CLK(n125), .C(n441) );
  CKNXD16 U1553 ( .I(n441), .ZN(AdrEna[523]) );
  CKBD0 U1554 ( .CLK(n184), .C(n443) );
  CKNXD16 U1555 ( .I(n443), .ZN(AdrEna[682]) );
  CKBD0 U1556 ( .CLK(n190), .C(n445) );
  CKNXD16 U1557 ( .I(n445), .ZN(AdrEna[698]) );
  CKBD0 U1558 ( .CLK(n196), .C(n447) );
  CKNXD16 U1559 ( .I(n447), .ZN(AdrEna[714]) );
  CKBD0 U1560 ( .CLK(n160), .C(n449) );
  CKNXD16 U1561 ( .I(n449), .ZN(AdrEna[618]) );
  CKBD0 U1562 ( .CLK(n166), .C(n451) );
  CKNXD16 U1563 ( .I(n451), .ZN(AdrEna[634]) );
  CKBD0 U1564 ( .CLK(n172), .C(n453) );
  CKNXD16 U1565 ( .I(n453), .ZN(AdrEna[650]) );
  CKBD0 U1566 ( .CLK(n178), .C(n455) );
  CKNXD16 U1567 ( .I(n455), .ZN(AdrEna[666]) );
  CKBD0 U1568 ( .CLK(n142), .C(n457) );
  CKNXD16 U1569 ( .I(n457), .ZN(AdrEna[570]) );
  CKBD0 U1570 ( .CLK(n148), .C(n459) );
  CKNXD16 U1571 ( .I(n459), .ZN(AdrEna[586]) );
  CKBD0 U1572 ( .CLK(n154), .C(n461) );
  CKNXD16 U1573 ( .I(n461), .ZN(AdrEna[602]) );
  CKBD0 U1574 ( .CLK(n222), .C(n463) );
  CKNXD16 U1575 ( .I(n463), .ZN(AdrEna[959]) );
  CKBD0 U1576 ( .CLK(n124), .C(n465) );
  CKNXD16 U1577 ( .I(n465), .ZN(AdrEna[522]) );
  CKBD0 U1578 ( .CLK(n130), .C(n467) );
  CKNXD16 U1579 ( .I(n467), .ZN(AdrEna[538]) );
  CKBD0 U1580 ( .CLK(n136), .C(n469) );
  CKNXD16 U1581 ( .I(n469), .ZN(AdrEna[554]) );
  CKBD0 U1582 ( .CLK(n123), .C(n471) );
  CKNXD16 U1583 ( .I(n471), .ZN(AdrEna[255]) );
  CKBD0 U1584 ( .CLK(n220), .C(n473) );
  CKNXD16 U1585 ( .I(n473), .ZN(AdrEna[927]) );
  CKBD0 U1586 ( .CLK(n221), .C(n475) );
  CKNXD16 U1587 ( .I(n475), .ZN(AdrEna[943]) );
  CKBD0 U1588 ( .CLK(n111), .C(n477) );
  CKNXD16 U1589 ( .I(n477), .ZN(AdrEna[191]) );
  CKBD0 U1590 ( .CLK(n114), .C(n479) );
  CKNXD16 U1591 ( .I(n479), .ZN(AdrEna[207]) );
  CKBD0 U1592 ( .CLK(n117), .C(n481) );
  CKNXD16 U1593 ( .I(n481), .ZN(AdrEna[223]) );
  CKBD0 U1594 ( .CLK(n120), .C(n483) );
  CKNXD16 U1595 ( .I(n483), .ZN(AdrEna[239]) );
  CKBD0 U1596 ( .CLK(n100), .C(n485) );
  CKNXD16 U1597 ( .I(n485), .ZN(AdrEna[143]) );
  CKBD0 U1598 ( .CLK(n104), .C(n487) );
  CKNXD16 U1599 ( .I(n487), .ZN(AdrEna[159]) );
  CKBD0 U1600 ( .CLK(n108), .C(n489) );
  CKNXD16 U1601 ( .I(n489), .ZN(AdrEna[175]) );
  CKBD0 U1602 ( .CLK(n84), .C(n491) );
  CKNXD16 U1603 ( .I(n491), .ZN(AdrEna[79]) );
  CKBD0 U1604 ( .CLK(n88), .C(n493) );
  CKNXD16 U1605 ( .I(n493), .ZN(AdrEna[95]) );
  CKBD0 U1606 ( .CLK(n92), .C(n495) );
  CKNXD16 U1607 ( .I(n495), .ZN(AdrEna[111]) );
  CKBD0 U1608 ( .CLK(n96), .C(n497) );
  CKNXD16 U1609 ( .I(n497), .ZN(AdrEna[127]) );
  CKBD0 U1610 ( .CLK(n72), .C(n499) );
  CKNXD16 U1611 ( .I(n499), .ZN(AdrEna[31]) );
  CKBD0 U1612 ( .CLK(n76), .C(n501) );
  CKNXD16 U1613 ( .I(n501), .ZN(AdrEna[47]) );
  CKBD0 U1614 ( .CLK(n80), .C(n503) );
  CKNXD16 U1615 ( .I(n503), .ZN(AdrEna[63]) );
  CKBD0 U1616 ( .CLK(n116), .C(n505) );
  CKNXD16 U1617 ( .I(n505), .ZN(AdrEna[222]) );
  CKBD0 U1618 ( .CLK(n119), .C(n507) );
  CKNXD16 U1619 ( .I(n507), .ZN(AdrEna[238]) );
  CKBD0 U1620 ( .CLK(n122), .C(n509) );
  CKNXD16 U1621 ( .I(n509), .ZN(AdrEna[254]) );
  CKBD0 U1622 ( .CLK(n68), .C(n511) );
  CKNXD16 U1623 ( .I(n511), .ZN(AdrEna[15]) );
  CKBD0 U1624 ( .CLK(n107), .C(n513) );
  CKNXD16 U1625 ( .I(n513), .ZN(AdrEna[174]) );
  CKBD0 U1626 ( .CLK(n110), .C(n515) );
  CKNXD16 U1627 ( .I(n515), .ZN(AdrEna[190]) );
  CKBD0 U1628 ( .CLK(n113), .C(n517) );
  CKNXD16 U1629 ( .I(n517), .ZN(AdrEna[206]) );
  CKBD0 U1630 ( .CLK(n91), .C(n519) );
  CKNXD16 U1631 ( .I(n519), .ZN(AdrEna[110]) );
  CKBD0 U1632 ( .CLK(n95), .C(n521) );
  CKNXD16 U1633 ( .I(n521), .ZN(AdrEna[126]) );
  CKBD0 U1634 ( .CLK(n99), .C(n523) );
  CKNXD16 U1635 ( .I(n523), .ZN(AdrEna[142]) );
  CKBD0 U1636 ( .CLK(n103), .C(n525) );
  CKNXD16 U1637 ( .I(n525), .ZN(AdrEna[158]) );
  CKBD0 U1638 ( .CLK(n79), .C(n527) );
  CKNXD16 U1639 ( .I(n527), .ZN(AdrEna[62]) );
  CKBD0 U1640 ( .CLK(n83), .C(n529) );
  CKNXD16 U1641 ( .I(n529), .ZN(AdrEna[78]) );
  CKBD0 U1642 ( .CLK(n87), .C(n531) );
  CKNXD16 U1643 ( .I(n531), .ZN(AdrEna[94]) );
  CKBD0 U1644 ( .CLK(n121), .C(n533) );
  CKNXD16 U1645 ( .I(n533), .ZN(AdrEna[253]) );
  CKBD0 U1646 ( .CLK(n67), .C(n535) );
  CKNXD16 U1647 ( .I(n535), .ZN(AdrEna[14]) );
  CKBD0 U1648 ( .CLK(n71), .C(n537) );
  CKNXD16 U1649 ( .I(n537), .ZN(AdrEna[30]) );
  CKBD0 U1650 ( .CLK(n75), .C(n539) );
  CKNXD16 U1651 ( .I(n539), .ZN(AdrEna[46]) );
  CKBD0 U1652 ( .CLK(n112), .C(n541) );
  CKNXD16 U1653 ( .I(n541), .ZN(AdrEna[205]) );
  CKBD0 U1654 ( .CLK(n115), .C(n543) );
  CKNXD16 U1655 ( .I(n543), .ZN(AdrEna[221]) );
  CKBD0 U1656 ( .CLK(n118), .C(n545) );
  CKNXD16 U1657 ( .I(n545), .ZN(AdrEna[237]) );
  CKBD0 U1658 ( .CLK(n98), .C(n547) );
  CKNXD16 U1659 ( .I(n547), .ZN(AdrEna[141]) );
  CKBD0 U1660 ( .CLK(n102), .C(n549) );
  CKNXD16 U1661 ( .I(n549), .ZN(AdrEna[157]) );
  CKBD0 U1662 ( .CLK(n106), .C(n551) );
  CKNXD16 U1663 ( .I(n551), .ZN(AdrEna[173]) );
  CKBD0 U1664 ( .CLK(n109), .C(n553) );
  CKNXD16 U1665 ( .I(n553), .ZN(AdrEna[189]) );
  CKBD0 U1666 ( .CLK(n86), .C(n555) );
  CKNXD16 U1667 ( .I(n555), .ZN(AdrEna[93]) );
  CKBD0 U1668 ( .CLK(n90), .C(n557) );
  CKNXD16 U1669 ( .I(n557), .ZN(AdrEna[109]) );
  CKBD0 U1670 ( .CLK(n94), .C(n559) );
  CKNXD16 U1671 ( .I(n559), .ZN(AdrEna[125]) );
  CKBD0 U1672 ( .CLK(n70), .C(n561) );
  CKNXD16 U1673 ( .I(n561), .ZN(AdrEna[29]) );
  CKBD0 U1674 ( .CLK(n74), .C(n563) );
  CKNXD16 U1675 ( .I(n563), .ZN(AdrEna[45]) );
  CKBD0 U1676 ( .CLK(n78), .C(n565) );
  CKNXD16 U1677 ( .I(n565), .ZN(AdrEna[61]) );
  CKBD0 U1678 ( .CLK(n82), .C(n567) );
  CKNXD16 U1679 ( .I(n567), .ZN(AdrEna[77]) );
  CKBD0 U1680 ( .CLK(n97), .C(n569) );
  CKNXD16 U1681 ( .I(n569), .ZN(AdrEna[139]) );
  CKBD0 U1682 ( .CLK(n101), .C(n571) );
  CKNXD16 U1683 ( .I(n571), .ZN(AdrEna[155]) );
  CKBD0 U1684 ( .CLK(n105), .C(n573) );
  CKNXD16 U1685 ( .I(n573), .ZN(AdrEna[171]) );
  CKBD0 U1686 ( .CLK(n81), .C(n575) );
  CKNXD16 U1687 ( .I(n575), .ZN(AdrEna[75]) );
  CKBD0 U1688 ( .CLK(n85), .C(n577) );
  CKNXD16 U1689 ( .I(n577), .ZN(AdrEna[91]) );
  CKBD0 U1690 ( .CLK(n89), .C(n579) );
  CKNXD16 U1691 ( .I(n579), .ZN(AdrEna[107]) );
  CKBD0 U1692 ( .CLK(n93), .C(n581) );
  CKNXD16 U1693 ( .I(n581), .ZN(AdrEna[123]) );
  CKBD0 U1694 ( .CLK(n219), .C(n583) );
  CKNXD16 U1695 ( .I(n583), .ZN(AdrEna[815]) );
  CKBD0 U1696 ( .CLK(n77), .C(n585) );
  CKNXD16 U1697 ( .I(n585), .ZN(AdrEna[59]) );
  CKND2D0 U1698 ( .A1(\DL3[40].tempL3[5] ), .A2(n28), .ZN(n587) );
  CKNXD16 U1699 ( .I(n587), .ZN(AdrEna[645]) );
  CKND2D0 U1700 ( .A1(\DL3[40].tempL3[6] ), .A2(n28), .ZN(n589) );
  CKNXD16 U1701 ( .I(n589), .ZN(AdrEna[646]) );
  CKND2D0 U1702 ( .A1(\DL3[31].tempL3[0] ), .A2(n38), .ZN(n591) );
  CKNXD16 U1703 ( .I(n591), .ZN(AdrEna[496]) );
  CKND2D0 U1704 ( .A1(\DL3[40].tempL3[7] ), .A2(n28), .ZN(n593) );
  CKNXD16 U1705 ( .I(n593), .ZN(AdrEna[647]) );
  CKND2D0 U1706 ( .A1(\DL3[31].tempL3[6] ), .A2(n38), .ZN(n595) );
  CKNXD16 U1707 ( .I(n595), .ZN(AdrEna[502]) );
  CKND2D0 U1708 ( .A1(\DL3[60].tempL3[15] ), .A2(n6), .ZN(n597) );
  CKNXD16 U1709 ( .I(n597), .ZN(AdrEna[975]) );
  CKND2D0 U1710 ( .A1(\DL3[63].tempL3[6] ), .A2(n65), .ZN(n599) );
  CKNXD16 U1711 ( .I(n599), .ZN(AdrEna[1014]) );
  CKND2D0 U1712 ( .A1(\DL3[47].tempL3[2] ), .A2(n21), .ZN(n601) );
  CKNXD16 U1713 ( .I(n601), .ZN(AdrEna[754]) );
  CKND2D0 U1714 ( .A1(\DL3[57].tempL3[9] ), .A2(n10), .ZN(n603) );
  CKNXD16 U1715 ( .I(n603), .ZN(AdrEna[921]) );
  CKND2D0 U1716 ( .A1(\DL3[31].tempL3[7] ), .A2(n38), .ZN(n605) );
  CKNXD16 U1717 ( .I(n605), .ZN(AdrEna[503]) );
  CKND2D0 U1718 ( .A1(\DL3[59].tempL3[8] ), .A2(n8), .ZN(n607) );
  CKNXD16 U1719 ( .I(n607), .ZN(AdrEna[952]) );
  CKND2D0 U1720 ( .A1(\DL3[31].tempL3[8] ), .A2(n38), .ZN(n609) );
  CKNXD16 U1721 ( .I(n609), .ZN(AdrEna[504]) );
  CKND2D0 U1722 ( .A1(\DL3[31].tempL3[10] ), .A2(n38), .ZN(n611) );
  CKNXD16 U1723 ( .I(n611), .ZN(AdrEna[506]) );
  CKND2D0 U1724 ( .A1(\DL3[63].tempL3[14] ), .A2(n65), .ZN(n613) );
  CKNXD16 U1725 ( .I(n613), .ZN(AdrEna[1022]) );
  CKND2D0 U1726 ( .A1(\DL3[55].tempL3[6] ), .A2(n12), .ZN(n615) );
  CKNXD16 U1727 ( .I(n615), .ZN(AdrEna[886]) );
  CKND2D0 U1728 ( .A1(\DL3[39].tempL3[7] ), .A2(n30), .ZN(n617) );
  CKNXD16 U1729 ( .I(n617), .ZN(AdrEna[631]) );
  CKND2D0 U1730 ( .A1(\DL3[39].tempL3[6] ), .A2(n30), .ZN(n619) );
  CKNXD16 U1731 ( .I(n619), .ZN(AdrEna[630]) );
  CKND2D0 U1732 ( .A1(\DL3[31].tempL3[11] ), .A2(n38), .ZN(n621) );
  CKNXD16 U1733 ( .I(n621), .ZN(AdrEna[507]) );
  CKND2D0 U1734 ( .A1(\DL3[30].tempL3[6] ), .A2(n39), .ZN(n623) );
  CKNXD16 U1735 ( .I(n623), .ZN(AdrEna[486]) );
  CKND2D0 U1736 ( .A1(\DL3[47].tempL3[6] ), .A2(n21), .ZN(n625) );
  CKNXD16 U1737 ( .I(n625), .ZN(AdrEna[758]) );
  CKND2D0 U1738 ( .A1(\DL3[31].tempL3[15] ), .A2(n38), .ZN(n627) );
  CKNXD16 U1739 ( .I(n627), .ZN(AdrEna[511]) );
  CKND2D0 U1740 ( .A1(\DL3[31].tempL3[14] ), .A2(n38), .ZN(n629) );
  CKNXD16 U1741 ( .I(n629), .ZN(AdrEna[510]) );
  CKND2D0 U1742 ( .A1(\DL3[46].tempL3[7] ), .A2(n22), .ZN(n631) );
  CKNXD16 U1743 ( .I(n631), .ZN(AdrEna[743]) );
  CKND2D0 U1744 ( .A1(\DL3[46].tempL3[5] ), .A2(n22), .ZN(n633) );
  CKNXD16 U1745 ( .I(n633), .ZN(AdrEna[741]) );
  CKND2D0 U1746 ( .A1(\DL3[39].tempL3[2] ), .A2(n30), .ZN(n635) );
  CKNXD16 U1747 ( .I(n635), .ZN(AdrEna[626]) );
  CKND2D0 U1748 ( .A1(\DL3[58].tempL3[2] ), .A2(n9), .ZN(n637) );
  CKNXD16 U1749 ( .I(n637), .ZN(AdrEna[930]) );
  CKND2D0 U1750 ( .A1(\DL3[57].tempL3[6] ), .A2(n10), .ZN(n639) );
  CKNXD16 U1751 ( .I(n639), .ZN(AdrEna[918]) );
  CKND2D0 U1752 ( .A1(\DL3[47].tempL3[9] ), .A2(n21), .ZN(n641) );
  CKNXD16 U1753 ( .I(n641), .ZN(AdrEna[761]) );
  CKND2D0 U1754 ( .A1(\DL3[41].tempL3[6] ), .A2(n27), .ZN(n643) );
  CKNXD16 U1755 ( .I(n643), .ZN(AdrEna[662]) );
  CKND2D0 U1756 ( .A1(\DL3[61].tempL3[15] ), .A2(n5), .ZN(n645) );
  CKNXD16 U1757 ( .I(n645), .ZN(AdrEna[991]) );
  CKND2D0 U1758 ( .A1(\DL3[59].tempL3[6] ), .A2(n8), .ZN(n647) );
  CKNXD16 U1759 ( .I(n647), .ZN(AdrEna[950]) );
  CKND2D0 U1760 ( .A1(\DL3[46].tempL3[6] ), .A2(n22), .ZN(n649) );
  CKNXD16 U1761 ( .I(n649), .ZN(AdrEna[742]) );
  CKND2D0 U1762 ( .A1(\DL3[38].tempL3[6] ), .A2(n31), .ZN(n651) );
  CKNXD16 U1763 ( .I(n651), .ZN(AdrEna[614]) );
  CKND2D0 U1764 ( .A1(\DL3[41].tempL3[5] ), .A2(n27), .ZN(n653) );
  CKNXD16 U1765 ( .I(n653), .ZN(AdrEna[661]) );
  AN2D1 U1766 ( .A1(\DL2[2].tempL2[6] ), .A2(DecodedL1[2]), .Z(n31) );
  CKND2D0 U1767 ( .A1(\DL3[38].tempL3[7] ), .A2(n31), .ZN(n655) );
  CKNXD16 U1768 ( .I(n655), .ZN(AdrEna[615]) );
  CKND2D0 U1769 ( .A1(\DL3[41].tempL3[7] ), .A2(n27), .ZN(n657) );
  CKNXD16 U1770 ( .I(n657), .ZN(AdrEna[663]) );
  CKND2D0 U1771 ( .A1(\DL3[53].tempL3[6] ), .A2(n14), .ZN(n659) );
  CKNXD16 U1772 ( .I(n659), .ZN(AdrEna[854]) );
  CKND2D0 U1773 ( .A1(\DL3[61].tempL3[7] ), .A2(n5), .ZN(n661) );
  CKNXD16 U1774 ( .I(n661), .ZN(AdrEna[983]) );
  CKND2D0 U1775 ( .A1(\DL3[38].tempL3[3] ), .A2(n31), .ZN(n663) );
  CKNXD16 U1776 ( .I(n663), .ZN(AdrEna[611]) );
  CKND2D0 U1777 ( .A1(\DL3[38].tempL3[5] ), .A2(n31), .ZN(n665) );
  CKNXD16 U1778 ( .I(n665), .ZN(AdrEna[613]) );
  CKND2D0 U1779 ( .A1(\DL3[29].tempL3[7] ), .A2(n41), .ZN(n667) );
  CKNXD16 U1780 ( .I(n667), .ZN(AdrEna[471]) );
  CKND2D0 U1781 ( .A1(\DL3[63].tempL3[7] ), .A2(n65), .ZN(n669) );
  CKNXD16 U1782 ( .I(n669), .ZN(AdrEna[1015]) );
  CKND2D0 U1783 ( .A1(\DL3[29].tempL3[6] ), .A2(n41), .ZN(n671) );
  CKNXD16 U1784 ( .I(n671), .ZN(AdrEna[470]) );
  CKND2D0 U1785 ( .A1(\DL3[63].tempL3[15] ), .A2(n65), .ZN(n673) );
  CKNXD16 U1786 ( .I(n673), .ZN(AdrEna[1023]) );
  CKND2D0 U1787 ( .A1(\DL3[61].tempL3[13] ), .A2(n5), .ZN(n675) );
  CKNXD16 U1788 ( .I(n675), .ZN(AdrEna[989]) );
  CKND2D0 U1789 ( .A1(\DL3[42].tempL3[2] ), .A2(n26), .ZN(n677) );
  CKNXD16 U1790 ( .I(n677), .ZN(AdrEna[674]) );
  CKND2D0 U1791 ( .A1(\DL3[38].tempL3[2] ), .A2(n31), .ZN(n679) );
  CKNXD16 U1792 ( .I(n679), .ZN(AdrEna[610]) );
  CKND2D0 U1793 ( .A1(\DL3[60].tempL3[13] ), .A2(n6), .ZN(n681) );
  CKNXD16 U1794 ( .I(n681), .ZN(AdrEna[973]) );
  CKND2D0 U1795 ( .A1(\DL3[59].tempL3[2] ), .A2(n8), .ZN(n683) );
  CKNXD16 U1796 ( .I(n683), .ZN(AdrEna[946]) );
  CKND2D0 U1797 ( .A1(\DL3[42].tempL3[7] ), .A2(n26), .ZN(n685) );
  CKNXD16 U1798 ( .I(n685), .ZN(AdrEna[679]) );
  CKND2D0 U1799 ( .A1(\DL3[52].tempL3[6] ), .A2(n15), .ZN(n687) );
  CKNXD16 U1800 ( .I(n687), .ZN(AdrEna[838]) );
  CKND2D0 U1801 ( .A1(\DL3[42].tempL3[6] ), .A2(n26), .ZN(n689) );
  CKNXD16 U1802 ( .I(n689), .ZN(AdrEna[678]) );
  CKND2D0 U1803 ( .A1(\DL3[58].tempL3[6] ), .A2(n9), .ZN(n691) );
  CKNXD16 U1804 ( .I(n691), .ZN(AdrEna[934]) );
  CKND2D0 U1805 ( .A1(\DL3[63].tempL3[11] ), .A2(n65), .ZN(n693) );
  CKNXD16 U1806 ( .I(n693), .ZN(AdrEna[1019]) );
  CKND2D0 U1807 ( .A1(\DL3[6].tempL3[9] ), .A2(n3), .ZN(n695) );
  CKNXD16 U1808 ( .I(n695), .ZN(AdrEna[105]) );
  CKND2D0 U1809 ( .A1(\DL3[26].tempL3[6] ), .A2(n44), .ZN(n697) );
  CKNXD16 U1810 ( .I(n697), .ZN(AdrEna[422]) );
  CKND2D0 U1811 ( .A1(\DL3[2].tempL3[9] ), .A2(n40), .ZN(n699) );
  CKNXD16 U1812 ( .I(n699), .ZN(AdrEna[41]) );
  CKND2D0 U1813 ( .A1(\DL3[42].tempL3[9] ), .A2(n26), .ZN(n701) );
  CKNXD16 U1814 ( .I(n701), .ZN(AdrEna[681]) );
  CKND2D0 U1815 ( .A1(\DL3[23].tempL3[13] ), .A2(n47), .ZN(n703) );
  CKNXD16 U1816 ( .I(n703), .ZN(AdrEna[381]) );
  CKND2D0 U1817 ( .A1(\DL3[62].tempL3[13] ), .A2(n4), .ZN(n705) );
  CKNXD16 U1818 ( .I(n705), .ZN(AdrEna[1005]) );
  CKND2D0 U1819 ( .A1(\DL3[58].tempL3[8] ), .A2(n9), .ZN(n707) );
  CKNXD16 U1820 ( .I(n707), .ZN(AdrEna[936]) );
  CKND2D0 U1821 ( .A1(\DL3[43].tempL3[5] ), .A2(n25), .ZN(n709) );
  CKNXD16 U1822 ( .I(n709), .ZN(AdrEna[693]) );
  CKND2D0 U1823 ( .A1(\DL3[8].tempL3[9] ), .A2(n63), .ZN(n711) );
  CKNXD16 U1824 ( .I(n711), .ZN(AdrEna[137]) );
  CKND2D0 U1825 ( .A1(\DL3[9].tempL3[9] ), .A2(n62), .ZN(n713) );
  CKNXD16 U1826 ( .I(n713), .ZN(AdrEna[153]) );
  CKND2D0 U1827 ( .A1(\DL3[15].tempL3[6] ), .A2(n56), .ZN(n715) );
  CKNXD16 U1828 ( .I(n715), .ZN(AdrEna[246]) );
  CKND2D0 U1829 ( .A1(\DL3[43].tempL3[6] ), .A2(n25), .ZN(n717) );
  CKNXD16 U1830 ( .I(n717), .ZN(AdrEna[694]) );
  CKND2D0 U1831 ( .A1(\DL3[28].tempL3[6] ), .A2(n42), .ZN(n719) );
  CKNXD16 U1832 ( .I(n719), .ZN(AdrEna[454]) );
  CKND2D0 U1833 ( .A1(\DL3[56].tempL3[6] ), .A2(n11), .ZN(n721) );
  CKNXD16 U1834 ( .I(n721), .ZN(AdrEna[902]) );
  CKND2D0 U1835 ( .A1(\DL3[56].tempL3[9] ), .A2(n11), .ZN(n723) );
  CKNXD16 U1836 ( .I(n723), .ZN(AdrEna[905]) );
  CKND2D0 U1837 ( .A1(\DL3[43].tempL3[7] ), .A2(n25), .ZN(n725) );
  CKNXD16 U1838 ( .I(n725), .ZN(AdrEna[695]) );
  CKND2D0 U1839 ( .A1(\DL3[13].tempL3[6] ), .A2(n58), .ZN(n727) );
  CKNXD16 U1840 ( .I(n727), .ZN(AdrEna[214]) );
  CKND2D0 U1841 ( .A1(\DL3[11].tempL3[9] ), .A2(n60), .ZN(n729) );
  CKNXD16 U1842 ( .I(n729), .ZN(AdrEna[185]) );
  CKND2D0 U1843 ( .A1(\DL3[21].tempL3[6] ), .A2(n49), .ZN(n731) );
  CKNXD16 U1844 ( .I(n731), .ZN(AdrEna[342]) );
  CKND2D0 U1845 ( .A1(\DL3[44].tempL3[2] ), .A2(n24), .ZN(n733) );
  CKNXD16 U1846 ( .I(n733), .ZN(AdrEna[706]) );
  CKND2D0 U1847 ( .A1(\DL3[25].tempL3[7] ), .A2(n45), .ZN(n735) );
  CKNXD16 U1848 ( .I(n735), .ZN(AdrEna[407]) );
  CKND2D0 U1849 ( .A1(\DL3[63].tempL3[10] ), .A2(n65), .ZN(n737) );
  CKNXD16 U1850 ( .I(n737), .ZN(AdrEna[1018]) );
  CKND2D0 U1851 ( .A1(\DL3[44].tempL3[5] ), .A2(n24), .ZN(n739) );
  CKNXD16 U1852 ( .I(n739), .ZN(AdrEna[709]) );
  CKND2D0 U1853 ( .A1(\DL3[44].tempL3[3] ), .A2(n24), .ZN(n741) );
  CKNXD16 U1854 ( .I(n741), .ZN(AdrEna[707]) );
  CKND2D0 U1855 ( .A1(\DL3[25].tempL3[6] ), .A2(n45), .ZN(n743) );
  CKNXD16 U1856 ( .I(n743), .ZN(AdrEna[406]) );
  CKND2D0 U1857 ( .A1(\DL3[23].tempL3[6] ), .A2(n47), .ZN(n745) );
  CKNXD16 U1858 ( .I(n745), .ZN(AdrEna[374]) );
  CKND2D0 U1859 ( .A1(\DL3[9].tempL3[5] ), .A2(n62), .ZN(n747) );
  CKNXD16 U1860 ( .I(n747), .ZN(AdrEna[149]) );
  CKND2D0 U1861 ( .A1(\DL3[51].tempL3[11] ), .A2(n16), .ZN(n749) );
  CKNXD16 U1862 ( .I(n749), .ZN(AdrEna[827]) );
  CKND2D0 U1863 ( .A1(\DL3[10].tempL3[9] ), .A2(n61), .ZN(n751) );
  CKNXD16 U1864 ( .I(n751), .ZN(AdrEna[169]) );
  CKND2D0 U1865 ( .A1(\DL3[44].tempL3[6] ), .A2(n24), .ZN(n753) );
  CKNXD16 U1866 ( .I(n753), .ZN(AdrEna[710]) );
  CKND2D0 U1867 ( .A1(\DL3[44].tempL3[7] ), .A2(n24), .ZN(n755) );
  CKNXD16 U1868 ( .I(n755), .ZN(AdrEna[711]) );
  CKND2D0 U1869 ( .A1(\DL3[61].tempL3[14] ), .A2(n5), .ZN(n757) );
  CKNXD16 U1870 ( .I(n757), .ZN(AdrEna[990]) );
  CKND2D0 U1871 ( .A1(\DL3[14].tempL3[6] ), .A2(n57), .ZN(n759) );
  CKNXD16 U1872 ( .I(n759), .ZN(AdrEna[230]) );
  CKND2D0 U1873 ( .A1(\DL3[1].tempL3[9] ), .A2(n51), .ZN(n761) );
  CKNXD16 U1874 ( .I(n761), .ZN(AdrEna[25]) );
  CKND2D0 U1875 ( .A1(\DL3[19].tempL3[6] ), .A2(n52), .ZN(n763) );
  CKNXD16 U1876 ( .I(n763), .ZN(AdrEna[310]) );
  CKND2D0 U1877 ( .A1(\DL3[60].tempL3[11] ), .A2(n6), .ZN(n765) );
  CKNXD16 U1878 ( .I(n765), .ZN(AdrEna[971]) );
  CKND2D0 U1879 ( .A1(\DL3[27].tempL3[7] ), .A2(n43), .ZN(n767) );
  CKNXD16 U1880 ( .I(n767), .ZN(AdrEna[439]) );
  CKND2D0 U1881 ( .A1(\DL3[60].tempL3[14] ), .A2(n6), .ZN(n769) );
  CKNXD16 U1882 ( .I(n769), .ZN(AdrEna[974]) );
  CKND2D0 U1883 ( .A1(\DL3[36].tempL3[6] ), .A2(n33), .ZN(n771) );
  CKNXD16 U1884 ( .I(n771), .ZN(AdrEna[582]) );
  CKND2D0 U1885 ( .A1(\DL3[36].tempL3[5] ), .A2(n33), .ZN(n773) );
  CKNXD16 U1886 ( .I(n773), .ZN(AdrEna[581]) );
  CKND2D0 U1887 ( .A1(\DL3[7].tempL3[9] ), .A2(n64), .ZN(n775) );
  CKNXD16 U1888 ( .I(n775), .ZN(AdrEna[121]) );
  CKND2D0 U1889 ( .A1(\DL3[27].tempL3[6] ), .A2(n43), .ZN(n777) );
  CKNXD16 U1890 ( .I(n777), .ZN(AdrEna[438]) );
  CKND2D0 U1891 ( .A1(\DL3[4].tempL3[9] ), .A2(n18), .ZN(n779) );
  CKNXD16 U1892 ( .I(n779), .ZN(AdrEna[73]) );
  CKND2D0 U1893 ( .A1(\DL3[36].tempL3[7] ), .A2(n33), .ZN(n781) );
  CKNXD16 U1894 ( .I(n781), .ZN(AdrEna[583]) );
  CKND2D0 U1895 ( .A1(\DL3[11].tempL3[8] ), .A2(n60), .ZN(n783) );
  CKNXD16 U1896 ( .I(n783), .ZN(AdrEna[184]) );
  CKND2D0 U1897 ( .A1(\DL3[54].tempL3[6] ), .A2(n13), .ZN(n785) );
  CKNXD16 U1898 ( .I(n785), .ZN(AdrEna[870]) );
  CKND2D0 U1899 ( .A1(\DL3[45].tempL3[6] ), .A2(n23), .ZN(n787) );
  CKNXD16 U1900 ( .I(n787), .ZN(AdrEna[726]) );
  CKND2D0 U1901 ( .A1(\DL3[62].tempL3[15] ), .A2(n4), .ZN(n789) );
  CKNXD16 U1902 ( .I(n789), .ZN(AdrEna[1007]) );
  CKND2D0 U1903 ( .A1(\DL3[12].tempL3[6] ), .A2(n59), .ZN(n791) );
  CKNXD16 U1904 ( .I(n791), .ZN(AdrEna[198]) );
  CKND2D0 U1905 ( .A1(\DL3[5].tempL3[9] ), .A2(n7), .ZN(n793) );
  CKNXD16 U1906 ( .I(n793), .ZN(AdrEna[89]) );
  CKND2D0 U1907 ( .A1(\DL3[17].tempL3[6] ), .A2(n54), .ZN(n795) );
  CKNXD16 U1908 ( .I(n795), .ZN(AdrEna[278]) );
  CKND2D0 U1909 ( .A1(\DL3[37].tempL3[2] ), .A2(n32), .ZN(n797) );
  CKNXD16 U1910 ( .I(n797), .ZN(AdrEna[594]) );
  CKND2D0 U1911 ( .A1(\DL3[22].tempL3[6] ), .A2(n48), .ZN(n799) );
  CKNXD16 U1912 ( .I(n799), .ZN(AdrEna[358]) );
  CKND2D0 U1913 ( .A1(\DL3[63].tempL3[2] ), .A2(n65), .ZN(n801) );
  CKNXD16 U1914 ( .I(n801), .ZN(AdrEna[1010]) );
  CKND2D0 U1915 ( .A1(\DL3[37].tempL3[6] ), .A2(n32), .ZN(n803) );
  CKNXD16 U1916 ( .I(n803), .ZN(AdrEna[598]) );
  CKND2D0 U1917 ( .A1(\DL3[45].tempL3[7] ), .A2(n23), .ZN(n805) );
  CKNXD16 U1918 ( .I(n805), .ZN(AdrEna[727]) );
  CKND2D0 U1919 ( .A1(\DL3[24].tempL3[6] ), .A2(n46), .ZN(n807) );
  CKNXD16 U1920 ( .I(n807), .ZN(AdrEna[390]) );
  CKND2D0 U1921 ( .A1(\DL3[20].tempL3[6] ), .A2(n50), .ZN(n809) );
  CKNXD16 U1922 ( .I(n809), .ZN(AdrEna[326]) );
  CKND2D0 U1923 ( .A1(\DL3[3].tempL3[9] ), .A2(n29), .ZN(n811) );
  CKNXD16 U1924 ( .I(n811), .ZN(AdrEna[57]) );
  CKND2D0 U1925 ( .A1(\DL3[37].tempL3[7] ), .A2(n32), .ZN(n813) );
  CKNXD16 U1926 ( .I(n813), .ZN(AdrEna[599]) );
  CKND2D0 U1927 ( .A1(\DL3[51].tempL3[3] ), .A2(n16), .ZN(n815) );
  CKNXD16 U1928 ( .I(n815), .ZN(AdrEna[819]) );
  CKND2D0 U1929 ( .A1(\DL3[51].tempL3[2] ), .A2(n16), .ZN(n817) );
  CKNXD16 U1930 ( .I(n817), .ZN(AdrEna[818]) );
  CKND2D0 U1931 ( .A1(\DL3[45].tempL3[9] ), .A2(n23), .ZN(n819) );
  CKNXD16 U1932 ( .I(n819), .ZN(AdrEna[729]) );
  CKND2D0 U1933 ( .A1(\DL3[18].tempL3[6] ), .A2(n53), .ZN(n821) );
  CKNXD16 U1934 ( .I(n821), .ZN(AdrEna[294]) );
  CKND2D0 U1935 ( .A1(\DL3[51].tempL3[5] ), .A2(n16), .ZN(n823) );
  CKNXD16 U1936 ( .I(n823), .ZN(AdrEna[821]) );
  CKND2D0 U1937 ( .A1(\DL3[41].tempL3[4] ), .A2(n27), .ZN(n825) );
  CKNXD16 U1938 ( .I(n825), .ZN(AdrEna[660]) );
  CKND2D0 U1939 ( .A1(\DL3[51].tempL3[7] ), .A2(n16), .ZN(n827) );
  CKNXD16 U1940 ( .I(n827), .ZN(AdrEna[823]) );
  CKND2D0 U1941 ( .A1(\DL3[30].tempL3[14] ), .A2(n39), .ZN(n829) );
  CKNXD16 U1942 ( .I(n829), .ZN(AdrEna[494]) );
  CKND2D0 U1943 ( .A1(\DL3[51].tempL3[4] ), .A2(n16), .ZN(n831) );
  CKNXD16 U1944 ( .I(n831), .ZN(AdrEna[820]) );
  CKND2D0 U1945 ( .A1(\DL3[51].tempL3[6] ), .A2(n16), .ZN(n833) );
  CKNXD16 U1946 ( .I(n833), .ZN(AdrEna[822]) );
  CKND2D0 U1947 ( .A1(\DL3[51].tempL3[13] ), .A2(n16), .ZN(n835) );
  CKNXD16 U1948 ( .I(n835), .ZN(AdrEna[829]) );
  CKND2D0 U1949 ( .A1(\DL3[51].tempL3[10] ), .A2(n16), .ZN(n837) );
  CKNXD16 U1950 ( .I(n837), .ZN(AdrEna[826]) );
  CKND2D0 U1951 ( .A1(\DL3[51].tempL3[12] ), .A2(n16), .ZN(n839) );
  CKNXD16 U1952 ( .I(n839), .ZN(AdrEna[828]) );
  CKND2D0 U1953 ( .A1(\DL3[51].tempL3[8] ), .A2(n16), .ZN(n841) );
  CKNXD16 U1954 ( .I(n841), .ZN(AdrEna[824]) );
  CKND2D0 U1955 ( .A1(\DL3[11].tempL3[10] ), .A2(n60), .ZN(n843) );
  CKNXD16 U1956 ( .I(n843), .ZN(AdrEna[186]) );
  CKND2D0 U1957 ( .A1(\DL3[51].tempL3[15] ), .A2(n16), .ZN(n845) );
  CKNXD16 U1958 ( .I(n845), .ZN(AdrEna[831]) );
  CKND2D0 U1959 ( .A1(\DL3[11].tempL3[11] ), .A2(n60), .ZN(n847) );
  CKNXD16 U1960 ( .I(n847), .ZN(AdrEna[187]) );
  CKND2D0 U1961 ( .A1(\DL3[51].tempL3[0] ), .A2(n16), .ZN(n849) );
  CKNXD16 U1962 ( .I(n849), .ZN(AdrEna[816]) );
  CKND2D0 U1963 ( .A1(\DL3[51].tempL3[14] ), .A2(n16), .ZN(n851) );
  CKNXD16 U1964 ( .I(n851), .ZN(AdrEna[830]) );
  CKND2D0 U1965 ( .A1(\DL3[51].tempL3[1] ), .A2(n16), .ZN(n853) );
  CKNXD16 U1966 ( .I(n853), .ZN(AdrEna[817]) );
  CKND2D0 U1967 ( .A1(\DL3[28].tempL3[9] ), .A2(n42), .ZN(n855) );
  CKNXD16 U1968 ( .I(n855), .ZN(AdrEna[457]) );
  CKND2D0 U1969 ( .A1(\DL3[28].tempL3[7] ), .A2(n42), .ZN(n857) );
  CKNXD16 U1970 ( .I(n857), .ZN(AdrEna[455]) );
  CKND2D0 U1971 ( .A1(\DL3[28].tempL3[8] ), .A2(n42), .ZN(n859) );
  CKNXD16 U1972 ( .I(n859), .ZN(AdrEna[456]) );
  CKND2D0 U1973 ( .A1(\DL3[51].tempL3[9] ), .A2(n16), .ZN(n861) );
  CKNXD16 U1974 ( .I(n861), .ZN(AdrEna[825]) );
  CKND2D0 U1975 ( .A1(\DL3[28].tempL3[4] ), .A2(n42), .ZN(n863) );
  CKNXD16 U1976 ( .I(n863), .ZN(AdrEna[452]) );
  CKND2D0 U1977 ( .A1(\DL3[28].tempL3[10] ), .A2(n42), .ZN(n865) );
  CKNXD16 U1978 ( .I(n865), .ZN(AdrEna[458]) );
  CKND2D0 U1979 ( .A1(\DL3[28].tempL3[12] ), .A2(n42), .ZN(n867) );
  CKNXD16 U1980 ( .I(n867), .ZN(AdrEna[460]) );
  CKND2D0 U1981 ( .A1(\DL3[28].tempL3[11] ), .A2(n42), .ZN(n869) );
  CKNXD16 U1982 ( .I(n869), .ZN(AdrEna[459]) );
  CKND2D0 U1983 ( .A1(\DL3[28].tempL3[13] ), .A2(n42), .ZN(n871) );
  CKNXD16 U1984 ( .I(n871), .ZN(AdrEna[461]) );
  CKND2D0 U1985 ( .A1(\DL3[28].tempL3[2] ), .A2(n42), .ZN(n873) );
  CKNXD16 U1986 ( .I(n873), .ZN(AdrEna[450]) );
  CKND2D0 U1987 ( .A1(\DL3[28].tempL3[3] ), .A2(n42), .ZN(n875) );
  CKNXD16 U1988 ( .I(n875), .ZN(AdrEna[451]) );
  CKND2D0 U1989 ( .A1(\DL3[28].tempL3[15] ), .A2(n42), .ZN(n877) );
  CKNXD16 U1990 ( .I(n877), .ZN(AdrEna[463]) );
  CKND2D0 U1991 ( .A1(\DL3[28].tempL3[0] ), .A2(n42), .ZN(n879) );
  CKNXD16 U1992 ( .I(n879), .ZN(AdrEna[448]) );
  CKND2D0 U1993 ( .A1(\DL3[28].tempL3[14] ), .A2(n42), .ZN(n881) );
  CKNXD16 U1994 ( .I(n881), .ZN(AdrEna[462]) );
  CKND2D0 U1995 ( .A1(\DL3[29].tempL3[0] ), .A2(n41), .ZN(n883) );
  CKNXD16 U1996 ( .I(n883), .ZN(AdrEna[464]) );
  CKND2D0 U1997 ( .A1(\DL3[28].tempL3[1] ), .A2(n42), .ZN(n885) );
  CKNXD16 U1998 ( .I(n885), .ZN(AdrEna[449]) );
  CKND2D0 U1999 ( .A1(\DL3[29].tempL3[1] ), .A2(n41), .ZN(n887) );
  CKNXD16 U2000 ( .I(n887), .ZN(AdrEna[465]) );
  CKND2D0 U2001 ( .A1(\DL3[27].tempL3[14] ), .A2(n43), .ZN(n889) );
  CKNXD16 U2002 ( .I(n889), .ZN(AdrEna[446]) );
  CKND2D0 U2003 ( .A1(\DL3[27].tempL3[15] ), .A2(n43), .ZN(n891) );
  CKNXD16 U2004 ( .I(n891), .ZN(AdrEna[447]) );
  CKND2D0 U2005 ( .A1(\DL3[29].tempL3[3] ), .A2(n41), .ZN(n893) );
  CKNXD16 U2006 ( .I(n893), .ZN(AdrEna[467]) );
  CKND2D0 U2007 ( .A1(\DL3[27].tempL3[12] ), .A2(n43), .ZN(n895) );
  CKNXD16 U2008 ( .I(n895), .ZN(AdrEna[444]) );
  CKND2D0 U2009 ( .A1(\DL3[29].tempL3[2] ), .A2(n41), .ZN(n897) );
  CKNXD16 U2010 ( .I(n897), .ZN(AdrEna[466]) );
  CKND2D0 U2011 ( .A1(\DL3[29].tempL3[4] ), .A2(n41), .ZN(n899) );
  CKNXD16 U2012 ( .I(n899), .ZN(AdrEna[468]) );
  CKND2D0 U2013 ( .A1(\DL3[27].tempL3[13] ), .A2(n43), .ZN(n901) );
  CKNXD16 U2014 ( .I(n901), .ZN(AdrEna[445]) );
  CKND2D0 U2015 ( .A1(\DL3[29].tempL3[5] ), .A2(n41), .ZN(n903) );
  CKNXD16 U2016 ( .I(n903), .ZN(AdrEna[469]) );
  CKND2D0 U2017 ( .A1(\DL3[27].tempL3[10] ), .A2(n43), .ZN(n905) );
  CKNXD16 U2018 ( .I(n905), .ZN(AdrEna[442]) );
  CKND2D0 U2019 ( .A1(\DL3[27].tempL3[11] ), .A2(n43), .ZN(n907) );
  CKNXD16 U2020 ( .I(n907), .ZN(AdrEna[443]) );
  CKND2D0 U2021 ( .A1(\DL3[29].tempL3[9] ), .A2(n41), .ZN(n909) );
  CKNXD16 U2022 ( .I(n909), .ZN(AdrEna[473]) );
  CKND2D0 U2023 ( .A1(\DL3[27].tempL3[8] ), .A2(n43), .ZN(n911) );
  CKNXD16 U2024 ( .I(n911), .ZN(AdrEna[440]) );
  CKND2D0 U2025 ( .A1(\DL3[29].tempL3[8] ), .A2(n41), .ZN(n913) );
  CKNXD16 U2026 ( .I(n913), .ZN(AdrEna[472]) );
  CKND2D0 U2027 ( .A1(\DL3[29].tempL3[10] ), .A2(n41), .ZN(n915) );
  CKNXD16 U2028 ( .I(n915), .ZN(AdrEna[474]) );
  CKND2D0 U2029 ( .A1(\DL3[27].tempL3[9] ), .A2(n43), .ZN(n917) );
  CKNXD16 U2030 ( .I(n917), .ZN(AdrEna[441]) );
  CKND2D0 U2031 ( .A1(\DL3[29].tempL3[11] ), .A2(n41), .ZN(n919) );
  CKNXD16 U2032 ( .I(n919), .ZN(AdrEna[475]) );
  CKND2D0 U2033 ( .A1(\DL3[27].tempL3[4] ), .A2(n43), .ZN(n921) );
  CKNXD16 U2034 ( .I(n921), .ZN(AdrEna[436]) );
  CKND2D0 U2035 ( .A1(\DL3[27].tempL3[5] ), .A2(n43), .ZN(n923) );
  CKNXD16 U2036 ( .I(n923), .ZN(AdrEna[437]) );
  CKND2D0 U2037 ( .A1(\DL3[29].tempL3[13] ), .A2(n41), .ZN(n925) );
  CKNXD16 U2038 ( .I(n925), .ZN(AdrEna[477]) );
  CKND2D0 U2039 ( .A1(\DL3[27].tempL3[2] ), .A2(n43), .ZN(n927) );
  CKNXD16 U2040 ( .I(n927), .ZN(AdrEna[434]) );
  CKND2D0 U2041 ( .A1(\DL3[29].tempL3[12] ), .A2(n41), .ZN(n929) );
  CKNXD16 U2042 ( .I(n929), .ZN(AdrEna[476]) );
  CKND2D0 U2043 ( .A1(\DL3[29].tempL3[14] ), .A2(n41), .ZN(n931) );
  CKNXD16 U2044 ( .I(n931), .ZN(AdrEna[478]) );
  CKND2D0 U2045 ( .A1(\DL3[27].tempL3[3] ), .A2(n43), .ZN(n933) );
  CKNXD16 U2046 ( .I(n933), .ZN(AdrEna[435]) );
  CKND2D0 U2047 ( .A1(\DL3[29].tempL3[15] ), .A2(n41), .ZN(n935) );
  CKNXD16 U2048 ( .I(n935), .ZN(AdrEna[479]) );
  CKND2D0 U2049 ( .A1(\DL3[27].tempL3[0] ), .A2(n43), .ZN(n937) );
  CKNXD16 U2050 ( .I(n937), .ZN(AdrEna[432]) );
  CKND2D0 U2051 ( .A1(\DL3[27].tempL3[1] ), .A2(n43), .ZN(n939) );
  CKNXD16 U2052 ( .I(n939), .ZN(AdrEna[433]) );
  CKND2D0 U2053 ( .A1(\DL3[30].tempL3[1] ), .A2(n39), .ZN(n941) );
  CKNXD16 U2054 ( .I(n941), .ZN(AdrEna[481]) );
  CKND2D0 U2055 ( .A1(\DL3[26].tempL3[14] ), .A2(n44), .ZN(n943) );
  CKNXD16 U2056 ( .I(n943), .ZN(AdrEna[430]) );
  CKND2D0 U2057 ( .A1(\DL3[30].tempL3[0] ), .A2(n39), .ZN(n945) );
  CKNXD16 U2058 ( .I(n945), .ZN(AdrEna[480]) );
  CKND2D0 U2059 ( .A1(\DL3[30].tempL3[2] ), .A2(n39), .ZN(n947) );
  CKNXD16 U2060 ( .I(n947), .ZN(AdrEna[482]) );
  CKND2D0 U2061 ( .A1(\DL3[26].tempL3[15] ), .A2(n44), .ZN(n949) );
  CKNXD16 U2062 ( .I(n949), .ZN(AdrEna[431]) );
  CKND2D0 U2063 ( .A1(\DL3[30].tempL3[3] ), .A2(n39), .ZN(n951) );
  CKNXD16 U2064 ( .I(n951), .ZN(AdrEna[483]) );
  CKND2D0 U2065 ( .A1(\DL3[26].tempL3[12] ), .A2(n44), .ZN(n953) );
  CKNXD16 U2066 ( .I(n953), .ZN(AdrEna[428]) );
  CKND2D0 U2067 ( .A1(\DL3[26].tempL3[13] ), .A2(n44), .ZN(n955) );
  CKNXD16 U2068 ( .I(n955), .ZN(AdrEna[429]) );
  CKND2D0 U2069 ( .A1(\DL3[28].tempL3[5] ), .A2(n42), .ZN(n957) );
  CKNXD16 U2070 ( .I(n957), .ZN(AdrEna[453]) );
  CKND2D0 U2071 ( .A1(\DL3[26].tempL3[10] ), .A2(n44), .ZN(n959) );
  CKNXD16 U2072 ( .I(n959), .ZN(AdrEna[426]) );
  CKND2D0 U2073 ( .A1(\DL3[30].tempL3[4] ), .A2(n39), .ZN(n961) );
  CKNXD16 U2074 ( .I(n961), .ZN(AdrEna[484]) );
  CKND2D0 U2075 ( .A1(\DL3[30].tempL3[7] ), .A2(n39), .ZN(n963) );
  CKNXD16 U2076 ( .I(n963), .ZN(AdrEna[487]) );
  CKND2D0 U2077 ( .A1(\DL3[26].tempL3[11] ), .A2(n44), .ZN(n965) );
  CKNXD16 U2078 ( .I(n965), .ZN(AdrEna[427]) );
  CKND2D0 U2079 ( .A1(\DL3[30].tempL3[10] ), .A2(n39), .ZN(n967) );
  CKNXD16 U2080 ( .I(n967), .ZN(AdrEna[490]) );
  CKND2D0 U2081 ( .A1(\DL3[26].tempL3[8] ), .A2(n44), .ZN(n969) );
  CKNXD16 U2082 ( .I(n969), .ZN(AdrEna[424]) );
  CKND2D0 U2083 ( .A1(\DL3[26].tempL3[9] ), .A2(n44), .ZN(n971) );
  CKNXD16 U2084 ( .I(n971), .ZN(AdrEna[425]) );
  CKND2D0 U2085 ( .A1(\DL3[30].tempL3[8] ), .A2(n39), .ZN(n973) );
  CKNXD16 U2086 ( .I(n973), .ZN(AdrEna[488]) );
  CKND2D0 U2087 ( .A1(\DL3[26].tempL3[5] ), .A2(n44), .ZN(n975) );
  CKNXD16 U2088 ( .I(n975), .ZN(AdrEna[421]) );
  CKND2D0 U2089 ( .A1(\DL3[30].tempL3[9] ), .A2(n39), .ZN(n977) );
  CKNXD16 U2090 ( .I(n977), .ZN(AdrEna[489]) );
  CKND2D0 U2091 ( .A1(\DL3[30].tempL3[11] ), .A2(n39), .ZN(n979) );
  CKNXD16 U2092 ( .I(n979), .ZN(AdrEna[491]) );
  CKND2D0 U2093 ( .A1(\DL3[26].tempL3[7] ), .A2(n44), .ZN(n981) );
  CKNXD16 U2094 ( .I(n981), .ZN(AdrEna[423]) );
  CKND2D0 U2095 ( .A1(\DL3[30].tempL3[13] ), .A2(n39), .ZN(n983) );
  CKNXD16 U2096 ( .I(n983), .ZN(AdrEna[493]) );
  CKND2D0 U2097 ( .A1(\DL3[26].tempL3[3] ), .A2(n44), .ZN(n985) );
  CKNXD16 U2098 ( .I(n985), .ZN(AdrEna[419]) );
  CKND2D0 U2099 ( .A1(\DL3[26].tempL3[4] ), .A2(n44), .ZN(n987) );
  CKNXD16 U2100 ( .I(n987), .ZN(AdrEna[420]) );
  CKND2D0 U2101 ( .A1(\DL3[30].tempL3[12] ), .A2(n39), .ZN(n989) );
  CKNXD16 U2102 ( .I(n989), .ZN(AdrEna[492]) );
  CKND2D0 U2103 ( .A1(\DL3[26].tempL3[2] ), .A2(n44), .ZN(n991) );
  CKNXD16 U2104 ( .I(n991), .ZN(AdrEna[418]) );
  CKND2D0 U2105 ( .A1(\DL3[30].tempL3[5] ), .A2(n39), .ZN(n993) );
  CKNXD16 U2106 ( .I(n993), .ZN(AdrEna[485]) );
  CKND2D0 U2107 ( .A1(\DL3[31].tempL3[1] ), .A2(n38), .ZN(n995) );
  CKNXD16 U2108 ( .I(n995), .ZN(AdrEna[497]) );
  CKND2D0 U2109 ( .A1(\DL3[26].tempL3[1] ), .A2(n44), .ZN(n997) );
  CKNXD16 U2110 ( .I(n997), .ZN(AdrEna[417]) );
  CKND2D0 U2111 ( .A1(\DL3[31].tempL3[4] ), .A2(n38), .ZN(n999) );
  CKNXD16 U2112 ( .I(n999), .ZN(AdrEna[500]) );
  CKND2D0 U2113 ( .A1(\DL3[25].tempL3[15] ), .A2(n45), .ZN(n1001) );
  CKNXD16 U2114 ( .I(n1001), .ZN(AdrEna[415]) );
  CKND2D0 U2115 ( .A1(\DL3[26].tempL3[0] ), .A2(n44), .ZN(n1003) );
  CKNXD16 U2116 ( .I(n1003), .ZN(AdrEna[416]) );
  CKND2D0 U2117 ( .A1(\DL3[31].tempL3[2] ), .A2(n38), .ZN(n1005) );
  CKNXD16 U2118 ( .I(n1005), .ZN(AdrEna[498]) );
  CKND2D0 U2119 ( .A1(\DL3[25].tempL3[14] ), .A2(n45), .ZN(n1007) );
  CKNXD16 U2120 ( .I(n1007), .ZN(AdrEna[414]) );
  CKND2D0 U2121 ( .A1(\DL3[31].tempL3[3] ), .A2(n38), .ZN(n1009) );
  CKNXD16 U2122 ( .I(n1009), .ZN(AdrEna[499]) );
  CKND2D0 U2123 ( .A1(\DL3[30].tempL3[15] ), .A2(n39), .ZN(n1011) );
  CKNXD16 U2124 ( .I(n1011), .ZN(AdrEna[495]) );
  CKND2D0 U2125 ( .A1(\DL3[25].tempL3[13] ), .A2(n45), .ZN(n1013) );
  CKNXD16 U2126 ( .I(n1013), .ZN(AdrEna[413]) );
  CKND2D0 U2127 ( .A1(\DL3[31].tempL3[9] ), .A2(n38), .ZN(n1015) );
  CKNXD16 U2128 ( .I(n1015), .ZN(AdrEna[505]) );
  CKND2D0 U2129 ( .A1(\DL3[25].tempL3[11] ), .A2(n45), .ZN(n1017) );
  CKNXD16 U2130 ( .I(n1017), .ZN(AdrEna[411]) );
  CKND2D0 U2131 ( .A1(\DL3[25].tempL3[12] ), .A2(n45), .ZN(n1019) );
  CKNXD16 U2132 ( .I(n1019), .ZN(AdrEna[412]) );
  CKND2D0 U2133 ( .A1(\DL3[31].tempL3[13] ), .A2(n38), .ZN(n1021) );
  CKNXD16 U2134 ( .I(n1021), .ZN(AdrEna[509]) );
  CKND2D0 U2135 ( .A1(\DL3[25].tempL3[10] ), .A2(n45), .ZN(n1023) );
  CKNXD16 U2136 ( .I(n1023), .ZN(AdrEna[410]) );
  CKND2D0 U2137 ( .A1(\DL3[31].tempL3[12] ), .A2(n38), .ZN(n1025) );
  CKNXD16 U2138 ( .I(n1025), .ZN(AdrEna[508]) );
  CKND2D0 U2139 ( .A1(\DL3[32].tempL3[0] ), .A2(n37), .ZN(n1027) );
  CKNXD16 U2140 ( .I(n1027), .ZN(AdrEna[512]) );
  CKND2D0 U2141 ( .A1(\DL3[25].tempL3[9] ), .A2(n45), .ZN(n1029) );
  CKNXD16 U2142 ( .I(n1029), .ZN(AdrEna[409]) );
  CKND2D0 U2143 ( .A1(\DL3[32].tempL3[1] ), .A2(n37), .ZN(n1031) );
  CKNXD16 U2144 ( .I(n1031), .ZN(AdrEna[513]) );
  CKND2D0 U2145 ( .A1(\DL3[25].tempL3[5] ), .A2(n45), .ZN(n1033) );
  CKNXD16 U2146 ( .I(n1033), .ZN(AdrEna[405]) );
  CKND2D0 U2147 ( .A1(\DL3[25].tempL3[8] ), .A2(n45), .ZN(n1035) );
  CKNXD16 U2148 ( .I(n1035), .ZN(AdrEna[408]) );
  CKND2D0 U2149 ( .A1(\DL3[32].tempL3[3] ), .A2(n37), .ZN(n1037) );
  CKNXD16 U2150 ( .I(n1037), .ZN(AdrEna[515]) );
  CKND2D0 U2151 ( .A1(\DL3[25].tempL3[4] ), .A2(n45), .ZN(n1039) );
  CKNXD16 U2152 ( .I(n1039), .ZN(AdrEna[404]) );
  CKND2D0 U2153 ( .A1(\DL3[32].tempL3[2] ), .A2(n37), .ZN(n1041) );
  CKNXD16 U2154 ( .I(n1041), .ZN(AdrEna[514]) );
  CKND2D0 U2155 ( .A1(\DL3[32].tempL3[4] ), .A2(n37), .ZN(n1043) );
  CKNXD16 U2156 ( .I(n1043), .ZN(AdrEna[516]) );
  CKND2D0 U2157 ( .A1(\DL3[25].tempL3[3] ), .A2(n45), .ZN(n1045) );
  CKNXD16 U2158 ( .I(n1045), .ZN(AdrEna[403]) );
  CKND2D0 U2159 ( .A1(\DL3[32].tempL3[5] ), .A2(n37), .ZN(n1047) );
  CKNXD16 U2160 ( .I(n1047), .ZN(AdrEna[517]) );
  CKND2D0 U2161 ( .A1(\DL3[25].tempL3[1] ), .A2(n45), .ZN(n1049) );
  CKNXD16 U2162 ( .I(n1049), .ZN(AdrEna[401]) );
  CKND2D0 U2163 ( .A1(\DL3[25].tempL3[2] ), .A2(n45), .ZN(n1051) );
  CKNXD16 U2164 ( .I(n1051), .ZN(AdrEna[402]) );
  CKND2D0 U2165 ( .A1(\DL3[32].tempL3[7] ), .A2(n37), .ZN(n1053) );
  CKNXD16 U2166 ( .I(n1053), .ZN(AdrEna[519]) );
  CKND2D0 U2167 ( .A1(\DL3[25].tempL3[0] ), .A2(n45), .ZN(n1055) );
  CKNXD16 U2168 ( .I(n1055), .ZN(AdrEna[400]) );
  CKND2D0 U2169 ( .A1(\DL3[32].tempL3[6] ), .A2(n37), .ZN(n1057) );
  CKNXD16 U2170 ( .I(n1057), .ZN(AdrEna[518]) );
  CKND2D0 U2171 ( .A1(\DL3[32].tempL3[8] ), .A2(n37), .ZN(n1059) );
  CKNXD16 U2172 ( .I(n1059), .ZN(AdrEna[520]) );
  CKND2D0 U2173 ( .A1(\DL3[24].tempL3[15] ), .A2(n46), .ZN(n1061) );
  CKNXD16 U2174 ( .I(n1061), .ZN(AdrEna[399]) );
  CKND2D0 U2175 ( .A1(\DL3[32].tempL3[9] ), .A2(n37), .ZN(n1063) );
  CKNXD16 U2176 ( .I(n1063), .ZN(AdrEna[521]) );
  CKND2D0 U2177 ( .A1(\DL3[24].tempL3[13] ), .A2(n46), .ZN(n1065) );
  CKNXD16 U2178 ( .I(n1065), .ZN(AdrEna[397]) );
  CKND2D0 U2179 ( .A1(\DL3[24].tempL3[14] ), .A2(n46), .ZN(n1067) );
  CKNXD16 U2180 ( .I(n1067), .ZN(AdrEna[398]) );
  CKND2D0 U2181 ( .A1(\DL3[33].tempL3[1] ), .A2(n36), .ZN(n1069) );
  CKNXD16 U2182 ( .I(n1069), .ZN(AdrEna[529]) );
  CKND2D0 U2183 ( .A1(\DL3[24].tempL3[12] ), .A2(n46), .ZN(n1071) );
  CKNXD16 U2184 ( .I(n1071), .ZN(AdrEna[396]) );
  CKND2D0 U2185 ( .A1(\DL3[33].tempL3[0] ), .A2(n36), .ZN(n1073) );
  CKNXD16 U2186 ( .I(n1073), .ZN(AdrEna[528]) );
  CKND2D0 U2187 ( .A1(\DL3[33].tempL3[2] ), .A2(n36), .ZN(n1075) );
  CKNXD16 U2188 ( .I(n1075), .ZN(AdrEna[530]) );
  CKND2D0 U2189 ( .A1(\DL3[24].tempL3[11] ), .A2(n46), .ZN(n1077) );
  CKNXD16 U2190 ( .I(n1077), .ZN(AdrEna[395]) );
  CKND2D0 U2191 ( .A1(\DL3[24].tempL3[9] ), .A2(n46), .ZN(n1079) );
  CKNXD16 U2192 ( .I(n1079), .ZN(AdrEna[393]) );
  CKND2D0 U2193 ( .A1(\DL3[24].tempL3[10] ), .A2(n46), .ZN(n1081) );
  CKNXD16 U2194 ( .I(n1081), .ZN(AdrEna[394]) );
  CKND2D0 U2195 ( .A1(\DL3[33].tempL3[3] ), .A2(n36), .ZN(n1083) );
  CKNXD16 U2196 ( .I(n1083), .ZN(AdrEna[531]) );
  CKND2D0 U2197 ( .A1(\DL3[24].tempL3[8] ), .A2(n46), .ZN(n1085) );
  CKNXD16 U2198 ( .I(n1085), .ZN(AdrEna[392]) );
  CKND2D0 U2199 ( .A1(\DL3[33].tempL3[4] ), .A2(n36), .ZN(n1087) );
  CKNXD16 U2200 ( .I(n1087), .ZN(AdrEna[532]) );
  CKND2D0 U2201 ( .A1(\DL3[33].tempL3[6] ), .A2(n36), .ZN(n1089) );
  CKNXD16 U2202 ( .I(n1089), .ZN(AdrEna[534]) );
  CKND2D0 U2203 ( .A1(\DL3[24].tempL3[7] ), .A2(n46), .ZN(n1091) );
  CKNXD16 U2204 ( .I(n1091), .ZN(AdrEna[391]) );
  CKND2D0 U2205 ( .A1(\DL3[33].tempL3[9] ), .A2(n36), .ZN(n1093) );
  CKNXD16 U2206 ( .I(n1093), .ZN(AdrEna[537]) );
  CKND2D0 U2207 ( .A1(\DL3[24].tempL3[4] ), .A2(n46), .ZN(n1095) );
  CKNXD16 U2208 ( .I(n1095), .ZN(AdrEna[388]) );
  CKND2D0 U2209 ( .A1(\DL3[24].tempL3[5] ), .A2(n46), .ZN(n1097) );
  CKNXD16 U2210 ( .I(n1097), .ZN(AdrEna[389]) );
  CKND2D0 U2211 ( .A1(\DL3[33].tempL3[7] ), .A2(n36), .ZN(n1099) );
  CKNXD16 U2212 ( .I(n1099), .ZN(AdrEna[535]) );
  CKND2D0 U2213 ( .A1(\DL3[24].tempL3[2] ), .A2(n46), .ZN(n1101) );
  CKNXD16 U2214 ( .I(n1101), .ZN(AdrEna[386]) );
  CKND2D0 U2215 ( .A1(\DL3[33].tempL3[8] ), .A2(n36), .ZN(n1103) );
  CKNXD16 U2216 ( .I(n1103), .ZN(AdrEna[536]) );
  CKND2D0 U2217 ( .A1(\DL3[34].tempL3[0] ), .A2(n35), .ZN(n1105) );
  CKNXD16 U2218 ( .I(n1105), .ZN(AdrEna[544]) );
  CKND2D0 U2219 ( .A1(\DL3[24].tempL3[3] ), .A2(n46), .ZN(n1107) );
  CKNXD16 U2220 ( .I(n1107), .ZN(AdrEna[387]) );
  CKND2D0 U2221 ( .A1(\DL3[34].tempL3[3] ), .A2(n35), .ZN(n1109) );
  CKNXD16 U2222 ( .I(n1109), .ZN(AdrEna[547]) );
  CKND2D0 U2223 ( .A1(\DL3[24].tempL3[0] ), .A2(n46), .ZN(n1111) );
  CKNXD16 U2224 ( .I(n1111), .ZN(AdrEna[384]) );
  CKND2D0 U2225 ( .A1(\DL3[24].tempL3[1] ), .A2(n46), .ZN(n1113) );
  CKNXD16 U2226 ( .I(n1113), .ZN(AdrEna[385]) );
  CKND2D0 U2227 ( .A1(\DL3[34].tempL3[1] ), .A2(n35), .ZN(n1115) );
  CKNXD16 U2228 ( .I(n1115), .ZN(AdrEna[545]) );
  CKND2D0 U2229 ( .A1(\DL3[23].tempL3[14] ), .A2(n47), .ZN(n1117) );
  CKNXD16 U2230 ( .I(n1117), .ZN(AdrEna[382]) );
  CKND2D0 U2231 ( .A1(\DL3[34].tempL3[2] ), .A2(n35), .ZN(n1119) );
  CKNXD16 U2232 ( .I(n1119), .ZN(AdrEna[546]) );
  CKND2D0 U2233 ( .A1(\DL3[34].tempL3[4] ), .A2(n35), .ZN(n1121) );
  CKNXD16 U2234 ( .I(n1121), .ZN(AdrEna[548]) );
  CKND2D0 U2235 ( .A1(\DL3[23].tempL3[15] ), .A2(n47), .ZN(n1123) );
  CKNXD16 U2236 ( .I(n1123), .ZN(AdrEna[383]) );
  CKND2D0 U2237 ( .A1(\DL3[34].tempL3[7] ), .A2(n35), .ZN(n1125) );
  CKNXD16 U2238 ( .I(n1125), .ZN(AdrEna[551]) );
  CKND2D0 U2239 ( .A1(\DL3[23].tempL3[11] ), .A2(n47), .ZN(n1127) );
  CKNXD16 U2240 ( .I(n1127), .ZN(AdrEna[379]) );
  CKND2D0 U2241 ( .A1(\DL3[23].tempL3[12] ), .A2(n47), .ZN(n1129) );
  CKNXD16 U2242 ( .I(n1129), .ZN(AdrEna[380]) );
  CKND2D0 U2243 ( .A1(\DL3[34].tempL3[5] ), .A2(n35), .ZN(n1131) );
  CKNXD16 U2244 ( .I(n1131), .ZN(AdrEna[549]) );
  CKND2D0 U2245 ( .A1(\DL3[23].tempL3[10] ), .A2(n47), .ZN(n1133) );
  CKNXD16 U2246 ( .I(n1133), .ZN(AdrEna[378]) );
  CKND2D0 U2247 ( .A1(\DL3[34].tempL3[6] ), .A2(n35), .ZN(n1135) );
  CKNXD16 U2248 ( .I(n1135), .ZN(AdrEna[550]) );
  CKND2D0 U2249 ( .A1(\DL3[34].tempL3[8] ), .A2(n35), .ZN(n1137) );
  CKNXD16 U2250 ( .I(n1137), .ZN(AdrEna[552]) );
  CKND2D0 U2251 ( .A1(\DL3[23].tempL3[9] ), .A2(n47), .ZN(n1139) );
  CKNXD16 U2252 ( .I(n1139), .ZN(AdrEna[377]) );
  CKND2D0 U2253 ( .A1(\DL3[35].tempL3[1] ), .A2(n34), .ZN(n1141) );
  CKNXD16 U2254 ( .I(n1141), .ZN(AdrEna[561]) );
  CKND2D0 U2255 ( .A1(\DL3[23].tempL3[7] ), .A2(n47), .ZN(n1143) );
  CKNXD16 U2256 ( .I(n1143), .ZN(AdrEna[375]) );
  CKND2D0 U2257 ( .A1(\DL3[23].tempL3[8] ), .A2(n47), .ZN(n1145) );
  CKNXD16 U2258 ( .I(n1145), .ZN(AdrEna[376]) );
  CKND2D0 U2259 ( .A1(\DL3[34].tempL3[9] ), .A2(n35), .ZN(n1147) );
  CKNXD16 U2260 ( .I(n1147), .ZN(AdrEna[553]) );
  CKND2D0 U2261 ( .A1(\DL3[23].tempL3[4] ), .A2(n47), .ZN(n1149) );
  CKNXD16 U2262 ( .I(n1149), .ZN(AdrEna[372]) );
  CKND2D0 U2263 ( .A1(\DL3[35].tempL3[0] ), .A2(n34), .ZN(n1151) );
  CKNXD16 U2264 ( .I(n1151), .ZN(AdrEna[560]) );
  CKND2D0 U2265 ( .A1(\DL3[35].tempL3[2] ), .A2(n34), .ZN(n1153) );
  CKNXD16 U2266 ( .I(n1153), .ZN(AdrEna[562]) );
  CKND2D0 U2267 ( .A1(\DL3[23].tempL3[5] ), .A2(n47), .ZN(n1155) );
  CKNXD16 U2268 ( .I(n1155), .ZN(AdrEna[373]) );
  CKND2D0 U2269 ( .A1(\DL3[35].tempL3[5] ), .A2(n34), .ZN(n1157) );
  CKNXD16 U2270 ( .I(n1157), .ZN(AdrEna[565]) );
  CKND2D0 U2271 ( .A1(\DL3[23].tempL3[2] ), .A2(n47), .ZN(n1159) );
  CKNXD16 U2272 ( .I(n1159), .ZN(AdrEna[370]) );
  CKND2D0 U2273 ( .A1(\DL3[23].tempL3[3] ), .A2(n47), .ZN(n1161) );
  CKNXD16 U2274 ( .I(n1161), .ZN(AdrEna[371]) );
  CKND2D0 U2275 ( .A1(\DL3[35].tempL3[3] ), .A2(n34), .ZN(n1163) );
  CKNXD16 U2276 ( .I(n1163), .ZN(AdrEna[563]) );
  CKND2D0 U2277 ( .A1(\DL3[23].tempL3[0] ), .A2(n47), .ZN(n1165) );
  CKNXD16 U2278 ( .I(n1165), .ZN(AdrEna[368]) );
  CKND2D0 U2279 ( .A1(\DL3[35].tempL3[4] ), .A2(n34), .ZN(n1167) );
  CKNXD16 U2280 ( .I(n1167), .ZN(AdrEna[564]) );
  CKND2D0 U2281 ( .A1(\DL3[35].tempL3[6] ), .A2(n34), .ZN(n1169) );
  CKNXD16 U2282 ( .I(n1169), .ZN(AdrEna[566]) );
  CKND2D0 U2283 ( .A1(\DL3[23].tempL3[1] ), .A2(n47), .ZN(n1171) );
  CKNXD16 U2284 ( .I(n1171), .ZN(AdrEna[369]) );
  CKND2D0 U2285 ( .A1(\DL3[35].tempL3[9] ), .A2(n34), .ZN(n1173) );
  CKNXD16 U2286 ( .I(n1173), .ZN(AdrEna[569]) );
  CKND2D0 U2287 ( .A1(\DL3[22].tempL3[14] ), .A2(n48), .ZN(n1175) );
  CKNXD16 U2288 ( .I(n1175), .ZN(AdrEna[366]) );
  CKND2D0 U2289 ( .A1(\DL3[22].tempL3[15] ), .A2(n48), .ZN(n1177) );
  CKNXD16 U2290 ( .I(n1177), .ZN(AdrEna[367]) );
  CKND2D0 U2291 ( .A1(\DL3[35].tempL3[7] ), .A2(n34), .ZN(n1179) );
  CKNXD16 U2292 ( .I(n1179), .ZN(AdrEna[567]) );
  CKND2D0 U2293 ( .A1(\DL3[22].tempL3[12] ), .A2(n48), .ZN(n1181) );
  CKNXD16 U2294 ( .I(n1181), .ZN(AdrEna[364]) );
  CKND2D0 U2295 ( .A1(\DL3[35].tempL3[8] ), .A2(n34), .ZN(n1183) );
  CKNXD16 U2296 ( .I(n1183), .ZN(AdrEna[568]) );
  CKND2D0 U2297 ( .A1(\DL3[36].tempL3[0] ), .A2(n33), .ZN(n1185) );
  CKNXD16 U2298 ( .I(n1185), .ZN(AdrEna[576]) );
  CKND2D0 U2299 ( .A1(\DL3[22].tempL3[13] ), .A2(n48), .ZN(n1187) );
  CKNXD16 U2300 ( .I(n1187), .ZN(AdrEna[365]) );
  CKND2D0 U2301 ( .A1(\DL3[36].tempL3[3] ), .A2(n33), .ZN(n1189) );
  CKNXD16 U2302 ( .I(n1189), .ZN(AdrEna[579]) );
  CKND2D0 U2303 ( .A1(\DL3[22].tempL3[10] ), .A2(n48), .ZN(n1191) );
  CKNXD16 U2304 ( .I(n1191), .ZN(AdrEna[362]) );
  CKND2D0 U2305 ( .A1(\DL3[22].tempL3[11] ), .A2(n48), .ZN(n1193) );
  CKNXD16 U2306 ( .I(n1193), .ZN(AdrEna[363]) );
  CKND2D0 U2307 ( .A1(\DL3[36].tempL3[1] ), .A2(n33), .ZN(n1195) );
  CKNXD16 U2308 ( .I(n1195), .ZN(AdrEna[577]) );
  CKND2D0 U2309 ( .A1(\DL3[22].tempL3[8] ), .A2(n48), .ZN(n1197) );
  CKNXD16 U2310 ( .I(n1197), .ZN(AdrEna[360]) );
  CKND2D0 U2311 ( .A1(\DL3[36].tempL3[2] ), .A2(n33), .ZN(n1199) );
  CKNXD16 U2312 ( .I(n1199), .ZN(AdrEna[578]) );
  CKND2D0 U2313 ( .A1(\DL3[31].tempL3[5] ), .A2(n38), .ZN(n1201) );
  CKNXD16 U2314 ( .I(n1201), .ZN(AdrEna[501]) );
  CKND2D0 U2315 ( .A1(\DL3[22].tempL3[9] ), .A2(n48), .ZN(n1203) );
  CKNXD16 U2316 ( .I(n1203), .ZN(AdrEna[361]) );
  CKND2D0 U2317 ( .A1(\DL3[36].tempL3[8] ), .A2(n33), .ZN(n1205) );
  CKNXD16 U2318 ( .I(n1205), .ZN(AdrEna[584]) );
  CKND2D0 U2319 ( .A1(\DL3[22].tempL3[5] ), .A2(n48), .ZN(n1207) );
  CKNXD16 U2320 ( .I(n1207), .ZN(AdrEna[357]) );
  CKND2D0 U2321 ( .A1(\DL3[22].tempL3[7] ), .A2(n48), .ZN(n1209) );
  CKNXD16 U2322 ( .I(n1209), .ZN(AdrEna[359]) );
  CKND2D0 U2323 ( .A1(\DL3[37].tempL3[0] ), .A2(n32), .ZN(n1211) );
  CKNXD16 U2324 ( .I(n1211), .ZN(AdrEna[592]) );
  CKND2D0 U2325 ( .A1(\DL3[22].tempL3[4] ), .A2(n48), .ZN(n1213) );
  CKNXD16 U2326 ( .I(n1213), .ZN(AdrEna[356]) );
  CKND2D0 U2327 ( .A1(\DL3[36].tempL3[9] ), .A2(n33), .ZN(n1215) );
  CKNXD16 U2328 ( .I(n1215), .ZN(AdrEna[585]) );
  CKND2D0 U2329 ( .A1(\DL3[36].tempL3[4] ), .A2(n33), .ZN(n1217) );
  CKNXD16 U2330 ( .I(n1217), .ZN(AdrEna[580]) );
  CKND2D0 U2331 ( .A1(\DL3[22].tempL3[3] ), .A2(n48), .ZN(n1219) );
  CKNXD16 U2332 ( .I(n1219), .ZN(AdrEna[355]) );
  CKND2D0 U2333 ( .A1(\DL3[37].tempL3[5] ), .A2(n32), .ZN(n1221) );
  CKNXD16 U2334 ( .I(n1221), .ZN(AdrEna[597]) );
  CKND2D0 U2335 ( .A1(\DL3[22].tempL3[1] ), .A2(n48), .ZN(n1223) );
  CKNXD16 U2336 ( .I(n1223), .ZN(AdrEna[353]) );
  CKND2D0 U2337 ( .A1(\DL3[22].tempL3[2] ), .A2(n48), .ZN(n1225) );
  CKNXD16 U2338 ( .I(n1225), .ZN(AdrEna[354]) );
  CKND2D0 U2339 ( .A1(\DL3[37].tempL3[3] ), .A2(n32), .ZN(n1227) );
  CKNXD16 U2340 ( .I(n1227), .ZN(AdrEna[595]) );
  CKND2D0 U2341 ( .A1(\DL3[22].tempL3[0] ), .A2(n48), .ZN(n1229) );
  CKNXD16 U2342 ( .I(n1229), .ZN(AdrEna[352]) );
  CKND2D0 U2343 ( .A1(\DL3[37].tempL3[4] ), .A2(n32), .ZN(n1231) );
  CKNXD16 U2344 ( .I(n1231), .ZN(AdrEna[596]) );
  CKND2D0 U2345 ( .A1(\DL3[37].tempL3[8] ), .A2(n32), .ZN(n1233) );
  CKNXD16 U2346 ( .I(n1233), .ZN(AdrEna[600]) );
  CKND2D0 U2347 ( .A1(\DL3[21].tempL3[15] ), .A2(n49), .ZN(n1235) );
  CKNXD16 U2348 ( .I(n1235), .ZN(AdrEna[351]) );
  CKND2D0 U2349 ( .A1(\DL3[38].tempL3[1] ), .A2(n31), .ZN(n1237) );
  CKNXD16 U2350 ( .I(n1237), .ZN(AdrEna[609]) );
  CKND2D0 U2351 ( .A1(\DL3[21].tempL3[13] ), .A2(n49), .ZN(n1239) );
  CKNXD16 U2352 ( .I(n1239), .ZN(AdrEna[349]) );
  CKND2D0 U2353 ( .A1(\DL3[21].tempL3[14] ), .A2(n49), .ZN(n1241) );
  CKNXD16 U2354 ( .I(n1241), .ZN(AdrEna[350]) );
  CKND2D0 U2355 ( .A1(\DL3[37].tempL3[9] ), .A2(n32), .ZN(n1243) );
  CKNXD16 U2356 ( .I(n1243), .ZN(AdrEna[601]) );
  CKND2D0 U2357 ( .A1(\DL3[21].tempL3[12] ), .A2(n49), .ZN(n1245) );
  CKNXD16 U2358 ( .I(n1245), .ZN(AdrEna[348]) );
  CKND2D0 U2359 ( .A1(\DL3[38].tempL3[0] ), .A2(n31), .ZN(n1247) );
  CKNXD16 U2360 ( .I(n1247), .ZN(AdrEna[608]) );
  CKND2D0 U2361 ( .A1(\DL3[37].tempL3[1] ), .A2(n32), .ZN(n1249) );
  CKNXD16 U2362 ( .I(n1249), .ZN(AdrEna[593]) );
  CKND2D0 U2363 ( .A1(\DL3[21].tempL3[11] ), .A2(n49), .ZN(n1251) );
  CKNXD16 U2364 ( .I(n1251), .ZN(AdrEna[347]) );
  CKND2D0 U2365 ( .A1(\DL3[38].tempL3[8] ), .A2(n31), .ZN(n1253) );
  CKNXD16 U2366 ( .I(n1253), .ZN(AdrEna[616]) );
  CKND2D0 U2367 ( .A1(\DL3[21].tempL3[9] ), .A2(n49), .ZN(n1255) );
  CKNXD16 U2368 ( .I(n1255), .ZN(AdrEna[345]) );
  CKND2D0 U2369 ( .A1(\DL3[21].tempL3[10] ), .A2(n49), .ZN(n1257) );
  CKNXD16 U2370 ( .I(n1257), .ZN(AdrEna[346]) );
  CKND2D0 U2371 ( .A1(\DL3[39].tempL3[0] ), .A2(n30), .ZN(n1259) );
  CKNXD16 U2372 ( .I(n1259), .ZN(AdrEna[624]) );
  CKND2D0 U2373 ( .A1(\DL3[21].tempL3[8] ), .A2(n49), .ZN(n1261) );
  CKNXD16 U2374 ( .I(n1261), .ZN(AdrEna[344]) );
  CKND2D0 U2375 ( .A1(\DL3[38].tempL3[9] ), .A2(n31), .ZN(n1263) );
  CKNXD16 U2376 ( .I(n1263), .ZN(AdrEna[617]) );
  CKND2D0 U2377 ( .A1(\DL3[38].tempL3[4] ), .A2(n31), .ZN(n1265) );
  CKNXD16 U2378 ( .I(n1265), .ZN(AdrEna[612]) );
  CKND2D0 U2379 ( .A1(\DL3[21].tempL3[7] ), .A2(n49), .ZN(n1267) );
  CKNXD16 U2380 ( .I(n1267), .ZN(AdrEna[343]) );
  CKND2D0 U2381 ( .A1(\DL3[39].tempL3[5] ), .A2(n30), .ZN(n1269) );
  CKNXD16 U2382 ( .I(n1269), .ZN(AdrEna[629]) );
  CKND2D0 U2383 ( .A1(\DL3[21].tempL3[4] ), .A2(n49), .ZN(n1271) );
  CKNXD16 U2384 ( .I(n1271), .ZN(AdrEna[340]) );
  CKND2D0 U2385 ( .A1(\DL3[21].tempL3[5] ), .A2(n49), .ZN(n1273) );
  CKNXD16 U2386 ( .I(n1273), .ZN(AdrEna[341]) );
  CKND2D0 U2387 ( .A1(\DL3[39].tempL3[3] ), .A2(n30), .ZN(n1275) );
  CKNXD16 U2388 ( .I(n1275), .ZN(AdrEna[627]) );
  CKND2D0 U2389 ( .A1(\DL3[21].tempL3[2] ), .A2(n49), .ZN(n1277) );
  CKNXD16 U2390 ( .I(n1277), .ZN(AdrEna[338]) );
  CKND2D0 U2391 ( .A1(\DL3[39].tempL3[4] ), .A2(n30), .ZN(n1279) );
  CKNXD16 U2392 ( .I(n1279), .ZN(AdrEna[628]) );
  CKND2D0 U2393 ( .A1(\DL3[39].tempL3[8] ), .A2(n30), .ZN(n1281) );
  CKNXD16 U2394 ( .I(n1281), .ZN(AdrEna[632]) );
  CKND2D0 U2395 ( .A1(\DL3[21].tempL3[3] ), .A2(n49), .ZN(n1283) );
  CKNXD16 U2396 ( .I(n1283), .ZN(AdrEna[339]) );
  CKND2D0 U2397 ( .A1(\DL3[40].tempL3[1] ), .A2(n28), .ZN(n1285) );
  CKNXD16 U2398 ( .I(n1285), .ZN(AdrEna[641]) );
  CKND2D0 U2399 ( .A1(\DL3[21].tempL3[0] ), .A2(n49), .ZN(n1287) );
  CKNXD16 U2400 ( .I(n1287), .ZN(AdrEna[336]) );
  CKND2D0 U2401 ( .A1(\DL3[21].tempL3[1] ), .A2(n49), .ZN(n1289) );
  CKNXD16 U2402 ( .I(n1289), .ZN(AdrEna[337]) );
  CKND2D0 U2403 ( .A1(\DL3[39].tempL3[9] ), .A2(n30), .ZN(n1291) );
  CKNXD16 U2404 ( .I(n1291), .ZN(AdrEna[633]) );
  CKND2D0 U2405 ( .A1(\DL3[20].tempL3[14] ), .A2(n50), .ZN(n1293) );
  CKNXD16 U2406 ( .I(n1293), .ZN(AdrEna[334]) );
  CKND2D0 U2407 ( .A1(\DL3[40].tempL3[0] ), .A2(n28), .ZN(n1295) );
  CKNXD16 U2408 ( .I(n1295), .ZN(AdrEna[640]) );
  CKND2D0 U2409 ( .A1(\DL3[40].tempL3[2] ), .A2(n28), .ZN(n1297) );
  CKNXD16 U2410 ( .I(n1297), .ZN(AdrEna[642]) );
  CKND2D0 U2411 ( .A1(\DL3[20].tempL3[15] ), .A2(n50), .ZN(n1299) );
  CKNXD16 U2412 ( .I(n1299), .ZN(AdrEna[335]) );
  CKND2D0 U2413 ( .A1(\DL3[40].tempL3[8] ), .A2(n28), .ZN(n1301) );
  CKNXD16 U2414 ( .I(n1301), .ZN(AdrEna[648]) );
  CKND2D0 U2415 ( .A1(\DL3[20].tempL3[12] ), .A2(n50), .ZN(n1303) );
  CKNXD16 U2416 ( .I(n1303), .ZN(AdrEna[332]) );
  CKND2D0 U2417 ( .A1(\DL3[20].tempL3[13] ), .A2(n50), .ZN(n1305) );
  CKNXD16 U2418 ( .I(n1305), .ZN(AdrEna[333]) );
  CKND2D0 U2419 ( .A1(\DL3[40].tempL3[3] ), .A2(n28), .ZN(n1307) );
  CKNXD16 U2420 ( .I(n1307), .ZN(AdrEna[643]) );
  CKND2D0 U2421 ( .A1(\DL3[20].tempL3[10] ), .A2(n50), .ZN(n1309) );
  CKNXD16 U2422 ( .I(n1309), .ZN(AdrEna[330]) );
  CKND2D0 U2423 ( .A1(\DL3[39].tempL3[1] ), .A2(n30), .ZN(n1311) );
  CKNXD16 U2424 ( .I(n1311), .ZN(AdrEna[625]) );
  CKND2D0 U2425 ( .A1(\DL3[40].tempL3[9] ), .A2(n28), .ZN(n1313) );
  CKNXD16 U2426 ( .I(n1313), .ZN(AdrEna[649]) );
  CKND2D0 U2427 ( .A1(\DL3[20].tempL3[11] ), .A2(n50), .ZN(n1315) );
  CKNXD16 U2428 ( .I(n1315), .ZN(AdrEna[331]) );
  CKND2D0 U2429 ( .A1(\DL3[41].tempL3[0] ), .A2(n27), .ZN(n1317) );
  CKNXD16 U2430 ( .I(n1317), .ZN(AdrEna[656]) );
  CKND2D0 U2431 ( .A1(\DL3[20].tempL3[8] ), .A2(n50), .ZN(n1319) );
  CKNXD16 U2432 ( .I(n1319), .ZN(AdrEna[328]) );
  CKND2D0 U2433 ( .A1(\DL3[20].tempL3[9] ), .A2(n50), .ZN(n1321) );
  CKNXD16 U2434 ( .I(n1321), .ZN(AdrEna[329]) );
  CKND2D0 U2435 ( .A1(\DL3[41].tempL3[2] ), .A2(n27), .ZN(n1323) );
  CKNXD16 U2436 ( .I(n1323), .ZN(AdrEna[658]) );
  CKND2D0 U2437 ( .A1(\DL3[20].tempL3[5] ), .A2(n50), .ZN(n1325) );
  CKNXD16 U2438 ( .I(n1325), .ZN(AdrEna[325]) );
  CKND2D0 U2439 ( .A1(\DL3[41].tempL3[1] ), .A2(n27), .ZN(n1327) );
  CKNXD16 U2440 ( .I(n1327), .ZN(AdrEna[657]) );
  CKND2D0 U2441 ( .A1(\DL3[41].tempL3[3] ), .A2(n27), .ZN(n1329) );
  CKNXD16 U2442 ( .I(n1329), .ZN(AdrEna[659]) );
  CKND2D0 U2443 ( .A1(\DL3[20].tempL3[7] ), .A2(n50), .ZN(n1331) );
  CKNXD16 U2444 ( .I(n1331), .ZN(AdrEna[327]) );
  CKND2D0 U2445 ( .A1(\DL3[41].tempL3[8] ), .A2(n27), .ZN(n1333) );
  CKNXD16 U2446 ( .I(n1333), .ZN(AdrEna[664]) );
  CKND2D0 U2447 ( .A1(\DL3[20].tempL3[3] ), .A2(n50), .ZN(n1335) );
  CKNXD16 U2448 ( .I(n1335), .ZN(AdrEna[323]) );
  CKND2D0 U2449 ( .A1(\DL3[20].tempL3[4] ), .A2(n50), .ZN(n1337) );
  CKNXD16 U2450 ( .I(n1337), .ZN(AdrEna[324]) );
  CKND2D0 U2451 ( .A1(\DL3[42].tempL3[0] ), .A2(n26), .ZN(n1339) );
  CKNXD16 U2452 ( .I(n1339), .ZN(AdrEna[672]) );
  CKND2D0 U2453 ( .A1(\DL3[20].tempL3[2] ), .A2(n50), .ZN(n1341) );
  CKNXD16 U2454 ( .I(n1341), .ZN(AdrEna[322]) );
  CKND2D0 U2455 ( .A1(\DL3[41].tempL3[9] ), .A2(n27), .ZN(n1343) );
  CKNXD16 U2456 ( .I(n1343), .ZN(AdrEna[665]) );
  CKND2D0 U2457 ( .A1(\DL3[40].tempL3[4] ), .A2(n28), .ZN(n1345) );
  CKNXD16 U2458 ( .I(n1345), .ZN(AdrEna[644]) );
  CKND2D0 U2459 ( .A1(\DL3[20].tempL3[1] ), .A2(n50), .ZN(n1347) );
  CKNXD16 U2460 ( .I(n1347), .ZN(AdrEna[321]) );
  CKND2D0 U2461 ( .A1(\DL3[42].tempL3[5] ), .A2(n26), .ZN(n1349) );
  CKNXD16 U2462 ( .I(n1349), .ZN(AdrEna[677]) );
  CKND2D0 U2463 ( .A1(\DL3[19].tempL3[15] ), .A2(n52), .ZN(n1351) );
  CKNXD16 U2464 ( .I(n1351), .ZN(AdrEna[319]) );
  CKND2D0 U2465 ( .A1(\DL3[20].tempL3[0] ), .A2(n50), .ZN(n1353) );
  CKNXD16 U2466 ( .I(n1353), .ZN(AdrEna[320]) );
  CKND2D0 U2467 ( .A1(\DL3[42].tempL3[3] ), .A2(n26), .ZN(n1355) );
  CKNXD16 U2468 ( .I(n1355), .ZN(AdrEna[675]) );
  CKND2D0 U2469 ( .A1(\DL3[19].tempL3[14] ), .A2(n52), .ZN(n1357) );
  CKNXD16 U2470 ( .I(n1357), .ZN(AdrEna[318]) );
  CKND2D0 U2471 ( .A1(\DL3[42].tempL3[4] ), .A2(n26), .ZN(n1359) );
  CKNXD16 U2472 ( .I(n1359), .ZN(AdrEna[676]) );
  CKND2D0 U2473 ( .A1(\DL3[42].tempL3[1] ), .A2(n26), .ZN(n1361) );
  CKNXD16 U2474 ( .I(n1361), .ZN(AdrEna[673]) );
  CKND2D0 U2475 ( .A1(\DL3[19].tempL3[13] ), .A2(n52), .ZN(n1363) );
  CKNXD16 U2476 ( .I(n1363), .ZN(AdrEna[317]) );
  CKND2D0 U2477 ( .A1(\DL3[43].tempL3[0] ), .A2(n25), .ZN(n1365) );
  CKNXD16 U2478 ( .I(n1365), .ZN(AdrEna[688]) );
  CKND2D0 U2479 ( .A1(\DL3[19].tempL3[11] ), .A2(n52), .ZN(n1367) );
  CKNXD16 U2480 ( .I(n1367), .ZN(AdrEna[315]) );
  CKND2D0 U2481 ( .A1(\DL3[19].tempL3[12] ), .A2(n52), .ZN(n1369) );
  CKNXD16 U2482 ( .I(n1369), .ZN(AdrEna[316]) );
  CKND2D0 U2483 ( .A1(\DL3[43].tempL3[2] ), .A2(n25), .ZN(n1371) );
  CKNXD16 U2484 ( .I(n1371), .ZN(AdrEna[690]) );
  CKND2D0 U2485 ( .A1(\DL3[19].tempL3[10] ), .A2(n52), .ZN(n1373) );
  CKNXD16 U2486 ( .I(n1373), .ZN(AdrEna[314]) );
  CKND2D0 U2487 ( .A1(\DL3[43].tempL3[1] ), .A2(n25), .ZN(n1375) );
  CKNXD16 U2488 ( .I(n1375), .ZN(AdrEna[689]) );
  CKND2D0 U2489 ( .A1(\DL3[43].tempL3[3] ), .A2(n25), .ZN(n1377) );
  CKNXD16 U2490 ( .I(n1377), .ZN(AdrEna[691]) );
  CKND2D0 U2491 ( .A1(\DL3[19].tempL3[9] ), .A2(n52), .ZN(n1379) );
  CKNXD16 U2492 ( .I(n1379), .ZN(AdrEna[313]) );
  CKND2D0 U2493 ( .A1(\DL3[43].tempL3[9] ), .A2(n25), .ZN(n1381) );
  CKNXD16 U2494 ( .I(n1381), .ZN(AdrEna[697]) );
  CKND2D0 U2495 ( .A1(\DL3[19].tempL3[7] ), .A2(n52), .ZN(n1383) );
  CKNXD16 U2496 ( .I(n1383), .ZN(AdrEna[311]) );
  CKND2D0 U2497 ( .A1(\DL3[19].tempL3[8] ), .A2(n52), .ZN(n1385) );
  CKNXD16 U2498 ( .I(n1385), .ZN(AdrEna[312]) );
  CKND2D0 U2499 ( .A1(\DL3[42].tempL3[8] ), .A2(n26), .ZN(n1387) );
  CKNXD16 U2500 ( .I(n1387), .ZN(AdrEna[680]) );
  CKND2D0 U2501 ( .A1(\DL3[19].tempL3[4] ), .A2(n52), .ZN(n1389) );
  CKNXD16 U2502 ( .I(n1389), .ZN(AdrEna[308]) );
  CKND2D0 U2503 ( .A1(\DL3[43].tempL3[8] ), .A2(n25), .ZN(n1391) );
  CKNXD16 U2504 ( .I(n1391), .ZN(AdrEna[696]) );
  CKND2D0 U2505 ( .A1(\DL3[44].tempL3[0] ), .A2(n24), .ZN(n1393) );
  CKNXD16 U2506 ( .I(n1393), .ZN(AdrEna[704]) );
  CKND2D0 U2507 ( .A1(\DL3[19].tempL3[5] ), .A2(n52), .ZN(n1395) );
  CKNXD16 U2508 ( .I(n1395), .ZN(AdrEna[309]) );
  CKND2D0 U2509 ( .A1(\DL3[44].tempL3[8] ), .A2(n24), .ZN(n1397) );
  CKNXD16 U2510 ( .I(n1397), .ZN(AdrEna[712]) );
  CKND2D0 U2511 ( .A1(\DL3[19].tempL3[2] ), .A2(n52), .ZN(n1399) );
  CKNXD16 U2512 ( .I(n1399), .ZN(AdrEna[306]) );
  CKND2D0 U2513 ( .A1(\DL3[19].tempL3[3] ), .A2(n52), .ZN(n1401) );
  CKNXD16 U2514 ( .I(n1401), .ZN(AdrEna[307]) );
  CKND2D0 U2515 ( .A1(\DL3[44].tempL3[1] ), .A2(n24), .ZN(n1403) );
  CKNXD16 U2516 ( .I(n1403), .ZN(AdrEna[705]) );
  CKND2D0 U2517 ( .A1(\DL3[19].tempL3[0] ), .A2(n52), .ZN(n1405) );
  CKNXD16 U2518 ( .I(n1405), .ZN(AdrEna[304]) );
  CKND2D0 U2519 ( .A1(\DL3[43].tempL3[4] ), .A2(n25), .ZN(n1407) );
  CKNXD16 U2520 ( .I(n1407), .ZN(AdrEna[692]) );
  CKND2D0 U2521 ( .A1(\DL3[44].tempL3[9] ), .A2(n24), .ZN(n1409) );
  CKNXD16 U2522 ( .I(n1409), .ZN(AdrEna[713]) );
  CKND2D0 U2523 ( .A1(\DL3[19].tempL3[1] ), .A2(n52), .ZN(n1411) );
  CKNXD16 U2524 ( .I(n1411), .ZN(AdrEna[305]) );
  CKND2D0 U2525 ( .A1(\DL3[45].tempL3[0] ), .A2(n23), .ZN(n1413) );
  CKNXD16 U2526 ( .I(n1413), .ZN(AdrEna[720]) );
  CKND2D0 U2527 ( .A1(\DL3[18].tempL3[14] ), .A2(n53), .ZN(n1415) );
  CKNXD16 U2528 ( .I(n1415), .ZN(AdrEna[302]) );
  CKND2D0 U2529 ( .A1(\DL3[18].tempL3[15] ), .A2(n53), .ZN(n1417) );
  CKNXD16 U2530 ( .I(n1417), .ZN(AdrEna[303]) );
  CKND2D0 U2531 ( .A1(\DL3[45].tempL3[2] ), .A2(n23), .ZN(n1419) );
  CKNXD16 U2532 ( .I(n1419), .ZN(AdrEna[722]) );
  CKND2D0 U2533 ( .A1(\DL3[18].tempL3[12] ), .A2(n53), .ZN(n1421) );
  CKNXD16 U2534 ( .I(n1421), .ZN(AdrEna[300]) );
  CKND2D0 U2535 ( .A1(\DL3[45].tempL3[1] ), .A2(n23), .ZN(n1423) );
  CKNXD16 U2536 ( .I(n1423), .ZN(AdrEna[721]) );
  CKND2D0 U2537 ( .A1(\DL3[45].tempL3[3] ), .A2(n23), .ZN(n1425) );
  CKNXD16 U2538 ( .I(n1425), .ZN(AdrEna[723]) );
  CKND2D0 U2539 ( .A1(\DL3[18].tempL3[13] ), .A2(n53), .ZN(n1427) );
  CKNXD16 U2540 ( .I(n1427), .ZN(AdrEna[301]) );
  CKND2D0 U2541 ( .A1(\DL3[45].tempL3[4] ), .A2(n23), .ZN(n1429) );
  CKNXD16 U2542 ( .I(n1429), .ZN(AdrEna[724]) );
  CKND2D0 U2543 ( .A1(\DL3[18].tempL3[10] ), .A2(n53), .ZN(n1431) );
  CKNXD16 U2544 ( .I(n1431), .ZN(AdrEna[298]) );
  CKND2D0 U2545 ( .A1(\DL3[18].tempL3[11] ), .A2(n53), .ZN(n1433) );
  CKNXD16 U2546 ( .I(n1433), .ZN(AdrEna[299]) );
  CKND2D0 U2547 ( .A1(\DL3[44].tempL3[4] ), .A2(n24), .ZN(n1435) );
  CKNXD16 U2548 ( .I(n1435), .ZN(AdrEna[708]) );
  CKND2D0 U2549 ( .A1(\DL3[18].tempL3[8] ), .A2(n53), .ZN(n1437) );
  CKNXD16 U2550 ( .I(n1437), .ZN(AdrEna[296]) );
  CKND2D0 U2551 ( .A1(\DL3[45].tempL3[5] ), .A2(n23), .ZN(n1439) );
  CKNXD16 U2552 ( .I(n1439), .ZN(AdrEna[725]) );
  CKND2D0 U2553 ( .A1(\DL3[46].tempL3[0] ), .A2(n22), .ZN(n1441) );
  CKNXD16 U2554 ( .I(n1441), .ZN(AdrEna[736]) );
  CKND2D0 U2555 ( .A1(\DL3[18].tempL3[9] ), .A2(n53), .ZN(n1443) );
  CKNXD16 U2556 ( .I(n1443), .ZN(AdrEna[297]) );
  CKND2D0 U2557 ( .A1(\DL3[46].tempL3[3] ), .A2(n22), .ZN(n1445) );
  CKNXD16 U2558 ( .I(n1445), .ZN(AdrEna[739]) );
  CKND2D0 U2559 ( .A1(\DL3[18].tempL3[5] ), .A2(n53), .ZN(n1447) );
  CKNXD16 U2560 ( .I(n1447), .ZN(AdrEna[293]) );
  CKND2D0 U2561 ( .A1(\DL3[18].tempL3[7] ), .A2(n53), .ZN(n1449) );
  CKNXD16 U2562 ( .I(n1449), .ZN(AdrEna[295]) );
  CKND2D0 U2563 ( .A1(\DL3[46].tempL3[1] ), .A2(n22), .ZN(n1451) );
  CKNXD16 U2564 ( .I(n1451), .ZN(AdrEna[737]) );
  CKND2D0 U2565 ( .A1(\DL3[18].tempL3[3] ), .A2(n53), .ZN(n1453) );
  CKNXD16 U2566 ( .I(n1453), .ZN(AdrEna[291]) );
  CKND2D0 U2567 ( .A1(\DL3[45].tempL3[8] ), .A2(n23), .ZN(n1455) );
  CKNXD16 U2568 ( .I(n1455), .ZN(AdrEna[728]) );
  CKND2D0 U2569 ( .A1(\DL3[18].tempL3[4] ), .A2(n53), .ZN(n1457) );
  CKNXD16 U2570 ( .I(n1457), .ZN(AdrEna[292]) );
  CKND2D0 U2571 ( .A1(\DL3[46].tempL3[8] ), .A2(n22), .ZN(n1459) );
  CKNXD16 U2572 ( .I(n1459), .ZN(AdrEna[744]) );
  CKND2D0 U2573 ( .A1(\DL3[18].tempL3[1] ), .A2(n53), .ZN(n1461) );
  CKNXD16 U2574 ( .I(n1461), .ZN(AdrEna[289]) );
  CKND2D0 U2575 ( .A1(\DL3[18].tempL3[2] ), .A2(n53), .ZN(n1463) );
  CKNXD16 U2576 ( .I(n1463), .ZN(AdrEna[290]) );
  CKND2D0 U2577 ( .A1(\DL3[47].tempL3[0] ), .A2(n21), .ZN(n1465) );
  CKNXD16 U2578 ( .I(n1465), .ZN(AdrEna[752]) );
  CKND2D0 U2579 ( .A1(\DL3[17].tempL3[15] ), .A2(n54), .ZN(n1467) );
  CKNXD16 U2580 ( .I(n1467), .ZN(AdrEna[287]) );
  CKND2D0 U2581 ( .A1(\DL3[46].tempL3[9] ), .A2(n22), .ZN(n1469) );
  CKNXD16 U2582 ( .I(n1469), .ZN(AdrEna[745]) );
  CKND2D0 U2583 ( .A1(\DL3[46].tempL3[4] ), .A2(n22), .ZN(n1471) );
  CKNXD16 U2584 ( .I(n1471), .ZN(AdrEna[740]) );
  CKND2D0 U2585 ( .A1(\DL3[18].tempL3[0] ), .A2(n53), .ZN(n1473) );
  CKNXD16 U2586 ( .I(n1473), .ZN(AdrEna[288]) );
  CKND2D0 U2587 ( .A1(\DL3[47].tempL3[1] ), .A2(n21), .ZN(n1475) );
  CKNXD16 U2588 ( .I(n1475), .ZN(AdrEna[753]) );
  CKND2D0 U2589 ( .A1(\DL3[17].tempL3[13] ), .A2(n54), .ZN(n1477) );
  CKNXD16 U2590 ( .I(n1477), .ZN(AdrEna[285]) );
  CKND2D0 U2591 ( .A1(\DL3[17].tempL3[14] ), .A2(n54), .ZN(n1479) );
  CKNXD16 U2592 ( .I(n1479), .ZN(AdrEna[286]) );
  CKND2D0 U2593 ( .A1(\DL3[47].tempL3[3] ), .A2(n21), .ZN(n1481) );
  CKNXD16 U2594 ( .I(n1481), .ZN(AdrEna[755]) );
  CKND2D0 U2595 ( .A1(\DL3[17].tempL3[11] ), .A2(n54), .ZN(n1483) );
  CKNXD16 U2596 ( .I(n1483), .ZN(AdrEna[283]) );
  CKND2D0 U2597 ( .A1(\DL3[47].tempL3[4] ), .A2(n21), .ZN(n1485) );
  CKNXD16 U2598 ( .I(n1485), .ZN(AdrEna[756]) );
  CKND2D0 U2599 ( .A1(\DL3[47].tempL3[7] ), .A2(n21), .ZN(n1487) );
  CKNXD16 U2600 ( .I(n1487), .ZN(AdrEna[759]) );
  CKND2D0 U2601 ( .A1(\DL3[17].tempL3[12] ), .A2(n54), .ZN(n1489) );
  CKNXD16 U2602 ( .I(n1489), .ZN(AdrEna[284]) );
  CKND2D0 U2603 ( .A1(\DL3[48].tempL3[0] ), .A2(n20), .ZN(n1491) );
  CKNXD16 U2604 ( .I(n1491), .ZN(AdrEna[768]) );
  CKND2D0 U2605 ( .A1(\DL3[17].tempL3[9] ), .A2(n54), .ZN(n1493) );
  CKNXD16 U2606 ( .I(n1493), .ZN(AdrEna[281]) );
  CKND2D0 U2607 ( .A1(\DL3[17].tempL3[10] ), .A2(n54), .ZN(n1495) );
  CKNXD16 U2608 ( .I(n1495), .ZN(AdrEna[282]) );
  CKND2D0 U2609 ( .A1(\DL3[47].tempL3[5] ), .A2(n21), .ZN(n1497) );
  CKNXD16 U2610 ( .I(n1497), .ZN(AdrEna[757]) );
  CKND2D0 U2611 ( .A1(\DL3[17].tempL3[7] ), .A2(n54), .ZN(n1499) );
  CKNXD16 U2612 ( .I(n1499), .ZN(AdrEna[279]) );
  CKND2D0 U2613 ( .A1(\DL3[47].tempL3[10] ), .A2(n21), .ZN(n1501) );
  CKNXD16 U2614 ( .I(n1501), .ZN(AdrEna[762]) );
  CKND2D0 U2615 ( .A1(\DL3[48].tempL3[1] ), .A2(n20), .ZN(n1503) );
  CKNXD16 U2616 ( .I(n1503), .ZN(AdrEna[769]) );
  CKND2D0 U2617 ( .A1(\DL3[17].tempL3[8] ), .A2(n54), .ZN(n1505) );
  CKNXD16 U2618 ( .I(n1505), .ZN(AdrEna[280]) );
  CKND2D0 U2619 ( .A1(\DL3[48].tempL3[4] ), .A2(n20), .ZN(n1507) );
  CKNXD16 U2620 ( .I(n1507), .ZN(AdrEna[772]) );
  CKND2D0 U2621 ( .A1(\DL3[17].tempL3[4] ), .A2(n54), .ZN(n1509) );
  CKNXD16 U2622 ( .I(n1509), .ZN(AdrEna[276]) );
  CKND2D0 U2623 ( .A1(\DL3[17].tempL3[5] ), .A2(n54), .ZN(n1511) );
  CKNXD16 U2624 ( .I(n1511), .ZN(AdrEna[277]) );
  CKND2D0 U2625 ( .A1(\DL3[48].tempL3[2] ), .A2(n20), .ZN(n1513) );
  CKNXD16 U2626 ( .I(n1513), .ZN(AdrEna[770]) );
  CKND2D0 U2627 ( .A1(\DL3[17].tempL3[3] ), .A2(n54), .ZN(n1515) );
  CKNXD16 U2628 ( .I(n1515), .ZN(AdrEna[275]) );
  CKND2D0 U2629 ( .A1(\DL3[48].tempL3[3] ), .A2(n20), .ZN(n1517) );
  CKNXD16 U2630 ( .I(n1517), .ZN(AdrEna[771]) );
  CKND2D0 U2631 ( .A1(\DL3[48].tempL3[5] ), .A2(n20), .ZN(n1519) );
  CKNXD16 U2632 ( .I(n1519), .ZN(AdrEna[773]) );
  CKND2D0 U2633 ( .A1(\DL3[17].tempL3[2] ), .A2(n54), .ZN(n1521) );
  CKNXD16 U2634 ( .I(n1521), .ZN(AdrEna[274]) );
  CKND2D0 U2635 ( .A1(\DL3[48].tempL3[8] ), .A2(n20), .ZN(n1523) );
  CKNXD16 U2636 ( .I(n1523), .ZN(AdrEna[776]) );
  CKND2D0 U2637 ( .A1(\DL3[17].tempL3[0] ), .A2(n54), .ZN(n1525) );
  CKNXD16 U2638 ( .I(n1525), .ZN(AdrEna[272]) );
  CKND2D0 U2639 ( .A1(\DL3[17].tempL3[1] ), .A2(n54), .ZN(n1527) );
  CKNXD16 U2640 ( .I(n1527), .ZN(AdrEna[273]) );
  CKND2D0 U2641 ( .A1(\DL3[48].tempL3[6] ), .A2(n20), .ZN(n1529) );
  CKNXD16 U2642 ( .I(n1529), .ZN(AdrEna[774]) );
  CKND2D0 U2643 ( .A1(\DL3[16].tempL3[15] ), .A2(n55), .ZN(n1531) );
  CKNXD16 U2644 ( .I(n1531), .ZN(AdrEna[271]) );
  CKND2D0 U2645 ( .A1(\DL3[48].tempL3[7] ), .A2(n20), .ZN(n1533) );
  CKNXD16 U2646 ( .I(n1533), .ZN(AdrEna[775]) );
  CKND2D0 U2647 ( .A1(\DL3[48].tempL3[9] ), .A2(n20), .ZN(n1535) );
  CKNXD16 U2648 ( .I(n1535), .ZN(AdrEna[777]) );
  CKND2D0 U2649 ( .A1(\DL3[16].tempL3[14] ), .A2(n55), .ZN(n1537) );
  CKNXD16 U2650 ( .I(n1537), .ZN(AdrEna[270]) );
  CKAN2D0 U2651 ( .A1(\DL2[1].tempL2[0] ), .A2(DecodedL1[1]), .Z(n55) );
  CKND2D0 U2652 ( .A1(\DL3[48].tempL3[12] ), .A2(n20), .ZN(n1539) );
  CKNXD16 U2653 ( .I(n1539), .ZN(AdrEna[780]) );
  CKND2D0 U2654 ( .A1(\DL3[16].tempL3[12] ), .A2(n55), .ZN(n1541) );
  CKNXD16 U2655 ( .I(n1541), .ZN(AdrEna[268]) );
  CKND2D0 U2656 ( .A1(\DL3[16].tempL3[13] ), .A2(n55), .ZN(n1543) );
  CKNXD16 U2657 ( .I(n1543), .ZN(AdrEna[269]) );
  CKND2D0 U2658 ( .A1(\DL3[48].tempL3[10] ), .A2(n20), .ZN(n1545) );
  CKNXD16 U2659 ( .I(n1545), .ZN(AdrEna[778]) );
  CKND2D0 U2660 ( .A1(\DL3[16].tempL3[11] ), .A2(n55), .ZN(n1547) );
  CKNXD16 U2661 ( .I(n1547), .ZN(AdrEna[267]) );
  CKND2D0 U2662 ( .A1(\DL3[48].tempL3[11] ), .A2(n20), .ZN(n1549) );
  CKNXD16 U2663 ( .I(n1549), .ZN(AdrEna[779]) );
  CKND2D0 U2664 ( .A1(\DL3[48].tempL3[13] ), .A2(n20), .ZN(n1551) );
  CKNXD16 U2665 ( .I(n1551), .ZN(AdrEna[781]) );
  CKND2D0 U2666 ( .A1(\DL3[16].tempL3[10] ), .A2(n55), .ZN(n1553) );
  CKNXD16 U2667 ( .I(n1553), .ZN(AdrEna[266]) );
  CKND2D0 U2668 ( .A1(\DL3[49].tempL3[0] ), .A2(n19), .ZN(n1555) );
  CKNXD16 U2669 ( .I(n1555), .ZN(AdrEna[784]) );
  CKND2D0 U2670 ( .A1(\DL3[16].tempL3[8] ), .A2(n55), .ZN(n1557) );
  CKNXD16 U2671 ( .I(n1557), .ZN(AdrEna[264]) );
  CKND2D0 U2672 ( .A1(\DL3[16].tempL3[9] ), .A2(n55), .ZN(n1559) );
  CKNXD16 U2673 ( .I(n1559), .ZN(AdrEna[265]) );
  CKND2D0 U2674 ( .A1(\DL3[48].tempL3[14] ), .A2(n20), .ZN(n1561) );
  CKNXD16 U2675 ( .I(n1561), .ZN(AdrEna[782]) );
  CKND2D0 U2676 ( .A1(\DL3[16].tempL3[7] ), .A2(n55), .ZN(n1563) );
  CKNXD16 U2677 ( .I(n1563), .ZN(AdrEna[263]) );
  CKND2D0 U2678 ( .A1(\DL3[48].tempL3[15] ), .A2(n20), .ZN(n1565) );
  CKNXD16 U2679 ( .I(n1565), .ZN(AdrEna[783]) );
  CKND2D0 U2680 ( .A1(\DL3[49].tempL3[1] ), .A2(n19), .ZN(n1567) );
  CKNXD16 U2681 ( .I(n1567), .ZN(AdrEna[785]) );
  CKND2D0 U2682 ( .A1(\DL3[16].tempL3[6] ), .A2(n55), .ZN(n1569) );
  CKNXD16 U2683 ( .I(n1569), .ZN(AdrEna[262]) );
  CKND2D0 U2684 ( .A1(\DL3[49].tempL3[4] ), .A2(n19), .ZN(n1571) );
  CKNXD16 U2685 ( .I(n1571), .ZN(AdrEna[788]) );
  CKND2D0 U2686 ( .A1(\DL3[16].tempL3[4] ), .A2(n55), .ZN(n1573) );
  CKNXD16 U2687 ( .I(n1573), .ZN(AdrEna[260]) );
  CKND2D0 U2688 ( .A1(\DL3[16].tempL3[5] ), .A2(n55), .ZN(n1575) );
  CKNXD16 U2689 ( .I(n1575), .ZN(AdrEna[261]) );
  CKND2D0 U2690 ( .A1(\DL3[49].tempL3[2] ), .A2(n19), .ZN(n1577) );
  CKNXD16 U2691 ( .I(n1577), .ZN(AdrEna[786]) );
  CKND2D0 U2692 ( .A1(\DL3[16].tempL3[3] ), .A2(n55), .ZN(n1579) );
  CKNXD16 U2693 ( .I(n1579), .ZN(AdrEna[259]) );
  CKND2D0 U2694 ( .A1(\DL3[49].tempL3[3] ), .A2(n19), .ZN(n1581) );
  CKNXD16 U2695 ( .I(n1581), .ZN(AdrEna[787]) );
  CKND2D0 U2696 ( .A1(\DL3[49].tempL3[5] ), .A2(n19), .ZN(n1583) );
  CKNXD16 U2697 ( .I(n1583), .ZN(AdrEna[789]) );
  CKND2D0 U2698 ( .A1(\DL3[16].tempL3[2] ), .A2(n55), .ZN(n1585) );
  CKNXD16 U2699 ( .I(n1585), .ZN(AdrEna[258]) );
  CKND2D0 U2700 ( .A1(\DL3[49].tempL3[8] ), .A2(n19), .ZN(n1587) );
  CKNXD16 U2701 ( .I(n1587), .ZN(AdrEna[792]) );
  CKND2D0 U2702 ( .A1(\DL3[16].tempL3[0] ), .A2(n55), .ZN(n1589) );
  CKNXD16 U2703 ( .I(n1589), .ZN(AdrEna[256]) );
  CKND2D0 U2704 ( .A1(\DL3[16].tempL3[1] ), .A2(n55), .ZN(n1591) );
  CKNXD16 U2705 ( .I(n1591), .ZN(AdrEna[257]) );
  CKND2D0 U2706 ( .A1(\DL3[49].tempL3[6] ), .A2(n19), .ZN(n1593) );
  CKNXD16 U2707 ( .I(n1593), .ZN(AdrEna[790]) );
  CKND2D0 U2708 ( .A1(\DL3[15].tempL3[12] ), .A2(n56), .ZN(n1595) );
  CKNXD16 U2709 ( .I(n1595), .ZN(AdrEna[252]) );
  CKND2D0 U2710 ( .A1(\DL3[49].tempL3[7] ), .A2(n19), .ZN(n1597) );
  CKNXD16 U2711 ( .I(n1597), .ZN(AdrEna[791]) );
  CKND2D0 U2712 ( .A1(\DL3[49].tempL3[9] ), .A2(n19), .ZN(n1599) );
  CKNXD16 U2713 ( .I(n1599), .ZN(AdrEna[793]) );
  CKND2D0 U2714 ( .A1(\DL3[15].tempL3[11] ), .A2(n56), .ZN(n1601) );
  CKNXD16 U2715 ( .I(n1601), .ZN(AdrEna[251]) );
  CKND2D0 U2716 ( .A1(\DL3[49].tempL3[12] ), .A2(n19), .ZN(n1603) );
  CKNXD16 U2717 ( .I(n1603), .ZN(AdrEna[796]) );
  CKND2D0 U2718 ( .A1(\DL3[15].tempL3[9] ), .A2(n56), .ZN(n1605) );
  CKNXD16 U2719 ( .I(n1605), .ZN(AdrEna[249]) );
  CKND2D0 U2720 ( .A1(\DL3[15].tempL3[10] ), .A2(n56), .ZN(n1607) );
  CKNXD16 U2721 ( .I(n1607), .ZN(AdrEna[250]) );
  CKND2D0 U2722 ( .A1(\DL3[49].tempL3[10] ), .A2(n19), .ZN(n1609) );
  CKNXD16 U2723 ( .I(n1609), .ZN(AdrEna[794]) );
  CKND2D0 U2724 ( .A1(\DL3[15].tempL3[8] ), .A2(n56), .ZN(n1611) );
  CKNXD16 U2725 ( .I(n1611), .ZN(AdrEna[248]) );
  CKND2D0 U2726 ( .A1(\DL3[49].tempL3[11] ), .A2(n19), .ZN(n1613) );
  CKNXD16 U2727 ( .I(n1613), .ZN(AdrEna[795]) );
  CKND2D0 U2728 ( .A1(\DL3[49].tempL3[13] ), .A2(n19), .ZN(n1615) );
  CKNXD16 U2729 ( .I(n1615), .ZN(AdrEna[797]) );
  CKND2D0 U2730 ( .A1(\DL3[15].tempL3[7] ), .A2(n56), .ZN(n1617) );
  CKNXD16 U2731 ( .I(n1617), .ZN(AdrEna[247]) );
  CKND2D0 U2732 ( .A1(\DL3[50].tempL3[0] ), .A2(n17), .ZN(n1619) );
  CKNXD16 U2733 ( .I(n1619), .ZN(AdrEna[800]) );
  CKND2D0 U2734 ( .A1(\DL3[15].tempL3[4] ), .A2(n56), .ZN(n1621) );
  CKNXD16 U2735 ( .I(n1621), .ZN(AdrEna[244]) );
  CKND2D0 U2736 ( .A1(\DL3[15].tempL3[5] ), .A2(n56), .ZN(n1623) );
  CKNXD16 U2737 ( .I(n1623), .ZN(AdrEna[245]) );
  CKND2D0 U2738 ( .A1(\DL3[49].tempL3[14] ), .A2(n19), .ZN(n1625) );
  CKNXD16 U2739 ( .I(n1625), .ZN(AdrEna[798]) );
  CKND2D0 U2740 ( .A1(\DL3[15].tempL3[2] ), .A2(n56), .ZN(n1627) );
  CKNXD16 U2741 ( .I(n1627), .ZN(AdrEna[242]) );
  CKND2D0 U2742 ( .A1(\DL3[49].tempL3[15] ), .A2(n19), .ZN(n1629) );
  CKNXD16 U2743 ( .I(n1629), .ZN(AdrEna[799]) );
  CKND2D0 U2744 ( .A1(\DL3[50].tempL3[1] ), .A2(n17), .ZN(n1631) );
  CKNXD16 U2745 ( .I(n1631), .ZN(AdrEna[801]) );
  CKND2D0 U2746 ( .A1(\DL3[15].tempL3[3] ), .A2(n56), .ZN(n1633) );
  CKNXD16 U2747 ( .I(n1633), .ZN(AdrEna[243]) );
  CKND2D0 U2748 ( .A1(\DL3[50].tempL3[4] ), .A2(n17), .ZN(n1635) );
  CKNXD16 U2749 ( .I(n1635), .ZN(AdrEna[804]) );
  CKND2D0 U2750 ( .A1(\DL3[15].tempL3[0] ), .A2(n56), .ZN(n1637) );
  CKNXD16 U2751 ( .I(n1637), .ZN(AdrEna[240]) );
  CKND2D0 U2752 ( .A1(\DL3[15].tempL3[1] ), .A2(n56), .ZN(n1639) );
  CKNXD16 U2753 ( .I(n1639), .ZN(AdrEna[241]) );
  CKND2D0 U2754 ( .A1(\DL3[50].tempL3[2] ), .A2(n17), .ZN(n1641) );
  CKNXD16 U2755 ( .I(n1641), .ZN(AdrEna[802]) );
  CKND2D0 U2756 ( .A1(\DL3[14].tempL3[11] ), .A2(n57), .ZN(n1643) );
  CKNXD16 U2757 ( .I(n1643), .ZN(AdrEna[235]) );
  CKND2D0 U2758 ( .A1(\DL3[50].tempL3[3] ), .A2(n17), .ZN(n1645) );
  CKNXD16 U2759 ( .I(n1645), .ZN(AdrEna[803]) );
  CKND2D0 U2760 ( .A1(\DL3[50].tempL3[5] ), .A2(n17), .ZN(n1647) );
  CKNXD16 U2761 ( .I(n1647), .ZN(AdrEna[805]) );
  CKND2D0 U2762 ( .A1(\DL3[14].tempL3[12] ), .A2(n57), .ZN(n1649) );
  CKNXD16 U2763 ( .I(n1649), .ZN(AdrEna[236]) );
  CKND2D0 U2764 ( .A1(\DL3[50].tempL3[8] ), .A2(n17), .ZN(n1651) );
  CKNXD16 U2765 ( .I(n1651), .ZN(AdrEna[808]) );
  CKND2D0 U2766 ( .A1(\DL3[14].tempL3[9] ), .A2(n57), .ZN(n1653) );
  CKNXD16 U2767 ( .I(n1653), .ZN(AdrEna[233]) );
  CKND2D0 U2768 ( .A1(\DL3[14].tempL3[10] ), .A2(n57), .ZN(n1655) );
  CKNXD16 U2769 ( .I(n1655), .ZN(AdrEna[234]) );
  CKND2D0 U2770 ( .A1(\DL3[50].tempL3[6] ), .A2(n17), .ZN(n1657) );
  CKNXD16 U2771 ( .I(n1657), .ZN(AdrEna[806]) );
  CKND2D0 U2772 ( .A1(\DL3[14].tempL3[7] ), .A2(n57), .ZN(n1659) );
  CKNXD16 U2773 ( .I(n1659), .ZN(AdrEna[231]) );
  CKND2D0 U2774 ( .A1(\DL3[50].tempL3[7] ), .A2(n17), .ZN(n1661) );
  CKNXD16 U2775 ( .I(n1661), .ZN(AdrEna[807]) );
  CKND2D0 U2776 ( .A1(\DL3[50].tempL3[9] ), .A2(n17), .ZN(n1663) );
  CKNXD16 U2777 ( .I(n1663), .ZN(AdrEna[809]) );
  CKND2D0 U2778 ( .A1(\DL3[14].tempL3[8] ), .A2(n57), .ZN(n1665) );
  CKNXD16 U2779 ( .I(n1665), .ZN(AdrEna[232]) );
  CKND2D0 U2780 ( .A1(\DL3[50].tempL3[12] ), .A2(n17), .ZN(n1667) );
  CKNXD16 U2781 ( .I(n1667), .ZN(AdrEna[812]) );
  CKND2D0 U2782 ( .A1(\DL3[14].tempL3[4] ), .A2(n57), .ZN(n1669) );
  CKNXD16 U2783 ( .I(n1669), .ZN(AdrEna[228]) );
  CKND2D0 U2784 ( .A1(\DL3[14].tempL3[5] ), .A2(n57), .ZN(n1671) );
  CKNXD16 U2785 ( .I(n1671), .ZN(AdrEna[229]) );
  CKND2D0 U2786 ( .A1(\DL3[50].tempL3[10] ), .A2(n17), .ZN(n1673) );
  CKNXD16 U2787 ( .I(n1673), .ZN(AdrEna[810]) );
  CKND2D0 U2788 ( .A1(\DL3[14].tempL3[3] ), .A2(n57), .ZN(n1675) );
  CKNXD16 U2789 ( .I(n1675), .ZN(AdrEna[227]) );
  CKND2D0 U2790 ( .A1(\DL3[50].tempL3[11] ), .A2(n17), .ZN(n1677) );
  CKNXD16 U2791 ( .I(n1677), .ZN(AdrEna[811]) );
  CKND2D0 U2792 ( .A1(\DL3[50].tempL3[13] ), .A2(n17), .ZN(n1679) );
  CKNXD16 U2793 ( .I(n1679), .ZN(AdrEna[813]) );
  CKND2D0 U2794 ( .A1(\DL3[14].tempL3[2] ), .A2(n57), .ZN(n1681) );
  CKNXD16 U2795 ( .I(n1681), .ZN(AdrEna[226]) );
  CKND2D0 U2796 ( .A1(\DL3[52].tempL3[1] ), .A2(n15), .ZN(n1683) );
  CKNXD16 U2797 ( .I(n1683), .ZN(AdrEna[833]) );
  CKND2D0 U2798 ( .A1(\DL3[14].tempL3[0] ), .A2(n57), .ZN(n1685) );
  CKNXD16 U2799 ( .I(n1685), .ZN(AdrEna[224]) );
  CKND2D0 U2800 ( .A1(\DL3[14].tempL3[1] ), .A2(n57), .ZN(n1687) );
  CKNXD16 U2801 ( .I(n1687), .ZN(AdrEna[225]) );
  CKND2D0 U2802 ( .A1(\DL3[50].tempL3[14] ), .A2(n17), .ZN(n1689) );
  CKNXD16 U2803 ( .I(n1689), .ZN(AdrEna[814]) );
  CKND2D0 U2804 ( .A1(\DL3[13].tempL3[12] ), .A2(n58), .ZN(n1691) );
  CKNXD16 U2805 ( .I(n1691), .ZN(AdrEna[220]) );
  CKND2D0 U2806 ( .A1(\DL3[52].tempL3[0] ), .A2(n15), .ZN(n1693) );
  CKNXD16 U2807 ( .I(n1693), .ZN(AdrEna[832]) );
  CKND2D0 U2808 ( .A1(\DL3[52].tempL3[2] ), .A2(n15), .ZN(n1695) );
  CKNXD16 U2809 ( .I(n1695), .ZN(AdrEna[834]) );
  CKND2D0 U2810 ( .A1(\DL3[13].tempL3[11] ), .A2(n58), .ZN(n1697) );
  CKNXD16 U2811 ( .I(n1697), .ZN(AdrEna[219]) );
  CKND2D0 U2812 ( .A1(\DL3[47].tempL3[8] ), .A2(n21), .ZN(n1699) );
  CKNXD16 U2813 ( .I(n1699), .ZN(AdrEna[760]) );
  CKND2D0 U2814 ( .A1(\DL3[13].tempL3[9] ), .A2(n58), .ZN(n1701) );
  CKNXD16 U2815 ( .I(n1701), .ZN(AdrEna[217]) );
  CKND2D0 U2816 ( .A1(\DL3[13].tempL3[10] ), .A2(n58), .ZN(n1703) );
  CKNXD16 U2817 ( .I(n1703), .ZN(AdrEna[218]) );
  CKND2D0 U2818 ( .A1(\DL3[52].tempL3[3] ), .A2(n15), .ZN(n1705) );
  CKNXD16 U2819 ( .I(n1705), .ZN(AdrEna[835]) );
  CKND2D0 U2820 ( .A1(\DL3[13].tempL3[8] ), .A2(n58), .ZN(n1707) );
  CKNXD16 U2821 ( .I(n1707), .ZN(AdrEna[216]) );
  CKND2D0 U2822 ( .A1(\DL3[52].tempL3[4] ), .A2(n15), .ZN(n1709) );
  CKNXD16 U2823 ( .I(n1709), .ZN(AdrEna[836]) );
  CKND2D0 U2824 ( .A1(\DL3[52].tempL3[7] ), .A2(n15), .ZN(n1711) );
  CKNXD16 U2825 ( .I(n1711), .ZN(AdrEna[839]) );
  CKND2D0 U2826 ( .A1(\DL3[13].tempL3[7] ), .A2(n58), .ZN(n1713) );
  CKNXD16 U2827 ( .I(n1713), .ZN(AdrEna[215]) );
  CKND2D0 U2828 ( .A1(\DL3[52].tempL3[8] ), .A2(n15), .ZN(n1715) );
  CKNXD16 U2829 ( .I(n1715), .ZN(AdrEna[840]) );
  CKND2D0 U2830 ( .A1(\DL3[13].tempL3[4] ), .A2(n58), .ZN(n1717) );
  CKNXD16 U2831 ( .I(n1717), .ZN(AdrEna[212]) );
  CKND2D0 U2832 ( .A1(\DL3[13].tempL3[5] ), .A2(n58), .ZN(n1719) );
  CKNXD16 U2833 ( .I(n1719), .ZN(AdrEna[213]) );
  CKND2D0 U2834 ( .A1(\DL3[52].tempL3[10] ), .A2(n15), .ZN(n1721) );
  CKNXD16 U2835 ( .I(n1721), .ZN(AdrEna[842]) );
  CKND2D0 U2836 ( .A1(\DL3[13].tempL3[2] ), .A2(n58), .ZN(n1723) );
  CKNXD16 U2837 ( .I(n1723), .ZN(AdrEna[210]) );
  CKND2D0 U2838 ( .A1(\DL3[52].tempL3[9] ), .A2(n15), .ZN(n1725) );
  CKNXD16 U2839 ( .I(n1725), .ZN(AdrEna[841]) );
  CKND2D0 U2840 ( .A1(\DL3[52].tempL3[11] ), .A2(n15), .ZN(n1727) );
  CKNXD16 U2841 ( .I(n1727), .ZN(AdrEna[843]) );
  CKND2D0 U2842 ( .A1(\DL3[13].tempL3[3] ), .A2(n58), .ZN(n1729) );
  CKNXD16 U2843 ( .I(n1729), .ZN(AdrEna[211]) );
  CKND2D0 U2844 ( .A1(\DL3[52].tempL3[12] ), .A2(n15), .ZN(n1731) );
  CKNXD16 U2845 ( .I(n1731), .ZN(AdrEna[844]) );
  CKND2D0 U2846 ( .A1(\DL3[13].tempL3[0] ), .A2(n58), .ZN(n1733) );
  CKNXD16 U2847 ( .I(n1733), .ZN(AdrEna[208]) );
  CKND2D0 U2848 ( .A1(\DL3[13].tempL3[1] ), .A2(n58), .ZN(n1735) );
  CKNXD16 U2849 ( .I(n1735), .ZN(AdrEna[209]) );
  CKND2D0 U2850 ( .A1(\DL3[52].tempL3[14] ), .A2(n15), .ZN(n1737) );
  CKNXD16 U2851 ( .I(n1737), .ZN(AdrEna[846]) );
  CKND2D0 U2852 ( .A1(\DL3[12].tempL3[11] ), .A2(n59), .ZN(n1739) );
  CKNXD16 U2853 ( .I(n1739), .ZN(AdrEna[203]) );
  CKND2D0 U2854 ( .A1(\DL3[52].tempL3[13] ), .A2(n15), .ZN(n1741) );
  CKNXD16 U2855 ( .I(n1741), .ZN(AdrEna[845]) );
  CKND2D0 U2856 ( .A1(\DL3[52].tempL3[15] ), .A2(n15), .ZN(n1743) );
  CKNXD16 U2857 ( .I(n1743), .ZN(AdrEna[847]) );
  CKND2D0 U2858 ( .A1(\DL3[12].tempL3[12] ), .A2(n59), .ZN(n1745) );
  CKNXD16 U2859 ( .I(n1745), .ZN(AdrEna[204]) );
  CKND2D0 U2860 ( .A1(\DL3[53].tempL3[0] ), .A2(n14), .ZN(n1747) );
  CKNXD16 U2861 ( .I(n1747), .ZN(AdrEna[848]) );
  CKND2D0 U2862 ( .A1(\DL3[12].tempL3[9] ), .A2(n59), .ZN(n1749) );
  CKNXD16 U2863 ( .I(n1749), .ZN(AdrEna[201]) );
  CKND2D0 U2864 ( .A1(\DL3[12].tempL3[10] ), .A2(n59), .ZN(n1751) );
  CKNXD16 U2865 ( .I(n1751), .ZN(AdrEna[202]) );
  CKND2D0 U2866 ( .A1(\DL3[53].tempL3[2] ), .A2(n14), .ZN(n1753) );
  CKNXD16 U2867 ( .I(n1753), .ZN(AdrEna[850]) );
  CKND2D0 U2868 ( .A1(\DL3[12].tempL3[7] ), .A2(n59), .ZN(n1755) );
  CKNXD16 U2869 ( .I(n1755), .ZN(AdrEna[199]) );
  CKND2D0 U2870 ( .A1(\DL3[53].tempL3[1] ), .A2(n14), .ZN(n1757) );
  CKNXD16 U2871 ( .I(n1757), .ZN(AdrEna[849]) );
  CKND2D0 U2872 ( .A1(\DL3[53].tempL3[3] ), .A2(n14), .ZN(n1759) );
  CKNXD16 U2873 ( .I(n1759), .ZN(AdrEna[851]) );
  CKND2D0 U2874 ( .A1(\DL3[12].tempL3[8] ), .A2(n59), .ZN(n1761) );
  CKNXD16 U2875 ( .I(n1761), .ZN(AdrEna[200]) );
  CKND2D0 U2876 ( .A1(\DL3[53].tempL3[4] ), .A2(n14), .ZN(n1763) );
  CKNXD16 U2877 ( .I(n1763), .ZN(AdrEna[852]) );
  CKND2D0 U2878 ( .A1(\DL3[12].tempL3[4] ), .A2(n59), .ZN(n1765) );
  CKNXD16 U2879 ( .I(n1765), .ZN(AdrEna[196]) );
  CKND2D0 U2880 ( .A1(\DL3[12].tempL3[5] ), .A2(n59), .ZN(n1767) );
  CKNXD16 U2881 ( .I(n1767), .ZN(AdrEna[197]) );
  CKND2D0 U2882 ( .A1(\DL3[53].tempL3[7] ), .A2(n14), .ZN(n1769) );
  CKNXD16 U2883 ( .I(n1769), .ZN(AdrEna[855]) );
  CKND2D0 U2884 ( .A1(\DL3[12].tempL3[3] ), .A2(n59), .ZN(n1771) );
  CKNXD16 U2885 ( .I(n1771), .ZN(AdrEna[195]) );
  CKND2D0 U2886 ( .A1(\DL3[52].tempL3[5] ), .A2(n15), .ZN(n1773) );
  CKNXD16 U2887 ( .I(n1773), .ZN(AdrEna[837]) );
  CKND2D0 U2888 ( .A1(\DL3[53].tempL3[8] ), .A2(n14), .ZN(n1775) );
  CKNXD16 U2889 ( .I(n1775), .ZN(AdrEna[856]) );
  CKND2D0 U2890 ( .A1(\DL3[12].tempL3[2] ), .A2(n59), .ZN(n1777) );
  CKNXD16 U2891 ( .I(n1777), .ZN(AdrEna[194]) );
  CKND2D0 U2892 ( .A1(\DL3[53].tempL3[11] ), .A2(n14), .ZN(n1779) );
  CKNXD16 U2893 ( .I(n1779), .ZN(AdrEna[859]) );
  CKND2D0 U2894 ( .A1(\DL3[12].tempL3[0] ), .A2(n59), .ZN(n1781) );
  CKNXD16 U2895 ( .I(n1781), .ZN(AdrEna[192]) );
  CKND2D0 U2896 ( .A1(\DL3[12].tempL3[1] ), .A2(n59), .ZN(n1783) );
  CKNXD16 U2897 ( .I(n1783), .ZN(AdrEna[193]) );
  CKND2D0 U2898 ( .A1(\DL3[53].tempL3[9] ), .A2(n14), .ZN(n1785) );
  CKNXD16 U2899 ( .I(n1785), .ZN(AdrEna[857]) );
  CKND2D0 U2900 ( .A1(\DL3[11].tempL3[12] ), .A2(n60), .ZN(n1787) );
  CKNXD16 U2901 ( .I(n1787), .ZN(AdrEna[188]) );
  CKND2D0 U2902 ( .A1(\DL3[53].tempL3[10] ), .A2(n14), .ZN(n1789) );
  CKNXD16 U2903 ( .I(n1789), .ZN(AdrEna[858]) );
  CKND2D0 U2904 ( .A1(\DL3[53].tempL3[12] ), .A2(n14), .ZN(n1791) );
  CKNXD16 U2905 ( .I(n1791), .ZN(AdrEna[860]) );
  CKND2D0 U2906 ( .A1(\DL3[11].tempL3[6] ), .A2(n60), .ZN(n1793) );
  CKNXD16 U2907 ( .I(n1793), .ZN(AdrEna[182]) );
  CKND2D0 U2908 ( .A1(\DL3[53].tempL3[15] ), .A2(n14), .ZN(n1795) );
  CKNXD16 U2909 ( .I(n1795), .ZN(AdrEna[863]) );
  CKND2D0 U2910 ( .A1(\DL3[11].tempL3[7] ), .A2(n60), .ZN(n1797) );
  CKNXD16 U2911 ( .I(n1797), .ZN(AdrEna[183]) );
  CKND2D0 U2912 ( .A1(\DL3[11].tempL3[5] ), .A2(n60), .ZN(n1799) );
  CKNXD16 U2913 ( .I(n1799), .ZN(AdrEna[181]) );
  CKND2D0 U2914 ( .A1(\DL3[53].tempL3[13] ), .A2(n14), .ZN(n1801) );
  CKNXD16 U2915 ( .I(n1801), .ZN(AdrEna[861]) );
  CKND2D0 U2916 ( .A1(\DL3[11].tempL3[4] ), .A2(n60), .ZN(n1803) );
  CKNXD16 U2917 ( .I(n1803), .ZN(AdrEna[180]) );
  CKND2D0 U2918 ( .A1(\DL3[53].tempL3[14] ), .A2(n14), .ZN(n1805) );
  CKNXD16 U2919 ( .I(n1805), .ZN(AdrEna[862]) );
  CKND2D0 U2920 ( .A1(\DL3[54].tempL3[0] ), .A2(n13), .ZN(n1807) );
  CKNXD16 U2921 ( .I(n1807), .ZN(AdrEna[864]) );
  CKND2D0 U2922 ( .A1(\DL3[11].tempL3[2] ), .A2(n60), .ZN(n1809) );
  CKNXD16 U2923 ( .I(n1809), .ZN(AdrEna[178]) );
  CKND2D0 U2924 ( .A1(\DL3[54].tempL3[3] ), .A2(n13), .ZN(n1811) );
  CKNXD16 U2925 ( .I(n1811), .ZN(AdrEna[867]) );
  CKND2D0 U2926 ( .A1(\DL3[11].tempL3[3] ), .A2(n60), .ZN(n1813) );
  CKNXD16 U2927 ( .I(n1813), .ZN(AdrEna[179]) );
  CKND2D0 U2928 ( .A1(\DL3[11].tempL3[1] ), .A2(n60), .ZN(n1815) );
  CKNXD16 U2929 ( .I(n1815), .ZN(AdrEna[177]) );
  CKND2D0 U2930 ( .A1(\DL3[54].tempL3[1] ), .A2(n13), .ZN(n1817) );
  CKNXD16 U2931 ( .I(n1817), .ZN(AdrEna[865]) );
  CKND2D0 U2932 ( .A1(\DL3[54].tempL3[2] ), .A2(n13), .ZN(n1819) );
  CKNXD16 U2933 ( .I(n1819), .ZN(AdrEna[866]) );
  CKND2D0 U2934 ( .A1(\DL3[54].tempL3[4] ), .A2(n13), .ZN(n1821) );
  CKNXD16 U2935 ( .I(n1821), .ZN(AdrEna[868]) );
  CKND2D0 U2936 ( .A1(\DL3[11].tempL3[0] ), .A2(n60), .ZN(n1823) );
  CKNXD16 U2937 ( .I(n1823), .ZN(AdrEna[176]) );
  CKND2D0 U2938 ( .A1(\DL3[53].tempL3[5] ), .A2(n14), .ZN(n1825) );
  CKNXD16 U2939 ( .I(n1825), .ZN(AdrEna[853]) );
  CKND2D0 U2940 ( .A1(\DL3[10].tempL3[12] ), .A2(n61), .ZN(n1827) );
  CKNXD16 U2941 ( .I(n1827), .ZN(AdrEna[172]) );
  CKND2D0 U2942 ( .A1(\DL3[10].tempL3[8] ), .A2(n61), .ZN(n1829) );
  CKNXD16 U2943 ( .I(n1829), .ZN(AdrEna[168]) );
  CKND2D0 U2944 ( .A1(\DL3[54].tempL3[8] ), .A2(n13), .ZN(n1831) );
  CKNXD16 U2945 ( .I(n1831), .ZN(AdrEna[872]) );
  CKND2D0 U2946 ( .A1(\DL3[10].tempL3[7] ), .A2(n61), .ZN(n1833) );
  CKNXD16 U2947 ( .I(n1833), .ZN(AdrEna[167]) );
  CKND2D0 U2948 ( .A1(\DL3[54].tempL3[7] ), .A2(n13), .ZN(n1835) );
  CKNXD16 U2949 ( .I(n1835), .ZN(AdrEna[871]) );
  CKND2D0 U2950 ( .A1(\DL3[54].tempL3[9] ), .A2(n13), .ZN(n1837) );
  CKNXD16 U2951 ( .I(n1837), .ZN(AdrEna[873]) );
  CKND2D0 U2952 ( .A1(\DL3[10].tempL3[5] ), .A2(n61), .ZN(n1839) );
  CKNXD16 U2953 ( .I(n1839), .ZN(AdrEna[165]) );
  CKND2D0 U2954 ( .A1(\DL3[54].tempL3[10] ), .A2(n13), .ZN(n1841) );
  CKNXD16 U2955 ( .I(n1841), .ZN(AdrEna[874]) );
  CKND2D0 U2956 ( .A1(\DL3[10].tempL3[6] ), .A2(n61), .ZN(n1843) );
  CKNXD16 U2957 ( .I(n1843), .ZN(AdrEna[166]) );
  CKND2D0 U2958 ( .A1(\DL3[10].tempL3[4] ), .A2(n61), .ZN(n1845) );
  CKNXD16 U2959 ( .I(n1845), .ZN(AdrEna[164]) );
  CKND2D0 U2960 ( .A1(\DL3[54].tempL3[12] ), .A2(n13), .ZN(n1847) );
  CKNXD16 U2961 ( .I(n1847), .ZN(AdrEna[876]) );
  CKND2D0 U2962 ( .A1(\DL3[10].tempL3[3] ), .A2(n61), .ZN(n1849) );
  CKNXD16 U2963 ( .I(n1849), .ZN(AdrEna[163]) );
  CKND2D0 U2964 ( .A1(\DL3[54].tempL3[11] ), .A2(n13), .ZN(n1851) );
  CKNXD16 U2965 ( .I(n1851), .ZN(AdrEna[875]) );
  CKND2D0 U2966 ( .A1(\DL3[54].tempL3[13] ), .A2(n13), .ZN(n1853) );
  CKNXD16 U2967 ( .I(n1853), .ZN(AdrEna[877]) );
  CKND2D0 U2968 ( .A1(\DL3[10].tempL3[1] ), .A2(n61), .ZN(n1855) );
  CKNXD16 U2969 ( .I(n1855), .ZN(AdrEna[161]) );
  CKND2D0 U2970 ( .A1(\DL3[54].tempL3[14] ), .A2(n13), .ZN(n1857) );
  CKNXD16 U2971 ( .I(n1857), .ZN(AdrEna[878]) );
  CKND2D0 U2972 ( .A1(\DL3[10].tempL3[2] ), .A2(n61), .ZN(n1859) );
  CKNXD16 U2973 ( .I(n1859), .ZN(AdrEna[162]) );
  CKND2D0 U2974 ( .A1(\DL3[10].tempL3[0] ), .A2(n61), .ZN(n1861) );
  CKNXD16 U2975 ( .I(n1861), .ZN(AdrEna[160]) );
  CKND2D0 U2976 ( .A1(\DL3[55].tempL3[0] ), .A2(n12), .ZN(n1863) );
  CKNXD16 U2977 ( .I(n1863), .ZN(AdrEna[880]) );
  CKND2D0 U2978 ( .A1(\DL3[9].tempL3[12] ), .A2(n62), .ZN(n1865) );
  CKNXD16 U2979 ( .I(n1865), .ZN(AdrEna[156]) );
  CKND2D0 U2980 ( .A1(\DL3[54].tempL3[15] ), .A2(n13), .ZN(n1867) );
  CKNXD16 U2981 ( .I(n1867), .ZN(AdrEna[879]) );
  CKND2D0 U2982 ( .A1(\DL3[55].tempL3[1] ), .A2(n12), .ZN(n1869) );
  CKNXD16 U2983 ( .I(n1869), .ZN(AdrEna[881]) );
  CKND2D0 U2984 ( .A1(\DL3[9].tempL3[8] ), .A2(n62), .ZN(n1871) );
  CKNXD16 U2985 ( .I(n1871), .ZN(AdrEna[152]) );
  CKND2D0 U2986 ( .A1(\DL3[55].tempL3[2] ), .A2(n12), .ZN(n1873) );
  CKNXD16 U2987 ( .I(n1873), .ZN(AdrEna[882]) );
  CKND2D0 U2988 ( .A1(\DL3[9].tempL3[10] ), .A2(n62), .ZN(n1875) );
  CKNXD16 U2989 ( .I(n1875), .ZN(AdrEna[154]) );
  CKND2D0 U2990 ( .A1(\DL3[9].tempL3[7] ), .A2(n62), .ZN(n1877) );
  CKNXD16 U2991 ( .I(n1877), .ZN(AdrEna[151]) );
  CKND2D0 U2992 ( .A1(\DL3[55].tempL3[4] ), .A2(n12), .ZN(n1879) );
  CKNXD16 U2993 ( .I(n1879), .ZN(AdrEna[884]) );
  CKND2D0 U2994 ( .A1(\DL3[9].tempL3[3] ), .A2(n62), .ZN(n1881) );
  CKNXD16 U2995 ( .I(n1881), .ZN(AdrEna[147]) );
  CKND2D0 U2996 ( .A1(\DL3[55].tempL3[3] ), .A2(n12), .ZN(n1883) );
  CKNXD16 U2997 ( .I(n1883), .ZN(AdrEna[883]) );
  CKND2D0 U2998 ( .A1(\DL3[54].tempL3[5] ), .A2(n13), .ZN(n1885) );
  CKNXD16 U2999 ( .I(n1885), .ZN(AdrEna[869]) );
  CKND2D0 U3000 ( .A1(\DL3[9].tempL3[6] ), .A2(n62), .ZN(n1887) );
  CKNXD16 U3001 ( .I(n1887), .ZN(AdrEna[150]) );
  CKND2D0 U3002 ( .A1(\DL3[55].tempL3[9] ), .A2(n12), .ZN(n1889) );
  CKNXD16 U3003 ( .I(n1889), .ZN(AdrEna[889]) );
  CKND2D0 U3004 ( .A1(\DL3[9].tempL3[4] ), .A2(n62), .ZN(n1891) );
  CKNXD16 U3005 ( .I(n1891), .ZN(AdrEna[148]) );
  CKND2D0 U3006 ( .A1(\DL3[9].tempL3[2] ), .A2(n62), .ZN(n1893) );
  CKNXD16 U3007 ( .I(n1893), .ZN(AdrEna[146]) );
  CKND2D0 U3008 ( .A1(\DL3[55].tempL3[7] ), .A2(n12), .ZN(n1895) );
  CKNXD16 U3009 ( .I(n1895), .ZN(AdrEna[887]) );
  CKND2D0 U3010 ( .A1(\DL3[9].tempL3[1] ), .A2(n62), .ZN(n1897) );
  CKNXD16 U3011 ( .I(n1897), .ZN(AdrEna[145]) );
  CKND2D0 U3012 ( .A1(\DL3[55].tempL3[8] ), .A2(n12), .ZN(n1899) );
  CKNXD16 U3013 ( .I(n1899), .ZN(AdrEna[888]) );
  CKND2D0 U3014 ( .A1(\DL3[55].tempL3[10] ), .A2(n12), .ZN(n1901) );
  CKNXD16 U3015 ( .I(n1901), .ZN(AdrEna[890]) );
  CKND2D0 U3016 ( .A1(\DL3[8].tempL3[12] ), .A2(n63), .ZN(n1903) );
  CKNXD16 U3017 ( .I(n1903), .ZN(AdrEna[140]) );
  CKND2D0 U3018 ( .A1(\DL3[55].tempL3[13] ), .A2(n12), .ZN(n1905) );
  CKNXD16 U3019 ( .I(n1905), .ZN(AdrEna[893]) );
  CKND2D0 U3020 ( .A1(\DL3[9].tempL3[0] ), .A2(n62), .ZN(n1907) );
  CKNXD16 U3021 ( .I(n1907), .ZN(AdrEna[144]) );
  CKND2D0 U3022 ( .A1(\DL3[8].tempL3[10] ), .A2(n63), .ZN(n1909) );
  CKNXD16 U3023 ( .I(n1909), .ZN(AdrEna[138]) );
  CKND2D0 U3024 ( .A1(\DL3[55].tempL3[11] ), .A2(n12), .ZN(n1911) );
  CKNXD16 U3025 ( .I(n1911), .ZN(AdrEna[891]) );
  CKND2D0 U3026 ( .A1(\DL3[8].tempL3[6] ), .A2(n63), .ZN(n1913) );
  CKNXD16 U3027 ( .I(n1913), .ZN(AdrEna[134]) );
  CKND2D0 U3028 ( .A1(\DL3[55].tempL3[12] ), .A2(n12), .ZN(n1915) );
  CKNXD16 U3029 ( .I(n1915), .ZN(AdrEna[892]) );
  CKND2D0 U3030 ( .A1(\DL3[55].tempL3[14] ), .A2(n12), .ZN(n1917) );
  CKNXD16 U3031 ( .I(n1917), .ZN(AdrEna[894]) );
  CKND2D0 U3032 ( .A1(\DL3[8].tempL3[8] ), .A2(n63), .ZN(n1919) );
  CKNXD16 U3033 ( .I(n1919), .ZN(AdrEna[136]) );
  CKND2D0 U3034 ( .A1(\DL3[56].tempL3[1] ), .A2(n11), .ZN(n1921) );
  CKNXD16 U3035 ( .I(n1921), .ZN(AdrEna[897]) );
  CKND2D0 U3036 ( .A1(\DL3[8].tempL3[7] ), .A2(n63), .ZN(n1923) );
  CKNXD16 U3037 ( .I(n1923), .ZN(AdrEna[135]) );
  CKND2D0 U3038 ( .A1(\DL3[8].tempL3[5] ), .A2(n63), .ZN(n1925) );
  CKNXD16 U3039 ( .I(n1925), .ZN(AdrEna[133]) );
  CKND2D0 U3040 ( .A1(\DL3[55].tempL3[15] ), .A2(n12), .ZN(n1927) );
  CKNXD16 U3041 ( .I(n1927), .ZN(AdrEna[895]) );
  CKND2D0 U3042 ( .A1(\DL3[8].tempL3[2] ), .A2(n63), .ZN(n1929) );
  CKNXD16 U3043 ( .I(n1929), .ZN(AdrEna[130]) );
  CKND2D0 U3044 ( .A1(\DL3[56].tempL3[0] ), .A2(n11), .ZN(n1931) );
  CKNXD16 U3045 ( .I(n1931), .ZN(AdrEna[896]) );
  CKND2D0 U3046 ( .A1(\DL3[56].tempL3[2] ), .A2(n11), .ZN(n1933) );
  CKNXD16 U3047 ( .I(n1933), .ZN(AdrEna[898]) );
  CKND2D0 U3048 ( .A1(\DL3[8].tempL3[4] ), .A2(n63), .ZN(n1935) );
  CKNXD16 U3049 ( .I(n1935), .ZN(AdrEna[132]) );
  CKND2D0 U3050 ( .A1(\DL3[55].tempL3[5] ), .A2(n12), .ZN(n1937) );
  CKNXD16 U3051 ( .I(n1937), .ZN(AdrEna[885]) );
  CKND2D0 U3052 ( .A1(\DL3[8].tempL3[3] ), .A2(n63), .ZN(n1939) );
  CKNXD16 U3053 ( .I(n1939), .ZN(AdrEna[131]) );
  CKND2D0 U3054 ( .A1(\DL3[8].tempL3[1] ), .A2(n63), .ZN(n1941) );
  CKNXD16 U3055 ( .I(n1941), .ZN(AdrEna[129]) );
  CKND2D0 U3056 ( .A1(\DL3[56].tempL3[3] ), .A2(n11), .ZN(n1943) );
  CKNXD16 U3057 ( .I(n1943), .ZN(AdrEna[899]) );
  CKND2D0 U3058 ( .A1(\DL3[7].tempL3[10] ), .A2(n64), .ZN(n1945) );
  CKNXD16 U3059 ( .I(n1945), .ZN(AdrEna[122]) );
  CKND2D0 U3060 ( .A1(\DL3[56].tempL3[4] ), .A2(n11), .ZN(n1947) );
  CKNXD16 U3061 ( .I(n1947), .ZN(AdrEna[900]) );
  CKND2D0 U3062 ( .A1(\DL3[56].tempL3[7] ), .A2(n11), .ZN(n1949) );
  CKNXD16 U3063 ( .I(n1949), .ZN(AdrEna[903]) );
  CKND2D0 U3064 ( .A1(\DL3[8].tempL3[0] ), .A2(n63), .ZN(n1951) );
  CKNXD16 U3065 ( .I(n1951), .ZN(AdrEna[128]) );
  CKND2D0 U3066 ( .A1(\DL3[56].tempL3[11] ), .A2(n11), .ZN(n1953) );
  CKNXD16 U3067 ( .I(n1953), .ZN(AdrEna[907]) );
  CKND2D0 U3068 ( .A1(\DL3[7].tempL3[12] ), .A2(n64), .ZN(n1955) );
  CKNXD16 U3069 ( .I(n1955), .ZN(AdrEna[124]) );
  CKND2D0 U3070 ( .A1(\DL3[7].tempL3[8] ), .A2(n64), .ZN(n1957) );
  CKNXD16 U3071 ( .I(n1957), .ZN(AdrEna[120]) );
  CKND2D0 U3072 ( .A1(\DL3[56].tempL3[5] ), .A2(n11), .ZN(n1959) );
  CKNXD16 U3073 ( .I(n1959), .ZN(AdrEna[901]) );
  CKND2D0 U3074 ( .A1(\DL3[7].tempL3[7] ), .A2(n64), .ZN(n1961) );
  CKNXD16 U3075 ( .I(n1961), .ZN(AdrEna[119]) );
  CKND2D0 U3076 ( .A1(\DL3[56].tempL3[10] ), .A2(n11), .ZN(n1963) );
  CKNXD16 U3077 ( .I(n1963), .ZN(AdrEna[906]) );
  CKND2D0 U3078 ( .A1(\DL3[56].tempL3[12] ), .A2(n11), .ZN(n1965) );
  CKNXD16 U3079 ( .I(n1965), .ZN(AdrEna[908]) );
  CKND2D0 U3080 ( .A1(\DL3[7].tempL3[5] ), .A2(n64), .ZN(n1967) );
  CKNXD16 U3081 ( .I(n1967), .ZN(AdrEna[117]) );
  CKND2D0 U3082 ( .A1(\DL3[56].tempL3[15] ), .A2(n11), .ZN(n1969) );
  CKNXD16 U3083 ( .I(n1969), .ZN(AdrEna[911]) );
  CKND2D0 U3084 ( .A1(\DL3[7].tempL3[6] ), .A2(n64), .ZN(n1971) );
  CKNXD16 U3085 ( .I(n1971), .ZN(AdrEna[118]) );
  CKND2D0 U3086 ( .A1(\DL3[7].tempL3[4] ), .A2(n64), .ZN(n1973) );
  CKNXD16 U3087 ( .I(n1973), .ZN(AdrEna[116]) );
  CKND2D0 U3088 ( .A1(\DL3[56].tempL3[13] ), .A2(n11), .ZN(n1975) );
  CKNXD16 U3089 ( .I(n1975), .ZN(AdrEna[909]) );
  CKND2D0 U3090 ( .A1(\DL3[7].tempL3[3] ), .A2(n64), .ZN(n1977) );
  CKNXD16 U3091 ( .I(n1977), .ZN(AdrEna[115]) );
  CKND2D0 U3092 ( .A1(\DL3[56].tempL3[14] ), .A2(n11), .ZN(n1979) );
  CKNXD16 U3093 ( .I(n1979), .ZN(AdrEna[910]) );
  CKND2D0 U3094 ( .A1(\DL3[57].tempL3[0] ), .A2(n10), .ZN(n1981) );
  CKNXD16 U3095 ( .I(n1981), .ZN(AdrEna[912]) );
  CKND2D0 U3096 ( .A1(\DL3[7].tempL3[1] ), .A2(n64), .ZN(n1983) );
  CKNXD16 U3097 ( .I(n1983), .ZN(AdrEna[113]) );
  CKND2D0 U3098 ( .A1(\DL3[57].tempL3[3] ), .A2(n10), .ZN(n1985) );
  CKNXD16 U3099 ( .I(n1985), .ZN(AdrEna[915]) );
  CKND2D0 U3100 ( .A1(\DL3[7].tempL3[2] ), .A2(n64), .ZN(n1987) );
  CKNXD16 U3101 ( .I(n1987), .ZN(AdrEna[114]) );
  CKND2D0 U3102 ( .A1(\DL3[7].tempL3[0] ), .A2(n64), .ZN(n1989) );
  CKNXD16 U3103 ( .I(n1989), .ZN(AdrEna[112]) );
  CKND2D0 U3104 ( .A1(\DL3[57].tempL3[1] ), .A2(n10), .ZN(n1991) );
  CKNXD16 U3105 ( .I(n1991), .ZN(AdrEna[913]) );
  CKND2D0 U3106 ( .A1(\DL3[6].tempL3[12] ), .A2(n3), .ZN(n1993) );
  CKNXD16 U3107 ( .I(n1993), .ZN(AdrEna[108]) );
  CKND2D0 U3108 ( .A1(\DL3[57].tempL3[2] ), .A2(n10), .ZN(n1995) );
  CKNXD16 U3109 ( .I(n1995), .ZN(AdrEna[914]) );
  CKND2D0 U3110 ( .A1(\DL3[57].tempL3[4] ), .A2(n10), .ZN(n1997) );
  CKNXD16 U3111 ( .I(n1997), .ZN(AdrEna[916]) );
  CKND2D0 U3112 ( .A1(\DL3[6].tempL3[8] ), .A2(n3), .ZN(n1999) );
  CKNXD16 U3113 ( .I(n1999), .ZN(AdrEna[104]) );
  CKND2D0 U3114 ( .A1(\DL3[56].tempL3[8] ), .A2(n11), .ZN(n2001) );
  CKNXD16 U3115 ( .I(n2001), .ZN(AdrEna[904]) );
  CKND2D0 U3116 ( .A1(\DL3[6].tempL3[10] ), .A2(n3), .ZN(n2003) );
  CKNXD16 U3117 ( .I(n2003), .ZN(AdrEna[106]) );
  CKND2D0 U3118 ( .A1(\DL3[6].tempL3[7] ), .A2(n3), .ZN(n2005) );
  CKNXD16 U3119 ( .I(n2005), .ZN(AdrEna[103]) );
  CKND2D0 U3120 ( .A1(\DL3[57].tempL3[5] ), .A2(n10), .ZN(n2007) );
  CKNXD16 U3121 ( .I(n2007), .ZN(AdrEna[917]) );
  CKND2D0 U3122 ( .A1(\DL3[6].tempL3[4] ), .A2(n3), .ZN(n2009) );
  CKNXD16 U3123 ( .I(n2009), .ZN(AdrEna[100]) );
  CKND2D0 U3124 ( .A1(\DL3[57].tempL3[7] ), .A2(n10), .ZN(n2011) );
  CKNXD16 U3125 ( .I(n2011), .ZN(AdrEna[919]) );
  CKND2D0 U3126 ( .A1(\DL3[57].tempL3[10] ), .A2(n10), .ZN(n2013) );
  CKNXD16 U3127 ( .I(n2013), .ZN(AdrEna[922]) );
  CKND2D0 U3128 ( .A1(\DL3[6].tempL3[6] ), .A2(n3), .ZN(n2015) );
  CKNXD16 U3129 ( .I(n2015), .ZN(AdrEna[102]) );
  CKND2D0 U3130 ( .A1(\DL3[57].tempL3[13] ), .A2(n10), .ZN(n2017) );
  CKNXD16 U3131 ( .I(n2017), .ZN(AdrEna[925]) );
  CKND2D0 U3132 ( .A1(\DL3[6].tempL3[5] ), .A2(n3), .ZN(n2019) );
  CKNXD16 U3133 ( .I(n2019), .ZN(AdrEna[101]) );
  CKND2D0 U3134 ( .A1(\DL3[6].tempL3[3] ), .A2(n3), .ZN(n2021) );
  CKNXD16 U3135 ( .I(n2021), .ZN(AdrEna[99]) );
  CKND2D0 U3136 ( .A1(\DL3[57].tempL3[11] ), .A2(n10), .ZN(n2023) );
  CKNXD16 U3137 ( .I(n2023), .ZN(AdrEna[923]) );
  CKND2D0 U3138 ( .A1(\DL3[6].tempL3[0] ), .A2(n3), .ZN(n2025) );
  CKNXD16 U3139 ( .I(n2025), .ZN(AdrEna[96]) );
  CKND2D0 U3140 ( .A1(\DL3[57].tempL3[12] ), .A2(n10), .ZN(n2027) );
  CKNXD16 U3141 ( .I(n2027), .ZN(AdrEna[924]) );
  CKND2D0 U3142 ( .A1(\DL3[57].tempL3[14] ), .A2(n10), .ZN(n2029) );
  CKNXD16 U3143 ( .I(n2029), .ZN(AdrEna[926]) );
  CKND2D0 U3144 ( .A1(\DL3[6].tempL3[2] ), .A2(n3), .ZN(n2031) );
  CKNXD16 U3145 ( .I(n2031), .ZN(AdrEna[98]) );
  CKND2D0 U3146 ( .A1(\DL3[58].tempL3[3] ), .A2(n9), .ZN(n2033) );
  CKNXD16 U3147 ( .I(n2033), .ZN(AdrEna[931]) );
  CKND2D0 U3148 ( .A1(\DL3[6].tempL3[1] ), .A2(n3), .ZN(n2035) );
  CKNXD16 U3149 ( .I(n2035), .ZN(AdrEna[97]) );
  CKND2D0 U3150 ( .A1(\DL3[5].tempL3[12] ), .A2(n7), .ZN(n2037) );
  CKNXD16 U3151 ( .I(n2037), .ZN(AdrEna[92]) );
  CKND2D0 U3152 ( .A1(\DL3[58].tempL3[0] ), .A2(n9), .ZN(n2039) );
  CKNXD16 U3153 ( .I(n2039), .ZN(AdrEna[928]) );
  CKND2D0 U3154 ( .A1(\DL3[5].tempL3[7] ), .A2(n7), .ZN(n2041) );
  CKNXD16 U3155 ( .I(n2041), .ZN(AdrEna[87]) );
  CKND2D0 U3156 ( .A1(\DL3[57].tempL3[8] ), .A2(n10), .ZN(n2043) );
  CKNXD16 U3157 ( .I(n2043), .ZN(AdrEna[920]) );
  CKND2D0 U3158 ( .A1(\DL3[58].tempL3[4] ), .A2(n9), .ZN(n2045) );
  CKNXD16 U3159 ( .I(n2045), .ZN(AdrEna[932]) );
  CKND2D0 U3160 ( .A1(\DL3[5].tempL3[10] ), .A2(n7), .ZN(n2047) );
  CKNXD16 U3161 ( .I(n2047), .ZN(AdrEna[90]) );
  CKND2D0 U3162 ( .A1(\DL3[58].tempL3[9] ), .A2(n9), .ZN(n2049) );
  CKNXD16 U3163 ( .I(n2049), .ZN(AdrEna[937]) );
  CKND2D0 U3164 ( .A1(\DL3[5].tempL3[8] ), .A2(n7), .ZN(n2051) );
  CKNXD16 U3165 ( .I(n2051), .ZN(AdrEna[88]) );
  CKND2D0 U3166 ( .A1(\DL3[5].tempL3[6] ), .A2(n7), .ZN(n2053) );
  CKNXD16 U3167 ( .I(n2053), .ZN(AdrEna[86]) );
  CKND2D0 U3168 ( .A1(\DL3[58].tempL3[1] ), .A2(n9), .ZN(n2055) );
  CKNXD16 U3169 ( .I(n2055), .ZN(AdrEna[929]) );
  CKND2D0 U3170 ( .A1(\DL3[5].tempL3[5] ), .A2(n7), .ZN(n2057) );
  CKNXD16 U3171 ( .I(n2057), .ZN(AdrEna[85]) );
  CKND2D0 U3172 ( .A1(\DL3[58].tempL3[5] ), .A2(n9), .ZN(n2059) );
  CKNXD16 U3173 ( .I(n2059), .ZN(AdrEna[933]) );
  CKND2D0 U3174 ( .A1(\DL3[58].tempL3[10] ), .A2(n9), .ZN(n2061) );
  CKNXD16 U3175 ( .I(n2061), .ZN(AdrEna[938]) );
  CKND2D0 U3176 ( .A1(\DL3[5].tempL3[3] ), .A2(n7), .ZN(n2063) );
  CKNXD16 U3177 ( .I(n2063), .ZN(AdrEna[83]) );
  CKND2D0 U3178 ( .A1(\DL3[58].tempL3[13] ), .A2(n9), .ZN(n2065) );
  CKNXD16 U3179 ( .I(n2065), .ZN(AdrEna[941]) );
  CKND2D0 U3180 ( .A1(\DL3[5].tempL3[4] ), .A2(n7), .ZN(n2067) );
  CKNXD16 U3181 ( .I(n2067), .ZN(AdrEna[84]) );
  CKND2D0 U3182 ( .A1(\DL3[58].tempL3[11] ), .A2(n9), .ZN(n2069) );
  CKNXD16 U3183 ( .I(n2069), .ZN(AdrEna[939]) );
  CKND2D0 U3184 ( .A1(\DL3[5].tempL3[1] ), .A2(n7), .ZN(n2071) );
  CKNXD16 U3185 ( .I(n2071), .ZN(AdrEna[81]) );
  CKND2D0 U3186 ( .A1(\DL3[58].tempL3[12] ), .A2(n9), .ZN(n2073) );
  CKNXD16 U3187 ( .I(n2073), .ZN(AdrEna[940]) );
  CKND2D0 U3188 ( .A1(\DL3[58].tempL3[14] ), .A2(n9), .ZN(n2075) );
  CKNXD16 U3189 ( .I(n2075), .ZN(AdrEna[942]) );
  CKND2D0 U3190 ( .A1(\DL3[4].tempL3[12] ), .A2(n18), .ZN(n2077) );
  CKNXD16 U3191 ( .I(n2077), .ZN(AdrEna[76]) );
  CKND2D0 U3192 ( .A1(\DL3[59].tempL3[3] ), .A2(n8), .ZN(n2079) );
  CKNXD16 U3193 ( .I(n2079), .ZN(AdrEna[947]) );
  CKND2D0 U3194 ( .A1(\DL3[5].tempL3[0] ), .A2(n7), .ZN(n2081) );
  CKNXD16 U3195 ( .I(n2081), .ZN(AdrEna[80]) );
  CKND2D0 U3196 ( .A1(\DL3[4].tempL3[10] ), .A2(n18), .ZN(n2083) );
  CKNXD16 U3197 ( .I(n2083), .ZN(AdrEna[74]) );
  CKND2D0 U3198 ( .A1(\DL3[59].tempL3[0] ), .A2(n8), .ZN(n2085) );
  CKNXD16 U3199 ( .I(n2085), .ZN(AdrEna[944]) );
  CKND2D0 U3200 ( .A1(\DL3[4].tempL3[6] ), .A2(n18), .ZN(n2087) );
  CKNXD16 U3201 ( .I(n2087), .ZN(AdrEna[70]) );
  CKND2D0 U3202 ( .A1(\DL3[58].tempL3[7] ), .A2(n9), .ZN(n2089) );
  CKNXD16 U3203 ( .I(n2089), .ZN(AdrEna[935]) );
  CKND2D0 U3204 ( .A1(\DL3[59].tempL3[4] ), .A2(n8), .ZN(n2091) );
  CKNXD16 U3205 ( .I(n2091), .ZN(AdrEna[948]) );
  CKND2D0 U3206 ( .A1(\DL3[4].tempL3[8] ), .A2(n18), .ZN(n2093) );
  CKNXD16 U3207 ( .I(n2093), .ZN(AdrEna[72]) );
  CKND2D0 U3208 ( .A1(\DL3[59].tempL3[9] ), .A2(n8), .ZN(n2095) );
  CKNXD16 U3209 ( .I(n2095), .ZN(AdrEna[953]) );
  CKND2D0 U3210 ( .A1(\DL3[4].tempL3[7] ), .A2(n18), .ZN(n2097) );
  CKNXD16 U3211 ( .I(n2097), .ZN(AdrEna[71]) );
  CKND2D0 U3212 ( .A1(\DL3[4].tempL3[5] ), .A2(n18), .ZN(n2099) );
  CKNXD16 U3213 ( .I(n2099), .ZN(AdrEna[69]) );
  CKND2D0 U3214 ( .A1(\DL3[59].tempL3[1] ), .A2(n8), .ZN(n2101) );
  CKNXD16 U3215 ( .I(n2101), .ZN(AdrEna[945]) );
  CKND2D0 U3216 ( .A1(\DL3[4].tempL3[2] ), .A2(n18), .ZN(n2103) );
  CKNXD16 U3217 ( .I(n2103), .ZN(AdrEna[66]) );
  CKND2D0 U3218 ( .A1(\DL3[59].tempL3[5] ), .A2(n8), .ZN(n2105) );
  CKNXD16 U3219 ( .I(n2105), .ZN(AdrEna[949]) );
  CKND2D0 U3220 ( .A1(\DL3[59].tempL3[10] ), .A2(n8), .ZN(n2107) );
  CKNXD16 U3221 ( .I(n2107), .ZN(AdrEna[954]) );
  CKND2D0 U3222 ( .A1(\DL3[4].tempL3[4] ), .A2(n18), .ZN(n2109) );
  CKNXD16 U3223 ( .I(n2109), .ZN(AdrEna[68]) );
  CKND2D0 U3224 ( .A1(\DL3[59].tempL3[11] ), .A2(n8), .ZN(n2111) );
  CKNXD16 U3225 ( .I(n2111), .ZN(AdrEna[955]) );
  CKND2D0 U3226 ( .A1(\DL3[4].tempL3[3] ), .A2(n18), .ZN(n2113) );
  CKNXD16 U3227 ( .I(n2113), .ZN(AdrEna[67]) );
  CKND2D0 U3228 ( .A1(\DL3[4].tempL3[1] ), .A2(n18), .ZN(n2115) );
  CKNXD16 U3229 ( .I(n2115), .ZN(AdrEna[65]) );
  CKND2D0 U3230 ( .A1(\DL3[59].tempL3[13] ), .A2(n8), .ZN(n2117) );
  CKNXD16 U3231 ( .I(n2117), .ZN(AdrEna[957]) );
  CKND2D0 U3232 ( .A1(\DL3[3].tempL3[12] ), .A2(n29), .ZN(n2119) );
  CKNXD16 U3233 ( .I(n2119), .ZN(AdrEna[60]) );
  CKND2D0 U3234 ( .A1(\DL3[59].tempL3[12] ), .A2(n8), .ZN(n2121) );
  CKNXD16 U3235 ( .I(n2121), .ZN(AdrEna[956]) );
  CKND2D0 U3236 ( .A1(\DL3[59].tempL3[14] ), .A2(n8), .ZN(n2123) );
  CKNXD16 U3237 ( .I(n2123), .ZN(AdrEna[958]) );
  CKND2D0 U3238 ( .A1(\DL3[4].tempL3[0] ), .A2(n18), .ZN(n2125) );
  CKNXD16 U3239 ( .I(n2125), .ZN(AdrEna[64]) );
  CKND2D0 U3240 ( .A1(\DL3[60].tempL3[0] ), .A2(n6), .ZN(n2127) );
  CKNXD16 U3241 ( .I(n2127), .ZN(AdrEna[960]) );
  CKND2D0 U3242 ( .A1(\DL3[3].tempL3[8] ), .A2(n29), .ZN(n2129) );
  CKNXD16 U3243 ( .I(n2129), .ZN(AdrEna[56]) );
  CKND2D0 U3244 ( .A1(\DL3[3].tempL3[10] ), .A2(n29), .ZN(n2131) );
  CKNXD16 U3245 ( .I(n2131), .ZN(AdrEna[58]) );
  CKND2D0 U3246 ( .A1(\DL3[60].tempL3[2] ), .A2(n6), .ZN(n2133) );
  CKNXD16 U3247 ( .I(n2133), .ZN(AdrEna[962]) );
  CKND2D0 U3248 ( .A1(\DL3[3].tempL3[7] ), .A2(n29), .ZN(n2135) );
  CKNXD16 U3249 ( .I(n2135), .ZN(AdrEna[55]) );
  CKND2D0 U3250 ( .A1(\DL3[60].tempL3[1] ), .A2(n6), .ZN(n2137) );
  CKNXD16 U3251 ( .I(n2137), .ZN(AdrEna[961]) );
  CKND2D0 U3252 ( .A1(\DL3[60].tempL3[3] ), .A2(n6), .ZN(n2139) );
  CKNXD16 U3253 ( .I(n2139), .ZN(AdrEna[963]) );
  CKND2D0 U3254 ( .A1(\DL3[3].tempL3[6] ), .A2(n29), .ZN(n2141) );
  CKNXD16 U3255 ( .I(n2141), .ZN(AdrEna[54]) );
  CKND2D0 U3256 ( .A1(\DL3[60].tempL3[4] ), .A2(n6), .ZN(n2143) );
  CKNXD16 U3257 ( .I(n2143), .ZN(AdrEna[964]) );
  CKND2D0 U3258 ( .A1(\DL3[3].tempL3[4] ), .A2(n29), .ZN(n2145) );
  CKNXD16 U3259 ( .I(n2145), .ZN(AdrEna[52]) );
  CKND2D0 U3260 ( .A1(\DL3[3].tempL3[5] ), .A2(n29), .ZN(n2147) );
  CKNXD16 U3261 ( .I(n2147), .ZN(AdrEna[53]) );
  CKND2D0 U3262 ( .A1(\DL3[60].tempL3[6] ), .A2(n6), .ZN(n2149) );
  CKNXD16 U3263 ( .I(n2149), .ZN(AdrEna[966]) );
  CKND2D0 U3264 ( .A1(\DL3[3].tempL3[3] ), .A2(n29), .ZN(n2151) );
  CKNXD16 U3265 ( .I(n2151), .ZN(AdrEna[51]) );
  CKND2D0 U3266 ( .A1(\DL3[60].tempL3[5] ), .A2(n6), .ZN(n2153) );
  CKNXD16 U3267 ( .I(n2153), .ZN(AdrEna[965]) );
  CKND2D0 U3268 ( .A1(\DL3[60].tempL3[7] ), .A2(n6), .ZN(n2155) );
  CKNXD16 U3269 ( .I(n2155), .ZN(AdrEna[967]) );
  CKND2D0 U3270 ( .A1(\DL3[3].tempL3[2] ), .A2(n29), .ZN(n2157) );
  CKNXD16 U3271 ( .I(n2157), .ZN(AdrEna[50]) );
  CKND2D0 U3272 ( .A1(\DL3[60].tempL3[8] ), .A2(n6), .ZN(n2159) );
  CKNXD16 U3273 ( .I(n2159), .ZN(AdrEna[968]) );
  CKND2D0 U3274 ( .A1(\DL3[3].tempL3[0] ), .A2(n29), .ZN(n2161) );
  CKNXD16 U3275 ( .I(n2161), .ZN(AdrEna[48]) );
  CKND2D0 U3276 ( .A1(\DL3[3].tempL3[1] ), .A2(n29), .ZN(n2163) );
  CKNXD16 U3277 ( .I(n2163), .ZN(AdrEna[49]) );
  CKND2D0 U3278 ( .A1(\DL3[59].tempL3[7] ), .A2(n8), .ZN(n2165) );
  CKNXD16 U3279 ( .I(n2165), .ZN(AdrEna[951]) );
  CKND2D0 U3280 ( .A1(\DL3[2].tempL3[12] ), .A2(n40), .ZN(n2167) );
  CKNXD16 U3281 ( .I(n2167), .ZN(AdrEna[44]) );
  CKND2D0 U3282 ( .A1(\DL3[60].tempL3[9] ), .A2(n6), .ZN(n2169) );
  CKNXD16 U3283 ( .I(n2169), .ZN(AdrEna[969]) );
  CKND2D0 U3284 ( .A1(\DL3[60].tempL3[10] ), .A2(n6), .ZN(n2171) );
  CKNXD16 U3285 ( .I(n2171), .ZN(AdrEna[970]) );
  CKND2D0 U3286 ( .A1(\DL3[2].tempL3[10] ), .A2(n40), .ZN(n2173) );
  CKNXD16 U3287 ( .I(n2173), .ZN(AdrEna[42]) );
  CKND2D0 U3288 ( .A1(\DL3[61].tempL3[0] ), .A2(n5), .ZN(n2175) );
  CKNXD16 U3289 ( .I(n2175), .ZN(AdrEna[976]) );
  CKND2D0 U3290 ( .A1(\DL3[2].tempL3[8] ), .A2(n40), .ZN(n2177) );
  CKNXD16 U3291 ( .I(n2177), .ZN(AdrEna[40]) );
  CKND2D0 U3292 ( .A1(\DL3[2].tempL3[7] ), .A2(n40), .ZN(n2179) );
  CKNXD16 U3293 ( .I(n2179), .ZN(AdrEna[39]) );
  CKND2D0 U3294 ( .A1(\DL3[61].tempL3[2] ), .A2(n5), .ZN(n2181) );
  CKNXD16 U3295 ( .I(n2181), .ZN(AdrEna[978]) );
  CKND2D0 U3296 ( .A1(\DL3[2].tempL3[5] ), .A2(n40), .ZN(n2183) );
  CKNXD16 U3297 ( .I(n2183), .ZN(AdrEna[37]) );
  CKND2D0 U3298 ( .A1(\DL3[61].tempL3[1] ), .A2(n5), .ZN(n2185) );
  CKNXD16 U3299 ( .I(n2185), .ZN(AdrEna[977]) );
  CKND2D0 U3300 ( .A1(\DL3[61].tempL3[3] ), .A2(n5), .ZN(n2187) );
  CKNXD16 U3301 ( .I(n2187), .ZN(AdrEna[979]) );
  CKND2D0 U3302 ( .A1(\DL3[2].tempL3[6] ), .A2(n40), .ZN(n2189) );
  CKNXD16 U3303 ( .I(n2189), .ZN(AdrEna[38]) );
  CKND2D0 U3304 ( .A1(\DL3[61].tempL3[4] ), .A2(n5), .ZN(n2191) );
  CKNXD16 U3305 ( .I(n2191), .ZN(AdrEna[980]) );
  CKND2D0 U3306 ( .A1(\DL3[2].tempL3[4] ), .A2(n40), .ZN(n2193) );
  CKNXD16 U3307 ( .I(n2193), .ZN(AdrEna[36]) );
  CKND2D0 U3308 ( .A1(\DL3[2].tempL3[3] ), .A2(n40), .ZN(n2195) );
  CKNXD16 U3309 ( .I(n2195), .ZN(AdrEna[35]) );
  CKND2D0 U3310 ( .A1(\DL3[60].tempL3[12] ), .A2(n6), .ZN(n2197) );
  CKNXD16 U3311 ( .I(n2197), .ZN(AdrEna[972]) );
  CKND2D0 U3312 ( .A1(\DL3[61].tempL3[10] ), .A2(n5), .ZN(n2199) );
  CKNXD16 U3313 ( .I(n2199), .ZN(AdrEna[986]) );
  CKND2D0 U3314 ( .A1(\DL3[61].tempL3[5] ), .A2(n5), .ZN(n2201) );
  CKNXD16 U3315 ( .I(n2201), .ZN(AdrEna[981]) );
  CKND2D0 U3316 ( .A1(\DL3[61].tempL3[8] ), .A2(n5), .ZN(n2203) );
  CKNXD16 U3317 ( .I(n2203), .ZN(AdrEna[984]) );
  CKND2D0 U3318 ( .A1(\DL3[2].tempL3[2] ), .A2(n40), .ZN(n2205) );
  CKNXD16 U3319 ( .I(n2205), .ZN(AdrEna[34]) );
  CKND2D0 U3320 ( .A1(\DL3[61].tempL3[11] ), .A2(n5), .ZN(n2207) );
  CKNXD16 U3321 ( .I(n2207), .ZN(AdrEna[987]) );
  CKND2D0 U3322 ( .A1(\DL3[2].tempL3[1] ), .A2(n40), .ZN(n2209) );
  CKNXD16 U3323 ( .I(n2209), .ZN(AdrEna[33]) );
  CKND2D0 U3324 ( .A1(\DL3[61].tempL3[6] ), .A2(n5), .ZN(n2211) );
  CKNXD16 U3325 ( .I(n2211), .ZN(AdrEna[982]) );
  CKND2D0 U3326 ( .A1(\DL3[61].tempL3[9] ), .A2(n5), .ZN(n2213) );
  CKNXD16 U3327 ( .I(n2213), .ZN(AdrEna[985]) );
  CKND2D0 U3328 ( .A1(\DL3[62].tempL3[0] ), .A2(n4), .ZN(n2215) );
  CKNXD16 U3329 ( .I(n2215), .ZN(AdrEna[992]) );
  CKND2D0 U3330 ( .A1(\DL3[2].tempL3[0] ), .A2(n40), .ZN(n2217) );
  CKNXD16 U3331 ( .I(n2217), .ZN(AdrEna[32]) );
  CKND2D0 U3332 ( .A1(\DL3[1].tempL3[8] ), .A2(n51), .ZN(n2219) );
  CKNXD16 U3333 ( .I(n2219), .ZN(AdrEna[24]) );
  CKND2D0 U3334 ( .A1(\DL3[1].tempL3[10] ), .A2(n51), .ZN(n2221) );
  CKNXD16 U3335 ( .I(n2221), .ZN(AdrEna[26]) );
  CKND2D0 U3336 ( .A1(\DL3[1].tempL3[7] ), .A2(n51), .ZN(n2223) );
  CKNXD16 U3337 ( .I(n2223), .ZN(AdrEna[23]) );
  CKND2D0 U3338 ( .A1(\DL3[62].tempL3[4] ), .A2(n4), .ZN(n2225) );
  CKNXD16 U3339 ( .I(n2225), .ZN(AdrEna[996]) );
  CKND2D0 U3340 ( .A1(\DL3[62].tempL3[5] ), .A2(n4), .ZN(n2227) );
  CKNXD16 U3341 ( .I(n2227), .ZN(AdrEna[997]) );
  CKND2D0 U3342 ( .A1(\DL3[62].tempL3[3] ), .A2(n4), .ZN(n2229) );
  CKNXD16 U3343 ( .I(n2229), .ZN(AdrEna[995]) );
  CKND2D0 U3344 ( .A1(\DL3[62].tempL3[6] ), .A2(n4), .ZN(n2231) );
  CKNXD16 U3345 ( .I(n2231), .ZN(AdrEna[998]) );
  CKND2D0 U3346 ( .A1(\DL3[1].tempL3[3] ), .A2(n51), .ZN(n2233) );
  CKNXD16 U3347 ( .I(n2233), .ZN(AdrEna[19]) );
  CKND2D0 U3348 ( .A1(\DL3[1].tempL3[2] ), .A2(n51), .ZN(n2235) );
  CKNXD16 U3349 ( .I(n2235), .ZN(AdrEna[18]) );
  CKND2D0 U3350 ( .A1(\DL3[1].tempL3[4] ), .A2(n51), .ZN(n2237) );
  CKNXD16 U3351 ( .I(n2237), .ZN(AdrEna[20]) );
  CKND2D0 U3352 ( .A1(\DL3[1].tempL3[1] ), .A2(n51), .ZN(n2239) );
  CKNXD16 U3353 ( .I(n2239), .ZN(AdrEna[17]) );
  CKND2D0 U3354 ( .A1(\DL3[62].tempL3[10] ), .A2(n4), .ZN(n2241) );
  CKNXD16 U3355 ( .I(n2241), .ZN(AdrEna[1002]) );
  CKND2D0 U3356 ( .A1(\DL3[62].tempL3[11] ), .A2(n4), .ZN(n2243) );
  CKNXD16 U3357 ( .I(n2243), .ZN(AdrEna[1003]) );
  CKND2D0 U3358 ( .A1(\DL3[62].tempL3[9] ), .A2(n4), .ZN(n2245) );
  CKNXD16 U3359 ( .I(n2245), .ZN(AdrEna[1001]) );
  CKND2D0 U3360 ( .A1(\DL3[0].tempL3[12] ), .A2(n2), .ZN(n2247) );
  CKNXD16 U3361 ( .I(n2247), .ZN(AdrEna[12]) );
  CKND2D0 U3362 ( .A1(\DL3[0].tempL3[10] ), .A2(n2), .ZN(n2249) );
  CKNXD16 U3363 ( .I(n2249), .ZN(AdrEna[10]) );
  CKND2D0 U3364 ( .A1(\DL3[0].tempL3[9] ), .A2(n2), .ZN(n2251) );
  CKNXD16 U3365 ( .I(n2251), .ZN(AdrEna[9]) );
  CKND2D0 U3366 ( .A1(\DL3[61].tempL3[12] ), .A2(n5), .ZN(n2253) );
  CKNXD16 U3367 ( .I(n2253), .ZN(AdrEna[988]) );
  CKND2D0 U3368 ( .A1(\DL3[0].tempL3[8] ), .A2(n2), .ZN(n2255) );
  CKNXD16 U3369 ( .I(n2255), .ZN(AdrEna[8]) );
  CKND2D0 U3370 ( .A1(\DL3[63].tempL3[4] ), .A2(n65), .ZN(n2257) );
  CKNXD16 U3371 ( .I(n2257), .ZN(AdrEna[1012]) );
  CKND2D0 U3372 ( .A1(\DL3[63].tempL3[8] ), .A2(n65), .ZN(n2259) );
  CKNXD16 U3373 ( .I(n2259), .ZN(AdrEna[1016]) );
  CKND2D0 U3374 ( .A1(\DL3[62].tempL3[14] ), .A2(n4), .ZN(n2261) );
  CKNXD16 U3375 ( .I(n2261), .ZN(AdrEna[1006]) );
  CKND2D0 U3376 ( .A1(\DL3[0].tempL3[2] ), .A2(n2), .ZN(n2263) );
  CKNXD16 U3377 ( .I(n2263), .ZN(AdrEna[2]) );
  CKND2D0 U3378 ( .A1(\DL3[0].tempL3[1] ), .A2(n2), .ZN(n2265) );
  CKNXD16 U3379 ( .I(n2265), .ZN(AdrEna[1]) );
  CKND2D0 U3380 ( .A1(\DL3[0].tempL3[0] ), .A2(n2), .ZN(n2267) );
  CKNXD16 U3381 ( .I(n2267), .ZN(AdrEna[0]) );
  CKND2D0 U3382 ( .A1(\DL3[63].tempL3[12] ), .A2(n65), .ZN(n2269) );
  CKNXD16 U3383 ( .I(n2269), .ZN(AdrEna[1020]) );
  INVD0 U3384 ( .I(n2286), .ZN(n2273) );
  CKAN2D0 U3385 ( .A1(\DL2[3].tempL2[3] ), .A2(DecodedL1[3]), .Z(n16) );
  TIEL U3386 ( .ZN(\*Logic0* ) );
endmodule


module Dec4_16_0 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n5, n6, n8, n9, n11, n12, n13, n14, n15, n16, n1, n2;

  NR2D1 U1 ( .A1(n1), .A2(n12), .ZN(Hot[0]) );
  NR2D1 U2 ( .A1(n5), .A2(n12), .ZN(Hot[1]) );
  NR2D1 U3 ( .A1(n2), .A2(n12), .ZN(Hot[2]) );
  NR2D1 U4 ( .A1(n8), .A2(n12), .ZN(Hot[3]) );
  OR2D1 U5 ( .A1(n14), .A2(n15), .Z(n8) );
  ND2D1 U6 ( .A1(n14), .A2(n15), .ZN(n1) );
  ND2D1 U7 ( .A1(Sel[1]), .A2(n15), .ZN(n2) );
  ND2D1 U8 ( .A1(Sel[0]), .A2(n14), .ZN(n5) );
  CKND0 U9 ( .CLK(Sel[1]), .CN(n14) );
  NR2D1 U10 ( .A1(n6), .A2(n2), .ZN(Hot[10]) );
  NR2D1 U11 ( .A1(n9), .A2(n2), .ZN(Hot[6]) );
  NR2D1 U12 ( .A1(n6), .A2(n1), .ZN(Hot[8]) );
  NR2D1 U13 ( .A1(n2), .A2(n13), .ZN(Hot[14]) );
  NR2D1 U14 ( .A1(n1), .A2(n13), .ZN(Hot[12]) );
  NR2D1 U15 ( .A1(n1), .A2(n9), .ZN(Hot[4]) );
  NR2D0 U16 ( .A1(n5), .A2(n13), .ZN(Hot[13]) );
  NR2D0 U17 ( .A1(n5), .A2(n9), .ZN(Hot[5]) );
  NR2D0 U18 ( .A1(n5), .A2(n6), .ZN(Hot[9]) );
  NR2D0 U19 ( .A1(n6), .A2(n8), .ZN(Hot[11]) );
  NR2D0 U20 ( .A1(n8), .A2(n13), .ZN(Hot[15]) );
  NR2D0 U21 ( .A1(n8), .A2(n9), .ZN(Hot[7]) );
  ND2D1 U22 ( .A1(n16), .A2(n11), .ZN(n12) );
  ND2D1 U23 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n13) );
  ND2D1 U24 ( .A1(Sel[2]), .A2(n11), .ZN(n9) );
  ND2D1 U25 ( .A1(Sel[3]), .A2(n16), .ZN(n6) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n16) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n15) );
endmodule


module Dec4_16_1 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2D0 U2 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2D0 U3 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D0 U4 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2D0 U5 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U6 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2D0 U7 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D0 U8 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  ND2D1 U9 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  NR2D0 U10 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  ND2D0 U11 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  NR2XD0 U12 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U13 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U14 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  CKND2D1 U15 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U16 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D0 U17 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U18 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U19 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U20 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2XD0 U21 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U22 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  INVD1 U25 ( .I(Sel[3]), .ZN(n4) );
  CKND0 U26 ( .CLK(Sel[2]), .CN(n3) );
  INVD1 U27 ( .I(Sel[0]), .ZN(n1) );
  CKND0 U28 ( .CLK(Sel[1]), .CN(n2) );
endmodule


module Dec4_16_2 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  ND2D1 U1 ( .A1(Sel[1]), .A2(n2), .ZN(n16) );
  ND2D1 U2 ( .A1(Sel[1]), .A2(n1), .ZN(n18) );
  NR2D1 U3 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D1 U4 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2D1 U5 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2D0 U6 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2D0 U7 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D1 U8 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  CKND2D1 U9 ( .A1(n2), .A2(n3), .ZN(n19) );
  CKND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n21) );
  ND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  ND2D1 U12 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  INVD1 U13 ( .I(n2), .ZN(n1) );
  ND2D0 U14 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  ND2D1 U15 ( .A1(n4), .A2(n11), .ZN(n15) );
  NR2XD0 U16 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U17 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U18 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U19 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U20 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U21 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U22 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U24 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U25 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n2) );
  CKND0 U29 ( .CLK(Sel[1]), .CN(n3) );
endmodule


module Dec4_16_3 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  ND2D1 U1 ( .A1(n1), .A2(n3), .ZN(n21) );
  ND2D1 U2 ( .A1(Sel[1]), .A2(n2), .ZN(n16) );
  NR2D1 U3 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U4 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2D0 U5 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2D1 U6 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D1 U7 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  CKND2D1 U8 ( .A1(n2), .A2(n3), .ZN(n19) );
  ND2D0 U9 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  ND2D1 U10 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  INVD1 U11 ( .I(n2), .ZN(n1) );
  ND2D0 U12 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  ND2D1 U13 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(n1), .ZN(n18) );
  NR2XD0 U15 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U16 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U17 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U18 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U19 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U20 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U21 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U22 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U24 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U25 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n2) );
  CKND0 U29 ( .CLK(Sel[1]), .CN(n3) );
endmodule


module Dec4_16_4 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  ND2D1 U1 ( .A1(Sel[1]), .A2(n1), .ZN(n18) );
  NR2D1 U2 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2D1 U3 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U4 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2D0 U5 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2D0 U6 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  CKND2D1 U7 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  ND2D1 U8 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD0 U9 ( .I(Sel[1]), .ZN(n3) );
  CKND2D1 U10 ( .A1(n2), .A2(n3), .ZN(n19) );
  INVD1 U11 ( .I(n2), .ZN(n1) );
  CKND0 U12 ( .CLK(Sel[3]), .CN(n11) );
  CKND2D0 U13 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(n2), .ZN(n16) );
  CKND0 U17 ( .CLK(Sel[2]), .CN(n4) );
  NR2XD0 U18 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U20 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U25 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2XD0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  INVD1 U29 ( .I(Sel[0]), .ZN(n2) );
endmodule


module Dec4_16_5 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D1 U2 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D1 U3 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U4 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  CKND2D1 U5 ( .A1(n1), .A2(n4), .ZN(n22) );
  INVD1 U6 ( .I(n4), .ZN(n3) );
  ND2D0 U7 ( .A1(n3), .A2(n1), .ZN(n19) );
  CKND2D0 U8 ( .A1(n11), .A2(n14), .ZN(n16) );
  CKND2D0 U9 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  CKND2D1 U10 ( .A1(n3), .A2(n2), .ZN(n17) );
  INVD0 U11 ( .I(Sel[3]), .ZN(n14) );
  CKND0 U12 ( .CLK(n2), .CN(n1) );
  INVD0 U13 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U14 ( .I(Sel[1]), .ZN(n4) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n15) );
  INVD0 U16 ( .I(Sel[2]), .ZN(n11) );
  ND2D1 U17 ( .A1(n2), .A2(n4), .ZN(n20) );
  CKND2D0 U18 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  NR2XD0 U19 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U20 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U21 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U23 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U24 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U25 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U26 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U27 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U28 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U29 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
endmodule


module Dec4_16_6 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  NR2D1 U2 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D1 U3 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D1 U4 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  CKND2D1 U5 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  INVD1 U6 ( .I(n3), .ZN(n2) );
  ND2D0 U7 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  CKND2D0 U8 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND2D0 U9 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND2D1 U10 ( .A1(n2), .A2(n1), .ZN(n17) );
  INVD0 U11 ( .I(Sel[3]), .ZN(n14) );
  INVD0 U12 ( .I(Sel[0]), .ZN(n1) );
  INVD0 U13 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  INVD0 U15 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U16 ( .I(n14), .ZN(n11) );
  ND2D1 U17 ( .A1(n1), .A2(n3), .ZN(n20) );
  NR2XD0 U18 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U21 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U22 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U23 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U25 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U26 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2XD0 U27 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U28 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U29 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
endmodule


module Dec4_16_7 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2D1 U2 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D1 U3 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U4 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  ND2D0 U5 ( .A1(n1), .A2(n3), .ZN(n19) );
  ND2D0 U6 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  INVD0 U7 ( .I(Sel[3]), .ZN(n11) );
  CKND2D0 U8 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  CKND2D0 U9 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  INVD0 U10 ( .I(Sel[2]), .ZN(n4) );
  ND2D0 U11 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U12 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  NR2D0 U13 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  INVD1 U14 ( .I(n3), .ZN(n2) );
  CKND0 U15 ( .CLK(Sel[1]), .CN(n3) );
  CKND0 U16 ( .CLK(Sel[0]), .CN(n1) );
  ND2D1 U17 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U18 ( .A1(n2), .A2(n1), .ZN(n16) );
  NR2XD0 U19 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U22 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U25 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U26 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2XD0 U28 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U29 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
endmodule


module Dec4_16_8 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D1 U2 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  CKND2D0 U4 ( .A1(n1), .A2(n3), .ZN(n19) );
  CKND2D0 U5 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U6 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  NR2XD0 U7 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  CKND2D0 U8 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  CKND2D0 U9 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U10 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  INVD1 U11 ( .I(n3), .ZN(n2) );
  CKND0 U12 ( .CLK(Sel[1]), .CN(n3) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U14 ( .A1(n2), .A2(n1), .ZN(n16) );
  CKND0 U15 ( .CLK(Sel[3]), .CN(n11) );
  NR2XD0 U16 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U17 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U18 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U19 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U25 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U26 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2XD0 U27 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n1) );
  CKND0 U29 ( .CLK(Sel[2]), .CN(n4) );
endmodule


module Dec4_16_9 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  CKND2D0 U3 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U4 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  ND2D1 U5 ( .A1(n2), .A2(n1), .ZN(n16) );
  INVD0 U6 ( .I(Sel[1]), .ZN(n3) );
  INVD0 U7 ( .I(Sel[0]), .ZN(n1) );
  INVD0 U8 ( .I(Sel[3]), .ZN(n11) );
  ND2D0 U9 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  ND2D0 U10 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  INVD0 U12 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U13 ( .I(n3), .ZN(n2) );
  ND2D1 U14 ( .A1(n1), .A2(n3), .ZN(n19) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  NR2XD0 U16 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U17 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U18 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U19 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U25 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U26 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2XD0 U28 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2XD0 U29 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
endmodule


module Dec4_16_10 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  ND2D1 U1 ( .A1(n4), .A2(n15), .ZN(n19) );
  NR2D0 U2 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2D0 U3 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2D0 U4 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U5 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D1 U6 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  CKND2D0 U7 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U8 ( .A1(n14), .A2(n11), .ZN(n22) );
  ND2D1 U9 ( .A1(n2), .A2(n1), .ZN(n18) );
  INVD0 U10 ( .I(Sel[1]), .ZN(n3) );
  INVD0 U11 ( .I(Sel[0]), .ZN(n1) );
  INVD0 U12 ( .I(Sel[3]), .ZN(n15) );
  ND2D0 U13 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  ND2D0 U14 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U15 ( .A1(n4), .A2(n14), .ZN(n16) );
  INVD1 U16 ( .I(n11), .ZN(n4) );
  INVD0 U17 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U18 ( .I(n15), .ZN(n14) );
  INVD1 U19 ( .I(n3), .ZN(n2) );
  ND2D1 U20 ( .A1(n1), .A2(n3), .ZN(n21) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U23 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U24 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U25 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U26 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U27 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2XD0 U28 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2XD0 U29 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2XD0 U30 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2XD0 U31 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
endmodule


module Dec4_16_11 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  CKND2D0 U4 ( .A1(n11), .A2(n14), .ZN(n16) );
  CKND2D0 U5 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  ND2D1 U6 ( .A1(n3), .A2(n2), .ZN(n17) );
  INVD0 U7 ( .I(Sel[1]), .ZN(n4) );
  INVD0 U8 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U9 ( .I(Sel[3]), .ZN(n14) );
  ND2D0 U10 ( .A1(n1), .A2(n4), .ZN(n22) );
  ND2D0 U11 ( .A1(n3), .A2(n1), .ZN(n19) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n15) );
  INVD0 U13 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U14 ( .I(n4), .ZN(n3) );
  INVD1 U15 ( .I(n2), .ZN(n1) );
  ND2D1 U16 ( .A1(n2), .A2(n4), .ZN(n20) );
  CKND2D0 U17 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  NR2XD0 U18 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U23 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U24 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U25 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U26 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2XD0 U27 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U28 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U29 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2XD0 U30 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
endmodule


module Dec4_16_12 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2XD0 U1 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2D0 U3 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D0 U4 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U5 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U6 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U7 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  ND2D1 U8 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  CKND2D0 U9 ( .A1(n11), .A2(n14), .ZN(n16) );
  CKND2D0 U10 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  ND2D1 U11 ( .A1(n3), .A2(n2), .ZN(n17) );
  INVD0 U12 ( .I(Sel[1]), .ZN(n4) );
  INVD0 U13 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U14 ( .I(Sel[3]), .ZN(n14) );
  ND2D0 U15 ( .A1(n1), .A2(n4), .ZN(n22) );
  ND2D0 U16 ( .A1(n3), .A2(n1), .ZN(n19) );
  CKND2D0 U17 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n15) );
  INVD0 U18 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U19 ( .I(n4), .ZN(n3) );
  INVD1 U20 ( .I(n2), .ZN(n1) );
  ND2D1 U21 ( .A1(n2), .A2(n4), .ZN(n20) );
  NR2XD0 U22 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U23 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U24 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U25 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U26 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U27 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U28 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U30 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
endmodule


module Dec4_16_13 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24;

  CKND2D0 U1 ( .A1(n2), .A2(n4), .ZN(n22) );
  CKND2D0 U2 ( .A1(n14), .A2(n16), .ZN(n18) );
  CKND2D0 U3 ( .A1(n1), .A2(n4), .ZN(n24) );
  CKND2D0 U4 ( .A1(n15), .A2(n14), .ZN(n23) );
  CKND2D0 U5 ( .A1(n11), .A2(n15), .ZN(n17) );
  INVD1 U6 ( .I(n16), .ZN(n15) );
  INVD1 U7 ( .I(n14), .ZN(n11) );
  INVD1 U8 ( .I(n4), .ZN(n3) );
  INVD1 U9 ( .I(n2), .ZN(n1) );
  CKND2D0 U10 ( .A1(n11), .A2(n16), .ZN(n20) );
  CKND2D0 U11 ( .A1(n3), .A2(n2), .ZN(n19) );
  CKND2D0 U12 ( .A1(n3), .A2(n1), .ZN(n21) );
  NR2XD0 U13 ( .A1(n22), .A2(n17), .ZN(Hot[12]) );
  NR2XD0 U14 ( .A1(n19), .A2(n17), .ZN(Hot[14]) );
  NR2XD0 U15 ( .A1(n24), .A2(n17), .ZN(Hot[13]) );
  NR2XD0 U16 ( .A1(n21), .A2(n17), .ZN(Hot[15]) );
  NR2XD0 U17 ( .A1(n22), .A2(n20), .ZN(Hot[4]) );
  NR2XD0 U18 ( .A1(n24), .A2(n20), .ZN(Hot[5]) );
  NR2XD0 U19 ( .A1(n21), .A2(n20), .ZN(Hot[7]) );
  NR2XD0 U20 ( .A1(n20), .A2(n19), .ZN(Hot[6]) );
  NR2XD0 U21 ( .A1(n23), .A2(n19), .ZN(Hot[10]) );
  NR2XD0 U22 ( .A1(n23), .A2(n22), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n24), .A2(n23), .ZN(Hot[9]) );
  NR2XD0 U24 ( .A1(n21), .A2(n18), .ZN(Hot[3]) );
  NR2XD0 U25 ( .A1(n19), .A2(n18), .ZN(Hot[2]) );
  NR2XD0 U26 ( .A1(n22), .A2(n18), .ZN(Hot[0]) );
  NR2XD0 U27 ( .A1(n24), .A2(n18), .ZN(Hot[1]) );
  INVD0 U28 ( .I(Sel[3]), .ZN(n16) );
  INVD0 U29 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U30 ( .I(Sel[2]), .ZN(n14) );
  INVD0 U31 ( .I(Sel[1]), .ZN(n4) );
  NR2D0 U32 ( .A1(n23), .A2(n21), .ZN(Hot[11]) );
endmodule


module Dec4_16_14 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2D1 U2 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2D1 U3 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D1 U4 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D1 U5 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2D1 U6 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D1 U7 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D1 U8 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2D1 U9 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D1 U10 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D1 U11 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D1 U12 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D1 U13 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D1 U14 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D1 U15 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  INVD0 U16 ( .I(Sel[1]), .ZN(n3) );
  CKND2D1 U17 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  CKND2D1 U18 ( .A1(Sel[1]), .A2(n1), .ZN(n19) );
  INVD1 U19 ( .I(n14), .ZN(n11) );
  INVD0 U20 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U21 ( .I(n2), .ZN(n1) );
  INVD0 U22 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U23 ( .I(Sel[2]), .ZN(n4) );
  ND2D1 U24 ( .A1(n4), .A2(n14), .ZN(n16) );
  ND2D1 U25 ( .A1(n2), .A2(n3), .ZN(n20) );
  ND2D1 U26 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  ND2D1 U27 ( .A1(Sel[1]), .A2(n2), .ZN(n17) );
  ND2D1 U28 ( .A1(n11), .A2(n4), .ZN(n21) );
  ND2D1 U29 ( .A1(n1), .A2(n3), .ZN(n22) );
  NR2D0 U30 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
endmodule


module Dec4_16_15 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24;

  ND2D1 U1 ( .A1(n11), .A2(n16), .ZN(n20) );
  ND2D1 U2 ( .A1(n15), .A2(n14), .ZN(n23) );
  ND2D1 U3 ( .A1(n2), .A2(n4), .ZN(n22) );
  ND2D1 U4 ( .A1(n1), .A2(n4), .ZN(n24) );
  ND2D1 U5 ( .A1(n3), .A2(n2), .ZN(n19) );
  ND2D1 U6 ( .A1(n3), .A2(n1), .ZN(n21) );
  ND2D1 U7 ( .A1(n11), .A2(n15), .ZN(n17) );
  NR2D1 U8 ( .A1(n22), .A2(n18), .ZN(Hot[0]) );
  NR2D1 U9 ( .A1(n21), .A2(n18), .ZN(Hot[3]) );
  NR2D1 U10 ( .A1(n22), .A2(n20), .ZN(Hot[4]) );
  NR2D1 U11 ( .A1(n24), .A2(n20), .ZN(Hot[5]) );
  NR2D1 U12 ( .A1(n20), .A2(n19), .ZN(Hot[6]) );
  NR2D1 U13 ( .A1(n21), .A2(n20), .ZN(Hot[7]) );
  NR2D1 U14 ( .A1(n23), .A2(n22), .ZN(Hot[8]) );
  NR2D1 U15 ( .A1(n24), .A2(n23), .ZN(Hot[9]) );
  NR2D1 U16 ( .A1(n23), .A2(n19), .ZN(Hot[10]) );
  NR2D1 U17 ( .A1(n23), .A2(n21), .ZN(Hot[11]) );
  NR2D1 U18 ( .A1(n22), .A2(n17), .ZN(Hot[12]) );
  NR2D1 U19 ( .A1(n24), .A2(n17), .ZN(Hot[13]) );
  NR2D1 U20 ( .A1(n19), .A2(n17), .ZN(Hot[14]) );
  NR2D1 U21 ( .A1(n21), .A2(n17), .ZN(Hot[15]) );
  INVD1 U22 ( .I(n4), .ZN(n3) );
  INVD1 U23 ( .I(n16), .ZN(n15) );
  INVD1 U24 ( .I(n2), .ZN(n1) );
  INVD1 U25 ( .I(n14), .ZN(n11) );
  NR2D1 U26 ( .A1(n24), .A2(n18), .ZN(Hot[1]) );
  NR2D1 U27 ( .A1(n19), .A2(n18), .ZN(Hot[2]) );
  INVD0 U28 ( .I(Sel[3]), .ZN(n16) );
  INVD0 U29 ( .I(Sel[0]), .ZN(n2) );
  INVD0 U30 ( .I(Sel[1]), .ZN(n4) );
  INVD0 U31 ( .I(Sel[2]), .ZN(n14) );
  ND2D1 U32 ( .A1(n14), .A2(n16), .ZN(n18) );
endmodule


module Dec4_16_16 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2D1 U2 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2D1 U3 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D1 U4 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D1 U5 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2D1 U6 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D1 U7 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D1 U8 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2D1 U9 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D1 U10 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D1 U11 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D1 U12 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D1 U13 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D1 U14 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D1 U15 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D1 U16 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  INVD1 U17 ( .I(n14), .ZN(n11) );
  INVD0 U18 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U19 ( .I(n3), .ZN(n2) );
  INVD0 U20 ( .I(Sel[0]), .ZN(n1) );
  INVD0 U21 ( .I(Sel[2]), .ZN(n4) );
  ND2D1 U22 ( .A1(n4), .A2(n14), .ZN(n16) );
  ND2D1 U23 ( .A1(n1), .A2(n3), .ZN(n20) );
  ND2D1 U24 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  ND2D1 U25 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  ND2D1 U26 ( .A1(n2), .A2(n1), .ZN(n17) );
  ND2D1 U27 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  ND2D1 U28 ( .A1(n11), .A2(n4), .ZN(n21) );
  ND2D1 U29 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  CKND0 U30 ( .CLK(Sel[1]), .CN(n3) );
endmodule


module Dec4_16_17 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2D1 U2 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2D0 U3 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  ND2D1 U4 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U6 ( .A1(n1), .A2(n2), .ZN(n17) );
  ND2D0 U7 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U8 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U9 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND2D0 U10 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U12 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U13 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U14 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2XD0 U15 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U16 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U17 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U18 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  INVD1 U20 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U21 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U22 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U23 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_18 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2D1 U2 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U3 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U4 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  NR2D0 U6 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  ND2D0 U7 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U8 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D0 U9 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U10 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U11 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U12 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND0 U13 ( .CLK(Sel[3]), .CN(n4) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U15 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U16 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U17 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U18 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2XD0 U19 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  INVD1 U20 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U21 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U22 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U23 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2D0 U27 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
endmodule


module Dec4_16_19 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  ND2D1 U1 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  ND2D1 U2 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D1 U3 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  ND2D0 U4 ( .A1(n1), .A2(n2), .ZN(n17) );
  ND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U6 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U7 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U8 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U9 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U10 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U11 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U12 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U13 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U14 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U15 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2XD0 U16 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U17 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U18 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  INVD1 U19 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U20 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U21 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U22 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U23 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2D0 U27 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
endmodule


module Dec4_16_20 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2D1 U2 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U3 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  ND2D1 U4 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  NR2XD0 U5 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  ND2D0 U6 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U7 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D0 U8 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U9 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U10 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U11 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U13 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U14 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U15 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U16 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2XD0 U17 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U18 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  INVD1 U19 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U20 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U21 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U22 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U23 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2D0 U27 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
endmodule


module Dec4_16_21 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  ND2D1 U1 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2D1 U2 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D1 U3 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  ND2D1 U4 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  ND2D0 U5 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U6 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D1 U7 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U8 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U9 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND0 U10 ( .CLK(Sel[3]), .CN(n4) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U12 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U13 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U14 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U15 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U16 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2XD0 U17 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U18 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  INVD1 U20 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U21 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U22 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U23 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2D0 U27 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
endmodule


module Dec4_16_22 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  ND2D1 U1 ( .A1(Sel[1]), .A2(n2), .ZN(n18) );
  NR2D1 U2 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2D1 U3 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U4 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  ND2D1 U5 ( .A1(n4), .A2(n15), .ZN(n19) );
  ND2D0 U6 ( .A1(n2), .A2(n3), .ZN(n21) );
  CKND2D0 U7 ( .A1(n1), .A2(n3), .ZN(n23) );
  CKND2D1 U8 ( .A1(n11), .A2(n15), .ZN(n17) );
  ND2D0 U9 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND0 U10 ( .CLK(n2), .CN(n1) );
  CKND0 U11 ( .CLK(n11), .CN(n4) );
  CKND0 U12 ( .CLK(n15), .CN(n14) );
  INVD1 U13 ( .I(Sel[3]), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(n1), .ZN(n20) );
  CKND2D0 U15 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U16 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U17 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U18 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U19 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  INVD1 U23 ( .I(Sel[0]), .ZN(n2) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U25 ( .I(Sel[2]), .ZN(n11) );
  NR2D0 U26 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U27 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U29 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_23 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2D0 U3 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D0 U4 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U5 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  ND2D0 U6 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U7 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D1 U8 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U9 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  INVD1 U10 ( .I(Sel[3]), .ZN(n4) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U12 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U13 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2XD0 U15 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2XD0 U16 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2XD0 U17 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U18 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U19 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  INVD1 U20 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U21 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U22 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U23 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U24 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2D0 U27 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
endmodule


module Dec4_16_24 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  NR2D1 U2 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D1 U3 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  INVD1 U4 ( .I(n3), .ZN(n2) );
  NR2D1 U5 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  ND2D1 U6 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  ND2D0 U7 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND2D0 U8 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D1 U9 ( .A1(n4), .A2(n14), .ZN(n16) );
  INVD1 U10 ( .I(n14), .ZN(n11) );
  CKND2D1 U11 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND2D0 U12 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  NR2XD0 U14 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U15 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U16 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U17 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U18 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U20 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  INVD1 U21 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U23 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n4) );
  NR2D0 U25 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U26 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U30 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
endmodule


module Dec4_16_25 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  ND2D1 U2 ( .A1(n4), .A2(n15), .ZN(n19) );
  ND2D0 U3 ( .A1(n1), .A2(n3), .ZN(n21) );
  CKND2D0 U4 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  ND2D1 U5 ( .A1(n11), .A2(n15), .ZN(n17) );
  INVD1 U6 ( .I(n15), .ZN(n14) );
  CKND2D1 U7 ( .A1(n14), .A2(n11), .ZN(n22) );
  INVD1 U8 ( .I(n3), .ZN(n2) );
  CKND0 U9 ( .CLK(n11), .CN(n4) );
  CKND2D0 U10 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U11 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U12 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U13 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U14 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U15 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U16 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U17 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U18 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U19 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U21 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  INVD1 U22 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U25 ( .I(Sel[2]), .ZN(n11) );
  NR2D0 U26 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U27 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U29 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_26 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(n4), .A2(n14), .ZN(n18) );
  NR2D1 U2 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D1 U3 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  ND2D1 U4 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  ND2D0 U5 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND2D0 U6 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D1 U7 ( .A1(n11), .A2(n14), .ZN(n16) );
  CKND2D1 U8 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  INVD1 U9 ( .I(n3), .ZN(n2) );
  CKND0 U10 ( .CLK(n11), .CN(n4) );
  CKND2D0 U11 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U12 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  NR2XD0 U13 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U14 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U15 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U16 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U17 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U18 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  INVD1 U21 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U23 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n11) );
  NR2D0 U25 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U26 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U30 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
endmodule


module Dec4_16_27 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D1 U2 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  ND2D0 U3 ( .A1(n2), .A2(n1), .ZN(n17) );
  ND2D1 U4 ( .A1(n4), .A2(n14), .ZN(n18) );
  ND2D0 U5 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND2D0 U6 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D1 U7 ( .A1(n11), .A2(n14), .ZN(n16) );
  CKND2D1 U8 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  INVD1 U9 ( .I(n3), .ZN(n2) );
  CKND0 U10 ( .CLK(n11), .CN(n4) );
  CKND2D0 U11 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  CKND0 U12 ( .CLK(Sel[3]), .CN(n14) );
  CKND2D0 U13 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  NR2XD0 U14 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U15 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U16 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U17 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U18 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U19 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U21 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  INVD1 U22 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U23 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n11) );
  NR2D0 U25 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U26 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U30 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
endmodule


module Dec4_16_28 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n19) );
  NR2D1 U2 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D1 U3 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  ND2D1 U4 ( .A1(n3), .A2(n14), .ZN(n18) );
  ND2D0 U5 ( .A1(n1), .A2(n2), .ZN(n20) );
  CKND2D0 U6 ( .A1(Sel[0]), .A2(n2), .ZN(n22) );
  ND2D1 U7 ( .A1(n4), .A2(n14), .ZN(n16) );
  INVD1 U8 ( .I(n14), .ZN(n11) );
  CKND2D1 U9 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND0 U10 ( .CLK(n4), .CN(n3) );
  CKND2D0 U11 ( .A1(Sel[1]), .A2(n1), .ZN(n17) );
  CKND2D0 U12 ( .A1(n3), .A2(n11), .ZN(n15) );
  NR2XD0 U13 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U14 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U15 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U16 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U17 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U18 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U19 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U20 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  INVD1 U21 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U23 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n4) );
  NR2D0 U25 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U26 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U30 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
endmodule


module Dec4_16_29 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D0 U1 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U2 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  ND2D0 U3 ( .A1(n1), .A2(n3), .ZN(n21) );
  CKND2D0 U4 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  ND2D1 U5 ( .A1(n14), .A2(n11), .ZN(n22) );
  ND2D0 U6 ( .A1(n4), .A2(n15), .ZN(n19) );
  INVD1 U7 ( .I(n3), .ZN(n2) );
  INVD0 U8 ( .I(Sel[1]), .ZN(n3) );
  CKND0 U9 ( .CLK(n11), .CN(n4) );
  INVD0 U10 ( .I(Sel[2]), .ZN(n11) );
  INVD0 U11 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U12 ( .I(n15), .ZN(n14) );
  ND2D1 U13 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U14 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U15 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U16 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U17 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U18 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U19 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U20 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U21 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U23 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U24 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  CKND0 U25 ( .CLK(Sel[3]), .CN(n15) );
  NR2D0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_30 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2D0 U2 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  ND2D0 U3 ( .A1(n1), .A2(n3), .ZN(n21) );
  CKND2D0 U4 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  ND2D1 U5 ( .A1(n14), .A2(n11), .ZN(n22) );
  ND2D0 U6 ( .A1(n4), .A2(n15), .ZN(n19) );
  INVD1 U7 ( .I(n3), .ZN(n2) );
  INVD0 U8 ( .I(Sel[1]), .ZN(n3) );
  CKND0 U9 ( .CLK(n11), .CN(n4) );
  INVD0 U10 ( .I(Sel[2]), .ZN(n11) );
  INVD0 U11 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U12 ( .I(n15), .ZN(n14) );
  ND2D1 U13 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U14 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U15 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U16 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U17 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U18 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U19 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U20 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U21 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U22 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U23 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  CKNXD0 U25 ( .I(Sel[3]), .ZN(n15) );
  NR2D0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_31 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2D0 U2 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2D0 U3 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2D0 U4 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U5 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  ND2D0 U6 ( .A1(n1), .A2(n3), .ZN(n21) );
  CKND2D0 U7 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  INVD1 U8 ( .I(n15), .ZN(n14) );
  ND2D1 U9 ( .A1(n14), .A2(n11), .ZN(n22) );
  INVD0 U10 ( .I(Sel[3]), .ZN(n15) );
  CKND0 U11 ( .CLK(n3), .CN(n2) );
  INVD0 U12 ( .I(Sel[1]), .ZN(n3) );
  ND2D0 U13 ( .A1(n4), .A2(n15), .ZN(n19) );
  CKND0 U14 ( .CLK(n11), .CN(n4) );
  INVD0 U15 ( .I(Sel[2]), .ZN(n11) );
  INVD0 U16 ( .I(Sel[0]), .ZN(n1) );
  ND2D1 U17 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U18 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U19 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U20 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U22 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U24 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U25 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_32 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D0 U1 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2D0 U2 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2D0 U3 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U4 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  ND2D0 U5 ( .A1(n1), .A2(n3), .ZN(n21) );
  CKND2D0 U6 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  ND2D1 U7 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND0 U8 ( .CLK(n3), .CN(n2) );
  INVD0 U9 ( .I(Sel[1]), .ZN(n3) );
  ND2D0 U10 ( .A1(n4), .A2(n15), .ZN(n19) );
  CKND0 U11 ( .CLK(n11), .CN(n4) );
  INVD0 U12 ( .I(Sel[2]), .ZN(n11) );
  INVD0 U13 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U14 ( .I(n15), .ZN(n14) );
  ND2D1 U15 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U16 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U17 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U18 ( .A1(n4), .A2(n14), .ZN(n16) );
  NR2XD0 U19 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U20 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U22 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U24 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  CKNXD0 U25 ( .I(Sel[3]), .ZN(n15) );
  NR2D0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U27 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U28 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U30 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U31 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
endmodule


module Dec4_16_33 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(n4), .A2(n14), .ZN(n18) );
  NR2D1 U2 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2D1 U3 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U4 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U5 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2XD0 U6 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2XD0 U7 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U8 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D0 U9 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U10 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U11 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  ND2D0 U12 ( .A1(n1), .A2(n3), .ZN(n20) );
  ND2D0 U13 ( .A1(n11), .A2(n14), .ZN(n16) );
  INVD0 U14 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U15 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  CKND2D0 U16 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND0 U17 ( .CLK(Sel[0]), .CN(n1) );
  INVD1 U18 ( .I(n11), .ZN(n4) );
  INVD1 U19 ( .I(n3), .ZN(n2) );
  CKND2D0 U20 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  CKND2D0 U21 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  CKND2D0 U22 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  CKND0 U23 ( .CLK(Sel[3]), .CN(n14) );
  NR2XD0 U24 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U25 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U26 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U27 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U28 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U29 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
endmodule


module Dec4_16_34 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U2 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U3 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  ND2D1 U5 ( .A1(n3), .A2(n11), .ZN(n17) );
  ND2D0 U6 ( .A1(n4), .A2(n11), .ZN(n15) );
  ND2D0 U7 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  NR2XD0 U8 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  CKND0 U9 ( .CLK(Sel[0]), .CN(n1) );
  ND2D0 U10 ( .A1(n3), .A2(Sel[3]), .ZN(n14) );
  INVD1 U11 ( .I(n4), .ZN(n3) );
  CKND2D0 U12 ( .A1(n1), .A2(n2), .ZN(n19) );
  CKND2D0 U13 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  CKND2D0 U15 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  CKND0 U16 ( .CLK(Sel[3]), .CN(n11) );
  NR2XD0 U17 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U18 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2XD0 U19 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U20 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U21 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U22 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U23 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U25 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U27 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  INVD1 U28 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U29 ( .I(Sel[1]), .ZN(n2) );
endmodule


module Dec4_16_35 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U2 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D0 U3 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D0 U4 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D0 U5 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U6 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U7 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U8 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U9 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  ND2D0 U10 ( .A1(n11), .A2(n14), .ZN(n16) );
  ND2D0 U11 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D0 U12 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  ND2D0 U13 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND0 U14 ( .CLK(n3), .CN(n2) );
  INVD0 U15 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U16 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  CKND0 U17 ( .CLK(n11), .CN(n4) );
  INVD0 U18 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U19 ( .A1(n4), .A2(n14), .ZN(n18) );
  CKND2D0 U20 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U21 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  NR2XD0 U22 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U23 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U24 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U25 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U27 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U28 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  INVD1 U29 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
endmodule


module Dec4_16_36 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U2 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U3 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U4 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D0 U5 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U6 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  ND2D1 U7 ( .A1(n4), .A2(n14), .ZN(n18) );
  ND2D0 U8 ( .A1(n11), .A2(n14), .ZN(n16) );
  ND2D0 U9 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D0 U10 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  ND2D0 U11 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND0 U12 ( .CLK(n3), .CN(n2) );
  INVD0 U13 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U14 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  CKND0 U15 ( .CLK(n11), .CN(n4) );
  INVD0 U16 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U17 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U18 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  NR2XD0 U19 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U20 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U23 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U25 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U27 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U28 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  INVD1 U29 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
endmodule


module Dec4_16_37 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  ND2D1 U1 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  NR2D1 U2 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D1 U3 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2D0 U4 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U5 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2D0 U6 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  ND2D0 U7 ( .A1(n4), .A2(n11), .ZN(n15) );
  ND2D0 U8 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  ND2D0 U9 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  ND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n19) );
  CKND0 U11 ( .CLK(n3), .CN(n2) );
  INVD0 U12 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  INVD0 U14 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U15 ( .A1(n2), .A2(n1), .ZN(n16) );
  CKND2D0 U16 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  NR2XD0 U17 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2XD0 U18 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U19 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U20 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U21 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U22 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U24 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U25 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2XD0 U27 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  INVD1 U28 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U29 ( .I(Sel[2]), .ZN(n4) );
endmodule


module Dec4_16_38 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U2 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U3 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U4 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U5 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2D0 U6 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  ND2D1 U7 ( .A1(n4), .A2(n14), .ZN(n18) );
  ND2D0 U8 ( .A1(n11), .A2(n14), .ZN(n16) );
  ND2D0 U9 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  ND2D0 U10 ( .A1(Sel[3]), .A2(n11), .ZN(n21) );
  ND2D0 U11 ( .A1(n1), .A2(n3), .ZN(n20) );
  CKND0 U12 ( .CLK(n3), .CN(n2) );
  INVD0 U13 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U14 ( .A1(n4), .A2(Sel[3]), .ZN(n15) );
  CKND0 U15 ( .CLK(n11), .CN(n4) );
  INVD0 U16 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U17 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U18 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  CKND0 U19 ( .CLK(Sel[3]), .CN(n14) );
  NR2XD0 U20 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2XD0 U21 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U22 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U24 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U25 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U27 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U28 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U29 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
endmodule


module Dec4_16_39 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U2 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2D0 U3 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U4 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  ND2D0 U5 ( .A1(n14), .A2(n15), .ZN(n17) );
  INVD1 U6 ( .I(n2), .ZN(n1) );
  ND2D0 U7 ( .A1(n1), .A2(n4), .ZN(n23) );
  ND2D0 U8 ( .A1(Sel[3]), .A2(n14), .ZN(n22) );
  ND2D0 U9 ( .A1(n2), .A2(n4), .ZN(n21) );
  CKND0 U10 ( .CLK(n4), .CN(n3) );
  INVD0 U11 ( .I(Sel[1]), .ZN(n4) );
  CKND2D0 U12 ( .A1(n11), .A2(Sel[3]), .ZN(n16) );
  CKND0 U13 ( .CLK(n14), .CN(n11) );
  INVD0 U14 ( .I(Sel[0]), .ZN(n2) );
  CKND2D0 U15 ( .A1(n11), .A2(n15), .ZN(n19) );
  CKND2D0 U16 ( .A1(n3), .A2(n2), .ZN(n18) );
  CKND2D0 U17 ( .A1(n3), .A2(n1), .ZN(n20) );
  NR2XD0 U18 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2XD0 U19 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2XD0 U20 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2XD0 U21 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2XD0 U23 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2XD0 U24 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2XD0 U25 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U27 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U28 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U29 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  INVD1 U30 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U31 ( .I(Sel[2]), .ZN(n14) );
endmodule


module Dec4_16_40 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D0 U1 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U2 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2D0 U3 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U4 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2D0 U5 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  ND2D1 U6 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  ND2D0 U7 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U8 ( .A1(n1), .A2(n3), .ZN(n19) );
  ND2D0 U9 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND0 U10 ( .CLK(n3), .CN(n2) );
  INVD0 U11 ( .I(Sel[1]), .ZN(n3) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  INVD0 U13 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U14 ( .A1(n2), .A2(n1), .ZN(n16) );
  CKND2D0 U15 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  CKND2D0 U16 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  NR2XD0 U17 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2XD0 U18 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2XD0 U19 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U25 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2XD0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U27 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  INVD1 U28 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U29 ( .I(Sel[2]), .ZN(n4) );
endmodule


module Dec4_16_41 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  ND2D1 U1 ( .A1(n3), .A2(n11), .ZN(n17) );
  NR2D1 U2 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D1 U3 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  INVD1 U4 ( .I(n4), .ZN(n3) );
  NR2D0 U5 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2D0 U6 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U7 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U8 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U9 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U10 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  ND2D1 U11 ( .A1(n3), .A2(Sel[3]), .ZN(n14) );
  CKND2D0 U12 ( .A1(n1), .A2(n2), .ZN(n19) );
  CKND2D0 U13 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U16 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U17 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  NR2XD0 U18 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U19 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2XD0 U20 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U21 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  NR2XD0 U25 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U27 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U28 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U29 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_42 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  ND2D1 U1 ( .A1(n3), .A2(n14), .ZN(n18) );
  INVD1 U2 ( .I(n4), .ZN(n3) );
  NR2D0 U3 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U4 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U5 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D0 U6 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U7 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U8 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U9 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D0 U10 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2D0 U11 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  CKND2D0 U12 ( .A1(n1), .A2(n2), .ZN(n20) );
  CKND2D0 U13 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n19) );
  CKND2D0 U15 ( .A1(n3), .A2(n11), .ZN(n15) );
  CKND0 U16 ( .CLK(n14), .CN(n11) );
  CKND2D0 U17 ( .A1(Sel[1]), .A2(n1), .ZN(n17) );
  CKND2D0 U18 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND2D0 U19 ( .A1(Sel[0]), .A2(n2), .ZN(n22) );
  NR2XD0 U20 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U21 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U22 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U23 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U24 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U25 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2XD0 U26 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  INVD1 U27 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U28 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U29 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U30 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_43 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U3 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U4 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2D0 U5 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U6 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2D0 U7 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2D0 U8 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  CKND2D0 U9 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U10 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U11 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U15 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U16 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND0 U17 ( .CLK(Sel[1]), .CN(n2) );
  NR2XD0 U18 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U19 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  NR2XD0 U24 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2XD0 U25 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_44 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  ND2D1 U1 ( .A1(n4), .A2(n15), .ZN(n19) );
  INVD1 U2 ( .I(n11), .ZN(n4) );
  NR2D0 U3 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U4 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U5 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U6 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2D0 U7 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2D0 U8 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  CKND2D0 U9 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD1 U10 ( .I(n3), .ZN(n2) );
  CKND2D0 U11 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U12 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U13 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND0 U14 ( .CLK(n15), .CN(n14) );
  CKND2D0 U15 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U16 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND2D0 U17 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  NR2XD0 U18 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U19 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U21 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U22 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2XD0 U24 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2XD0 U25 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2XD0 U26 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2XD0 U27 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  INVD1 U28 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U29 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U31 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_45 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2D0 U3 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U5 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U6 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U7 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2D0 U8 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U9 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  CKND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n19) );
  INVD1 U11 ( .I(n3), .ZN(n2) );
  CKND2D0 U12 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U13 ( .A1(n2), .A2(Sel[0]), .ZN(n18) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n14) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U16 ( .A1(n2), .A2(n1), .ZN(n16) );
  CKND2D0 U17 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U18 ( .A1(Sel[0]), .A2(n3), .ZN(n21) );
  NR2XD0 U19 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2XD0 U20 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2XD0 U21 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2XD0 U24 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U25 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U27 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U28 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U29 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_46 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D0 U1 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2D0 U2 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
  NR2D0 U3 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U5 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U6 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2D0 U7 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2D0 U8 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  ND2D1 U9 ( .A1(n4), .A2(n15), .ZN(n19) );
  CKND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD1 U11 ( .I(n11), .ZN(n4) );
  INVD1 U12 ( .I(n3), .ZN(n2) );
  CKND2D0 U13 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U14 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U15 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND0 U16 ( .CLK(n15), .CN(n14) );
  CKND2D0 U17 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U18 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND2D0 U19 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  NR2XD0 U20 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2XD0 U21 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U22 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2XD0 U23 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U24 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2XD0 U25 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U27 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  INVD1 U28 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U29 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U30 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U31 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_47 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D0 U3 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U4 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U5 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U6 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2D0 U7 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D0 U8 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D0 U9 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  CKND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n20) );
  INVD1 U11 ( .I(n3), .ZN(n2) );
  CKND2D0 U12 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND2D0 U13 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  CKND0 U15 ( .CLK(n14), .CN(n11) );
  CKND2D0 U16 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  CKND2D0 U17 ( .A1(n2), .A2(n1), .ZN(n17) );
  CKND2D0 U18 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND2D0 U19 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  NR2XD0 U20 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2XD0 U21 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U22 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2XD0 U23 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U25 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U26 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  INVD1 U27 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U28 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U29 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U30 ( .I(Sel[0]), .ZN(n1) );
endmodule


module Dec4_16_48 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D1 U2 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D1 U3 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2D1 U4 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2D1 U5 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  INVD1 U6 ( .I(n14), .ZN(n11) );
  INVD0 U7 ( .I(Sel[1]), .ZN(n2) );
  INVD1 U8 ( .I(n4), .ZN(n3) );
  INVD0 U9 ( .I(Sel[2]), .ZN(n4) );
  INVD0 U10 ( .I(Sel[0]), .ZN(n1) );
  INVD0 U11 ( .I(Sel[3]), .ZN(n14) );
  ND2D1 U12 ( .A1(n4), .A2(n14), .ZN(n16) );
  ND2D1 U13 ( .A1(n1), .A2(n2), .ZN(n20) );
  NR2XD0 U14 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U15 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U16 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U17 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U18 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U19 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U20 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2XD0 U21 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U22 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U23 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U24 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  ND2D1 U25 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n19) );
  ND2D1 U26 ( .A1(n3), .A2(n11), .ZN(n15) );
  ND2D1 U27 ( .A1(n3), .A2(n14), .ZN(n18) );
  ND2D1 U28 ( .A1(Sel[1]), .A2(n1), .ZN(n17) );
  ND2D1 U29 ( .A1(n11), .A2(n4), .ZN(n21) );
  ND2D1 U30 ( .A1(Sel[0]), .A2(n2), .ZN(n22) );
endmodule


module Dec4_16_49 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D0 U1 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U2 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U3 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U4 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2D0 U5 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2D0 U6 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2D0 U7 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2D0 U8 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  ND2D1 U9 ( .A1(n4), .A2(n15), .ZN(n19) );
  ND2D0 U10 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD1 U11 ( .I(n11), .ZN(n4) );
  INVD1 U12 ( .I(n3), .ZN(n2) );
  CKND2D0 U13 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U14 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U15 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND0 U16 ( .CLK(n15), .CN(n14) );
  CKND2D0 U17 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U18 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND2D0 U19 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  CKND0 U20 ( .CLK(Sel[0]), .CN(n1) );
  NR2XD0 U21 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2XD0 U22 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U23 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2XD0 U25 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  INVD1 U26 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U27 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U28 ( .I(Sel[2]), .ZN(n11) );
  NR2D0 U29 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U31 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
endmodule


module Dec4_16_50 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  NR2D1 U1 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2D0 U5 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2D0 U6 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2D0 U7 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2D0 U8 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2D0 U9 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2D0 U10 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  ND2D0 U11 ( .A1(n1), .A2(n2), .ZN(n20) );
  INVD1 U12 ( .I(n4), .ZN(n3) );
  CKND2D0 U13 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n19) );
  CKND2D0 U15 ( .A1(n3), .A2(n11), .ZN(n15) );
  CKND0 U16 ( .CLK(n14), .CN(n11) );
  CKND2D0 U17 ( .A1(n3), .A2(n14), .ZN(n18) );
  CKND2D0 U18 ( .A1(Sel[1]), .A2(n1), .ZN(n17) );
  CKND2D0 U19 ( .A1(n11), .A2(n4), .ZN(n21) );
  CKND2D0 U20 ( .A1(Sel[0]), .A2(n2), .ZN(n22) );
  CKND0 U21 ( .CLK(Sel[1]), .CN(n2) );
  NR2XD0 U22 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U23 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U24 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  INVD1 U25 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U26 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U27 ( .I(Sel[0]), .ZN(n1) );
  NR2D0 U28 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U29 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
  NR2D0 U30 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
endmodule


module Dec4_16_51 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2D0 U2 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U5 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2D0 U6 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  NR2D0 U7 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  ND2D1 U8 ( .A1(n4), .A2(n15), .ZN(n19) );
  ND2D0 U9 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD1 U10 ( .I(n11), .ZN(n4) );
  INVD1 U11 ( .I(n3), .ZN(n2) );
  CKND2D0 U12 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U13 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U14 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND0 U15 ( .CLK(n15), .CN(n14) );
  CKND2D0 U16 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U17 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND2D0 U18 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  NR2XD0 U19 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2XD0 U20 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2XD0 U22 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2XD0 U24 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  INVD1 U25 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U26 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n1) );
  NR2D0 U29 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U31 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
endmodule


module Dec4_16_52 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
;

  NR2D1 U1 ( .A1(n19), .A2(n18), .ZN(Hot[6]) );
  NR2D0 U2 ( .A1(n23), .A2(n22), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n22), .A2(n18), .ZN(Hot[10]) );
  NR2D0 U4 ( .A1(n20), .A2(n19), .ZN(Hot[7]) );
  NR2D0 U5 ( .A1(n22), .A2(n21), .ZN(Hot[8]) );
  NR2D0 U6 ( .A1(n21), .A2(n19), .ZN(Hot[4]) );
  NR2D0 U7 ( .A1(n23), .A2(n19), .ZN(Hot[5]) );
  NR2D0 U8 ( .A1(n20), .A2(n17), .ZN(Hot[3]) );
  NR2D0 U9 ( .A1(n18), .A2(n17), .ZN(Hot[2]) );
  NR2D0 U10 ( .A1(n21), .A2(n17), .ZN(Hot[0]) );
  ND2D0 U11 ( .A1(n1), .A2(n3), .ZN(n21) );
  INVD1 U12 ( .I(n11), .ZN(n4) );
  INVD1 U13 ( .I(n3), .ZN(n2) );
  CKND2D0 U14 ( .A1(n11), .A2(n15), .ZN(n17) );
  CKND2D0 U15 ( .A1(n2), .A2(Sel[0]), .ZN(n20) );
  CKND2D0 U16 ( .A1(n4), .A2(n14), .ZN(n16) );
  CKND0 U17 ( .CLK(n15), .CN(n14) );
  CKND2D0 U18 ( .A1(n4), .A2(n15), .ZN(n19) );
  CKND2D0 U19 ( .A1(n2), .A2(n1), .ZN(n18) );
  CKND2D0 U20 ( .A1(n14), .A2(n11), .ZN(n22) );
  CKND2D0 U21 ( .A1(Sel[0]), .A2(n3), .ZN(n23) );
  NR2XD0 U22 ( .A1(n21), .A2(n16), .ZN(Hot[12]) );
  NR2XD0 U23 ( .A1(n22), .A2(n20), .ZN(Hot[11]) );
  NR2XD0 U24 ( .A1(n23), .A2(n17), .ZN(Hot[1]) );
  INVD1 U25 ( .I(Sel[3]), .ZN(n15) );
  INVD1 U26 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U27 ( .I(Sel[2]), .ZN(n11) );
  INVD1 U28 ( .I(Sel[0]), .ZN(n1) );
  NR2D0 U29 ( .A1(n18), .A2(n16), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n20), .A2(n16), .ZN(Hot[15]) );
  NR2D0 U31 ( .A1(n23), .A2(n16), .ZN(Hot[13]) );
endmodule


module Dec4_16_53 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  NR2D0 U2 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U3 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D0 U4 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D1 U5 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  CKND2D1 U6 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  NR2XD0 U7 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
  ND2D1 U8 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D1 U9 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D1 U10 ( .A1(n3), .A2(n4), .ZN(n13) );
  ND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  NR2D0 U12 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2D0 U13 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND0 U17 ( .CLK(Sel[0]), .CN(n1) );
  CKND0 U18 ( .CLK(Sel[2]), .CN(n3) );
  NR2XD0 U19 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U20 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2XD0 U21 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U22 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U23 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  INVD1 U24 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U25 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U28 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
endmodule


module Dec4_16_54 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U2 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2D0 U3 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2D0 U4 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U5 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D0 U6 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U7 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U8 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  INVD0 U9 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U10 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U12 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U13 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  CKND0 U14 ( .CLK(Sel[2]), .CN(n3) );
  NR2XD0 U15 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2XD0 U16 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U17 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U18 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U19 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U20 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U21 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U25 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_55 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D0 U1 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2D0 U2 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2D0 U3 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2D0 U4 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U5 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  NR2XD0 U6 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  ND2D0 U7 ( .A1(n1), .A2(n2), .ZN(n17) );
  CKND2D0 U8 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U9 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  INVD0 U10 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U11 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U13 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2XD0 U15 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2XD0 U16 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2XD0 U17 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2XD0 U18 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2XD0 U19 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U20 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U23 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U25 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_56 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D0 U1 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2D0 U2 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U3 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D0 U4 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D0 U5 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2D0 U6 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2D0 U7 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U8 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D0 U9 ( .A1(n1), .A2(n2), .ZN(n17) );
  INVD0 U10 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U11 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U12 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2XD0 U17 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2XD0 U18 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U19 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2XD0 U20 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U23 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U25 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_57 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U2 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U3 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2D0 U4 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U5 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2D0 U6 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2D0 U7 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U8 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  ND2D0 U9 ( .A1(n1), .A2(n2), .ZN(n19) );
  INVD0 U10 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U11 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U12 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U13 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  CKND2D0 U14 ( .A1(n3), .A2(Sel[3]), .ZN(n14) );
  CKND0 U15 ( .CLK(n4), .CN(n3) );
  CKND2D0 U16 ( .A1(n3), .A2(n11), .ZN(n17) );
  CKND2D0 U17 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U18 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  NR2XD0 U19 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U20 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2XD0 U22 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U25 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U26 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U29 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
endmodule


module Dec4_16_58 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D0 U1 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2D0 U2 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U3 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U4 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2D0 U5 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U6 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  ND2D1 U7 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  ND2D0 U8 ( .A1(n1), .A2(n2), .ZN(n19) );
  INVD0 U9 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U10 ( .A1(n3), .A2(n11), .ZN(n15) );
  CKND2D0 U11 ( .A1(n4), .A2(n3), .ZN(n20) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(n4), .ZN(n14) );
  INVD1 U13 ( .I(n11), .ZN(n4) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  NR2XD0 U17 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U18 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U19 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U20 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U21 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2XD0 U22 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U25 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U26 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U29 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
endmodule


module Dec4_16_59 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D1 U2 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U3 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U4 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U5 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2D0 U6 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2D0 U7 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U8 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  NR2D0 U9 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  ND2D0 U10 ( .A1(n1), .A2(n2), .ZN(n19) );
  INVD0 U11 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U12 ( .A1(n3), .A2(n11), .ZN(n15) );
  CKND2D0 U13 ( .A1(n4), .A2(n3), .ZN(n20) );
  CKND2D0 U14 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(n4), .ZN(n14) );
  INVD1 U16 ( .I(n11), .ZN(n4) );
  CKND2D0 U17 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U18 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U19 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  CKND0 U20 ( .CLK(Sel[1]), .CN(n2) );
  NR2XD0 U21 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U22 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U23 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  INVD1 U24 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U25 ( .I(Sel[2]), .ZN(n3) );
  NR2D0 U26 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U29 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
endmodule


module Dec4_16_60 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  INVD0 U1 ( .I(Sel[3]), .ZN(n4) );
  NR2D0 U2 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  NR2D0 U3 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U4 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D0 U5 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D0 U6 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2D0 U7 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2D0 U8 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U9 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  ND2D0 U10 ( .A1(n1), .A2(n2), .ZN(n17) );
  INVD0 U11 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U12 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U13 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U15 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U17 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2XD0 U18 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2XD0 U19 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U20 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2XD0 U21 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U22 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  INVD1 U23 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U25 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_61 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D1 U1 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  NR2D0 U2 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U3 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U4 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2D0 U5 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U6 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2D0 U7 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  ND2D0 U8 ( .A1(n1), .A2(n2), .ZN(n19) );
  INVD0 U9 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U10 ( .A1(n4), .A2(n11), .ZN(n15) );
  CKND2D0 U11 ( .A1(Sel[3]), .A2(n4), .ZN(n20) );
  CKND2D0 U12 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  CKND2D0 U13 ( .A1(n3), .A2(Sel[3]), .ZN(n14) );
  CKND0 U14 ( .CLK(n4), .CN(n3) );
  CKND2D0 U15 ( .A1(n3), .A2(n11), .ZN(n17) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U17 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  NR2XD0 U18 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U19 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2XD0 U20 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U21 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U22 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n4) );
  INVD1 U25 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U26 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U29 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
endmodule


module Dec4_16_62 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21;

  NR2D0 U1 ( .A1(n20), .A2(n19), .ZN(Hot[8]) );
  NR2D0 U2 ( .A1(n21), .A2(n17), .ZN(Hot[5]) );
  NR2D0 U3 ( .A1(n17), .A2(n16), .ZN(Hot[6]) );
  NR2D0 U4 ( .A1(n19), .A2(n17), .ZN(Hot[4]) );
  NR2D0 U5 ( .A1(n16), .A2(n15), .ZN(Hot[2]) );
  NR2D0 U6 ( .A1(n21), .A2(n15), .ZN(Hot[1]) );
  ND2D1 U7 ( .A1(Sel[0]), .A2(n2), .ZN(n21) );
  ND2D0 U8 ( .A1(n1), .A2(n2), .ZN(n19) );
  INVD0 U9 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U10 ( .A1(n3), .A2(n11), .ZN(n15) );
  CKND2D0 U11 ( .A1(n4), .A2(n3), .ZN(n20) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(n4), .ZN(n14) );
  INVD1 U13 ( .I(n11), .ZN(n4) );
  CKND2D0 U14 ( .A1(Sel[2]), .A2(n11), .ZN(n17) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(n1), .ZN(n16) );
  CKND2D0 U16 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n18) );
  NR2XD0 U17 ( .A1(n19), .A2(n14), .ZN(Hot[12]) );
  NR2XD0 U18 ( .A1(n18), .A2(n17), .ZN(Hot[7]) );
  NR2XD0 U19 ( .A1(n20), .A2(n16), .ZN(Hot[10]) );
  NR2XD0 U20 ( .A1(n19), .A2(n15), .ZN(Hot[0]) );
  NR2XD0 U21 ( .A1(n18), .A2(n15), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n21), .A2(n20), .ZN(Hot[9]) );
  INVD1 U23 ( .I(Sel[3]), .ZN(n11) );
  INVD1 U24 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U25 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U26 ( .A1(n16), .A2(n14), .ZN(Hot[14]) );
  NR2D0 U27 ( .A1(n21), .A2(n14), .ZN(Hot[13]) );
  NR2D0 U28 ( .A1(n18), .A2(n14), .ZN(Hot[15]) );
  NR2D0 U29 ( .A1(n20), .A2(n18), .ZN(Hot[11]) );
endmodule


module Dec4_16_63 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n13, n14, n15, n16, n17, n18, n19;

  NR2D1 U1 ( .A1(n17), .A2(n11), .ZN(Hot[12]) );
  NR2D0 U2 ( .A1(n19), .A2(n15), .ZN(Hot[5]) );
  NR2D0 U3 ( .A1(n16), .A2(n15), .ZN(Hot[7]) );
  NR2D0 U4 ( .A1(n17), .A2(n15), .ZN(Hot[4]) );
  NR2D0 U5 ( .A1(n19), .A2(n13), .ZN(Hot[1]) );
  NR2D0 U6 ( .A1(n19), .A2(n18), .ZN(Hot[9]) );
  ND2D0 U7 ( .A1(n1), .A2(n2), .ZN(n17) );
  INVD0 U8 ( .I(Sel[0]), .ZN(n1) );
  CKND2D0 U9 ( .A1(n3), .A2(n4), .ZN(n13) );
  CKND2D0 U10 ( .A1(Sel[3]), .A2(n3), .ZN(n18) );
  CKND2D0 U11 ( .A1(Sel[0]), .A2(n2), .ZN(n19) );
  CKND2D0 U12 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n11) );
  CKND2D0 U13 ( .A1(Sel[2]), .A2(n4), .ZN(n15) );
  CKND2D0 U14 ( .A1(Sel[1]), .A2(n1), .ZN(n14) );
  CKND2D0 U15 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n16) );
  NR2XD0 U16 ( .A1(n15), .A2(n14), .ZN(Hot[6]) );
  NR2XD0 U17 ( .A1(n18), .A2(n14), .ZN(Hot[10]) );
  NR2XD0 U18 ( .A1(n17), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n14), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U20 ( .A1(n16), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U21 ( .A1(n18), .A2(n17), .ZN(Hot[8]) );
  INVD1 U22 ( .I(Sel[3]), .ZN(n4) );
  INVD1 U23 ( .I(Sel[2]), .ZN(n3) );
  INVD1 U24 ( .I(Sel[1]), .ZN(n2) );
  NR2D0 U25 ( .A1(n14), .A2(n11), .ZN(Hot[14]) );
  NR2D0 U26 ( .A1(n19), .A2(n11), .ZN(Hot[13]) );
  NR2D0 U27 ( .A1(n16), .A2(n11), .ZN(Hot[15]) );
  NR2D0 U28 ( .A1(n18), .A2(n16), .ZN(Hot[11]) );
endmodule


module Dec4_16_64 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n11, n14, n15, n16, n17, n18, n19, n20, n21, n22;

  CKND2D1 U1 ( .A1(Sel[0]), .A2(n3), .ZN(n22) );
  CKND2D1 U2 ( .A1(n2), .A2(Sel[0]), .ZN(n19) );
  INVD1 U3 ( .I(n3), .ZN(n2) );
  INVD0 U4 ( .I(Sel[1]), .ZN(n3) );
  INVD0 U5 ( .I(Sel[2]), .ZN(n4) );
  INVD0 U6 ( .I(Sel[0]), .ZN(n1) );
  INVD1 U7 ( .I(n14), .ZN(n11) );
  INVD0 U8 ( .I(Sel[3]), .ZN(n14) );
  ND2D1 U9 ( .A1(n4), .A2(n14), .ZN(n16) );
  ND2D1 U10 ( .A1(n1), .A2(n3), .ZN(n20) );
  NR2XD0 U11 ( .A1(n20), .A2(n15), .ZN(Hot[12]) );
  NR2XD0 U12 ( .A1(n22), .A2(n15), .ZN(Hot[13]) );
  NR2XD0 U13 ( .A1(n20), .A2(n18), .ZN(Hot[4]) );
  NR2XD0 U14 ( .A1(n22), .A2(n18), .ZN(Hot[5]) );
  NR2XD0 U15 ( .A1(n18), .A2(n17), .ZN(Hot[6]) );
  NR2XD0 U16 ( .A1(n19), .A2(n18), .ZN(Hot[7]) );
  NR2XD0 U17 ( .A1(n21), .A2(n17), .ZN(Hot[10]) );
  NR2XD0 U18 ( .A1(n20), .A2(n16), .ZN(Hot[0]) );
  NR2XD0 U19 ( .A1(n22), .A2(n16), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n17), .A2(n16), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n19), .A2(n16), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n21), .A2(n20), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n22), .A2(n21), .ZN(Hot[9]) );
  ND2D1 U24 ( .A1(Sel[2]), .A2(n11), .ZN(n15) );
  ND2D1 U25 ( .A1(Sel[2]), .A2(n14), .ZN(n18) );
  ND2D1 U26 ( .A1(n2), .A2(n1), .ZN(n17) );
  ND2D1 U27 ( .A1(n11), .A2(n4), .ZN(n21) );
  NR2D0 U28 ( .A1(n21), .A2(n19), .ZN(Hot[11]) );
  NR2D0 U29 ( .A1(n17), .A2(n15), .ZN(Hot[14]) );
  NR2D0 U30 ( .A1(n19), .A2(n15), .ZN(Hot[15]) );
endmodule


module Dec4_16_65 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n13, n14, n15, n16, n17, n18, n19, n20;

  INVD1 U1 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U2 ( .I(Sel[2]), .ZN(n1) );
  INVD1 U3 ( .I(Sel[1]), .ZN(n3) );
  ND2D1 U4 ( .A1(n1), .A2(n14), .ZN(n13) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(n14), .ZN(n16) );
  ND2D1 U6 ( .A1(Sel[3]), .A2(n1), .ZN(n19) );
  ND2D1 U7 ( .A1(Sel[0]), .A2(n3), .ZN(n20) );
  ND2D1 U8 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n4) );
  NR2D1 U9 ( .A1(n18), .A2(n13), .ZN(Hot[0]) );
  NR2D1 U10 ( .A1(n20), .A2(n13), .ZN(Hot[1]) );
  NR2D1 U11 ( .A1(n15), .A2(n13), .ZN(Hot[2]) );
  ND2D1 U12 ( .A1(n2), .A2(n3), .ZN(n18) );
  NR2XD0 U13 ( .A1(n19), .A2(n15), .ZN(Hot[10]) );
  NR2XD0 U14 ( .A1(n20), .A2(n19), .ZN(Hot[9]) );
  NR2XD0 U15 ( .A1(n18), .A2(n4), .ZN(Hot[12]) );
  NR2XD0 U16 ( .A1(n15), .A2(n4), .ZN(Hot[14]) );
  NR2XD0 U17 ( .A1(n20), .A2(n16), .ZN(Hot[5]) );
  NR2XD0 U18 ( .A1(n17), .A2(n16), .ZN(Hot[7]) );
  NR2XD0 U19 ( .A1(n16), .A2(n15), .ZN(Hot[6]) );
  NR2XD0 U20 ( .A1(n18), .A2(n16), .ZN(Hot[4]) );
  NR2XD0 U21 ( .A1(n17), .A2(n4), .ZN(Hot[15]) );
  NR2XD0 U22 ( .A1(n19), .A2(n18), .ZN(Hot[8]) );
  NR2XD0 U23 ( .A1(n19), .A2(n17), .ZN(Hot[11]) );
  NR2XD0 U24 ( .A1(n20), .A2(n4), .ZN(Hot[13]) );
  NR2D0 U25 ( .A1(n17), .A2(n13), .ZN(Hot[3]) );
  ND2D1 U26 ( .A1(Sel[1]), .A2(n2), .ZN(n15) );
  CKND0 U27 ( .CLK(Sel[0]), .CN(n2) );
  ND2D1 U28 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n17) );
endmodule


module Dec4_16_66 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n13, n14, n15, n16, n17, n18, n19, n20;

  INVD1 U1 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U2 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U3 ( .I(Sel[0]), .ZN(n2) );
  ND2D1 U4 ( .A1(Sel[3]), .A2(n1), .ZN(n19) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n4) );
  ND2D0 U6 ( .A1(Sel[2]), .A2(n14), .ZN(n16) );
  ND2D1 U7 ( .A1(n1), .A2(n14), .ZN(n13) );
  CKND2D1 U8 ( .A1(Sel[0]), .A2(n3), .ZN(n20) );
  ND2D0 U9 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n17) );
  CKND2D1 U10 ( .A1(Sel[1]), .A2(n2), .ZN(n15) );
  ND2D1 U11 ( .A1(n2), .A2(n3), .ZN(n18) );
  NR2XD0 U12 ( .A1(n18), .A2(n13), .ZN(Hot[0]) );
  NR2XD0 U13 ( .A1(n15), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U14 ( .A1(n17), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U15 ( .A1(n18), .A2(n16), .ZN(Hot[4]) );
  NR2XD0 U16 ( .A1(n17), .A2(n16), .ZN(Hot[7]) );
  NR2XD0 U17 ( .A1(n19), .A2(n18), .ZN(Hot[8]) );
  NR2XD0 U18 ( .A1(n16), .A2(n15), .ZN(Hot[6]) );
  NR2XD0 U19 ( .A1(n19), .A2(n15), .ZN(Hot[10]) );
  NR2XD0 U20 ( .A1(n20), .A2(n19), .ZN(Hot[9]) );
  NR2XD0 U21 ( .A1(n18), .A2(n4), .ZN(Hot[12]) );
  NR2XD0 U22 ( .A1(n20), .A2(n4), .ZN(Hot[13]) );
  NR2XD0 U23 ( .A1(n15), .A2(n4), .ZN(Hot[14]) );
  NR2XD0 U24 ( .A1(n19), .A2(n17), .ZN(Hot[11]) );
  NR2XD0 U25 ( .A1(n20), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U26 ( .A1(n20), .A2(n16), .ZN(Hot[5]) );
  NR2XD0 U27 ( .A1(n17), .A2(n4), .ZN(Hot[15]) );
  CKND0 U28 ( .CLK(Sel[2]), .CN(n1) );
endmodule


module Dec4_16_67 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n13, n14, n15, n16, n17, n18, n19, n20;

  INVD1 U1 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U2 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U3 ( .I(Sel[0]), .ZN(n2) );
  ND2D1 U4 ( .A1(Sel[3]), .A2(n1), .ZN(n19) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n4) );
  ND2D0 U6 ( .A1(Sel[2]), .A2(n14), .ZN(n16) );
  CKND2D1 U7 ( .A1(Sel[0]), .A2(n3), .ZN(n20) );
  CKND2D1 U8 ( .A1(Sel[1]), .A2(n2), .ZN(n15) );
  INVD0 U9 ( .I(Sel[2]), .ZN(n1) );
  NR2XD0 U10 ( .A1(n18), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U11 ( .A1(n1), .A2(n14), .ZN(n13) );
  ND2D1 U12 ( .A1(n2), .A2(n3), .ZN(n18) );
  NR2XD0 U13 ( .A1(n17), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U14 ( .A1(n18), .A2(n16), .ZN(Hot[4]) );
  NR2XD0 U15 ( .A1(n20), .A2(n16), .ZN(Hot[5]) );
  NR2XD0 U16 ( .A1(n19), .A2(n18), .ZN(Hot[8]) );
  NR2XD0 U17 ( .A1(n16), .A2(n15), .ZN(Hot[6]) );
  NR2XD0 U18 ( .A1(n19), .A2(n15), .ZN(Hot[10]) );
  NR2XD0 U19 ( .A1(n20), .A2(n19), .ZN(Hot[9]) );
  NR2XD0 U20 ( .A1(n18), .A2(n4), .ZN(Hot[12]) );
  NR2XD0 U21 ( .A1(n20), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U22 ( .A1(n20), .A2(n4), .ZN(Hot[13]) );
  NR2XD0 U23 ( .A1(n19), .A2(n17), .ZN(Hot[11]) );
  NR2XD0 U24 ( .A1(n15), .A2(n4), .ZN(Hot[14]) );
  NR2XD0 U25 ( .A1(n15), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U26 ( .A1(n17), .A2(n16), .ZN(Hot[7]) );
  NR2XD0 U27 ( .A1(n17), .A2(n4), .ZN(Hot[15]) );
  ND2D1 U28 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n17) );
endmodule


module Dec4_16_68 ( Hot, Sel );
  output [15:0] Hot;
  input [3:0] Sel;
  wire   n1, n2, n3, n4, n13, n14, n15, n16, n17, n18, n19, n20;

  INVD1 U1 ( .I(Sel[3]), .ZN(n14) );
  INVD1 U2 ( .I(Sel[1]), .ZN(n3) );
  INVD1 U3 ( .I(Sel[0]), .ZN(n2) );
  ND2D1 U4 ( .A1(Sel[3]), .A2(n1), .ZN(n19) );
  ND2D1 U5 ( .A1(Sel[2]), .A2(Sel[3]), .ZN(n4) );
  ND2D1 U6 ( .A1(Sel[1]), .A2(Sel[0]), .ZN(n17) );
  ND2D0 U7 ( .A1(Sel[2]), .A2(n14), .ZN(n16) );
  CKND2D1 U8 ( .A1(Sel[0]), .A2(n3), .ZN(n20) );
  CKND2D1 U9 ( .A1(Sel[1]), .A2(n2), .ZN(n15) );
  INVD0 U10 ( .I(Sel[2]), .ZN(n1) );
  NR2XD0 U11 ( .A1(n18), .A2(n13), .ZN(Hot[0]) );
  ND2D1 U12 ( .A1(n1), .A2(n14), .ZN(n13) );
  ND2D1 U13 ( .A1(n2), .A2(n3), .ZN(n18) );
  NR2XD0 U14 ( .A1(n18), .A2(n4), .ZN(Hot[12]) );
  NR2XD0 U15 ( .A1(n20), .A2(n4), .ZN(Hot[13]) );
  NR2XD0 U16 ( .A1(n15), .A2(n4), .ZN(Hot[14]) );
  NR2XD0 U17 ( .A1(n17), .A2(n4), .ZN(Hot[15]) );
  NR2XD0 U18 ( .A1(n19), .A2(n17), .ZN(Hot[11]) );
  NR2XD0 U19 ( .A1(n20), .A2(n13), .ZN(Hot[1]) );
  NR2XD0 U20 ( .A1(n15), .A2(n13), .ZN(Hot[2]) );
  NR2XD0 U21 ( .A1(n17), .A2(n13), .ZN(Hot[3]) );
  NR2XD0 U22 ( .A1(n18), .A2(n16), .ZN(Hot[4]) );
  NR2XD0 U23 ( .A1(n20), .A2(n16), .ZN(Hot[5]) );
  NR2XD0 U24 ( .A1(n17), .A2(n16), .ZN(Hot[7]) );
  NR2XD0 U25 ( .A1(n19), .A2(n18), .ZN(Hot[8]) );
  NR2XD0 U26 ( .A1(n16), .A2(n15), .ZN(Hot[6]) );
  NR2XD0 U27 ( .A1(n19), .A2(n15), .ZN(Hot[10]) );
  NR2XD0 U28 ( .A1(n20), .A2(n19), .ZN(Hot[9]) );
endmodule

