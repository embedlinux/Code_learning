library verilog;
use verilog.vl_types.all;
entity tlv5618_tb is
end tlv5618_tb;
