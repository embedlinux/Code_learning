`timescale 1ns/1ns

module tlv5618(
	Clk,
	Rst_n,
	
	DAC_DATA,
	Start,
	Set_Done,
	DIV_PARAM,
	
	CS_N,
	DIN,
	SCLK,
	DAC_State
);

	input Clk;
	input Rst_n;
	input [15:0]DAC_DATA;
	input Start;
	output Set_Done;
	input [7:0]DIV_PARAM;
	
	output reg CS_N;
	output reg DIN;
	output reg SCLK;
	output DAC_State;
	
	assign DAC_State = CS_N;
	
	reg [15:0]r_DAC_DATA;
	
	reg [7:0]DIV_CNT;//分频计数器
	reg SCLK2X;//2倍SCLK的采样时钟
	
	reg [5:0]SCLK_GEN_CNT;//SCLK生成暨序列机计数器
	
	reg en;//转换使能信号
	
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		en  <= 1'b0;
	else if(Start)
		en  <= 1'b1;
	else if(Set_Done)
		en  <= 1'b0;
	else
		en  <= en;

	//生成2倍SCLK使能时钟计数器
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		DIV_CNT  <= 8'd0;
	else if(en)begin
		if(DIV_CNT == (DIV_PARAM - 1'b1))
			DIV_CNT  <= 8'd0;
		else 
			DIV_CNT  <= DIV_CNT + 1'b1;
	end else	
		DIV_CNT  <= 8'd0;

	//生成2倍SCLK使能时钟计数器
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		SCLK2X  <= 1'b0;
	else if(en && (DIV_CNT == (DIV_PARAM - 1'b1)))
		SCLK2X  <= 1'b1;
	else
		SCLK2X  <= 1'b0;
		
	//生成序列计数器
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		SCLK_GEN_CNT  <= 6'd0;
	else if(SCLK2X && en)begin
		if(SCLK_GEN_CNT == 6'd32)
			SCLK_GEN_CNT  <= 6'd0;
		else
			SCLK_GEN_CNT  <= SCLK_GEN_CNT + 1'd1;
	end else
		SCLK_GEN_CNT  <= SCLK_GEN_CNT;

	//依次将数据移出到DAC芯片		
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)begin
		DIN  <= 1'b1;
		SCLK  <= 1'b0;
		r_DAC_DATA  <= 16'd0;
	end else begin
		if(Start)//收到开始发送命令时，寄存DAC_DATA值	
			r_DAC_DATA  <= DAC_DATA;
		if(!Set_Done && SCLK2X) begin
			if(!SCLK_GEN_CNT[0])begin	//偶数，0,2,4,6,8,10,12,14,16,18,20,22,24,26,28,30:
				SCLK  <= 1'b1; 
				DIN  <= r_DAC_DATA[15]; 
				r_DAC_DATA  <= r_DAC_DATA << 1;
			end else	 //奇数，1,3,5,7,9,11,13,15,17,19,21,23,25,27,29,31:
				SCLK  <= 1'b0;
		end
	end
	
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		CS_N  <= 1'b1;
	else if(en && SCLK2X)
		CS_N  <= SCLK_GEN_CNT[5];
	else 
		CS_N  <= CS_N;
		
	assign Set_Done = SCLK_GEN_CNT[5] && SCLK2X;
	
endmodule
