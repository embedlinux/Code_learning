// *****************************************************************
// Specman Elite Verilog stubs file: specman.v
// Topmost e module: test_cpu.e
// Generated using seed = 1
// Date: Tue May 10 13:30:33 2005
// Specman Elite version: 4.3.1
// *****************************************************************



//               Verilog time                
// ================================================================

`timescale 1ns/1ns


module specman;


    //               Stub attributes section               
    // ================================================================

    parameter sn_version_id = 658186680;   /* Stub checksum */
    parameter sn_version_date = 131102; /* Stub version */
    parameter sn_use_wave = 1; /* specman_wave module existance*/
    parameter sn_declarations_num = 1; /* The number of reflected HDL declarations */


    //               General section               
    // ================================================================

    event sn_never_happens;
    always @sn_never_happens begin
         $sn();
    end
    reg sn_register_memory;
    event sn_register_memory_event;
    initial begin
        sn_register_memory=0;
    end
    always @(sn_register_memory_event) begin
        sn_register_memory=1;
    end
    initial begin

        ->sn_register_memory_event;
    end



    event require_specman_tick;
    event emit_specman_tick;
    always @(require_specman_tick) begin
        #0 ->emit_specman_tick ;
    end

    reg finish_test;
    always @(posedge finish_test) begin
        $finish;
    end

    //               Verilog time attributes
    parameter sn_declaration1_id = 658186681;
    parameter sn_declaration1_desc = "verilog time: ";



    //               Verilog code section               
    // ================================================================

    //         *** No Verilog code to reflect *** 


    //               Verilog variable section               
    // ================================================================

    //         *** No Verilog variable to reflect *** 


    //               Verilog subprogram section               
    // ================================================================

    //         *** No Verilog subprogram to reflect *** 


    //               Verilog ports section               
    // ================================================================

    //         *** No Verilog ports to reflect *** 


    //               Event ports (hdl_expression) section               
    // ================================================================

    //         *** No Event ports (hdl_expression) to reflect *** 


endmodule /* specman */





module specman_wave;



     /* Errors */

    parameter sn_error_num = 1;
    parameter sn_error_len = 80;
    reg [647:0] sn_err_str1;

     /* Output */

    parameter sn_message_num = 3;
    parameter sn_message_len = 80;
    reg [647:0] sn_msg_str1;
    reg [647:0] sn_msg_str2;
    reg [647:0] sn_msg_str3;

     /* Events */

    parameter sn_event_num = 100;
    reg  sn_emit_event1;
    event  sn_event1;
    always @sn_emit_event1 begin
        ->sn_event1;
    end
    reg  sn_emit_event2;
    event  sn_event2;
    always @sn_emit_event2 begin
        ->sn_event2;
    end
    reg  sn_emit_event3;
    event  sn_event3;
    always @sn_emit_event3 begin
        ->sn_event3;
    end
    reg  sn_emit_event4;
    event  sn_event4;
    always @sn_emit_event4 begin
        ->sn_event4;
    end
    reg  sn_emit_event5;
    event  sn_event5;
    always @sn_emit_event5 begin
        ->sn_event5;
    end
    reg  sn_emit_event6;
    event  sn_event6;
    always @sn_emit_event6 begin
        ->sn_event6;
    end
    reg  sn_emit_event7;
    event  sn_event7;
    always @sn_emit_event7 begin
        ->sn_event7;
    end
    reg  sn_emit_event8;
    event  sn_event8;
    always @sn_emit_event8 begin
        ->sn_event8;
    end
    reg  sn_emit_event9;
    event  sn_event9;
    always @sn_emit_event9 begin
        ->sn_event9;
    end
    reg  sn_emit_event10;
    event  sn_event10;
    always @sn_emit_event10 begin
        ->sn_event10;
    end
    reg  sn_emit_event11;
    event  sn_event11;
    always @sn_emit_event11 begin
        ->sn_event11;
    end
    reg  sn_emit_event12;
    event  sn_event12;
    always @sn_emit_event12 begin
        ->sn_event12;
    end
    reg  sn_emit_event13;
    event  sn_event13;
    always @sn_emit_event13 begin
        ->sn_event13;
    end
    reg  sn_emit_event14;
    event  sn_event14;
    always @sn_emit_event14 begin
        ->sn_event14;
    end
    reg  sn_emit_event15;
    event  sn_event15;
    always @sn_emit_event15 begin
        ->sn_event15;
    end
    reg  sn_emit_event16;
    event  sn_event16;
    always @sn_emit_event16 begin
        ->sn_event16;
    end
    reg  sn_emit_event17;
    event  sn_event17;
    always @sn_emit_event17 begin
        ->sn_event17;
    end
    reg  sn_emit_event18;
    event  sn_event18;
    always @sn_emit_event18 begin
        ->sn_event18;
    end
    reg  sn_emit_event19;
    event  sn_event19;
    always @sn_emit_event19 begin
        ->sn_event19;
    end
    reg  sn_emit_event20;
    event  sn_event20;
    always @sn_emit_event20 begin
        ->sn_event20;
    end
    reg  sn_emit_event21;
    event  sn_event21;
    always @sn_emit_event21 begin
        ->sn_event21;
    end
    reg  sn_emit_event22;
    event  sn_event22;
    always @sn_emit_event22 begin
        ->sn_event22;
    end
    reg  sn_emit_event23;
    event  sn_event23;
    always @sn_emit_event23 begin
        ->sn_event23;
    end
    reg  sn_emit_event24;
    event  sn_event24;
    always @sn_emit_event24 begin
        ->sn_event24;
    end
    reg  sn_emit_event25;
    event  sn_event25;
    always @sn_emit_event25 begin
        ->sn_event25;
    end
    reg  sn_emit_event26;
    event  sn_event26;
    always @sn_emit_event26 begin
        ->sn_event26;
    end
    reg  sn_emit_event27;
    event  sn_event27;
    always @sn_emit_event27 begin
        ->sn_event27;
    end
    reg  sn_emit_event28;
    event  sn_event28;
    always @sn_emit_event28 begin
        ->sn_event28;
    end
    reg  sn_emit_event29;
    event  sn_event29;
    always @sn_emit_event29 begin
        ->sn_event29;
    end
    reg  sn_emit_event30;
    event  sn_event30;
    always @sn_emit_event30 begin
        ->sn_event30;
    end
    reg  sn_emit_event31;
    event  sn_event31;
    always @sn_emit_event31 begin
        ->sn_event31;
    end
    reg  sn_emit_event32;
    event  sn_event32;
    always @sn_emit_event32 begin
        ->sn_event32;
    end
    reg  sn_emit_event33;
    event  sn_event33;
    always @sn_emit_event33 begin
        ->sn_event33;
    end
    reg  sn_emit_event34;
    event  sn_event34;
    always @sn_emit_event34 begin
        ->sn_event34;
    end
    reg  sn_emit_event35;
    event  sn_event35;
    always @sn_emit_event35 begin
        ->sn_event35;
    end
    reg  sn_emit_event36;
    event  sn_event36;
    always @sn_emit_event36 begin
        ->sn_event36;
    end
    reg  sn_emit_event37;
    event  sn_event37;
    always @sn_emit_event37 begin
        ->sn_event37;
    end
    reg  sn_emit_event38;
    event  sn_event38;
    always @sn_emit_event38 begin
        ->sn_event38;
    end
    reg  sn_emit_event39;
    event  sn_event39;
    always @sn_emit_event39 begin
        ->sn_event39;
    end
    reg  sn_emit_event40;
    event  sn_event40;
    always @sn_emit_event40 begin
        ->sn_event40;
    end
    reg  sn_emit_event41;
    event  sn_event41;
    always @sn_emit_event41 begin
        ->sn_event41;
    end
    reg  sn_emit_event42;
    event  sn_event42;
    always @sn_emit_event42 begin
        ->sn_event42;
    end
    reg  sn_emit_event43;
    event  sn_event43;
    always @sn_emit_event43 begin
        ->sn_event43;
    end
    reg  sn_emit_event44;
    event  sn_event44;
    always @sn_emit_event44 begin
        ->sn_event44;
    end
    reg  sn_emit_event45;
    event  sn_event45;
    always @sn_emit_event45 begin
        ->sn_event45;
    end
    reg  sn_emit_event46;
    event  sn_event46;
    always @sn_emit_event46 begin
        ->sn_event46;
    end
    reg  sn_emit_event47;
    event  sn_event47;
    always @sn_emit_event47 begin
        ->sn_event47;
    end
    reg  sn_emit_event48;
    event  sn_event48;
    always @sn_emit_event48 begin
        ->sn_event48;
    end
    reg  sn_emit_event49;
    event  sn_event49;
    always @sn_emit_event49 begin
        ->sn_event49;
    end
    reg  sn_emit_event50;
    event  sn_event50;
    always @sn_emit_event50 begin
        ->sn_event50;
    end
    reg  sn_emit_event51;
    event  sn_event51;
    always @sn_emit_event51 begin
        ->sn_event51;
    end
    reg  sn_emit_event52;
    event  sn_event52;
    always @sn_emit_event52 begin
        ->sn_event52;
    end
    reg  sn_emit_event53;
    event  sn_event53;
    always @sn_emit_event53 begin
        ->sn_event53;
    end
    reg  sn_emit_event54;
    event  sn_event54;
    always @sn_emit_event54 begin
        ->sn_event54;
    end
    reg  sn_emit_event55;
    event  sn_event55;
    always @sn_emit_event55 begin
        ->sn_event55;
    end
    reg  sn_emit_event56;
    event  sn_event56;
    always @sn_emit_event56 begin
        ->sn_event56;
    end
    reg  sn_emit_event57;
    event  sn_event57;
    always @sn_emit_event57 begin
        ->sn_event57;
    end
    reg  sn_emit_event58;
    event  sn_event58;
    always @sn_emit_event58 begin
        ->sn_event58;
    end
    reg  sn_emit_event59;
    event  sn_event59;
    always @sn_emit_event59 begin
        ->sn_event59;
    end
    reg  sn_emit_event60;
    event  sn_event60;
    always @sn_emit_event60 begin
        ->sn_event60;
    end
    reg  sn_emit_event61;
    event  sn_event61;
    always @sn_emit_event61 begin
        ->sn_event61;
    end
    reg  sn_emit_event62;
    event  sn_event62;
    always @sn_emit_event62 begin
        ->sn_event62;
    end
    reg  sn_emit_event63;
    event  sn_event63;
    always @sn_emit_event63 begin
        ->sn_event63;
    end
    reg  sn_emit_event64;
    event  sn_event64;
    always @sn_emit_event64 begin
        ->sn_event64;
    end
    reg  sn_emit_event65;
    event  sn_event65;
    always @sn_emit_event65 begin
        ->sn_event65;
    end
    reg  sn_emit_event66;
    event  sn_event66;
    always @sn_emit_event66 begin
        ->sn_event66;
    end
    reg  sn_emit_event67;
    event  sn_event67;
    always @sn_emit_event67 begin
        ->sn_event67;
    end
    reg  sn_emit_event68;
    event  sn_event68;
    always @sn_emit_event68 begin
        ->sn_event68;
    end
    reg  sn_emit_event69;
    event  sn_event69;
    always @sn_emit_event69 begin
        ->sn_event69;
    end
    reg  sn_emit_event70;
    event  sn_event70;
    always @sn_emit_event70 begin
        ->sn_event70;
    end
    reg  sn_emit_event71;
    event  sn_event71;
    always @sn_emit_event71 begin
        ->sn_event71;
    end
    reg  sn_emit_event72;
    event  sn_event72;
    always @sn_emit_event72 begin
        ->sn_event72;
    end
    reg  sn_emit_event73;
    event  sn_event73;
    always @sn_emit_event73 begin
        ->sn_event73;
    end
    reg  sn_emit_event74;
    event  sn_event74;
    always @sn_emit_event74 begin
        ->sn_event74;
    end
    reg  sn_emit_event75;
    event  sn_event75;
    always @sn_emit_event75 begin
        ->sn_event75;
    end
    reg  sn_emit_event76;
    event  sn_event76;
    always @sn_emit_event76 begin
        ->sn_event76;
    end
    reg  sn_emit_event77;
    event  sn_event77;
    always @sn_emit_event77 begin
        ->sn_event77;
    end
    reg  sn_emit_event78;
    event  sn_event78;
    always @sn_emit_event78 begin
        ->sn_event78;
    end
    reg  sn_emit_event79;
    event  sn_event79;
    always @sn_emit_event79 begin
        ->sn_event79;
    end
    reg  sn_emit_event80;
    event  sn_event80;
    always @sn_emit_event80 begin
        ->sn_event80;
    end
    reg  sn_emit_event81;
    event  sn_event81;
    always @sn_emit_event81 begin
        ->sn_event81;
    end
    reg  sn_emit_event82;
    event  sn_event82;
    always @sn_emit_event82 begin
        ->sn_event82;
    end
    reg  sn_emit_event83;
    event  sn_event83;
    always @sn_emit_event83 begin
        ->sn_event83;
    end
    reg  sn_emit_event84;
    event  sn_event84;
    always @sn_emit_event84 begin
        ->sn_event84;
    end
    reg  sn_emit_event85;
    event  sn_event85;
    always @sn_emit_event85 begin
        ->sn_event85;
    end
    reg  sn_emit_event86;
    event  sn_event86;
    always @sn_emit_event86 begin
        ->sn_event86;
    end
    reg  sn_emit_event87;
    event  sn_event87;
    always @sn_emit_event87 begin
        ->sn_event87;
    end
    reg  sn_emit_event88;
    event  sn_event88;
    always @sn_emit_event88 begin
        ->sn_event88;
    end
    reg  sn_emit_event89;
    event  sn_event89;
    always @sn_emit_event89 begin
        ->sn_event89;
    end
    reg  sn_emit_event90;
    event  sn_event90;
    always @sn_emit_event90 begin
        ->sn_event90;
    end
    reg  sn_emit_event91;
    event  sn_event91;
    always @sn_emit_event91 begin
        ->sn_event91;
    end
    reg  sn_emit_event92;
    event  sn_event92;
    always @sn_emit_event92 begin
        ->sn_event92;
    end
    reg  sn_emit_event93;
    event  sn_event93;
    always @sn_emit_event93 begin
        ->sn_event93;
    end
    reg  sn_emit_event94;
    event  sn_event94;
    always @sn_emit_event94 begin
        ->sn_event94;
    end
    reg  sn_emit_event95;
    event  sn_event95;
    always @sn_emit_event95 begin
        ->sn_event95;
    end
    reg  sn_emit_event96;
    event  sn_event96;
    always @sn_emit_event96 begin
        ->sn_event96;
    end
    reg  sn_emit_event97;
    event  sn_event97;
    always @sn_emit_event97 begin
        ->sn_event97;
    end
    reg  sn_emit_event98;
    event  sn_event98;
    always @sn_emit_event98 begin
        ->sn_event98;
    end
    reg  sn_emit_event99;
    event  sn_event99;
    always @sn_emit_event99 begin
        ->sn_event99;
    end
    reg  sn_emit_event100;
    event  sn_event100;
    always @sn_emit_event100 begin
        ->sn_event100;
    end

     /* Bits */

    parameter sn_boolean_num = 100;
    reg  sn_bool1;
    reg  sn_bool2;
    reg  sn_bool3;
    reg  sn_bool4;
    reg  sn_bool5;
    reg  sn_bool6;
    reg  sn_bool7;
    reg  sn_bool8;
    reg  sn_bool9;
    reg  sn_bool10;
    reg  sn_bool11;
    reg  sn_bool12;
    reg  sn_bool13;
    reg  sn_bool14;
    reg  sn_bool15;
    reg  sn_bool16;
    reg  sn_bool17;
    reg  sn_bool18;
    reg  sn_bool19;
    reg  sn_bool20;
    reg  sn_bool21;
    reg  sn_bool22;
    reg  sn_bool23;
    reg  sn_bool24;
    reg  sn_bool25;
    reg  sn_bool26;
    reg  sn_bool27;
    reg  sn_bool28;
    reg  sn_bool29;
    reg  sn_bool30;
    reg  sn_bool31;
    reg  sn_bool32;
    reg  sn_bool33;
    reg  sn_bool34;
    reg  sn_bool35;
    reg  sn_bool36;
    reg  sn_bool37;
    reg  sn_bool38;
    reg  sn_bool39;
    reg  sn_bool40;
    reg  sn_bool41;
    reg  sn_bool42;
    reg  sn_bool43;
    reg  sn_bool44;
    reg  sn_bool45;
    reg  sn_bool46;
    reg  sn_bool47;
    reg  sn_bool48;
    reg  sn_bool49;
    reg  sn_bool50;
    reg  sn_bool51;
    reg  sn_bool52;
    reg  sn_bool53;
    reg  sn_bool54;
    reg  sn_bool55;
    reg  sn_bool56;
    reg  sn_bool57;
    reg  sn_bool58;
    reg  sn_bool59;
    reg  sn_bool60;
    reg  sn_bool61;
    reg  sn_bool62;
    reg  sn_bool63;
    reg  sn_bool64;
    reg  sn_bool65;
    reg  sn_bool66;
    reg  sn_bool67;
    reg  sn_bool68;
    reg  sn_bool69;
    reg  sn_bool70;
    reg  sn_bool71;
    reg  sn_bool72;
    reg  sn_bool73;
    reg  sn_bool74;
    reg  sn_bool75;
    reg  sn_bool76;
    reg  sn_bool77;
    reg  sn_bool78;
    reg  sn_bool79;
    reg  sn_bool80;
    reg  sn_bool81;
    reg  sn_bool82;
    reg  sn_bool83;
    reg  sn_bool84;
    reg  sn_bool85;
    reg  sn_bool86;
    reg  sn_bool87;
    reg  sn_bool88;
    reg  sn_bool89;
    reg  sn_bool90;
    reg  sn_bool91;
    reg  sn_bool92;
    reg  sn_bool93;
    reg  sn_bool94;
    reg  sn_bool95;
    reg  sn_bool96;
    reg  sn_bool97;
    reg  sn_bool98;
    reg  sn_bool99;
    reg  sn_bool100;

     /* scalars */

    parameter sn_integer_num = 100;
    reg [31:0] sn_intg1;
    reg [31:0] sn_intg2;
    reg [31:0] sn_intg3;
    reg [31:0] sn_intg4;
    reg [31:0] sn_intg5;
    reg [31:0] sn_intg6;
    reg [31:0] sn_intg7;
    reg [31:0] sn_intg8;
    reg [31:0] sn_intg9;
    reg [31:0] sn_intg10;
    reg [31:0] sn_intg11;
    reg [31:0] sn_intg12;
    reg [31:0] sn_intg13;
    reg [31:0] sn_intg14;
    reg [31:0] sn_intg15;
    reg [31:0] sn_intg16;
    reg [31:0] sn_intg17;
    reg [31:0] sn_intg18;
    reg [31:0] sn_intg19;
    reg [31:0] sn_intg20;
    reg [31:0] sn_intg21;
    reg [31:0] sn_intg22;
    reg [31:0] sn_intg23;
    reg [31:0] sn_intg24;
    reg [31:0] sn_intg25;
    reg [31:0] sn_intg26;
    reg [31:0] sn_intg27;
    reg [31:0] sn_intg28;
    reg [31:0] sn_intg29;
    reg [31:0] sn_intg30;
    reg [31:0] sn_intg31;
    reg [31:0] sn_intg32;
    reg [31:0] sn_intg33;
    reg [31:0] sn_intg34;
    reg [31:0] sn_intg35;
    reg [31:0] sn_intg36;
    reg [31:0] sn_intg37;
    reg [31:0] sn_intg38;
    reg [31:0] sn_intg39;
    reg [31:0] sn_intg40;
    reg [31:0] sn_intg41;
    reg [31:0] sn_intg42;
    reg [31:0] sn_intg43;
    reg [31:0] sn_intg44;
    reg [31:0] sn_intg45;
    reg [31:0] sn_intg46;
    reg [31:0] sn_intg47;
    reg [31:0] sn_intg48;
    reg [31:0] sn_intg49;
    reg [31:0] sn_intg50;
    reg [31:0] sn_intg51;
    reg [31:0] sn_intg52;
    reg [31:0] sn_intg53;
    reg [31:0] sn_intg54;
    reg [31:0] sn_intg55;
    reg [31:0] sn_intg56;
    reg [31:0] sn_intg57;
    reg [31:0] sn_intg58;
    reg [31:0] sn_intg59;
    reg [31:0] sn_intg60;
    reg [31:0] sn_intg61;
    reg [31:0] sn_intg62;
    reg [31:0] sn_intg63;
    reg [31:0] sn_intg64;
    reg [31:0] sn_intg65;
    reg [31:0] sn_intg66;
    reg [31:0] sn_intg67;
    reg [31:0] sn_intg68;
    reg [31:0] sn_intg69;
    reg [31:0] sn_intg70;
    reg [31:0] sn_intg71;
    reg [31:0] sn_intg72;
    reg [31:0] sn_intg73;
    reg [31:0] sn_intg74;
    reg [31:0] sn_intg75;
    reg [31:0] sn_intg76;
    reg [31:0] sn_intg77;
    reg [31:0] sn_intg78;
    reg [31:0] sn_intg79;
    reg [31:0] sn_intg80;
    reg [31:0] sn_intg81;
    reg [31:0] sn_intg82;
    reg [31:0] sn_intg83;
    reg [31:0] sn_intg84;
    reg [31:0] sn_intg85;
    reg [31:0] sn_intg86;
    reg [31:0] sn_intg87;
    reg [31:0] sn_intg88;
    reg [31:0] sn_intg89;
    reg [31:0] sn_intg90;
    reg [31:0] sn_intg91;
    reg [31:0] sn_intg92;
    reg [31:0] sn_intg93;
    reg [31:0] sn_intg94;
    reg [31:0] sn_intg95;
    reg [31:0] sn_intg96;
    reg [31:0] sn_intg97;
    reg [31:0] sn_intg98;
    reg [31:0] sn_intg99;
    reg [31:0] sn_intg100;

     /* Strings */

    parameter sn_string_num = 200;
    parameter sn_string_len = 80;
    reg [647:0] sn_str1;
    reg [647:0] sn_str2;
    reg [647:0] sn_str3;
    reg [647:0] sn_str4;
    reg [647:0] sn_str5;
    reg [647:0] sn_str6;
    reg [647:0] sn_str7;
    reg [647:0] sn_str8;
    reg [647:0] sn_str9;
    reg [647:0] sn_str10;
    reg [647:0] sn_str11;
    reg [647:0] sn_str12;
    reg [647:0] sn_str13;
    reg [647:0] sn_str14;
    reg [647:0] sn_str15;
    reg [647:0] sn_str16;
    reg [647:0] sn_str17;
    reg [647:0] sn_str18;
    reg [647:0] sn_str19;
    reg [647:0] sn_str20;
    reg [647:0] sn_str21;
    reg [647:0] sn_str22;
    reg [647:0] sn_str23;
    reg [647:0] sn_str24;
    reg [647:0] sn_str25;
    reg [647:0] sn_str26;
    reg [647:0] sn_str27;
    reg [647:0] sn_str28;
    reg [647:0] sn_str29;
    reg [647:0] sn_str30;
    reg [647:0] sn_str31;
    reg [647:0] sn_str32;
    reg [647:0] sn_str33;
    reg [647:0] sn_str34;
    reg [647:0] sn_str35;
    reg [647:0] sn_str36;
    reg [647:0] sn_str37;
    reg [647:0] sn_str38;
    reg [647:0] sn_str39;
    reg [647:0] sn_str40;
    reg [647:0] sn_str41;
    reg [647:0] sn_str42;
    reg [647:0] sn_str43;
    reg [647:0] sn_str44;
    reg [647:0] sn_str45;
    reg [647:0] sn_str46;
    reg [647:0] sn_str47;
    reg [647:0] sn_str48;
    reg [647:0] sn_str49;
    reg [647:0] sn_str50;
    reg [647:0] sn_str51;
    reg [647:0] sn_str52;
    reg [647:0] sn_str53;
    reg [647:0] sn_str54;
    reg [647:0] sn_str55;
    reg [647:0] sn_str56;
    reg [647:0] sn_str57;
    reg [647:0] sn_str58;
    reg [647:0] sn_str59;
    reg [647:0] sn_str60;
    reg [647:0] sn_str61;
    reg [647:0] sn_str62;
    reg [647:0] sn_str63;
    reg [647:0] sn_str64;
    reg [647:0] sn_str65;
    reg [647:0] sn_str66;
    reg [647:0] sn_str67;
    reg [647:0] sn_str68;
    reg [647:0] sn_str69;
    reg [647:0] sn_str70;
    reg [647:0] sn_str71;
    reg [647:0] sn_str72;
    reg [647:0] sn_str73;
    reg [647:0] sn_str74;
    reg [647:0] sn_str75;
    reg [647:0] sn_str76;
    reg [647:0] sn_str77;
    reg [647:0] sn_str78;
    reg [647:0] sn_str79;
    reg [647:0] sn_str80;
    reg [647:0] sn_str81;
    reg [647:0] sn_str82;
    reg [647:0] sn_str83;
    reg [647:0] sn_str84;
    reg [647:0] sn_str85;
    reg [647:0] sn_str86;
    reg [647:0] sn_str87;
    reg [647:0] sn_str88;
    reg [647:0] sn_str89;
    reg [647:0] sn_str90;
    reg [647:0] sn_str91;
    reg [647:0] sn_str92;
    reg [647:0] sn_str93;
    reg [647:0] sn_str94;
    reg [647:0] sn_str95;
    reg [647:0] sn_str96;
    reg [647:0] sn_str97;
    reg [647:0] sn_str98;
    reg [647:0] sn_str99;
    reg [647:0] sn_str100;
    reg [647:0] sn_str101;
    reg [647:0] sn_str102;
    reg [647:0] sn_str103;
    reg [647:0] sn_str104;
    reg [647:0] sn_str105;
    reg [647:0] sn_str106;
    reg [647:0] sn_str107;
    reg [647:0] sn_str108;
    reg [647:0] sn_str109;
    reg [647:0] sn_str110;
    reg [647:0] sn_str111;
    reg [647:0] sn_str112;
    reg [647:0] sn_str113;
    reg [647:0] sn_str114;
    reg [647:0] sn_str115;
    reg [647:0] sn_str116;
    reg [647:0] sn_str117;
    reg [647:0] sn_str118;
    reg [647:0] sn_str119;
    reg [647:0] sn_str120;
    reg [647:0] sn_str121;
    reg [647:0] sn_str122;
    reg [647:0] sn_str123;
    reg [647:0] sn_str124;
    reg [647:0] sn_str125;
    reg [647:0] sn_str126;
    reg [647:0] sn_str127;
    reg [647:0] sn_str128;
    reg [647:0] sn_str129;
    reg [647:0] sn_str130;
    reg [647:0] sn_str131;
    reg [647:0] sn_str132;
    reg [647:0] sn_str133;
    reg [647:0] sn_str134;
    reg [647:0] sn_str135;
    reg [647:0] sn_str136;
    reg [647:0] sn_str137;
    reg [647:0] sn_str138;
    reg [647:0] sn_str139;
    reg [647:0] sn_str140;
    reg [647:0] sn_str141;
    reg [647:0] sn_str142;
    reg [647:0] sn_str143;
    reg [647:0] sn_str144;
    reg [647:0] sn_str145;
    reg [647:0] sn_str146;
    reg [647:0] sn_str147;
    reg [647:0] sn_str148;
    reg [647:0] sn_str149;
    reg [647:0] sn_str150;
    reg [647:0] sn_str151;
    reg [647:0] sn_str152;
    reg [647:0] sn_str153;
    reg [647:0] sn_str154;
    reg [647:0] sn_str155;
    reg [647:0] sn_str156;
    reg [647:0] sn_str157;
    reg [647:0] sn_str158;
    reg [647:0] sn_str159;
    reg [647:0] sn_str160;
    reg [647:0] sn_str161;
    reg [647:0] sn_str162;
    reg [647:0] sn_str163;
    reg [647:0] sn_str164;
    reg [647:0] sn_str165;
    reg [647:0] sn_str166;
    reg [647:0] sn_str167;
    reg [647:0] sn_str168;
    reg [647:0] sn_str169;
    reg [647:0] sn_str170;
    reg [647:0] sn_str171;
    reg [647:0] sn_str172;
    reg [647:0] sn_str173;
    reg [647:0] sn_str174;
    reg [647:0] sn_str175;
    reg [647:0] sn_str176;
    reg [647:0] sn_str177;
    reg [647:0] sn_str178;
    reg [647:0] sn_str179;
    reg [647:0] sn_str180;
    reg [647:0] sn_str181;
    reg [647:0] sn_str182;
    reg [647:0] sn_str183;
    reg [647:0] sn_str184;
    reg [647:0] sn_str185;
    reg [647:0] sn_str186;
    reg [647:0] sn_str187;
    reg [647:0] sn_str188;
    reg [647:0] sn_str189;
    reg [647:0] sn_str190;
    reg [647:0] sn_str191;
    reg [647:0] sn_str192;
    reg [647:0] sn_str193;
    reg [647:0] sn_str194;
    reg [647:0] sn_str195;
    reg [647:0] sn_str196;
    reg [647:0] sn_str197;
    reg [647:0] sn_str198;
    reg [647:0] sn_str199;
    reg [647:0] sn_str200;

    initial begin

       sn_str1=1'bz;
       sn_str2=1'bz;
       sn_str3=1'bz;
       sn_str4=1'bz;
       sn_str5=1'bz;
       sn_str6=1'bz;
       sn_str7=1'bz;
       sn_str8=1'bz;
       sn_str9=1'bz;
       sn_str10=1'bz;
       sn_str11=1'bz;
       sn_str12=1'bz;
       sn_str13=1'bz;
       sn_str14=1'bz;
       sn_str15=1'bz;
       sn_str16=1'bz;
       sn_str17=1'bz;
       sn_str18=1'bz;
       sn_str19=1'bz;
       sn_str20=1'bz;
       sn_str21=1'bz;
       sn_str22=1'bz;
       sn_str23=1'bz;
       sn_str24=1'bz;
       sn_str25=1'bz;
       sn_str26=1'bz;
       sn_str27=1'bz;
       sn_str28=1'bz;
       sn_str29=1'bz;
       sn_str30=1'bz;
       sn_str31=1'bz;
       sn_str32=1'bz;
       sn_str33=1'bz;
       sn_str34=1'bz;
       sn_str35=1'bz;
       sn_str36=1'bz;
       sn_str37=1'bz;
       sn_str38=1'bz;
       sn_str39=1'bz;
       sn_str40=1'bz;
       sn_str41=1'bz;
       sn_str42=1'bz;
       sn_str43=1'bz;
       sn_str44=1'bz;
       sn_str45=1'bz;
       sn_str46=1'bz;
       sn_str47=1'bz;
       sn_str48=1'bz;
       sn_str49=1'bz;
       sn_str50=1'bz;
       sn_str51=1'bz;
       sn_str52=1'bz;
       sn_str53=1'bz;
       sn_str54=1'bz;
       sn_str55=1'bz;
       sn_str56=1'bz;
       sn_str57=1'bz;
       sn_str58=1'bz;
       sn_str59=1'bz;
       sn_str60=1'bz;
       sn_str61=1'bz;
       sn_str62=1'bz;
       sn_str63=1'bz;
       sn_str64=1'bz;
       sn_str65=1'bz;
       sn_str66=1'bz;
       sn_str67=1'bz;
       sn_str68=1'bz;
       sn_str69=1'bz;
       sn_str70=1'bz;
       sn_str71=1'bz;
       sn_str72=1'bz;
       sn_str73=1'bz;
       sn_str74=1'bz;
       sn_str75=1'bz;
       sn_str76=1'bz;
       sn_str77=1'bz;
       sn_str78=1'bz;
       sn_str79=1'bz;
       sn_str80=1'bz;
       sn_str81=1'bz;
       sn_str82=1'bz;
       sn_str83=1'bz;
       sn_str84=1'bz;
       sn_str85=1'bz;
       sn_str86=1'bz;
       sn_str87=1'bz;
       sn_str88=1'bz;
       sn_str89=1'bz;
       sn_str90=1'bz;
       sn_str91=1'bz;
       sn_str92=1'bz;
       sn_str93=1'bz;
       sn_str94=1'bz;
       sn_str95=1'bz;
       sn_str96=1'bz;
       sn_str97=1'bz;
       sn_str98=1'bz;
       sn_str99=1'bz;
       sn_str100=1'bz;
       sn_str101=1'bz;
       sn_str102=1'bz;
       sn_str103=1'bz;
       sn_str104=1'bz;
       sn_str105=1'bz;
       sn_str106=1'bz;
       sn_str107=1'bz;
       sn_str108=1'bz;
       sn_str109=1'bz;
       sn_str110=1'bz;
       sn_str111=1'bz;
       sn_str112=1'bz;
       sn_str113=1'bz;
       sn_str114=1'bz;
       sn_str115=1'bz;
       sn_str116=1'bz;
       sn_str117=1'bz;
       sn_str118=1'bz;
       sn_str119=1'bz;
       sn_str120=1'bz;
       sn_str121=1'bz;
       sn_str122=1'bz;
       sn_str123=1'bz;
       sn_str124=1'bz;
       sn_str125=1'bz;
       sn_str126=1'bz;
       sn_str127=1'bz;
       sn_str128=1'bz;
       sn_str129=1'bz;
       sn_str130=1'bz;
       sn_str131=1'bz;
       sn_str132=1'bz;
       sn_str133=1'bz;
       sn_str134=1'bz;
       sn_str135=1'bz;
       sn_str136=1'bz;
       sn_str137=1'bz;
       sn_str138=1'bz;
       sn_str139=1'bz;
       sn_str140=1'bz;
       sn_str141=1'bz;
       sn_str142=1'bz;
       sn_str143=1'bz;
       sn_str144=1'bz;
       sn_str145=1'bz;
       sn_str146=1'bz;
       sn_str147=1'bz;
       sn_str148=1'bz;
       sn_str149=1'bz;
       sn_str150=1'bz;
       sn_str151=1'bz;
       sn_str152=1'bz;
       sn_str153=1'bz;
       sn_str154=1'bz;
       sn_str155=1'bz;
       sn_str156=1'bz;
       sn_str157=1'bz;
       sn_str158=1'bz;
       sn_str159=1'bz;
       sn_str160=1'bz;
       sn_str161=1'bz;
       sn_str162=1'bz;
       sn_str163=1'bz;
       sn_str164=1'bz;
       sn_str165=1'bz;
       sn_str166=1'bz;
       sn_str167=1'bz;
       sn_str168=1'bz;
       sn_str169=1'bz;
       sn_str170=1'bz;
       sn_str171=1'bz;
       sn_str172=1'bz;
       sn_str173=1'bz;
       sn_str174=1'bz;
       sn_str175=1'bz;
       sn_str176=1'bz;
       sn_str177=1'bz;
       sn_str178=1'bz;
       sn_str179=1'bz;
       sn_str180=1'bz;
       sn_str181=1'bz;
       sn_str182=1'bz;
       sn_str183=1'bz;
       sn_str184=1'bz;
       sn_str185=1'bz;
       sn_str186=1'bz;
       sn_str187=1'bz;
       sn_str188=1'bz;
       sn_str189=1'bz;
       sn_str190=1'bz;
       sn_str191=1'bz;
       sn_str192=1'bz;
       sn_str193=1'bz;
       sn_str194=1'bz;
       sn_str195=1'bz;
       sn_str196=1'bz;
       sn_str197=1'bz;
       sn_str198=1'bz;
       sn_str199=1'bz;
       sn_str200=1'bz;
    end

endmodule /* specman_wave */
