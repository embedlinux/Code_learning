library verilog;
use verilog.vl_types.all;
entity key_model is
    port(
        key             : out    vl_logic
    );
end key_model;
