library verilog;
use verilog.vl_types.all;
entity dut_interface is
    port(
        clk             : in     vl_logic
    );
end dut_interface;
