library verilog;
use verilog.vl_types.all;
entity pwm_generator_tb is
end pwm_generator_tb;
