library verilog;
use verilog.vl_types.all;
entity Hello_tb is
end Hello_tb;
