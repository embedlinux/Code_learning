
module FullDup ( OutParDataA, OutParDataB, InParDataA, InParDataB, InParValidA, 
        InParValidB, ClockA, ClockB, Reset );
  output [31:0] OutParDataA;
  output [31:0] OutParDataB;
  input [31:0] InParDataA;
  input [31:0] InParDataB;
  input InParValidA, InParValidB, ClockA, ClockB, Reset;
  wire   \*Logic1* , SerLine1, SerLine2, n1, n2, n3, n4, n5;

  SerDes_DWid32_RxLogDepth4_TxLogDepth3 SerDes_U1 ( .ParOutRxClk(OutParDataB), 
        .SerLineXfer(SerLine1), .ParDataIn(InParDataA), .InParClk(n3), 
        .InParValid(InParValidA), .OutParClk(n2), .RxRequest(\*Logic1* ), 
        .TxRequest(InParValidA), .Reset(n4) );
  SerDes_DWid32_RxLogDepth3_TxLogDepth4 SerDes_U2 ( .ParOutRxClk(OutParDataA), 
        .SerLineXfer(SerLine2), .ParDataIn(InParDataB), .InParClk(n2), 
        .InParValid(InParValidB), .OutParClk(n3), .RxRequest(\*Logic1* ), 
        .TxRequest(InParValidB), .Reset(n4) );
  INVD1 U2 ( .I(n5), .ZN(n4) );
  INVD1 U3 ( .I(n1), .ZN(n5) );
  BUFFD1 U4 ( .I(Reset), .Z(n1) );
  BUFFD1 U5 ( .I(ClockB), .Z(n2) );
  BUFFD1 U6 ( .I(ClockA), .Z(n3) );
  TIEH U7 ( .Z(\*Logic1* ) );
endmodule


module SerDes_DWid32_RxLogDepth4_TxLogDepth3 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4;

  Serializer_DWid32_AWid3 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n4), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid4_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n3), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD2 U1 ( .I(OutParClk), .Z(n3) );
  INVD1 U2 ( .I(n2), .ZN(n1) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  BUFFD1 U4 ( .I(InParClk), .Z(n4) );
endmodule


module SerDes_DWid32_RxLogDepth3_TxLogDepth4 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4;

  Serializer_DWid32_AWid4 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n3), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid3_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n4), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD2 U1 ( .I(OutParClk), .Z(n4) );
  INVD1 U2 ( .I(n2), .ZN(n1) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  BUFFD1 U4 ( .I(InParClk), .Z(n3) );
endmodule


module Serializer_DWid32_AWid3 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid3_DWid32_0 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(F_ReadReq), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n1) );
  SerEncoder_DWid32_0 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n1) );
  SerialTx_0 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n1) );
  INVD0 U1 ( .I(n3), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n3) );
  AN3D1 U3 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U4 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U5 ( .A1(n1), .A2(FIFOEmpty), .ZN(F_Valid) );
  INR2D1 U6 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
endmodule


module Deserializer_AWid4_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n4, n6,
         n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34,
         n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62,
         n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid4_DWid32_0 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n98)
         );
  DesDecoder_DWid32_0 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n98) );
  SerialRx_0 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n98) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n102), .Q(n104) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n101), .Q(n105) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n101), .Q(n106) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n101), .Q(n107) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n101), .Q(n108) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n101), .Q(n109) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n101), .Q(n110) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n101), .Q(n111) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n101), .Q(n112) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n101), .Q(n113) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n101), .Q(n114) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n101), .Q(n115) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n101), .Q(n116) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n101), .Q(n117) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n100), .Q(n118) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n100), .Q(n119) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n100), .Q(n120) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n100), .Q(n121) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n100), .Q(n122) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n100), .Q(n123) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n100), .Q(n124) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n100), .Q(n125) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n100), .Q(n126) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n100), .Q(n127) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n100), .Q(n128) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n100), .Q(n129) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n100), .Q(n130) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n99), .Q(n131) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n99), .Q(n132) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n99), .Q(n133) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n99), .Q(n134) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n99), .Q(n135) );
  DFCNQD1 ParValidr_reg ( .D(N35), .CP(ParOutClk), .CDN(n102), .Q(ParValid) );
  CKBD0 U3 ( .CLK(n97), .C(n1) );
  CKNXD16 U4 ( .I(n1), .ZN(ParOut[31]) );
  CKBD0 U5 ( .CLK(n96), .C(n4) );
  CKNXD16 U6 ( .I(n4), .ZN(ParOut[30]) );
  CKBD0 U7 ( .CLK(n95), .C(n6) );
  CKNXD16 U8 ( .I(n6), .ZN(ParOut[29]) );
  CKBD0 U9 ( .CLK(n94), .C(n8) );
  CKNXD16 U10 ( .I(n8), .ZN(ParOut[28]) );
  CKBD0 U11 ( .CLK(n93), .C(n10) );
  CKNXD16 U12 ( .I(n10), .ZN(ParOut[27]) );
  CKBD0 U13 ( .CLK(n92), .C(n12) );
  CKNXD16 U14 ( .I(n12), .ZN(ParOut[26]) );
  CKBD0 U15 ( .CLK(n91), .C(n14) );
  CKNXD16 U16 ( .I(n14), .ZN(ParOut[25]) );
  CKBD0 U17 ( .CLK(n90), .C(n16) );
  CKNXD16 U18 ( .I(n16), .ZN(ParOut[24]) );
  CKBD0 U19 ( .CLK(n89), .C(n18) );
  CKNXD16 U20 ( .I(n18), .ZN(ParOut[23]) );
  CKBD0 U21 ( .CLK(n88), .C(n20) );
  CKNXD16 U22 ( .I(n20), .ZN(ParOut[22]) );
  CKBD0 U23 ( .CLK(n87), .C(n22) );
  CKNXD16 U24 ( .I(n22), .ZN(ParOut[21]) );
  CKBD0 U25 ( .CLK(n86), .C(n24) );
  CKNXD16 U26 ( .I(n24), .ZN(ParOut[20]) );
  CKBD0 U27 ( .CLK(n85), .C(n26) );
  CKNXD16 U28 ( .I(n26), .ZN(ParOut[19]) );
  CKBD0 U29 ( .CLK(n84), .C(n28) );
  CKNXD16 U30 ( .I(n28), .ZN(ParOut[18]) );
  CKBD0 U31 ( .CLK(n83), .C(n30) );
  CKNXD16 U32 ( .I(n30), .ZN(ParOut[17]) );
  CKBD0 U33 ( .CLK(n82), .C(n32) );
  CKNXD16 U34 ( .I(n32), .ZN(ParOut[16]) );
  CKBD0 U35 ( .CLK(n81), .C(n34) );
  CKNXD16 U36 ( .I(n34), .ZN(ParOut[15]) );
  CKBD0 U37 ( .CLK(n80), .C(n36) );
  CKNXD16 U38 ( .I(n36), .ZN(ParOut[14]) );
  CKBD0 U39 ( .CLK(n79), .C(n38) );
  CKNXD16 U40 ( .I(n38), .ZN(ParOut[13]) );
  CKBD0 U41 ( .CLK(n78), .C(n40) );
  CKNXD16 U42 ( .I(n40), .ZN(ParOut[12]) );
  CKBD0 U43 ( .CLK(n77), .C(n42) );
  CKNXD16 U44 ( .I(n42), .ZN(ParOut[11]) );
  CKBD0 U45 ( .CLK(n76), .C(n44) );
  CKNXD16 U46 ( .I(n44), .ZN(ParOut[10]) );
  CKBD0 U47 ( .CLK(n75), .C(n46) );
  CKNXD16 U48 ( .I(n46), .ZN(ParOut[9]) );
  CKBD0 U49 ( .CLK(n74), .C(n48) );
  CKNXD16 U50 ( .I(n48), .ZN(ParOut[8]) );
  CKBD0 U51 ( .CLK(n73), .C(n50) );
  CKNXD16 U52 ( .I(n50), .ZN(ParOut[7]) );
  CKBD0 U53 ( .CLK(n72), .C(n52) );
  CKNXD16 U54 ( .I(n52), .ZN(ParOut[6]) );
  CKBD0 U55 ( .CLK(n71), .C(n54) );
  CKNXD16 U56 ( .I(n54), .ZN(ParOut[5]) );
  CKBD0 U57 ( .CLK(n70), .C(n56) );
  CKNXD16 U58 ( .I(n56), .ZN(ParOut[4]) );
  CKBD0 U59 ( .CLK(n69), .C(n58) );
  CKNXD16 U60 ( .I(n58), .ZN(ParOut[3]) );
  CKBD0 U61 ( .CLK(n68), .C(n60) );
  CKNXD16 U62 ( .I(n60), .ZN(ParOut[2]) );
  CKBD0 U63 ( .CLK(n67), .C(n62) );
  CKNXD16 U64 ( .I(n62), .ZN(ParOut[1]) );
  CKBD0 U65 ( .CLK(n66), .C(n64) );
  CKNXD16 U66 ( .I(n64), .ZN(ParOut[0]) );
  INVD1 U67 ( .I(n99), .ZN(n98) );
  BUFFD1 U68 ( .I(n103), .Z(n99) );
  BUFFD1 U69 ( .I(n103), .Z(n100) );
  BUFFD1 U70 ( .I(n103), .Z(n101) );
  BUFFD1 U71 ( .I(n103), .Z(n102) );
  INVD1 U72 ( .I(Reset), .ZN(n103) );
  NR2D1 U73 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  INVD0 U74 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U75 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U76 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U77 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U78 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U79 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U80 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U81 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U82 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U83 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U84 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U85 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U86 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U87 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U88 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U89 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U90 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U91 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U92 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U93 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U94 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U95 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U96 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U97 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U98 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U99 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U100 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U101 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U102 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U103 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U104 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U105 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U106 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U107 ( .CLK(n135), .CN(n66) );
  CKND0 U108 ( .CLK(n134), .CN(n67) );
  CKND0 U109 ( .CLK(n133), .CN(n68) );
  CKND0 U110 ( .CLK(n132), .CN(n69) );
  CKND0 U111 ( .CLK(n131), .CN(n70) );
  CKND0 U112 ( .CLK(n130), .CN(n71) );
  CKND0 U113 ( .CLK(n129), .CN(n72) );
  CKND0 U114 ( .CLK(n128), .CN(n73) );
  CKND0 U115 ( .CLK(n127), .CN(n74) );
  CKND0 U116 ( .CLK(n126), .CN(n75) );
  CKND0 U117 ( .CLK(n125), .CN(n76) );
  CKND0 U118 ( .CLK(n124), .CN(n77) );
  CKND0 U119 ( .CLK(n123), .CN(n78) );
  CKND0 U120 ( .CLK(n122), .CN(n79) );
  CKND0 U121 ( .CLK(n121), .CN(n80) );
  CKND0 U122 ( .CLK(n120), .CN(n81) );
  CKND0 U123 ( .CLK(n119), .CN(n82) );
  CKND0 U124 ( .CLK(n118), .CN(n83) );
  CKND0 U125 ( .CLK(n117), .CN(n84) );
  CKND0 U126 ( .CLK(n116), .CN(n85) );
  CKND0 U127 ( .CLK(n115), .CN(n86) );
  CKND0 U128 ( .CLK(n114), .CN(n87) );
  CKND0 U129 ( .CLK(n113), .CN(n88) );
  CKND0 U130 ( .CLK(n112), .CN(n89) );
  CKND0 U131 ( .CLK(n111), .CN(n90) );
  CKND0 U132 ( .CLK(n110), .CN(n91) );
  CKND0 U133 ( .CLK(n109), .CN(n92) );
  CKND0 U134 ( .CLK(n108), .CN(n93) );
  CKND0 U135 ( .CLK(n107), .CN(n94) );
  CKND0 U136 ( .CLK(n106), .CN(n95) );
  CKND0 U137 ( .CLK(n105), .CN(n96) );
  CKND0 U138 ( .CLK(n104), .CN(n97) );
endmodule


module Serializer_DWid32_AWid4 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid4_DWid32_1 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(F_ReadReq), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n1) );
  SerEncoder_DWid32_1 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n1) );
  SerialTx_1 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n1) );
  INVD0 U1 ( .I(n3), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n3) );
  AN3D1 U3 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U4 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U5 ( .A1(n1), .A2(FIFOEmpty), .ZN(F_Valid) );
  INR2D1 U6 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
endmodule


module Deserializer_AWid3_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n4, n6,
         n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34,
         n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62,
         n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid3_DWid32_1 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n98)
         );
  DesDecoder_DWid32_1 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n98) );
  SerialRx_1 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n98) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n102), .Q(n104) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n101), .Q(n105) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n101), .Q(n106) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n101), .Q(n107) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n101), .Q(n108) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n101), .Q(n109) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n101), .Q(n110) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n101), .Q(n111) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n101), .Q(n112) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n101), .Q(n113) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n101), .Q(n114) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n101), .Q(n115) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n101), .Q(n116) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n101), .Q(n117) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n100), .Q(n118) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n100), .Q(n119) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n100), .Q(n120) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n100), .Q(n121) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n100), .Q(n122) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n100), .Q(n123) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n100), .Q(n124) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n100), .Q(n125) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n100), .Q(n126) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n100), .Q(n127) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n100), .Q(n128) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n100), .Q(n129) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n100), .Q(n130) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n99), .Q(n131) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n99), .Q(n132) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n99), .Q(n133) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n99), .Q(n134) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n99), .Q(n135) );
  DFCNQD1 ParValidr_reg ( .D(N35), .CP(ParOutClk), .CDN(n102), .Q(ParValid) );
  CKBD0 U3 ( .CLK(n97), .C(n1) );
  CKNXD16 U4 ( .I(n1), .ZN(ParOut[31]) );
  CKBD0 U5 ( .CLK(n96), .C(n4) );
  CKNXD16 U6 ( .I(n4), .ZN(ParOut[30]) );
  CKBD0 U7 ( .CLK(n95), .C(n6) );
  CKNXD16 U8 ( .I(n6), .ZN(ParOut[29]) );
  CKBD0 U9 ( .CLK(n94), .C(n8) );
  CKNXD16 U10 ( .I(n8), .ZN(ParOut[28]) );
  CKBD0 U11 ( .CLK(n93), .C(n10) );
  CKNXD16 U12 ( .I(n10), .ZN(ParOut[27]) );
  CKBD0 U13 ( .CLK(n92), .C(n12) );
  CKNXD16 U14 ( .I(n12), .ZN(ParOut[26]) );
  CKBD0 U15 ( .CLK(n91), .C(n14) );
  CKNXD16 U16 ( .I(n14), .ZN(ParOut[25]) );
  CKBD0 U17 ( .CLK(n90), .C(n16) );
  CKNXD16 U18 ( .I(n16), .ZN(ParOut[24]) );
  CKBD0 U19 ( .CLK(n89), .C(n18) );
  CKNXD16 U20 ( .I(n18), .ZN(ParOut[23]) );
  CKBD0 U21 ( .CLK(n88), .C(n20) );
  CKNXD16 U22 ( .I(n20), .ZN(ParOut[22]) );
  CKBD0 U23 ( .CLK(n87), .C(n22) );
  CKNXD16 U24 ( .I(n22), .ZN(ParOut[21]) );
  CKBD0 U25 ( .CLK(n86), .C(n24) );
  CKNXD16 U26 ( .I(n24), .ZN(ParOut[20]) );
  CKBD0 U27 ( .CLK(n85), .C(n26) );
  CKNXD16 U28 ( .I(n26), .ZN(ParOut[19]) );
  CKBD0 U29 ( .CLK(n84), .C(n28) );
  CKNXD16 U30 ( .I(n28), .ZN(ParOut[18]) );
  CKBD0 U31 ( .CLK(n83), .C(n30) );
  CKNXD16 U32 ( .I(n30), .ZN(ParOut[17]) );
  CKBD0 U33 ( .CLK(n82), .C(n32) );
  CKNXD16 U34 ( .I(n32), .ZN(ParOut[16]) );
  CKBD0 U35 ( .CLK(n81), .C(n34) );
  CKNXD16 U36 ( .I(n34), .ZN(ParOut[15]) );
  CKBD0 U37 ( .CLK(n80), .C(n36) );
  CKNXD16 U38 ( .I(n36), .ZN(ParOut[14]) );
  CKBD0 U39 ( .CLK(n79), .C(n38) );
  CKNXD16 U40 ( .I(n38), .ZN(ParOut[13]) );
  CKBD0 U41 ( .CLK(n78), .C(n40) );
  CKNXD16 U42 ( .I(n40), .ZN(ParOut[12]) );
  CKBD0 U43 ( .CLK(n77), .C(n42) );
  CKNXD16 U44 ( .I(n42), .ZN(ParOut[11]) );
  CKBD0 U45 ( .CLK(n76), .C(n44) );
  CKNXD16 U46 ( .I(n44), .ZN(ParOut[10]) );
  CKBD0 U47 ( .CLK(n75), .C(n46) );
  CKNXD16 U48 ( .I(n46), .ZN(ParOut[9]) );
  CKBD0 U49 ( .CLK(n74), .C(n48) );
  CKNXD16 U50 ( .I(n48), .ZN(ParOut[8]) );
  CKBD0 U51 ( .CLK(n73), .C(n50) );
  CKNXD16 U52 ( .I(n50), .ZN(ParOut[7]) );
  CKBD0 U53 ( .CLK(n72), .C(n52) );
  CKNXD16 U54 ( .I(n52), .ZN(ParOut[6]) );
  CKBD0 U55 ( .CLK(n71), .C(n54) );
  CKNXD16 U56 ( .I(n54), .ZN(ParOut[5]) );
  CKBD0 U57 ( .CLK(n70), .C(n56) );
  CKNXD16 U58 ( .I(n56), .ZN(ParOut[4]) );
  CKBD0 U59 ( .CLK(n69), .C(n58) );
  CKNXD16 U60 ( .I(n58), .ZN(ParOut[3]) );
  CKBD0 U61 ( .CLK(n68), .C(n60) );
  CKNXD16 U62 ( .I(n60), .ZN(ParOut[2]) );
  CKBD0 U63 ( .CLK(n67), .C(n62) );
  CKNXD16 U64 ( .I(n62), .ZN(ParOut[1]) );
  CKBD0 U65 ( .CLK(n66), .C(n64) );
  CKNXD16 U66 ( .I(n64), .ZN(ParOut[0]) );
  INVD1 U67 ( .I(n99), .ZN(n98) );
  BUFFD1 U68 ( .I(n103), .Z(n99) );
  BUFFD1 U69 ( .I(n103), .Z(n100) );
  BUFFD1 U70 ( .I(n103), .Z(n101) );
  BUFFD1 U71 ( .I(n103), .Z(n102) );
  INVD1 U72 ( .I(Reset), .ZN(n103) );
  NR2D1 U73 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  INVD0 U74 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U75 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U76 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U77 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U78 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U79 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U80 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U81 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U82 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U83 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U84 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U85 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U86 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U87 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U88 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U89 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U90 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U91 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U92 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U93 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U94 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U95 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U96 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U97 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U98 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U99 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U100 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U101 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U102 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U103 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U104 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U105 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U106 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U107 ( .CLK(n135), .CN(n66) );
  CKND0 U108 ( .CLK(n134), .CN(n67) );
  CKND0 U109 ( .CLK(n133), .CN(n68) );
  CKND0 U110 ( .CLK(n132), .CN(n69) );
  CKND0 U111 ( .CLK(n131), .CN(n70) );
  CKND0 U112 ( .CLK(n130), .CN(n71) );
  CKND0 U113 ( .CLK(n129), .CN(n72) );
  CKND0 U114 ( .CLK(n128), .CN(n73) );
  CKND0 U115 ( .CLK(n127), .CN(n74) );
  CKND0 U116 ( .CLK(n126), .CN(n75) );
  CKND0 U117 ( .CLK(n125), .CN(n76) );
  CKND0 U118 ( .CLK(n124), .CN(n77) );
  CKND0 U119 ( .CLK(n123), .CN(n78) );
  CKND0 U120 ( .CLK(n122), .CN(n79) );
  CKND0 U121 ( .CLK(n121), .CN(n80) );
  CKND0 U122 ( .CLK(n120), .CN(n81) );
  CKND0 U123 ( .CLK(n119), .CN(n82) );
  CKND0 U124 ( .CLK(n118), .CN(n83) );
  CKND0 U125 ( .CLK(n117), .CN(n84) );
  CKND0 U126 ( .CLK(n116), .CN(n85) );
  CKND0 U127 ( .CLK(n115), .CN(n86) );
  CKND0 U128 ( .CLK(n114), .CN(n87) );
  CKND0 U129 ( .CLK(n113), .CN(n88) );
  CKND0 U130 ( .CLK(n112), .CN(n89) );
  CKND0 U131 ( .CLK(n111), .CN(n90) );
  CKND0 U132 ( .CLK(n110), .CN(n91) );
  CKND0 U133 ( .CLK(n109), .CN(n92) );
  CKND0 U134 ( .CLK(n108), .CN(n93) );
  CKND0 U135 ( .CLK(n107), .CN(n94) );
  CKND0 U136 ( .CLK(n106), .CN(n95) );
  CKND0 U137 ( .CLK(n105), .CN(n96) );
  CKND0 U138 ( .CLK(n104), .CN(n97) );
endmodule


module FIFOTop_AWid3_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid3_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD0 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_0 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_0_DW01_dec_0 \ShifterBlock/sub_132  ( .A({\Sh_N[5] , N6, 
        N5, N4, N3, N2}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n17), .CP(n23), .CDN(n29), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n24), .CP(ParClk), .CDN(n27), .Q(HalfParClkr)
         );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(n23), .CDN(n27), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n23), .CDN(n27), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n23), .CDN(n28), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n22), .CDN(n29), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n22), .CDN(n27), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(n22), .CDN(n29), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(n22), .CDN(n28), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(n22), .CDN(n28), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(n21), .CDN(n28), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n21), .CDN(n28), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n21), .CDN(n28), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(n21), .CDN(n28), .Q(InBuf[9]) );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n23), .CDN(n29), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(n23), .CDN(n29), .Q(InBuf[5]) );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n23), .CDN(n29), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(n22), .CDN(n29), .Q(InBuf[1]) );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(n23), .CDN(n27), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n23), .CDN(n28), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(n23), .CDN(n27), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(n22), .CDN(n29), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(n22), .CDN(n28), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n22), .CDN(n27), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n22), .CDN(n29), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(n21), .CDN(n28), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(n21), .CDN(n28), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(n21), .CDN(n28), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(n21), .CDN(n28), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(n21), .CDN(n29), .Q(InBuf[8]) );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n21), .CDN(n29), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(n23), .CDN(n29), .Q(InBuf[4]) );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n22), .CDN(n29), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(n21), .CDN(n29), .Q(InBuf[0]) );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n27), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n27), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n27), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n27), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n27), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n27), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(N31), .CP(SerClk), .CDN(n28), .Q(SerOut) );
  INR2D1 U3 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
  CKBD0 U4 ( .CLK(Reset), .C(n25) );
  CKBXD0 U5 ( .I(Reset), .Z(n26) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(N4), .ZN(n1) );
  MUX2ND0 U7 ( .I0(n7), .I1(n8), .S(N4), .ZN(n2) );
  INVD0 U8 ( .I(n19), .ZN(n24) );
  MUX2ND0 U9 ( .I0(n9), .I1(n10), .S(N4), .ZN(n3) );
  MUX2ND0 U10 ( .I0(n5), .I1(n6), .S(N4), .ZN(n4) );
  INVD0 U11 ( .I(n20), .ZN(n19) );
  INVD0 U12 ( .I(HalfParClkr), .ZN(n20) );
  INVD1 U13 ( .I(n25), .ZN(n29) );
  INVD1 U14 ( .I(n26), .ZN(n28) );
  INVD1 U15 ( .I(n26), .ZN(n27) );
  INVD1 U16 ( .I(n24), .ZN(n21) );
  INVD1 U17 ( .I(n20), .ZN(n22) );
  INVD1 U18 ( .I(n20), .ZN(n23) );
  INVD1 U19 ( .I(n18), .ZN(n17) );
  INVD1 U20 ( .I(n31), .ZN(n30) );
  ND2D1 U21 ( .A1(N3), .A2(N2), .ZN(n32) );
  AN2D1 U22 ( .A1(N4), .A2(n30), .Z(N26) );
  MUX4ND0 U23 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n5) );
  MUX4ND0 U24 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n6) );
  MUX4ND0 U25 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n7) );
  MUX4ND0 U26 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n8) );
  MUX4ND0 U27 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n9) );
  MUX4ND0 U28 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n10) );
  MUX4ND0 U29 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n11) );
  MUX4ND0 U30 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n12) );
  NR2D1 U31 ( .A1(n32), .A2(N4), .ZN(N24) );
  INVD1 U32 ( .I(N85), .ZN(n18) );
  MUX2ND0 U33 ( .I0(n13), .I1(n14), .S(N6), .ZN(N29) );
  MUX2ND0 U34 ( .I0(n15), .I1(n16), .S(N6), .ZN(N27) );
  MUX2ND0 U35 ( .I0(n14), .I1(n13), .S(N6), .ZN(N25) );
  MUX2ND0 U36 ( .I0(n16), .I1(n15), .S(N6), .ZN(N23) );
  MUX2ND0 U37 ( .I0(n2), .I1(n3), .S(N5), .ZN(n14) );
  MUX2ND0 U38 ( .I0(n1), .I1(n4), .S(N5), .ZN(n13) );
  MUX2ND0 U39 ( .I0(n3), .I1(n1), .S(N5), .ZN(n16) );
  MUX2ND0 U40 ( .I0(n4), .I1(n2), .S(N5), .ZN(n15) );
  OR2D1 U41 ( .A1(N2), .A2(N3), .Z(n31) );
  MUX2ND0 U42 ( .I0(n32), .I1(n31), .S(N4), .ZN(N28) );
  AN2D0 U43 ( .A1(ParIn[31]), .A2(n17), .Z(N84) );
  AN2D0 U44 ( .A1(ParIn[30]), .A2(n17), .Z(N83) );
  AN2D0 U45 ( .A1(ParIn[29]), .A2(n17), .Z(N82) );
  AN2D0 U46 ( .A1(ParIn[28]), .A2(n17), .Z(N81) );
  AN2D0 U47 ( .A1(ParIn[27]), .A2(N85), .Z(N80) );
  AN2D0 U48 ( .A1(ParIn[26]), .A2(N85), .Z(N79) );
  AN2D0 U49 ( .A1(ParIn[25]), .A2(N85), .Z(N78) );
  AN2D0 U50 ( .A1(ParIn[24]), .A2(N85), .Z(N77) );
  AN2D0 U51 ( .A1(ParIn[23]), .A2(N85), .Z(N76) );
  AN2D0 U52 ( .A1(ParIn[22]), .A2(N85), .Z(N75) );
  AN2D0 U53 ( .A1(ParIn[21]), .A2(N85), .Z(N74) );
  AN2D0 U54 ( .A1(ParIn[20]), .A2(N85), .Z(N73) );
  AN2D0 U55 ( .A1(ParIn[19]), .A2(N85), .Z(N72) );
  AN2D0 U56 ( .A1(ParIn[18]), .A2(N85), .Z(N71) );
  AN2D0 U57 ( .A1(ParIn[17]), .A2(n17), .Z(N70) );
  AN2D0 U58 ( .A1(ParIn[16]), .A2(n17), .Z(N69) );
  AN2D0 U59 ( .A1(ParIn[15]), .A2(n17), .Z(N68) );
  AN2D0 U60 ( .A1(ParIn[14]), .A2(n17), .Z(N67) );
  AN2D0 U61 ( .A1(ParIn[13]), .A2(n17), .Z(N66) );
  AN2D0 U62 ( .A1(ParIn[12]), .A2(n17), .Z(N65) );
  AN2D0 U63 ( .A1(ParIn[11]), .A2(n17), .Z(N64) );
  AN2D0 U64 ( .A1(ParIn[10]), .A2(n17), .Z(N63) );
  AN2D0 U65 ( .A1(ParIn[9]), .A2(N85), .Z(N62) );
  AN2D0 U66 ( .A1(ParIn[8]), .A2(N85), .Z(N61) );
  AN2D0 U67 ( .A1(ParIn[7]), .A2(n17), .Z(N60) );
  AN2D0 U68 ( .A1(ParIn[6]), .A2(n17), .Z(N59) );
  AN2D0 U69 ( .A1(ParIn[5]), .A2(n17), .Z(N58) );
  AN2D0 U70 ( .A1(ParIn[4]), .A2(n17), .Z(N57) );
  AN2D0 U71 ( .A1(ParIn[3]), .A2(n17), .Z(N56) );
  AN2D0 U72 ( .A1(ParIn[2]), .A2(N85), .Z(N55) );
  AN2D0 U73 ( .A1(ParIn[1]), .A2(n17), .Z(N54) );
  AN2D0 U74 ( .A1(ParIn[0]), .A2(n17), .Z(N53) );
  IND2D0 U75 ( .A1(n33), .B1(n34), .ZN(N31) );
  OAI21D0 U76 ( .A1(N23), .A2(n35), .B(n36), .ZN(n34) );
  MUX2ND0 U77 ( .I0(n37), .I1(n38), .S(n35), .ZN(n36) );
  MUX3ND0 U78 ( .I0(N25), .I1(n39), .I2(N24), .S0(\Sh_N[5] ), .S1(n40), .ZN(
        n38) );
  NR2D0 U79 ( .A1(\Sh_N[5] ), .A2(N5), .ZN(n40) );
  MUX2D0 U80 ( .I0(n41), .I1(N26), .S(n42), .Z(n39) );
  NR2D0 U81 ( .A1(N6), .A2(N5), .ZN(n42) );
  INR2D0 U82 ( .A1(N27), .B1(N6), .ZN(n41) );
  CKND0 U83 ( .CLK(N5), .CN(n37) );
  CKND2D0 U84 ( .A1(n43), .A2(n44), .ZN(n35) );
  MUX2ND0 U85 ( .I0(n45), .I1(n46), .S(N5), .ZN(n33) );
  CKND2D0 U86 ( .A1(N29), .A2(n47), .ZN(n46) );
  CKND2D0 U87 ( .A1(N28), .A2(n47), .ZN(n45) );
  NR2D0 U88 ( .A1(n44), .A2(n43), .ZN(n47) );
  CKND0 U89 ( .CLK(N6), .CN(n43) );
  CKND0 U90 ( .CLK(\Sh_N[5] ), .CN(n44) );
  INR3D0 U91 ( .A1(N85), .B1(Reset), .B2(n24), .ZN(FIFO_ReadReq) );
endmodule


module SerialTx_0 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_0 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(n1), .ClkW(ClkW), .Reset(n3) );
  DPMem1kx32_AWid4_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(n1), .ClkW(ClkW), .ChipEna(
        \*Logic1* ), .Read(n2), .Write(SM_MemWriteCmd), .Reset(n3) );
  INVD0 U2 ( .I(n4), .ZN(n3) );
  BUFFD0 U3 ( .I(ClkR), .Z(n1) );
  INVD1 U4 ( .I(Reseter), .ZN(n4) );
  BUFFD1 U5 ( .I(SM_MemReadCmd), .Z(n2) );
  TIEH U6 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_0 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n230, n231, n232, n1, n4, n5, n30, n31, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9027, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U39 ( .A1(n9127), .A2(n54), .B1(n9129), .B2(Decoder[9]), .ZN(n123)
         );
  MOAI22D1 U40 ( .A1(n9127), .A2(n55), .B1(n9129), .B2(Decoder[8]), .ZN(n124)
         );
  OR3D1 U92 ( .A1(n8960), .A2(n8963), .A3(n8972), .Z(n22) );
  OR3D1 U94 ( .A1(n8962), .A2(n8966), .A3(n8974), .Z(n23) );
  OR3D1 U96 ( .A1(n8964), .A2(n8970), .A3(n8973), .Z(n24) );
  OA21D1 U99 ( .A1(n26), .A2(n27), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n28) );
  DesDecoder_DWid32_0_DW01_inc_0 \ClkGen/add_206  ( .A({Count32[4:2], n6895, 
        n6903}), .SUM({N34, N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(n4), .CPN(n9135), .CDN(n9149), .Q(FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(n30), .CPN(n9132), .CDN(n9148), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(n227), .CPN(n9130), .CDN(n9148), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(n327), .CPN(n9130), .CDN(n9149), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(n423), .CPN(SerClock), .CDN(n9149), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(n520), .CPN(n9136), .CDN(n9151), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(n616), .CPN(n9134), .CDN(n9148), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(n713), .CPN(n9136), .CDN(n9149), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(n715), .CPN(n9134), .CDN(n9149), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(n812), .CPN(n9135), .CDN(n9152), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(n909), .CPN(n9145), .CDN(n9147), .Q(FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(n912), .CPN(n9145), .CDN(n9147), .Q(FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(n914), .CPN(n9145), .CDN(n9154), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(n916), .CPN(n9145), .CDN(n9152), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(n918), .CPN(n9145), .CDN(n9149), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(n920), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(n922), .CPN(n9145), .CDN(n9150), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(n924), .CPN(n9136), .CDN(n9151), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(n926), .CPN(n9131), .CDN(n9153), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(n1022), .CPN(n9131), .CDN(n9148), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(n1119), .CPN(n9135), .CDN(n9148), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(n1121), .CPN(n9133), .CDN(n9148), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(n1123), .CPN(SerClock), .CDN(n9148), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(n1125), .CPN(n9135), .CDN(n9148), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(n1127), .CPN(n9133), .CDN(n9148), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(n1129), .CPN(n9132), .CDN(n9149), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(n1131), .CPN(n9134), .CDN(n9149), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(n1133), .CPN(n9131), .CDN(n9150), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(n1230), .CPN(n9130), .CDN(n9150), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(n1232), .CPN(n9136), .CDN(n9150), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(n1234), .CPN(n9130), .CDN(n9150), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(n1236), .CPN(n9134), .CDN(n9150), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(n1238), .CPN(n9136), .CDN(n9150), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(n1240), .CPN(SerClock), .CDN(n9150), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(n1242), .CPN(n9136), .CDN(n9150), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(n1244), .CPN(n9134), .CDN(n9151), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(n1341), .CPN(n9146), .CDN(n9153), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(n1343), .CPN(n9132), .CDN(n9151), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(n1345), .CPN(n9136), .CDN(n9152), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(n1347), .CPN(SerClock), .CDN(n9147), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(n1349), .CPN(n9130), .CDN(n9152), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(n1351), .CPN(n9131), .CDN(n9154), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[0]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(n1353), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(n1355), .CPN(n9130), .CDN(n9148), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(n1451), .CPN(n9130), .CDN(n9149), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(n1547), .CPN(n9135), .CDN(n9150), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(n1643), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(n1646), .CPN(n9145), .CDN(n9147), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(n1650), .CPN(n9131), .CDN(n9152), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(n1746), .CPN(n9132), .CDN(n9149), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(n1843), .CPN(n9133), .CDN(n9150), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(n1845), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(n1848), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(n1851), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(n1854), .CPN(n9145), .CDN(n9147), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(n1858), .CPN(n9132), .CDN(n9148), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(n1954), .CPN(n9133), .CDN(n9149), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(n2050), .CPN(SerClock), .CDN(n9154), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(n2146), .CPN(n9135), .CDN(n9153), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(n2242), .CPN(n9131), .CDN(n9149), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(n2338), .CPN(SerClock), .CDN(n9152), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(n2434), .CPN(n9133), .CDN(n9154), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(n2530), .CPN(n9134), .CDN(n9147), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(n2532), .E(SerValid), .CP(n9137), .CDN(n9153), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n2533), .CPN(n9134), .CDN(n9153), .Q(
        Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n2667), .CPN(n9146), .CDN(n9151), .Q(
        Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n2803), .CPN(n9133), .CDN(n9152), .Q(
        Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n2939), .CPN(n9132), .CDN(n9150), .Q(
        Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n3075), .CPN(n9146), .CDN(n9151), .Q(
        Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n3211), .CPN(n9144), .CDN(n9151), .Q(
        Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n3347), .CPN(n9144), .CDN(n9150), .Q(
        Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n3483), .CPN(n9144), .CDN(n9149), .Q(
        Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n3619), .CPN(n9144), .CDN(n9147), .Q(
        Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n3755), .CPN(n9144), .CDN(n9154), .Q(
        Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n3891), .CPN(n9144), .CDN(n9153), .Q(
        Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n4027), .CPN(n9144), .CDN(n9151), .Q(
        Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n4163), .CPN(n9144), .CDN(n9152), .Q(
        Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n4299), .CPN(n9144), .CDN(n9150), .Q(
        Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n4435), .CPN(n9143), .CDN(n9153), .Q(
        Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n4571), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n4707), .CPN(n9143), .CDN(n9152), .Q(
        Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n4843), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n4979), .CPN(n9143), .CDN(n9148), .Q(
        Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n5115), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n5251), .CPN(n9143), .CDN(n9147), .Q(
        Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n5387), .CPN(n9143), .CDN(n9151), .Q(
        Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n5524), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[9]) );
  DFNCND1 \Decoder_reg[8]  ( .D(n5661), .CPN(n9142), .CDN(n9153), .Q(
        Decoder[8]) );
  DFNCND1 \Decoder_reg[7]  ( .D(n5797), .CPN(n9142), .CDN(n9151), .Q(
        Decoder[7]) );
  DFNCND1 \Decoder_reg[6]  ( .D(n5934), .CPN(n9142), .CDN(n9152), .Q(
        Decoder[6]) );
  DFNCND1 \Decoder_reg[5]  ( .D(n6070), .CPN(n9142), .CDN(n9153), .Q(
        Decoder[5]) );
  DFNCND1 \Decoder_reg[4]  ( .D(n6207), .CPN(n9142), .CDN(n9151), .Q(
        Decoder[4]) );
  DFNCND1 \Decoder_reg[3]  ( .D(n6344), .CPN(n9142), .CDN(n9152), .Q(
        Decoder[3]) );
  DFNCND1 \Decoder_reg[2]  ( .D(n6481), .CPN(n9142), .CDN(n9153), .Q(
        Decoder[2]) );
  DFNCND1 \Decoder_reg[1]  ( .D(n6618), .CPN(n9142), .CDN(n9150), .Q(
        Decoder[1]) );
  DFNCND1 \Decoder_reg[0]  ( .D(n6755), .CPN(n9142), .CDN(n9152), .Q(
        Decoder[0]) );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n6892), .CPN(n9138), .CDN(n9153), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(n6894), .E(SerValid), .CP(n9137), .CDN(n9153), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n6896), .CPN(n9138), .CDN(n9154), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(n6898), .E(SerValid), .CP(n9137), .CDN(n9151), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(n6900), .E(SerValid), .CP(n9137), .CDN(n9151), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(n6902), .E(SerValid), .CP(n9137), .CDN(n9149), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n6904), .CPN(n9141), .CDN(n9154), .Q(ParOut[0]), .QN(n63) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n6908), .CPN(n9141), .CDN(n9149), .Q(ParOut[1]), .QN(n62) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n6912), .CPN(n9141), .CDN(n9153), .Q(ParOut[2]), .QN(n61) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n6916), .CPN(n9141), .CDN(n9151), .Q(ParOut[3]), .QN(n60) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n6920), .CPN(n9141), .CDN(n9150), .Q(ParOut[4]), .QN(n59) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n6924), .CPN(n9141), .CDN(n9152), .Q(ParOut[5]), .QN(n58) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n6928), .CPN(n9141), .CDN(n9148), .Q(ParOut[6]), .QN(n57) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n6932), .CPN(n9140), .CDN(n9153), .Q(ParOut[7]), .QN(n56) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n6936), .CPN(n9140), .CDN(n9149), .Q(ParOut[8]), .QN(n55) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n6940), .CPN(n9140), .CDN(n9147), .Q(ParOut[9]), .QN(n54) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n6944), .CPN(n9140), .CDN(n9154), .Q(
        ParOut[10]), .QN(n53) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n6948), .CPN(n9140), .CDN(n9152), .Q(
        ParOut[11]), .QN(n52) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n6952), .CPN(n9140), .CDN(n9153), .Q(
        ParOut[12]), .QN(n51) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n6956), .CPN(n9140), .CDN(n9148), .Q(
        ParOut[13]), .QN(n50) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n6960), .CPN(n9140), .CDN(n9153), .Q(
        ParOut[14]), .QN(n49) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n6964), .CPN(n9140), .CDN(n9152), .Q(
        ParOut[15]), .QN(n48) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n6968), .CPN(n9139), .CDN(n9151), .Q(
        ParOut[16]), .QN(n47) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n6972), .CPN(n9139), .CDN(n9154), .Q(
        ParOut[17]), .QN(n46) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n6976), .CPN(n9139), .CDN(n9150), .Q(
        ParOut[18]), .QN(n45) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n6980), .CPN(n9139), .CDN(n9148), .Q(
        ParOut[19]), .QN(n44) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n6984), .CPN(n9139), .CDN(n9149), .Q(
        ParOut[20]), .QN(n43) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n6988), .CPN(n9139), .CDN(n9148), .Q(
        ParOut[21]), .QN(n42) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n6992), .CPN(n9139), .CDN(n9153), .Q(
        ParOut[22]), .QN(n41) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n6996), .CPN(n9139), .CDN(n9149), .Q(
        ParOut[23]), .QN(n40) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n7000), .CPN(n9139), .CDN(n9147), .Q(
        ParOut[24]), .QN(n39) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n7004), .CPN(n9138), .CDN(n9147), .Q(
        ParOut[25]), .QN(n38) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n7008), .CPN(n9138), .CDN(n9148), .Q(
        ParOut[26]), .QN(n37) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n7012), .CPN(n9138), .CDN(n9151), .Q(
        ParOut[27]), .QN(n36) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n7016), .CPN(n9138), .CDN(n9152), .Q(
        ParOut[28]), .QN(n35) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n7020), .CPN(n9138), .CDN(n9154), .Q(
        ParOut[29]), .QN(n34) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n7024), .CPN(n9138), .CDN(n9152), .Q(
        ParOut[30]), .QN(n33) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n7028), .CPN(n9138), .CDN(n9152), .Q(
        ParOut[31]), .QN(n32) );
  EDFCNQD1 ParClkr_reg ( .D(n7032), .E(n7034), .CP(n9137), .CDN(n9151), .Q(
        ParClk) );
  DFNCND1 ParValidr_reg ( .D(n7036), .CPN(n9137), .CDN(n9150), .Q(ParValid), 
        .QN(n29) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n9141), .CDN(n9154), .Q(n27), .QN(n2)
         );
  DFNCND1 UnLoad_reg ( .D(n9017), .CPN(n9141), .CDN(n9154), .Q(n1), .QN(n231)
         );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n9019), .CPN(n9137), .CDN(n9154), .QN(
        n232) );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n9022), .CPN(n9137), .CDN(n9154), .QN(
        n230) );
  IOA22D0 U3 ( .B1(n9128), .B2(n32), .A1(n1), .A2(Decoder[31]), .ZN(n101) );
  CKAN2D0 U4 ( .A1(N30), .A2(n2), .Z(N38) );
  INVD0 U5 ( .I(ParValidTimer[0]), .ZN(n6) );
  BUFFD0 U6 ( .I(n2802), .Z(n4) );
  CKBD0 U7 ( .CLK(FrameSR[62]), .C(n5) );
  BUFFD0 U8 ( .I(n8992), .Z(n30) );
  CKBD0 U9 ( .CLK(FrameSR[21]), .C(n31) );
  CKBD0 U10 ( .CLK(n31), .C(n64) );
  BUFFD0 U11 ( .I(n64), .Z(n65) );
  CKBD0 U12 ( .CLK(n65), .C(n66) );
  CKBD0 U13 ( .CLK(n66), .C(n67) );
  CKBD0 U14 ( .CLK(n67), .C(n68) );
  CKBD0 U15 ( .CLK(n68), .C(n69) );
  CKBD0 U16 ( .CLK(n69), .C(n70) );
  CKBD0 U17 ( .CLK(n70), .C(n71) );
  CKBD0 U18 ( .CLK(n71), .C(n72) );
  CKBD0 U19 ( .CLK(n72), .C(n73) );
  CKBD0 U20 ( .CLK(n73), .C(n74) );
  CKBD0 U21 ( .CLK(n74), .C(n75) );
  BUFFD0 U22 ( .I(n75), .Z(n76) );
  CKBD0 U23 ( .CLK(n76), .C(n77) );
  CKBD0 U24 ( .CLK(n77), .C(n78) );
  CKBD0 U25 ( .CLK(n78), .C(n79) );
  CKBD0 U26 ( .CLK(n79), .C(n80) );
  CKBD0 U27 ( .CLK(n80), .C(n81) );
  CKBD0 U28 ( .CLK(n81), .C(n82) );
  CKBD0 U29 ( .CLK(n82), .C(n83) );
  CKBD0 U30 ( .CLK(n83), .C(n84) );
  CKBD0 U31 ( .CLK(n84), .C(n85) );
  BUFFD0 U32 ( .I(n85), .Z(n86) );
  CKBD0 U33 ( .CLK(n86), .C(n87) );
  CKBD0 U34 ( .CLK(n87), .C(n88) );
  CKBD0 U35 ( .CLK(n88), .C(n89) );
  CKBD0 U36 ( .CLK(n89), .C(n90) );
  CKBD0 U37 ( .CLK(n90), .C(n91) );
  CKBD0 U38 ( .CLK(n91), .C(n92) );
  CKBD0 U41 ( .CLK(n92), .C(n93) );
  CKBD0 U42 ( .CLK(n93), .C(n94) );
  CKBD0 U43 ( .CLK(n94), .C(n95) );
  CKBD0 U44 ( .CLK(n95), .C(n165) );
  BUFFD0 U45 ( .I(n165), .Z(n166) );
  CKBD0 U46 ( .CLK(n166), .C(n167) );
  CKBD0 U47 ( .CLK(n167), .C(n168) );
  CKBD0 U48 ( .CLK(n168), .C(n169) );
  CKBD0 U49 ( .CLK(n169), .C(n170) );
  CKBD0 U50 ( .CLK(n170), .C(n171) );
  CKBD0 U51 ( .CLK(n171), .C(n172) );
  CKBD0 U52 ( .CLK(n172), .C(n173) );
  CKBD0 U53 ( .CLK(n173), .C(n174) );
  CKBD0 U54 ( .CLK(n174), .C(n175) );
  CKBD0 U55 ( .CLK(n175), .C(n176) );
  BUFFD0 U56 ( .I(n176), .Z(n177) );
  CKBD0 U57 ( .CLK(n177), .C(n178) );
  CKBD0 U58 ( .CLK(n178), .C(n179) );
  CKBD0 U59 ( .CLK(n179), .C(n180) );
  CKBD0 U60 ( .CLK(n180), .C(n181) );
  CKBD0 U61 ( .CLK(n181), .C(n182) );
  CKBD0 U62 ( .CLK(n182), .C(n183) );
  CKBD0 U63 ( .CLK(n183), .C(n184) );
  CKBD0 U64 ( .CLK(n184), .C(n185) );
  CKBD0 U65 ( .CLK(n185), .C(n186) );
  CKBD0 U66 ( .CLK(n186), .C(n187) );
  BUFFD0 U67 ( .I(n187), .Z(n188) );
  CKBD0 U68 ( .CLK(n188), .C(n189) );
  CKBD0 U69 ( .CLK(n189), .C(n190) );
  CKBD0 U70 ( .CLK(n190), .C(n191) );
  CKBD0 U71 ( .CLK(n191), .C(n192) );
  CKBD0 U72 ( .CLK(n192), .C(n193) );
  CKBD0 U73 ( .CLK(n193), .C(n194) );
  CKBD0 U74 ( .CLK(n194), .C(n195) );
  CKBD0 U75 ( .CLK(n195), .C(n196) );
  CKBD0 U76 ( .CLK(n196), .C(n197) );
  CKBD0 U77 ( .CLK(n197), .C(n198) );
  BUFFD0 U78 ( .I(n198), .Z(n199) );
  CKBD0 U79 ( .CLK(n199), .C(n200) );
  CKBD0 U80 ( .CLK(n200), .C(n201) );
  CKBD0 U81 ( .CLK(n201), .C(n202) );
  CKBD0 U82 ( .CLK(n202), .C(n203) );
  CKBD0 U83 ( .CLK(n203), .C(n204) );
  CKBD0 U84 ( .CLK(n204), .C(n205) );
  CKBD0 U85 ( .CLK(n205), .C(n206) );
  CKBD0 U86 ( .CLK(n206), .C(n207) );
  CKBD0 U87 ( .CLK(n207), .C(n208) );
  CKBD0 U88 ( .CLK(n208), .C(n209) );
  BUFFD0 U89 ( .I(n209), .Z(n210) );
  CKBD0 U90 ( .CLK(n210), .C(n211) );
  CKBD0 U91 ( .CLK(n211), .C(n212) );
  CKBD0 U93 ( .CLK(n212), .C(n213) );
  CKBD0 U95 ( .CLK(n213), .C(n214) );
  CKBD0 U97 ( .CLK(n214), .C(n215) );
  CKBD0 U98 ( .CLK(n215), .C(n216) );
  CKBD0 U100 ( .CLK(n216), .C(n217) );
  CKBD0 U102 ( .CLK(n217), .C(n218) );
  CKBD0 U103 ( .CLK(n218), .C(n219) );
  CKBD0 U104 ( .CLK(n219), .C(n220) );
  BUFFD0 U105 ( .I(n220), .Z(n221) );
  CKBD0 U106 ( .CLK(n221), .C(n222) );
  CKBD0 U107 ( .CLK(n222), .C(n223) );
  CKBD0 U108 ( .CLK(n223), .C(n224) );
  CKBD0 U109 ( .CLK(n224), .C(n225) );
  CKBD0 U110 ( .CLK(n225), .C(n226) );
  BUFFD0 U111 ( .I(n8973), .Z(n227) );
  CKBD0 U112 ( .CLK(FrameSR[22]), .C(n228) );
  BUFFD0 U113 ( .I(n228), .Z(n229) );
  CKBD0 U114 ( .CLK(n229), .C(n233) );
  CKBD0 U115 ( .CLK(n233), .C(n234) );
  CKBD0 U116 ( .CLK(n234), .C(n235) );
  CKBD0 U117 ( .CLK(n235), .C(n236) );
  CKBD0 U118 ( .CLK(n236), .C(n237) );
  CKBD0 U119 ( .CLK(n237), .C(n238) );
  CKBD0 U120 ( .CLK(n238), .C(n239) );
  CKBD0 U121 ( .CLK(n239), .C(n240) );
  CKBD0 U122 ( .CLK(n240), .C(n241) );
  CKBD0 U123 ( .CLK(n241), .C(n242) );
  BUFFD0 U124 ( .I(n242), .Z(n243) );
  CKBD0 U125 ( .CLK(n243), .C(n244) );
  CKBD0 U126 ( .CLK(n244), .C(n245) );
  CKBD0 U127 ( .CLK(n245), .C(n246) );
  CKBD0 U128 ( .CLK(n246), .C(n247) );
  CKBD0 U129 ( .CLK(n247), .C(n248) );
  CKBD0 U130 ( .CLK(n248), .C(n249) );
  CKBD0 U131 ( .CLK(n249), .C(n250) );
  CKBD0 U132 ( .CLK(n250), .C(n251) );
  CKBD0 U133 ( .CLK(n251), .C(n252) );
  CKBD0 U134 ( .CLK(n252), .C(n253) );
  BUFFD0 U135 ( .I(n253), .Z(n254) );
  CKBD0 U136 ( .CLK(n254), .C(n255) );
  CKBD0 U137 ( .CLK(n255), .C(n256) );
  CKBD0 U138 ( .CLK(n256), .C(n257) );
  CKBD0 U139 ( .CLK(n257), .C(n258) );
  CKBD0 U140 ( .CLK(n258), .C(n259) );
  CKBD0 U141 ( .CLK(n259), .C(n260) );
  CKBD0 U142 ( .CLK(n260), .C(n261) );
  CKBD0 U143 ( .CLK(n261), .C(n262) );
  CKBD0 U144 ( .CLK(n262), .C(n263) );
  CKBD0 U145 ( .CLK(n263), .C(n264) );
  BUFFD0 U146 ( .I(n264), .Z(n265) );
  CKBD0 U147 ( .CLK(n265), .C(n266) );
  CKBD0 U148 ( .CLK(n266), .C(n267) );
  CKBD0 U149 ( .CLK(n267), .C(n268) );
  CKBD0 U150 ( .CLK(n268), .C(n269) );
  CKBD0 U151 ( .CLK(n269), .C(n270) );
  CKBD0 U152 ( .CLK(n270), .C(n271) );
  CKBD0 U153 ( .CLK(n271), .C(n272) );
  CKBD0 U154 ( .CLK(n272), .C(n273) );
  CKBD0 U155 ( .CLK(n273), .C(n274) );
  BUFFD0 U156 ( .I(n274), .Z(n275) );
  CKBD0 U157 ( .CLK(n275), .C(n276) );
  CKBD0 U158 ( .CLK(n276), .C(n277) );
  CKBD0 U159 ( .CLK(n277), .C(n278) );
  CKBD0 U160 ( .CLK(n278), .C(n279) );
  CKBD0 U161 ( .CLK(n279), .C(n280) );
  CKBD0 U162 ( .CLK(n280), .C(n281) );
  CKBD0 U163 ( .CLK(n281), .C(n282) );
  CKBD0 U164 ( .CLK(n282), .C(n283) );
  CKBD0 U165 ( .CLK(n283), .C(n284) );
  CKBD0 U166 ( .CLK(n284), .C(n285) );
  BUFFD0 U167 ( .I(n285), .Z(n286) );
  CKBD0 U168 ( .CLK(n286), .C(n287) );
  CKBD0 U169 ( .CLK(n287), .C(n288) );
  CKBD0 U170 ( .CLK(n288), .C(n289) );
  CKBD0 U171 ( .CLK(n289), .C(n290) );
  CKBD0 U172 ( .CLK(n290), .C(n291) );
  CKBD0 U173 ( .CLK(n291), .C(n292) );
  CKBD0 U174 ( .CLK(n292), .C(n293) );
  CKBD0 U175 ( .CLK(n293), .C(n294) );
  CKBD0 U176 ( .CLK(n294), .C(n295) );
  CKBD0 U177 ( .CLK(n295), .C(n296) );
  BUFFD0 U178 ( .I(n296), .Z(n297) );
  CKBD0 U179 ( .CLK(n297), .C(n298) );
  CKBD0 U180 ( .CLK(n298), .C(n299) );
  CKBD0 U181 ( .CLK(n299), .C(n300) );
  CKBD0 U182 ( .CLK(n300), .C(n301) );
  CKBD0 U183 ( .CLK(n301), .C(n302) );
  CKBD0 U184 ( .CLK(n302), .C(n303) );
  CKBD0 U185 ( .CLK(n303), .C(n304) );
  CKBD0 U186 ( .CLK(n304), .C(n305) );
  CKBD0 U187 ( .CLK(n305), .C(n306) );
  CKBD0 U188 ( .CLK(n306), .C(n307) );
  BUFFD0 U189 ( .I(n307), .Z(n308) );
  CKBD0 U190 ( .CLK(n308), .C(n309) );
  CKBD0 U191 ( .CLK(n309), .C(n310) );
  CKBD0 U192 ( .CLK(n310), .C(n311) );
  CKBD0 U193 ( .CLK(n311), .C(n312) );
  CKBD0 U194 ( .CLK(n312), .C(n313) );
  CKBD0 U195 ( .CLK(n313), .C(n314) );
  CKBD0 U196 ( .CLK(n314), .C(n315) );
  CKBD0 U197 ( .CLK(n315), .C(n316) );
  CKBD0 U198 ( .CLK(n316), .C(n317) );
  CKBD0 U199 ( .CLK(n317), .C(n318) );
  BUFFD0 U200 ( .I(n318), .Z(n319) );
  CKBD0 U201 ( .CLK(n319), .C(n320) );
  CKBD0 U202 ( .CLK(n320), .C(n321) );
  CKBD0 U203 ( .CLK(n321), .C(n322) );
  CKBD0 U204 ( .CLK(n322), .C(n323) );
  CKBD0 U205 ( .CLK(n323), .C(n324) );
  CKBD0 U206 ( .CLK(n324), .C(n325) );
  CKBD0 U207 ( .CLK(n325), .C(n326) );
  BUFFD0 U208 ( .I(n8979), .Z(n327) );
  CKBD0 U209 ( .CLK(FrameSR[36]), .C(n328) );
  CKBD0 U210 ( .CLK(n328), .C(n329) );
  CKBD0 U211 ( .CLK(n329), .C(n330) );
  CKBD0 U212 ( .CLK(n330), .C(n331) );
  CKBD0 U213 ( .CLK(n331), .C(n332) );
  CKBD0 U214 ( .CLK(n332), .C(n333) );
  CKBD0 U215 ( .CLK(n333), .C(n334) );
  CKBD0 U216 ( .CLK(n334), .C(n335) );
  CKBD0 U217 ( .CLK(n335), .C(n336) );
  CKBD0 U218 ( .CLK(n336), .C(n337) );
  BUFFD0 U219 ( .I(n337), .Z(n338) );
  CKBD0 U220 ( .CLK(n338), .C(n339) );
  CKBD0 U221 ( .CLK(n339), .C(n340) );
  CKBD0 U222 ( .CLK(n340), .C(n341) );
  CKBD0 U223 ( .CLK(n341), .C(n342) );
  CKBD0 U224 ( .CLK(n342), .C(n343) );
  CKBD0 U225 ( .CLK(n343), .C(n344) );
  CKBD0 U226 ( .CLK(n344), .C(n345) );
  CKBD0 U227 ( .CLK(n345), .C(n346) );
  CKBD0 U228 ( .CLK(n346), .C(n347) );
  CKBD0 U229 ( .CLK(n347), .C(n348) );
  BUFFD0 U230 ( .I(n348), .Z(n349) );
  CKBD0 U231 ( .CLK(n349), .C(n350) );
  CKBD0 U232 ( .CLK(n350), .C(n351) );
  CKBD0 U233 ( .CLK(n351), .C(n352) );
  CKBD0 U234 ( .CLK(n352), .C(n353) );
  CKBD0 U235 ( .CLK(n353), .C(n354) );
  CKBD0 U236 ( .CLK(n354), .C(n355) );
  CKBD0 U237 ( .CLK(n355), .C(n356) );
  CKBD0 U238 ( .CLK(n356), .C(n357) );
  CKBD0 U239 ( .CLK(n357), .C(n358) );
  CKBD0 U240 ( .CLK(n358), .C(n359) );
  BUFFD0 U241 ( .I(n359), .Z(n360) );
  CKBD0 U242 ( .CLK(n360), .C(n361) );
  CKBD0 U243 ( .CLK(n361), .C(n362) );
  CKBD0 U244 ( .CLK(n362), .C(n363) );
  CKBD0 U245 ( .CLK(n363), .C(n364) );
  CKBD0 U246 ( .CLK(n364), .C(n365) );
  CKBD0 U247 ( .CLK(n365), .C(n366) );
  CKBD0 U248 ( .CLK(n366), .C(n367) );
  CKBD0 U249 ( .CLK(n367), .C(n368) );
  CKBD0 U250 ( .CLK(n368), .C(n369) );
  BUFFD0 U251 ( .I(n369), .Z(n370) );
  CKBD0 U252 ( .CLK(n370), .C(n371) );
  CKBD0 U253 ( .CLK(n371), .C(n372) );
  CKBD0 U254 ( .CLK(n372), .C(n373) );
  CKBD0 U255 ( .CLK(n373), .C(n374) );
  CKBD0 U256 ( .CLK(n374), .C(n375) );
  CKBD0 U257 ( .CLK(n375), .C(n376) );
  CKBD0 U258 ( .CLK(n376), .C(n377) );
  CKBD0 U259 ( .CLK(n377), .C(n378) );
  CKBD0 U260 ( .CLK(n378), .C(n379) );
  CKBD0 U261 ( .CLK(n379), .C(n380) );
  BUFFD0 U262 ( .I(n380), .Z(n381) );
  CKBD0 U263 ( .CLK(n381), .C(n382) );
  CKBD0 U264 ( .CLK(n382), .C(n383) );
  CKBD0 U265 ( .CLK(n383), .C(n384) );
  CKBD0 U266 ( .CLK(n384), .C(n385) );
  CKBD0 U267 ( .CLK(n385), .C(n386) );
  CKBD0 U268 ( .CLK(n386), .C(n387) );
  CKBD0 U269 ( .CLK(n387), .C(n388) );
  CKBD0 U270 ( .CLK(n388), .C(n389) );
  CKBD0 U271 ( .CLK(n389), .C(n390) );
  CKBD0 U272 ( .CLK(n390), .C(n391) );
  BUFFD0 U273 ( .I(n391), .Z(n392) );
  CKBD0 U274 ( .CLK(n392), .C(n393) );
  CKBD0 U275 ( .CLK(n393), .C(n394) );
  CKBD0 U276 ( .CLK(n394), .C(n395) );
  CKBD0 U277 ( .CLK(n395), .C(n396) );
  CKBD0 U278 ( .CLK(n396), .C(n397) );
  CKBD0 U279 ( .CLK(n397), .C(n398) );
  CKBD0 U280 ( .CLK(n398), .C(n399) );
  CKBD0 U281 ( .CLK(n399), .C(n400) );
  CKBD0 U282 ( .CLK(n400), .C(n401) );
  CKBD0 U283 ( .CLK(n401), .C(n402) );
  BUFFD0 U284 ( .I(n402), .Z(n403) );
  CKBD0 U285 ( .CLK(n403), .C(n404) );
  CKBD0 U286 ( .CLK(n404), .C(n405) );
  CKBD0 U287 ( .CLK(n405), .C(n406) );
  CKBD0 U288 ( .CLK(n406), .C(n407) );
  CKBD0 U289 ( .CLK(n407), .C(n408) );
  CKBD0 U290 ( .CLK(n408), .C(n409) );
  CKBD0 U291 ( .CLK(n409), .C(n410) );
  CKBD0 U292 ( .CLK(n410), .C(n411) );
  CKBD0 U293 ( .CLK(n411), .C(n412) );
  CKBD0 U294 ( .CLK(n412), .C(n413) );
  BUFFD0 U295 ( .I(n413), .Z(n414) );
  CKBD0 U296 ( .CLK(n414), .C(n415) );
  CKBD0 U297 ( .CLK(n415), .C(n416) );
  CKBD0 U298 ( .CLK(n416), .C(n417) );
  CKBD0 U299 ( .CLK(n417), .C(n418) );
  CKBD0 U300 ( .CLK(n418), .C(n419) );
  CKBD0 U301 ( .CLK(n419), .C(n420) );
  CKBD0 U302 ( .CLK(n420), .C(n421) );
  CKBD0 U303 ( .CLK(n421), .C(n422) );
  BUFFD0 U304 ( .I(n8974), .Z(n423) );
  CKBD0 U305 ( .CLK(FrameSR[37]), .C(n424) );
  BUFFD0 U306 ( .I(n424), .Z(n425) );
  CKBD0 U307 ( .CLK(n425), .C(n426) );
  CKBD0 U308 ( .CLK(n426), .C(n427) );
  CKBD0 U309 ( .CLK(n427), .C(n428) );
  CKBD0 U310 ( .CLK(n428), .C(n429) );
  CKBD0 U311 ( .CLK(n429), .C(n430) );
  CKBD0 U312 ( .CLK(n430), .C(n431) );
  CKBD0 U313 ( .CLK(n431), .C(n432) );
  CKBD0 U314 ( .CLK(n432), .C(n433) );
  CKBD0 U315 ( .CLK(n433), .C(n434) );
  CKBD0 U316 ( .CLK(n434), .C(n435) );
  BUFFD0 U317 ( .I(n435), .Z(n436) );
  CKBD0 U318 ( .CLK(n436), .C(n437) );
  CKBD0 U319 ( .CLK(n437), .C(n438) );
  CKBD0 U320 ( .CLK(n438), .C(n439) );
  CKBD0 U321 ( .CLK(n439), .C(n440) );
  CKBD0 U322 ( .CLK(n440), .C(n441) );
  CKBD0 U323 ( .CLK(n441), .C(n442) );
  CKBD0 U324 ( .CLK(n442), .C(n443) );
  CKBD0 U325 ( .CLK(n443), .C(n444) );
  CKBD0 U326 ( .CLK(n444), .C(n445) );
  CKBD0 U327 ( .CLK(n445), .C(n446) );
  BUFFD0 U328 ( .I(n446), .Z(n447) );
  CKBD0 U329 ( .CLK(n447), .C(n448) );
  CKBD0 U330 ( .CLK(n448), .C(n449) );
  CKBD0 U331 ( .CLK(n449), .C(n450) );
  CKBD0 U332 ( .CLK(n450), .C(n451) );
  CKBD0 U333 ( .CLK(n451), .C(n452) );
  CKBD0 U334 ( .CLK(n452), .C(n453) );
  CKBD0 U335 ( .CLK(n453), .C(n454) );
  CKBD0 U336 ( .CLK(n454), .C(n455) );
  CKBD0 U337 ( .CLK(n455), .C(n456) );
  CKBD0 U338 ( .CLK(n456), .C(n457) );
  BUFFD0 U339 ( .I(n457), .Z(n458) );
  CKBD0 U340 ( .CLK(n458), .C(n459) );
  CKBD0 U341 ( .CLK(n459), .C(n460) );
  CKBD0 U342 ( .CLK(n460), .C(n461) );
  CKBD0 U343 ( .CLK(n461), .C(n462) );
  CKBD0 U344 ( .CLK(n462), .C(n463) );
  CKBD0 U345 ( .CLK(n463), .C(n464) );
  CKBD0 U346 ( .CLK(n464), .C(n465) );
  CKBD0 U347 ( .CLK(n465), .C(n466) );
  CKBD0 U348 ( .CLK(n466), .C(n467) );
  BUFFD0 U349 ( .I(n467), .Z(n468) );
  CKBD0 U350 ( .CLK(n468), .C(n469) );
  CKBD0 U351 ( .CLK(n469), .C(n470) );
  CKBD0 U352 ( .CLK(n470), .C(n471) );
  CKBD0 U353 ( .CLK(n471), .C(n472) );
  CKBD0 U354 ( .CLK(n472), .C(n473) );
  CKBD0 U355 ( .CLK(n473), .C(n474) );
  CKBD0 U356 ( .CLK(n474), .C(n475) );
  CKBD0 U357 ( .CLK(n475), .C(n476) );
  CKBD0 U358 ( .CLK(n476), .C(n477) );
  CKBD0 U359 ( .CLK(n477), .C(n478) );
  BUFFD0 U360 ( .I(n478), .Z(n479) );
  CKBD0 U361 ( .CLK(n479), .C(n480) );
  CKBD0 U362 ( .CLK(n480), .C(n481) );
  CKBD0 U363 ( .CLK(n481), .C(n482) );
  CKBD0 U364 ( .CLK(n482), .C(n483) );
  CKBD0 U365 ( .CLK(n483), .C(n484) );
  CKBD0 U366 ( .CLK(n484), .C(n485) );
  CKBD0 U367 ( .CLK(n485), .C(n486) );
  CKBD0 U368 ( .CLK(n486), .C(n487) );
  CKBD0 U369 ( .CLK(n487), .C(n488) );
  CKBD0 U370 ( .CLK(n488), .C(n489) );
  BUFFD0 U371 ( .I(n489), .Z(n490) );
  CKBD0 U372 ( .CLK(n490), .C(n491) );
  CKBD0 U373 ( .CLK(n491), .C(n492) );
  CKBD0 U374 ( .CLK(n492), .C(n493) );
  CKBD0 U375 ( .CLK(n493), .C(n494) );
  CKBD0 U376 ( .CLK(n494), .C(n495) );
  CKBD0 U377 ( .CLK(n495), .C(n496) );
  CKBD0 U378 ( .CLK(n496), .C(n497) );
  CKBD0 U379 ( .CLK(n497), .C(n498) );
  CKBD0 U380 ( .CLK(n498), .C(n499) );
  CKBD0 U381 ( .CLK(n499), .C(n500) );
  BUFFD0 U382 ( .I(n500), .Z(n501) );
  CKBD0 U383 ( .CLK(n501), .C(n502) );
  CKBD0 U384 ( .CLK(n502), .C(n503) );
  CKBD0 U385 ( .CLK(n503), .C(n504) );
  CKBD0 U386 ( .CLK(n504), .C(n505) );
  CKBD0 U387 ( .CLK(n505), .C(n506) );
  CKBD0 U388 ( .CLK(n506), .C(n507) );
  CKBD0 U389 ( .CLK(n507), .C(n508) );
  CKBD0 U390 ( .CLK(n508), .C(n509) );
  CKBD0 U391 ( .CLK(n509), .C(n510) );
  CKBD0 U392 ( .CLK(n510), .C(n511) );
  BUFFD0 U393 ( .I(n511), .Z(n512) );
  CKBD0 U394 ( .CLK(n512), .C(n513) );
  CKBD0 U395 ( .CLK(n513), .C(n514) );
  CKBD0 U396 ( .CLK(n514), .C(n515) );
  CKBD0 U397 ( .CLK(n515), .C(n516) );
  CKBD0 U398 ( .CLK(n516), .C(n517) );
  CKBD0 U399 ( .CLK(n517), .C(n518) );
  CKBD0 U400 ( .CLK(n518), .C(n519) );
  BUFFD0 U401 ( .I(n8978), .Z(n520) );
  CKBD0 U402 ( .CLK(FrameSR[52]), .C(n521) );
  CKBD0 U403 ( .CLK(n521), .C(n522) );
  CKBD0 U404 ( .CLK(n522), .C(n523) );
  CKBD0 U405 ( .CLK(n523), .C(n524) );
  CKBD0 U406 ( .CLK(n524), .C(n525) );
  CKBD0 U407 ( .CLK(n525), .C(n526) );
  CKBD0 U408 ( .CLK(n526), .C(n527) );
  CKBD0 U409 ( .CLK(n527), .C(n528) );
  CKBD0 U410 ( .CLK(n528), .C(n529) );
  CKBD0 U411 ( .CLK(n529), .C(n530) );
  BUFFD0 U412 ( .I(n530), .Z(n531) );
  CKBD0 U413 ( .CLK(n531), .C(n532) );
  CKBD0 U414 ( .CLK(n532), .C(n533) );
  CKBD0 U415 ( .CLK(n533), .C(n534) );
  CKBD0 U416 ( .CLK(n534), .C(n535) );
  CKBD0 U417 ( .CLK(n535), .C(n536) );
  CKBD0 U418 ( .CLK(n536), .C(n537) );
  CKBD0 U419 ( .CLK(n537), .C(n538) );
  CKBD0 U420 ( .CLK(n538), .C(n539) );
  CKBD0 U421 ( .CLK(n539), .C(n540) );
  CKBD0 U422 ( .CLK(n540), .C(n541) );
  BUFFD0 U423 ( .I(n541), .Z(n542) );
  CKBD0 U424 ( .CLK(n542), .C(n543) );
  CKBD0 U425 ( .CLK(n543), .C(n544) );
  CKBD0 U426 ( .CLK(n544), .C(n545) );
  CKBD0 U427 ( .CLK(n545), .C(n546) );
  CKBD0 U428 ( .CLK(n546), .C(n547) );
  CKBD0 U429 ( .CLK(n547), .C(n548) );
  CKBD0 U430 ( .CLK(n548), .C(n549) );
  CKBD0 U431 ( .CLK(n549), .C(n550) );
  CKBD0 U432 ( .CLK(n550), .C(n551) );
  CKBD0 U433 ( .CLK(n551), .C(n552) );
  BUFFD0 U434 ( .I(n552), .Z(n553) );
  CKBD0 U435 ( .CLK(n553), .C(n554) );
  CKBD0 U436 ( .CLK(n554), .C(n555) );
  CKBD0 U437 ( .CLK(n555), .C(n556) );
  CKBD0 U438 ( .CLK(n556), .C(n557) );
  CKBD0 U439 ( .CLK(n557), .C(n558) );
  CKBD0 U440 ( .CLK(n558), .C(n559) );
  CKBD0 U441 ( .CLK(n559), .C(n560) );
  CKBD0 U442 ( .CLK(n560), .C(n561) );
  CKBD0 U443 ( .CLK(n561), .C(n562) );
  CKBD0 U444 ( .CLK(n562), .C(n563) );
  BUFFD0 U445 ( .I(n563), .Z(n564) );
  CKBD0 U446 ( .CLK(n564), .C(n565) );
  CKBD0 U447 ( .CLK(n565), .C(n566) );
  CKBD0 U448 ( .CLK(n566), .C(n567) );
  CKBD0 U449 ( .CLK(n567), .C(n568) );
  CKBD0 U450 ( .CLK(n568), .C(n569) );
  CKBD0 U451 ( .CLK(n569), .C(n570) );
  CKBD0 U452 ( .CLK(n570), .C(n571) );
  CKBD0 U453 ( .CLK(n571), .C(n572) );
  CKBD0 U454 ( .CLK(n572), .C(n573) );
  CKBD0 U455 ( .CLK(n573), .C(n574) );
  BUFFD0 U456 ( .I(n574), .Z(n575) );
  CKBD0 U457 ( .CLK(n575), .C(n576) );
  CKBD0 U458 ( .CLK(n576), .C(n577) );
  CKBD0 U459 ( .CLK(n577), .C(n578) );
  CKBD0 U460 ( .CLK(n578), .C(n579) );
  CKBD0 U461 ( .CLK(n579), .C(n580) );
  CKBD0 U462 ( .CLK(n580), .C(n581) );
  CKBD0 U463 ( .CLK(n581), .C(n582) );
  CKBD0 U464 ( .CLK(n582), .C(n583) );
  CKBD0 U465 ( .CLK(n583), .C(n584) );
  CKBD0 U466 ( .CLK(n584), .C(n585) );
  BUFFD0 U467 ( .I(n585), .Z(n586) );
  CKBD0 U468 ( .CLK(n586), .C(n587) );
  CKBD0 U469 ( .CLK(n587), .C(n588) );
  CKBD0 U470 ( .CLK(n588), .C(n589) );
  CKBD0 U471 ( .CLK(n589), .C(n590) );
  CKBD0 U472 ( .CLK(n590), .C(n591) );
  CKBD0 U473 ( .CLK(n591), .C(n592) );
  CKBD0 U474 ( .CLK(n592), .C(n593) );
  CKBD0 U475 ( .CLK(n593), .C(n594) );
  CKBD0 U476 ( .CLK(n594), .C(n595) );
  BUFFD0 U477 ( .I(n595), .Z(n596) );
  CKBD0 U478 ( .CLK(n596), .C(n597) );
  CKBD0 U479 ( .CLK(n597), .C(n598) );
  CKBD0 U480 ( .CLK(n598), .C(n599) );
  CKBD0 U481 ( .CLK(n599), .C(n600) );
  CKBD0 U482 ( .CLK(n600), .C(n601) );
  CKBD0 U483 ( .CLK(n601), .C(n602) );
  CKBD0 U484 ( .CLK(n602), .C(n603) );
  CKBD0 U485 ( .CLK(n603), .C(n604) );
  CKBD0 U486 ( .CLK(n604), .C(n605) );
  CKBD0 U487 ( .CLK(n605), .C(n606) );
  BUFFD0 U488 ( .I(n606), .Z(n607) );
  CKBD0 U489 ( .CLK(n607), .C(n608) );
  CKBD0 U490 ( .CLK(n608), .C(n609) );
  CKBD0 U491 ( .CLK(n609), .C(n610) );
  CKBD0 U492 ( .CLK(n610), .C(n611) );
  CKBD0 U493 ( .CLK(n611), .C(n612) );
  CKBD0 U494 ( .CLK(n612), .C(n613) );
  CKBD0 U495 ( .CLK(n613), .C(n614) );
  CKBD0 U496 ( .CLK(n614), .C(n615) );
  BUFFD0 U497 ( .I(n8972), .Z(n616) );
  CKBD0 U498 ( .CLK(FrameSR[53]), .C(n617) );
  BUFFD0 U499 ( .I(n617), .Z(n618) );
  CKBD0 U500 ( .CLK(n618), .C(n619) );
  CKBD0 U501 ( .CLK(n619), .C(n620) );
  CKBD0 U502 ( .CLK(n620), .C(n621) );
  CKBD0 U503 ( .CLK(n621), .C(n622) );
  CKBD0 U504 ( .CLK(n622), .C(n623) );
  CKBD0 U505 ( .CLK(n623), .C(n624) );
  CKBD0 U506 ( .CLK(n624), .C(n625) );
  CKBD0 U507 ( .CLK(n625), .C(n626) );
  CKBD0 U508 ( .CLK(n626), .C(n627) );
  CKBD0 U509 ( .CLK(n627), .C(n628) );
  BUFFD0 U510 ( .I(n628), .Z(n629) );
  CKBD0 U511 ( .CLK(n629), .C(n630) );
  CKBD0 U512 ( .CLK(n630), .C(n631) );
  CKBD0 U513 ( .CLK(n631), .C(n632) );
  CKBD0 U514 ( .CLK(n632), .C(n633) );
  CKBD0 U515 ( .CLK(n633), .C(n634) );
  CKBD0 U516 ( .CLK(n634), .C(n635) );
  CKBD0 U517 ( .CLK(n635), .C(n636) );
  CKBD0 U518 ( .CLK(n636), .C(n637) );
  CKBD0 U519 ( .CLK(n637), .C(n638) );
  CKBD0 U520 ( .CLK(n638), .C(n639) );
  BUFFD0 U521 ( .I(n639), .Z(n640) );
  CKBD0 U522 ( .CLK(n640), .C(n641) );
  CKBD0 U523 ( .CLK(n641), .C(n642) );
  CKBD0 U524 ( .CLK(n642), .C(n643) );
  CKBD0 U525 ( .CLK(n643), .C(n644) );
  CKBD0 U526 ( .CLK(n644), .C(n645) );
  CKBD0 U527 ( .CLK(n645), .C(n646) );
  CKBD0 U528 ( .CLK(n646), .C(n647) );
  CKBD0 U529 ( .CLK(n647), .C(n648) );
  CKBD0 U530 ( .CLK(n648), .C(n649) );
  CKBD0 U531 ( .CLK(n649), .C(n650) );
  BUFFD0 U532 ( .I(n650), .Z(n651) );
  CKBD0 U533 ( .CLK(n651), .C(n652) );
  CKBD0 U534 ( .CLK(n652), .C(n653) );
  CKBD0 U535 ( .CLK(n653), .C(n654) );
  CKBD0 U536 ( .CLK(n654), .C(n655) );
  CKBD0 U537 ( .CLK(n655), .C(n656) );
  CKBD0 U538 ( .CLK(n656), .C(n657) );
  CKBD0 U539 ( .CLK(n657), .C(n658) );
  CKBD0 U540 ( .CLK(n658), .C(n659) );
  CKBD0 U541 ( .CLK(n659), .C(n660) );
  BUFFD0 U542 ( .I(n660), .Z(n661) );
  CKBD0 U543 ( .CLK(n661), .C(n662) );
  CKBD0 U544 ( .CLK(n662), .C(n663) );
  CKBD0 U545 ( .CLK(n663), .C(n664) );
  CKBD0 U546 ( .CLK(n664), .C(n665) );
  CKBD0 U547 ( .CLK(n665), .C(n666) );
  CKBD0 U548 ( .CLK(n666), .C(n667) );
  CKBD0 U549 ( .CLK(n667), .C(n668) );
  CKBD0 U550 ( .CLK(n668), .C(n669) );
  CKBD0 U551 ( .CLK(n669), .C(n670) );
  CKBD0 U552 ( .CLK(n670), .C(n671) );
  BUFFD0 U553 ( .I(n671), .Z(n672) );
  CKBD0 U554 ( .CLK(n672), .C(n673) );
  CKBD0 U555 ( .CLK(n673), .C(n674) );
  CKBD0 U556 ( .CLK(n674), .C(n675) );
  CKBD0 U557 ( .CLK(n675), .C(n676) );
  CKBD0 U558 ( .CLK(n676), .C(n677) );
  CKBD0 U559 ( .CLK(n677), .C(n678) );
  CKBD0 U560 ( .CLK(n678), .C(n679) );
  CKBD0 U561 ( .CLK(n679), .C(n680) );
  CKBD0 U562 ( .CLK(n680), .C(n681) );
  CKBD0 U563 ( .CLK(n681), .C(n682) );
  BUFFD0 U564 ( .I(n682), .Z(n683) );
  CKBD0 U565 ( .CLK(n683), .C(n684) );
  CKBD0 U566 ( .CLK(n684), .C(n685) );
  CKBD0 U567 ( .CLK(n685), .C(n686) );
  CKBD0 U568 ( .CLK(n686), .C(n687) );
  CKBD0 U569 ( .CLK(n687), .C(n688) );
  CKBD0 U570 ( .CLK(n688), .C(n689) );
  CKBD0 U571 ( .CLK(n689), .C(n690) );
  CKBD0 U572 ( .CLK(n690), .C(n691) );
  CKBD0 U573 ( .CLK(n691), .C(n692) );
  CKBD0 U574 ( .CLK(n692), .C(n693) );
  BUFFD0 U575 ( .I(n693), .Z(n694) );
  CKBD0 U576 ( .CLK(n694), .C(n695) );
  CKBD0 U577 ( .CLK(n695), .C(n696) );
  CKBD0 U578 ( .CLK(n696), .C(n697) );
  CKBD0 U579 ( .CLK(n697), .C(n698) );
  CKBD0 U580 ( .CLK(n698), .C(n699) );
  CKBD0 U581 ( .CLK(n699), .C(n700) );
  CKBD0 U582 ( .CLK(n700), .C(n701) );
  CKBD0 U583 ( .CLK(n701), .C(n702) );
  CKBD0 U584 ( .CLK(n702), .C(n703) );
  CKBD0 U585 ( .CLK(n703), .C(n704) );
  BUFFD0 U586 ( .I(n704), .Z(n705) );
  CKBD0 U587 ( .CLK(n705), .C(n706) );
  CKBD0 U588 ( .CLK(n706), .C(n707) );
  CKBD0 U589 ( .CLK(n707), .C(n708) );
  CKBD0 U590 ( .CLK(n708), .C(n709) );
  CKBD0 U591 ( .CLK(n709), .C(n710) );
  CKBD0 U592 ( .CLK(n710), .C(n711) );
  CKBD0 U593 ( .CLK(n711), .C(n712) );
  BUFFD0 U594 ( .I(n4842), .Z(n713) );
  CKBD0 U595 ( .CLK(FrameSR[31]), .C(n714) );
  BUFFD0 U596 ( .I(n8966), .Z(n715) );
  CKBD0 U597 ( .CLK(FrameSR[38]), .C(n716) );
  BUFFD0 U598 ( .I(n716), .Z(n717) );
  CKBD0 U599 ( .CLK(n717), .C(n718) );
  CKBD0 U600 ( .CLK(n718), .C(n719) );
  CKBD0 U601 ( .CLK(n719), .C(n720) );
  CKBD0 U602 ( .CLK(n720), .C(n721) );
  CKBD0 U603 ( .CLK(n721), .C(n722) );
  CKBD0 U604 ( .CLK(n722), .C(n723) );
  CKBD0 U605 ( .CLK(n723), .C(n724) );
  CKBD0 U606 ( .CLK(n724), .C(n725) );
  CKBD0 U607 ( .CLK(n725), .C(n726) );
  CKBD0 U608 ( .CLK(n726), .C(n727) );
  BUFFD0 U609 ( .I(n727), .Z(n728) );
  CKBD0 U610 ( .CLK(n728), .C(n729) );
  CKBD0 U611 ( .CLK(n729), .C(n730) );
  CKBD0 U612 ( .CLK(n730), .C(n731) );
  CKBD0 U613 ( .CLK(n731), .C(n732) );
  CKBD0 U614 ( .CLK(n732), .C(n733) );
  CKBD0 U615 ( .CLK(n733), .C(n734) );
  CKBD0 U616 ( .CLK(n734), .C(n735) );
  CKBD0 U617 ( .CLK(n735), .C(n736) );
  CKBD0 U618 ( .CLK(n736), .C(n737) );
  CKBD0 U619 ( .CLK(n737), .C(n738) );
  BUFFD0 U620 ( .I(n738), .Z(n739) );
  CKBD0 U621 ( .CLK(n739), .C(n740) );
  CKBD0 U622 ( .CLK(n740), .C(n741) );
  CKBD0 U623 ( .CLK(n741), .C(n742) );
  CKBD0 U624 ( .CLK(n742), .C(n743) );
  CKBD0 U625 ( .CLK(n743), .C(n744) );
  CKBD0 U626 ( .CLK(n744), .C(n745) );
  CKBD0 U627 ( .CLK(n745), .C(n746) );
  CKBD0 U628 ( .CLK(n746), .C(n747) );
  CKBD0 U629 ( .CLK(n747), .C(n748) );
  CKBD0 U630 ( .CLK(n748), .C(n749) );
  BUFFD0 U631 ( .I(n749), .Z(n750) );
  CKBD0 U632 ( .CLK(n750), .C(n751) );
  CKBD0 U633 ( .CLK(n751), .C(n752) );
  CKBD0 U634 ( .CLK(n752), .C(n753) );
  CKBD0 U635 ( .CLK(n753), .C(n754) );
  CKBD0 U636 ( .CLK(n754), .C(n755) );
  CKBD0 U637 ( .CLK(n755), .C(n756) );
  CKBD0 U638 ( .CLK(n756), .C(n757) );
  CKBD0 U639 ( .CLK(n757), .C(n758) );
  CKBD0 U640 ( .CLK(n758), .C(n759) );
  BUFFD0 U641 ( .I(n759), .Z(n760) );
  CKBD0 U642 ( .CLK(n760), .C(n761) );
  CKBD0 U643 ( .CLK(n761), .C(n762) );
  CKBD0 U644 ( .CLK(n762), .C(n763) );
  CKBD0 U645 ( .CLK(n763), .C(n764) );
  CKBD0 U646 ( .CLK(n764), .C(n765) );
  CKBD0 U647 ( .CLK(n765), .C(n766) );
  CKBD0 U648 ( .CLK(n766), .C(n767) );
  CKBD0 U649 ( .CLK(n767), .C(n768) );
  CKBD0 U650 ( .CLK(n768), .C(n769) );
  CKBD0 U651 ( .CLK(n769), .C(n770) );
  BUFFD0 U652 ( .I(n770), .Z(n771) );
  CKBD0 U653 ( .CLK(n771), .C(n772) );
  CKBD0 U654 ( .CLK(n772), .C(n773) );
  CKBD0 U655 ( .CLK(n773), .C(n774) );
  CKBD0 U656 ( .CLK(n774), .C(n775) );
  CKBD0 U657 ( .CLK(n775), .C(n776) );
  CKBD0 U658 ( .CLK(n776), .C(n777) );
  CKBD0 U659 ( .CLK(n777), .C(n778) );
  CKBD0 U660 ( .CLK(n778), .C(n779) );
  CKBD0 U661 ( .CLK(n779), .C(n780) );
  CKBD0 U662 ( .CLK(n780), .C(n781) );
  BUFFD0 U663 ( .I(n781), .Z(n782) );
  CKBD0 U664 ( .CLK(n782), .C(n783) );
  CKBD0 U665 ( .CLK(n783), .C(n784) );
  CKBD0 U666 ( .CLK(n784), .C(n785) );
  CKBD0 U667 ( .CLK(n785), .C(n786) );
  CKBD0 U668 ( .CLK(n786), .C(n787) );
  CKBD0 U669 ( .CLK(n787), .C(n788) );
  CKBD0 U670 ( .CLK(n788), .C(n789) );
  CKBD0 U671 ( .CLK(n789), .C(n790) );
  CKBD0 U672 ( .CLK(n790), .C(n791) );
  CKBD0 U673 ( .CLK(n791), .C(n792) );
  BUFFD0 U674 ( .I(n792), .Z(n793) );
  CKBD0 U675 ( .CLK(n793), .C(n794) );
  CKBD0 U676 ( .CLK(n794), .C(n795) );
  CKBD0 U677 ( .CLK(n795), .C(n796) );
  CKBD0 U678 ( .CLK(n796), .C(n797) );
  CKBD0 U679 ( .CLK(n797), .C(n798) );
  CKBD0 U680 ( .CLK(n798), .C(n799) );
  CKBD0 U681 ( .CLK(n799), .C(n800) );
  CKBD0 U682 ( .CLK(n800), .C(n801) );
  CKBD0 U683 ( .CLK(n801), .C(n802) );
  CKBD0 U684 ( .CLK(n802), .C(n803) );
  BUFFD0 U685 ( .I(n803), .Z(n804) );
  CKBD0 U686 ( .CLK(n804), .C(n805) );
  CKBD0 U687 ( .CLK(n805), .C(n806) );
  CKBD0 U688 ( .CLK(n806), .C(n807) );
  CKBD0 U689 ( .CLK(n807), .C(n808) );
  CKBD0 U690 ( .CLK(n808), .C(n809) );
  CKBD0 U691 ( .CLK(n809), .C(n810) );
  CKBD0 U692 ( .CLK(n810), .C(n811) );
  BUFFD0 U693 ( .I(n8963), .Z(n812) );
  CKBD0 U694 ( .CLK(FrameSR[54]), .C(n813) );
  BUFFD0 U695 ( .I(n813), .Z(n814) );
  CKBD0 U696 ( .CLK(n814), .C(n815) );
  CKBD0 U697 ( .CLK(n815), .C(n816) );
  CKBD0 U698 ( .CLK(n816), .C(n817) );
  CKBD0 U699 ( .CLK(n817), .C(n818) );
  CKBD0 U700 ( .CLK(n818), .C(n819) );
  CKBD0 U701 ( .CLK(n819), .C(n820) );
  CKBD0 U702 ( .CLK(n820), .C(n821) );
  CKBD0 U703 ( .CLK(n821), .C(n822) );
  CKBD0 U704 ( .CLK(n822), .C(n823) );
  CKBD0 U705 ( .CLK(n823), .C(n824) );
  BUFFD0 U706 ( .I(n824), .Z(n825) );
  CKBD0 U707 ( .CLK(n825), .C(n826) );
  CKBD0 U708 ( .CLK(n826), .C(n827) );
  CKBD0 U709 ( .CLK(n827), .C(n828) );
  CKBD0 U710 ( .CLK(n828), .C(n829) );
  CKBD0 U711 ( .CLK(n829), .C(n830) );
  CKBD0 U712 ( .CLK(n830), .C(n831) );
  CKBD0 U713 ( .CLK(n831), .C(n832) );
  CKBD0 U714 ( .CLK(n832), .C(n833) );
  CKBD0 U715 ( .CLK(n833), .C(n834) );
  CKBD0 U716 ( .CLK(n834), .C(n835) );
  BUFFD0 U717 ( .I(n835), .Z(n836) );
  CKBD0 U718 ( .CLK(n836), .C(n837) );
  CKBD0 U719 ( .CLK(n837), .C(n838) );
  CKBD0 U720 ( .CLK(n838), .C(n839) );
  CKBD0 U721 ( .CLK(n839), .C(n840) );
  CKBD0 U722 ( .CLK(n840), .C(n841) );
  CKBD0 U723 ( .CLK(n841), .C(n842) );
  CKBD0 U724 ( .CLK(n842), .C(n843) );
  CKBD0 U725 ( .CLK(n843), .C(n844) );
  CKBD0 U726 ( .CLK(n844), .C(n845) );
  CKBD0 U727 ( .CLK(n845), .C(n846) );
  BUFFD0 U728 ( .I(n846), .Z(n847) );
  CKBD0 U729 ( .CLK(n847), .C(n848) );
  CKBD0 U730 ( .CLK(n848), .C(n849) );
  CKBD0 U731 ( .CLK(n849), .C(n850) );
  CKBD0 U732 ( .CLK(n850), .C(n851) );
  CKBD0 U733 ( .CLK(n851), .C(n852) );
  CKBD0 U734 ( .CLK(n852), .C(n853) );
  CKBD0 U735 ( .CLK(n853), .C(n854) );
  CKBD0 U736 ( .CLK(n854), .C(n855) );
  CKBD0 U737 ( .CLK(n855), .C(n856) );
  BUFFD0 U738 ( .I(n856), .Z(n857) );
  CKBD0 U739 ( .CLK(n857), .C(n858) );
  CKBD0 U740 ( .CLK(n858), .C(n859) );
  CKBD0 U741 ( .CLK(n859), .C(n860) );
  CKBD0 U742 ( .CLK(n860), .C(n861) );
  CKBD0 U743 ( .CLK(n861), .C(n862) );
  CKBD0 U744 ( .CLK(n862), .C(n863) );
  CKBD0 U745 ( .CLK(n863), .C(n864) );
  CKBD0 U746 ( .CLK(n864), .C(n865) );
  CKBD0 U747 ( .CLK(n865), .C(n866) );
  CKBD0 U748 ( .CLK(n866), .C(n867) );
  BUFFD0 U749 ( .I(n867), .Z(n868) );
  CKBD0 U750 ( .CLK(n868), .C(n869) );
  CKBD0 U751 ( .CLK(n869), .C(n870) );
  CKBD0 U752 ( .CLK(n870), .C(n871) );
  CKBD0 U753 ( .CLK(n871), .C(n872) );
  CKBD0 U754 ( .CLK(n872), .C(n873) );
  CKBD0 U755 ( .CLK(n873), .C(n874) );
  CKBD0 U756 ( .CLK(n874), .C(n875) );
  CKBD0 U757 ( .CLK(n875), .C(n876) );
  CKBD0 U758 ( .CLK(n876), .C(n877) );
  CKBD0 U759 ( .CLK(n877), .C(n878) );
  BUFFD0 U760 ( .I(n878), .Z(n879) );
  CKBD0 U761 ( .CLK(n879), .C(n880) );
  CKBD0 U762 ( .CLK(n880), .C(n881) );
  CKBD0 U763 ( .CLK(n881), .C(n882) );
  CKBD0 U764 ( .CLK(n882), .C(n883) );
  CKBD0 U765 ( .CLK(n883), .C(n884) );
  CKBD0 U766 ( .CLK(n884), .C(n885) );
  CKBD0 U767 ( .CLK(n885), .C(n886) );
  CKBD0 U768 ( .CLK(n886), .C(n887) );
  CKBD0 U769 ( .CLK(n887), .C(n888) );
  CKBD0 U770 ( .CLK(n888), .C(n889) );
  BUFFD0 U771 ( .I(n889), .Z(n890) );
  CKBD0 U772 ( .CLK(n890), .C(n891) );
  CKBD0 U773 ( .CLK(n891), .C(n892) );
  CKBD0 U774 ( .CLK(n892), .C(n893) );
  CKBD0 U775 ( .CLK(n893), .C(n894) );
  CKBD0 U776 ( .CLK(n894), .C(n895) );
  CKBD0 U777 ( .CLK(n895), .C(n896) );
  CKBD0 U778 ( .CLK(n896), .C(n897) );
  CKBD0 U779 ( .CLK(n897), .C(n898) );
  CKBD0 U780 ( .CLK(n898), .C(n899) );
  CKBD0 U781 ( .CLK(n899), .C(n900) );
  BUFFD0 U782 ( .I(n900), .Z(n901) );
  CKBD0 U783 ( .CLK(n901), .C(n902) );
  CKBD0 U784 ( .CLK(n902), .C(n903) );
  CKBD0 U785 ( .CLK(n903), .C(n904) );
  CKBD0 U786 ( .CLK(n904), .C(n905) );
  CKBD0 U787 ( .CLK(n905), .C(n906) );
  CKBD0 U788 ( .CLK(n906), .C(n907) );
  CKBD0 U789 ( .CLK(n907), .C(n908) );
  BUFFD0 U790 ( .I(n9016), .Z(n909) );
  CKBD0 U791 ( .CLK(FrameSR[7]), .C(n910) );
  BUFFD0 U792 ( .I(n910), .Z(n911) );
  BUFFD0 U793 ( .I(n6891), .Z(n912) );
  CKBD0 U794 ( .CLK(FrameSR[8]), .C(n913) );
  BUFFD0 U795 ( .I(n6754), .Z(n914) );
  CKBD0 U796 ( .CLK(FrameSR[9]), .C(n915) );
  BUFFD0 U797 ( .I(n6617), .Z(n916) );
  CKBD0 U798 ( .CLK(FrameSR[10]), .C(n917) );
  BUFFD0 U799 ( .I(n6480), .Z(n918) );
  CKBD0 U800 ( .CLK(FrameSR[11]), .C(n919) );
  BUFFD0 U801 ( .I(n6343), .Z(n920) );
  CKBD0 U802 ( .CLK(FrameSR[12]), .C(n921) );
  BUFFD0 U803 ( .I(n6206), .Z(n922) );
  CKBD0 U804 ( .CLK(FrameSR[13]), .C(n923) );
  BUFFD0 U805 ( .I(n6069), .Z(n924) );
  CKBD0 U806 ( .CLK(FrameSR[14]), .C(n925) );
  BUFFD0 U807 ( .I(n9007), .Z(n926) );
  CKBD0 U808 ( .CLK(FrameSR[18]), .C(n927) );
  CKBD0 U809 ( .CLK(n927), .C(n928) );
  BUFFD0 U810 ( .I(n928), .Z(n929) );
  CKBD0 U811 ( .CLK(n929), .C(n930) );
  CKBD0 U812 ( .CLK(n930), .C(n931) );
  CKBD0 U813 ( .CLK(n931), .C(n932) );
  CKBD0 U814 ( .CLK(n932), .C(n933) );
  CKBD0 U815 ( .CLK(n933), .C(n934) );
  CKBD0 U816 ( .CLK(n934), .C(n935) );
  CKBD0 U817 ( .CLK(n935), .C(n936) );
  CKBD0 U818 ( .CLK(n936), .C(n937) );
  CKBD0 U819 ( .CLK(n937), .C(n938) );
  CKBD0 U820 ( .CLK(n938), .C(n939) );
  BUFFD0 U821 ( .I(n939), .Z(n940) );
  CKBD0 U822 ( .CLK(n940), .C(n941) );
  CKBD0 U823 ( .CLK(n941), .C(n942) );
  CKBD0 U824 ( .CLK(n942), .C(n943) );
  CKBD0 U825 ( .CLK(n943), .C(n944) );
  CKBD0 U826 ( .CLK(n944), .C(n945) );
  CKBD0 U827 ( .CLK(n945), .C(n946) );
  CKBD0 U828 ( .CLK(n946), .C(n947) );
  CKBD0 U829 ( .CLK(n947), .C(n948) );
  CKBD0 U830 ( .CLK(n948), .C(n949) );
  BUFFD0 U831 ( .I(n949), .Z(n950) );
  CKBD0 U832 ( .CLK(n950), .C(n951) );
  CKBD0 U833 ( .CLK(n951), .C(n952) );
  CKBD0 U834 ( .CLK(n952), .C(n953) );
  CKBD0 U835 ( .CLK(n953), .C(n954) );
  CKBD0 U836 ( .CLK(n954), .C(n955) );
  CKBD0 U837 ( .CLK(n955), .C(n956) );
  CKBD0 U838 ( .CLK(n956), .C(n957) );
  CKBD0 U839 ( .CLK(n957), .C(n958) );
  CKBD0 U840 ( .CLK(n958), .C(n959) );
  CKBD0 U841 ( .CLK(n959), .C(n960) );
  BUFFD0 U842 ( .I(n960), .Z(n961) );
  CKBD0 U843 ( .CLK(n961), .C(n962) );
  CKBD0 U844 ( .CLK(n962), .C(n963) );
  CKBD0 U845 ( .CLK(n963), .C(n964) );
  CKBD0 U846 ( .CLK(n964), .C(n965) );
  CKBD0 U847 ( .CLK(n965), .C(n966) );
  CKBD0 U848 ( .CLK(n966), .C(n967) );
  CKBD0 U849 ( .CLK(n967), .C(n968) );
  CKBD0 U850 ( .CLK(n968), .C(n969) );
  CKBD0 U851 ( .CLK(n969), .C(n970) );
  CKBD0 U852 ( .CLK(n970), .C(n971) );
  BUFFD0 U853 ( .I(n971), .Z(n972) );
  CKBD0 U854 ( .CLK(n972), .C(n973) );
  CKBD0 U855 ( .CLK(n973), .C(n974) );
  CKBD0 U856 ( .CLK(n974), .C(n975) );
  CKBD0 U857 ( .CLK(n975), .C(n976) );
  CKBD0 U858 ( .CLK(n976), .C(n977) );
  CKBD0 U859 ( .CLK(n977), .C(n978) );
  CKBD0 U860 ( .CLK(n978), .C(n979) );
  CKBD0 U861 ( .CLK(n979), .C(n980) );
  CKBD0 U862 ( .CLK(n980), .C(n981) );
  CKBD0 U863 ( .CLK(n981), .C(n982) );
  BUFFD0 U864 ( .I(n982), .Z(n983) );
  CKBD0 U865 ( .CLK(n983), .C(n984) );
  CKBD0 U866 ( .CLK(n984), .C(n985) );
  CKBD0 U867 ( .CLK(n985), .C(n986) );
  CKBD0 U868 ( .CLK(n986), .C(n987) );
  CKBD0 U869 ( .CLK(n987), .C(n988) );
  CKBD0 U870 ( .CLK(n988), .C(n989) );
  CKBD0 U871 ( .CLK(n989), .C(n990) );
  CKBD0 U872 ( .CLK(n990), .C(n991) );
  CKBD0 U873 ( .CLK(n991), .C(n992) );
  CKBD0 U874 ( .CLK(n992), .C(n993) );
  BUFFD0 U875 ( .I(n993), .Z(n994) );
  CKBD0 U876 ( .CLK(n994), .C(n995) );
  CKBD0 U877 ( .CLK(n995), .C(n996) );
  CKBD0 U878 ( .CLK(n996), .C(n997) );
  CKBD0 U879 ( .CLK(n997), .C(n998) );
  CKBD0 U880 ( .CLK(n998), .C(n999) );
  CKBD0 U881 ( .CLK(n999), .C(n1000) );
  CKBD0 U882 ( .CLK(n1000), .C(n1001) );
  CKBD0 U883 ( .CLK(n1001), .C(n1002) );
  CKBD0 U884 ( .CLK(n1002), .C(n1003) );
  CKBD0 U885 ( .CLK(n1003), .C(n1004) );
  BUFFD0 U886 ( .I(n1004), .Z(n1005) );
  CKBD0 U887 ( .CLK(n1005), .C(n1006) );
  CKBD0 U888 ( .CLK(n1006), .C(n1007) );
  CKBD0 U889 ( .CLK(n1007), .C(n1008) );
  CKBD0 U890 ( .CLK(n1008), .C(n1009) );
  CKBD0 U891 ( .CLK(n1009), .C(n1010) );
  CKBD0 U892 ( .CLK(n1010), .C(n1011) );
  CKBD0 U893 ( .CLK(n1011), .C(n1012) );
  CKBD0 U894 ( .CLK(n1012), .C(n1013) );
  CKBD0 U895 ( .CLK(n1013), .C(n1014) );
  CKBD0 U896 ( .CLK(n1014), .C(n1015) );
  BUFFD0 U897 ( .I(n1015), .Z(n1016) );
  CKBD0 U898 ( .CLK(n1016), .C(n1017) );
  CKBD0 U899 ( .CLK(n1017), .C(n1018) );
  CKBD0 U900 ( .CLK(n1018), .C(n1019) );
  CKBD0 U901 ( .CLK(n1019), .C(n1020) );
  CKBD0 U902 ( .CLK(n1020), .C(n1021) );
  BUFFD0 U903 ( .I(n8970), .Z(n1022) );
  CKBD0 U904 ( .CLK(FrameSR[23]), .C(n1023) );
  BUFFD0 U905 ( .I(n1023), .Z(n1024) );
  CKBD0 U906 ( .CLK(n1024), .C(n1025) );
  CKBD0 U907 ( .CLK(n1025), .C(n1026) );
  CKBD0 U908 ( .CLK(n1026), .C(n1027) );
  CKBD0 U909 ( .CLK(n1027), .C(n1028) );
  CKBD0 U910 ( .CLK(n1028), .C(n1029) );
  CKBD0 U911 ( .CLK(n1029), .C(n1030) );
  CKBD0 U912 ( .CLK(n1030), .C(n1031) );
  CKBD0 U913 ( .CLK(n1031), .C(n1032) );
  CKBD0 U914 ( .CLK(n1032), .C(n1033) );
  CKBD0 U915 ( .CLK(n1033), .C(n1034) );
  BUFFD0 U916 ( .I(n1034), .Z(n1035) );
  CKBD0 U917 ( .CLK(n1035), .C(n1036) );
  CKBD0 U918 ( .CLK(n1036), .C(n1037) );
  CKBD0 U919 ( .CLK(n1037), .C(n1038) );
  CKBD0 U920 ( .CLK(n1038), .C(n1039) );
  CKBD0 U921 ( .CLK(n1039), .C(n1040) );
  CKBD0 U922 ( .CLK(n1040), .C(n1041) );
  CKBD0 U923 ( .CLK(n1041), .C(n1042) );
  CKBD0 U924 ( .CLK(n1042), .C(n1043) );
  CKBD0 U925 ( .CLK(n1043), .C(n1044) );
  CKBD0 U926 ( .CLK(n1044), .C(n1045) );
  BUFFD0 U927 ( .I(n1045), .Z(n1046) );
  CKBD0 U928 ( .CLK(n1046), .C(n1047) );
  CKBD0 U929 ( .CLK(n1047), .C(n1048) );
  CKBD0 U930 ( .CLK(n1048), .C(n1049) );
  CKBD0 U931 ( .CLK(n1049), .C(n1050) );
  CKBD0 U932 ( .CLK(n1050), .C(n1051) );
  CKBD0 U933 ( .CLK(n1051), .C(n1052) );
  CKBD0 U934 ( .CLK(n1052), .C(n1053) );
  CKBD0 U935 ( .CLK(n1053), .C(n1054) );
  CKBD0 U936 ( .CLK(n1054), .C(n1055) );
  CKBD0 U937 ( .CLK(n1055), .C(n1056) );
  BUFFD0 U938 ( .I(n1056), .Z(n1057) );
  CKBD0 U939 ( .CLK(n1057), .C(n1058) );
  CKBD0 U940 ( .CLK(n1058), .C(n1059) );
  CKBD0 U941 ( .CLK(n1059), .C(n1060) );
  CKBD0 U942 ( .CLK(n1060), .C(n1061) );
  CKBD0 U943 ( .CLK(n1061), .C(n1062) );
  CKBD0 U944 ( .CLK(n1062), .C(n1063) );
  CKBD0 U945 ( .CLK(n1063), .C(n1064) );
  CKBD0 U946 ( .CLK(n1064), .C(n1065) );
  CKBD0 U947 ( .CLK(n1065), .C(n1066) );
  BUFFD0 U948 ( .I(n1066), .Z(n1067) );
  CKBD0 U949 ( .CLK(n1067), .C(n1068) );
  CKBD0 U950 ( .CLK(n1068), .C(n1069) );
  CKBD0 U951 ( .CLK(n1069), .C(n1070) );
  CKBD0 U952 ( .CLK(n1070), .C(n1071) );
  CKBD0 U953 ( .CLK(n1071), .C(n1072) );
  CKBD0 U954 ( .CLK(n1072), .C(n1073) );
  CKBD0 U955 ( .CLK(n1073), .C(n1074) );
  CKBD0 U956 ( .CLK(n1074), .C(n1075) );
  CKBD0 U957 ( .CLK(n1075), .C(n1076) );
  CKBD0 U958 ( .CLK(n1076), .C(n1077) );
  BUFFD0 U959 ( .I(n1077), .Z(n1078) );
  CKBD0 U960 ( .CLK(n1078), .C(n1079) );
  CKBD0 U961 ( .CLK(n1079), .C(n1080) );
  CKBD0 U962 ( .CLK(n1080), .C(n1081) );
  CKBD0 U963 ( .CLK(n1081), .C(n1082) );
  CKBD0 U964 ( .CLK(n1082), .C(n1083) );
  CKBD0 U965 ( .CLK(n1083), .C(n1084) );
  CKBD0 U966 ( .CLK(n1084), .C(n1085) );
  CKBD0 U967 ( .CLK(n1085), .C(n1086) );
  CKBD0 U968 ( .CLK(n1086), .C(n1087) );
  CKBD0 U969 ( .CLK(n1087), .C(n1088) );
  BUFFD0 U970 ( .I(n1088), .Z(n1089) );
  CKBD0 U971 ( .CLK(n1089), .C(n1090) );
  CKBD0 U972 ( .CLK(n1090), .C(n1091) );
  CKBD0 U973 ( .CLK(n1091), .C(n1092) );
  CKBD0 U974 ( .CLK(n1092), .C(n1093) );
  CKBD0 U975 ( .CLK(n1093), .C(n1094) );
  CKBD0 U976 ( .CLK(n1094), .C(n1095) );
  CKBD0 U977 ( .CLK(n1095), .C(n1096) );
  CKBD0 U978 ( .CLK(n1096), .C(n1097) );
  CKBD0 U979 ( .CLK(n1097), .C(n1098) );
  CKBD0 U980 ( .CLK(n1098), .C(n1099) );
  BUFFD0 U981 ( .I(n1099), .Z(n1100) );
  CKBD0 U982 ( .CLK(n1100), .C(n1101) );
  CKBD0 U983 ( .CLK(n1101), .C(n1102) );
  CKBD0 U984 ( .CLK(n1102), .C(n1103) );
  CKBD0 U985 ( .CLK(n1103), .C(n1104) );
  CKBD0 U986 ( .CLK(n1104), .C(n1105) );
  CKBD0 U987 ( .CLK(n1105), .C(n1106) );
  CKBD0 U988 ( .CLK(n1106), .C(n1107) );
  CKBD0 U989 ( .CLK(n1107), .C(n1108) );
  CKBD0 U990 ( .CLK(n1108), .C(n1109) );
  CKBD0 U991 ( .CLK(n1109), .C(n1110) );
  BUFFD0 U992 ( .I(n1110), .Z(n1111) );
  CKBD0 U993 ( .CLK(n1111), .C(n1112) );
  CKBD0 U994 ( .CLK(n1112), .C(n1113) );
  CKBD0 U995 ( .CLK(n1113), .C(n1114) );
  CKBD0 U996 ( .CLK(n1114), .C(n1115) );
  CKBD0 U997 ( .CLK(n1115), .C(n1116) );
  CKBD0 U998 ( .CLK(n1116), .C(n1117) );
  CKBD0 U999 ( .CLK(n1117), .C(n1118) );
  BUFFD0 U1000 ( .I(n5796), .Z(n1119) );
  CKBD0 U1001 ( .CLK(FrameSR[24]), .C(n1120) );
  BUFFD0 U1002 ( .I(n5659), .Z(n1121) );
  CKBD0 U1003 ( .CLK(FrameSR[25]), .C(n1122) );
  BUFFD0 U1004 ( .I(n5522), .Z(n1123) );
  CKBD0 U1005 ( .CLK(FrameSR[26]), .C(n1124) );
  BUFFD0 U1006 ( .I(n5386), .Z(n1125) );
  CKBD0 U1007 ( .CLK(FrameSR[27]), .C(n1126) );
  BUFFD0 U1008 ( .I(n5250), .Z(n1127) );
  CKBD0 U1009 ( .CLK(FrameSR[28]), .C(n1128) );
  BUFFD0 U1010 ( .I(n5114), .Z(n1129) );
  CKBD0 U1011 ( .CLK(FrameSR[29]), .C(n1130) );
  BUFFD0 U1012 ( .I(n4978), .Z(n1131) );
  CKBD0 U1013 ( .CLK(FrameSR[30]), .C(n1132) );
  BUFFD0 U1014 ( .I(n8962), .Z(n1133) );
  CKBD0 U1015 ( .CLK(FrameSR[39]), .C(n1134) );
  BUFFD0 U1016 ( .I(n1134), .Z(n1135) );
  CKBD0 U1017 ( .CLK(n1135), .C(n1136) );
  CKBD0 U1018 ( .CLK(n1136), .C(n1137) );
  CKBD0 U1019 ( .CLK(n1137), .C(n1138) );
  CKBD0 U1020 ( .CLK(n1138), .C(n1139) );
  CKBD0 U1021 ( .CLK(n1139), .C(n1140) );
  CKBD0 U1022 ( .CLK(n1140), .C(n1141) );
  CKBD0 U1023 ( .CLK(n1141), .C(n1142) );
  CKBD0 U1024 ( .CLK(n1142), .C(n1143) );
  CKBD0 U1025 ( .CLK(n1143), .C(n1144) );
  BUFFD0 U1026 ( .I(n1144), .Z(n1145) );
  CKBD0 U1027 ( .CLK(n1145), .C(n1146) );
  CKBD0 U1028 ( .CLK(n1146), .C(n1147) );
  CKBD0 U1029 ( .CLK(n1147), .C(n1148) );
  CKBD0 U1030 ( .CLK(n1148), .C(n1149) );
  CKBD0 U1031 ( .CLK(n1149), .C(n1150) );
  CKBD0 U1032 ( .CLK(n1150), .C(n1151) );
  CKBD0 U1033 ( .CLK(n1151), .C(n1152) );
  CKBD0 U1034 ( .CLK(n1152), .C(n1153) );
  CKBD0 U1035 ( .CLK(n1153), .C(n1154) );
  CKBD0 U1036 ( .CLK(n1154), .C(n1155) );
  BUFFD0 U1037 ( .I(n1155), .Z(n1156) );
  CKBD0 U1038 ( .CLK(n1156), .C(n1157) );
  CKBD0 U1039 ( .CLK(n1157), .C(n1158) );
  CKBD0 U1040 ( .CLK(n1158), .C(n1159) );
  CKBD0 U1041 ( .CLK(n1159), .C(n1160) );
  CKBD0 U1042 ( .CLK(n1160), .C(n1161) );
  CKBD0 U1043 ( .CLK(n1161), .C(n1162) );
  CKBD0 U1044 ( .CLK(n1162), .C(n1163) );
  CKBD0 U1045 ( .CLK(n1163), .C(n1164) );
  CKBD0 U1046 ( .CLK(n1164), .C(n1165) );
  CKBD0 U1047 ( .CLK(n1165), .C(n1166) );
  BUFFD0 U1048 ( .I(n1166), .Z(n1167) );
  CKBD0 U1049 ( .CLK(n1167), .C(n1168) );
  CKBD0 U1050 ( .CLK(n1168), .C(n1169) );
  CKBD0 U1051 ( .CLK(n1169), .C(n1170) );
  CKBD0 U1052 ( .CLK(n1170), .C(n1171) );
  CKBD0 U1053 ( .CLK(n1171), .C(n1172) );
  CKBD0 U1054 ( .CLK(n1172), .C(n1173) );
  CKBD0 U1055 ( .CLK(n1173), .C(n1174) );
  CKBD0 U1056 ( .CLK(n1174), .C(n1175) );
  CKBD0 U1057 ( .CLK(n1175), .C(n1176) );
  CKBD0 U1058 ( .CLK(n1176), .C(n1177) );
  BUFFD0 U1059 ( .I(n1177), .Z(n1178) );
  CKBD0 U1060 ( .CLK(n1178), .C(n1179) );
  CKBD0 U1061 ( .CLK(n1179), .C(n1180) );
  CKBD0 U1062 ( .CLK(n1180), .C(n1181) );
  CKBD0 U1063 ( .CLK(n1181), .C(n1182) );
  CKBD0 U1064 ( .CLK(n1182), .C(n1183) );
  CKBD0 U1065 ( .CLK(n1183), .C(n1184) );
  CKBD0 U1066 ( .CLK(n1184), .C(n1185) );
  CKBD0 U1067 ( .CLK(n1185), .C(n1186) );
  CKBD0 U1068 ( .CLK(n1186), .C(n1187) );
  CKBD0 U1069 ( .CLK(n1187), .C(n1188) );
  BUFFD0 U1070 ( .I(n1188), .Z(n1189) );
  CKBD0 U1071 ( .CLK(n1189), .C(n1190) );
  CKBD0 U1072 ( .CLK(n1190), .C(n1191) );
  CKBD0 U1073 ( .CLK(n1191), .C(n1192) );
  CKBD0 U1074 ( .CLK(n1192), .C(n1193) );
  CKBD0 U1075 ( .CLK(n1193), .C(n1194) );
  CKBD0 U1076 ( .CLK(n1194), .C(n1195) );
  CKBD0 U1077 ( .CLK(n1195), .C(n1196) );
  CKBD0 U1078 ( .CLK(n1196), .C(n1197) );
  CKBD0 U1079 ( .CLK(n1197), .C(n1198) );
  CKBD0 U1080 ( .CLK(n1198), .C(n1199) );
  BUFFD0 U1081 ( .I(n1199), .Z(n1200) );
  CKBD0 U1082 ( .CLK(n1200), .C(n1201) );
  CKBD0 U1083 ( .CLK(n1201), .C(n1202) );
  CKBD0 U1084 ( .CLK(n1202), .C(n1203) );
  CKBD0 U1085 ( .CLK(n1203), .C(n1204) );
  CKBD0 U1086 ( .CLK(n1204), .C(n1205) );
  CKBD0 U1087 ( .CLK(n1205), .C(n1206) );
  CKBD0 U1088 ( .CLK(n1206), .C(n1207) );
  CKBD0 U1089 ( .CLK(n1207), .C(n1208) );
  CKBD0 U1090 ( .CLK(n1208), .C(n1209) );
  CKBD0 U1091 ( .CLK(n1209), .C(n1210) );
  BUFFD0 U1092 ( .I(n1210), .Z(n1211) );
  CKBD0 U1093 ( .CLK(n1211), .C(n1212) );
  CKBD0 U1094 ( .CLK(n1212), .C(n1213) );
  CKBD0 U1095 ( .CLK(n1213), .C(n1214) );
  CKBD0 U1096 ( .CLK(n1214), .C(n1215) );
  CKBD0 U1097 ( .CLK(n1215), .C(n1216) );
  CKBD0 U1098 ( .CLK(n1216), .C(n1217) );
  CKBD0 U1099 ( .CLK(n1217), .C(n1218) );
  CKBD0 U1100 ( .CLK(n1218), .C(n1219) );
  CKBD0 U1101 ( .CLK(n1219), .C(n1220) );
  BUFFD0 U1102 ( .I(n1220), .Z(n1221) );
  CKBD0 U1103 ( .CLK(n1221), .C(n1222) );
  CKBD0 U1104 ( .CLK(n1222), .C(n1223) );
  CKBD0 U1105 ( .CLK(n1223), .C(n1224) );
  CKBD0 U1106 ( .CLK(n1224), .C(n1225) );
  CKBD0 U1107 ( .CLK(n1225), .C(n1226) );
  CKBD0 U1108 ( .CLK(n1226), .C(n1227) );
  CKBD0 U1109 ( .CLK(n1227), .C(n1228) );
  CKBD0 U1110 ( .CLK(n1228), .C(n1229) );
  BUFFD0 U1111 ( .I(n4706), .Z(n1230) );
  CKBD0 U1112 ( .CLK(FrameSR[40]), .C(n1231) );
  BUFFD0 U1113 ( .I(n4570), .Z(n1232) );
  CKBD0 U1114 ( .CLK(FrameSR[41]), .C(n1233) );
  BUFFD0 U1115 ( .I(n4434), .Z(n1234) );
  CKBD0 U1116 ( .CLK(FrameSR[42]), .C(n1235) );
  BUFFD0 U1117 ( .I(n4298), .Z(n1236) );
  CKBD0 U1118 ( .CLK(FrameSR[43]), .C(n1237) );
  BUFFD0 U1119 ( .I(n4162), .Z(n1238) );
  CKBD0 U1120 ( .CLK(FrameSR[44]), .C(n1239) );
  BUFFD0 U1121 ( .I(n4026), .Z(n1240) );
  CKBD0 U1122 ( .CLK(FrameSR[45]), .C(n1241) );
  BUFFD0 U1123 ( .I(n3890), .Z(n1242) );
  CKBD0 U1124 ( .CLK(FrameSR[46]), .C(n1243) );
  BUFFD0 U1125 ( .I(n8960), .Z(n1244) );
  CKBD0 U1126 ( .CLK(FrameSR[55]), .C(n1245) );
  BUFFD0 U1127 ( .I(n1245), .Z(n1246) );
  CKBD0 U1128 ( .CLK(n1246), .C(n1247) );
  CKBD0 U1129 ( .CLK(n1247), .C(n1248) );
  CKBD0 U1130 ( .CLK(n1248), .C(n1249) );
  CKBD0 U1131 ( .CLK(n1249), .C(n1250) );
  CKBD0 U1132 ( .CLK(n1250), .C(n1251) );
  CKBD0 U1133 ( .CLK(n1251), .C(n1252) );
  CKBD0 U1134 ( .CLK(n1252), .C(n1253) );
  CKBD0 U1135 ( .CLK(n1253), .C(n1254) );
  CKBD0 U1136 ( .CLK(n1254), .C(n1255) );
  BUFFD0 U1137 ( .I(n1255), .Z(n1256) );
  CKBD0 U1138 ( .CLK(n1256), .C(n1257) );
  CKBD0 U1139 ( .CLK(n1257), .C(n1258) );
  CKBD0 U1140 ( .CLK(n1258), .C(n1259) );
  CKBD0 U1141 ( .CLK(n1259), .C(n1260) );
  CKBD0 U1142 ( .CLK(n1260), .C(n1261) );
  CKBD0 U1143 ( .CLK(n1261), .C(n1262) );
  CKBD0 U1144 ( .CLK(n1262), .C(n1263) );
  CKBD0 U1145 ( .CLK(n1263), .C(n1264) );
  CKBD0 U1146 ( .CLK(n1264), .C(n1265) );
  CKBD0 U1147 ( .CLK(n1265), .C(n1266) );
  BUFFD0 U1148 ( .I(n1266), .Z(n1267) );
  CKBD0 U1149 ( .CLK(n1267), .C(n1268) );
  CKBD0 U1150 ( .CLK(n1268), .C(n1269) );
  CKBD0 U1151 ( .CLK(n1269), .C(n1270) );
  CKBD0 U1152 ( .CLK(n1270), .C(n1271) );
  CKBD0 U1153 ( .CLK(n1271), .C(n1272) );
  CKBD0 U1154 ( .CLK(n1272), .C(n1273) );
  CKBD0 U1155 ( .CLK(n1273), .C(n1274) );
  CKBD0 U1156 ( .CLK(n1274), .C(n1275) );
  CKBD0 U1157 ( .CLK(n1275), .C(n1276) );
  CKBD0 U1158 ( .CLK(n1276), .C(n1277) );
  BUFFD0 U1159 ( .I(n1277), .Z(n1278) );
  CKBD0 U1160 ( .CLK(n1278), .C(n1279) );
  CKBD0 U1161 ( .CLK(n1279), .C(n1280) );
  CKBD0 U1162 ( .CLK(n1280), .C(n1281) );
  CKBD0 U1163 ( .CLK(n1281), .C(n1282) );
  CKBD0 U1164 ( .CLK(n1282), .C(n1283) );
  CKBD0 U1165 ( .CLK(n1283), .C(n1284) );
  CKBD0 U1166 ( .CLK(n1284), .C(n1285) );
  CKBD0 U1167 ( .CLK(n1285), .C(n1286) );
  CKBD0 U1168 ( .CLK(n1286), .C(n1287) );
  CKBD0 U1169 ( .CLK(n1287), .C(n1288) );
  BUFFD0 U1170 ( .I(n1288), .Z(n1289) );
  CKBD0 U1171 ( .CLK(n1289), .C(n1290) );
  CKBD0 U1172 ( .CLK(n1290), .C(n1291) );
  CKBD0 U1173 ( .CLK(n1291), .C(n1292) );
  CKBD0 U1174 ( .CLK(n1292), .C(n1293) );
  CKBD0 U1175 ( .CLK(n1293), .C(n1294) );
  CKBD0 U1176 ( .CLK(n1294), .C(n1295) );
  CKBD0 U1177 ( .CLK(n1295), .C(n1296) );
  CKBD0 U1178 ( .CLK(n1296), .C(n1297) );
  CKBD0 U1179 ( .CLK(n1297), .C(n1298) );
  CKBD0 U1180 ( .CLK(n1298), .C(n1299) );
  BUFFD0 U1181 ( .I(n1299), .Z(n1300) );
  CKBD0 U1182 ( .CLK(n1300), .C(n1301) );
  CKBD0 U1183 ( .CLK(n1301), .C(n1302) );
  CKBD0 U1184 ( .CLK(n1302), .C(n1303) );
  CKBD0 U1185 ( .CLK(n1303), .C(n1304) );
  CKBD0 U1186 ( .CLK(n1304), .C(n1305) );
  CKBD0 U1187 ( .CLK(n1305), .C(n1306) );
  CKBD0 U1188 ( .CLK(n1306), .C(n1307) );
  CKBD0 U1189 ( .CLK(n1307), .C(n1308) );
  CKBD0 U1190 ( .CLK(n1308), .C(n1309) );
  CKBD0 U1191 ( .CLK(n1309), .C(n1310) );
  BUFFD0 U1192 ( .I(n1310), .Z(n1311) );
  CKBD0 U1193 ( .CLK(n1311), .C(n1312) );
  CKBD0 U1194 ( .CLK(n1312), .C(n1313) );
  CKBD0 U1195 ( .CLK(n1313), .C(n1314) );
  CKBD0 U1196 ( .CLK(n1314), .C(n1315) );
  CKBD0 U1197 ( .CLK(n1315), .C(n1316) );
  CKBD0 U1198 ( .CLK(n1316), .C(n1317) );
  CKBD0 U1199 ( .CLK(n1317), .C(n1318) );
  CKBD0 U1200 ( .CLK(n1318), .C(n1319) );
  CKBD0 U1201 ( .CLK(n1319), .C(n1320) );
  CKBD0 U1202 ( .CLK(n1320), .C(n1321) );
  BUFFD0 U1203 ( .I(n1321), .Z(n1322) );
  CKBD0 U1204 ( .CLK(n1322), .C(n1323) );
  CKBD0 U1205 ( .CLK(n1323), .C(n1324) );
  CKBD0 U1206 ( .CLK(n1324), .C(n1325) );
  CKBD0 U1207 ( .CLK(n1325), .C(n1326) );
  CKBD0 U1208 ( .CLK(n1326), .C(n1327) );
  CKBD0 U1209 ( .CLK(n1327), .C(n1328) );
  CKBD0 U1210 ( .CLK(n1328), .C(n1329) );
  CKBD0 U1211 ( .CLK(n1329), .C(n1330) );
  CKBD0 U1212 ( .CLK(n1330), .C(n1331) );
  BUFFD0 U1213 ( .I(n1331), .Z(n1332) );
  CKBD0 U1214 ( .CLK(n1332), .C(n1333) );
  CKBD0 U1215 ( .CLK(n1333), .C(n1334) );
  CKBD0 U1216 ( .CLK(n1334), .C(n1335) );
  CKBD0 U1217 ( .CLK(n1335), .C(n1336) );
  CKBD0 U1218 ( .CLK(n1336), .C(n1337) );
  CKBD0 U1219 ( .CLK(n1337), .C(n1338) );
  CKBD0 U1220 ( .CLK(n1338), .C(n1339) );
  CKBD0 U1221 ( .CLK(n1339), .C(n1340) );
  BUFFD0 U1222 ( .I(n3618), .Z(n1341) );
  CKBD0 U1223 ( .CLK(FrameSR[56]), .C(n1342) );
  BUFFD0 U1224 ( .I(n3482), .Z(n1343) );
  CKBD0 U1225 ( .CLK(FrameSR[57]), .C(n1344) );
  BUFFD0 U1226 ( .I(n3346), .Z(n1345) );
  CKBD0 U1227 ( .CLK(FrameSR[58]), .C(n1346) );
  BUFFD0 U1228 ( .I(n3210), .Z(n1347) );
  CKBD0 U1229 ( .CLK(FrameSR[59]), .C(n1348) );
  BUFFD0 U1230 ( .I(n3074), .Z(n1349) );
  CKBD0 U1231 ( .CLK(FrameSR[60]), .C(n1350) );
  BUFFD0 U1232 ( .I(n2938), .Z(n1351) );
  CKBD0 U1233 ( .CLK(FrameSR[61]), .C(n1352) );
  BUFFD0 U1234 ( .I(n9015), .Z(n1353) );
  CKBD0 U1235 ( .CLK(FrameSR[3]), .C(n1354) );
  BUFFD0 U1236 ( .I(n8982), .Z(n1355) );
  CKBD0 U1237 ( .CLK(FrameSR[19]), .C(n1356) );
  CKBD0 U1238 ( .CLK(n1356), .C(n1357) );
  BUFFD0 U1239 ( .I(n1357), .Z(n1358) );
  CKBD0 U1240 ( .CLK(n1358), .C(n1359) );
  CKBD0 U1241 ( .CLK(n1359), .C(n1360) );
  CKBD0 U1242 ( .CLK(n1360), .C(n1361) );
  CKBD0 U1243 ( .CLK(n1361), .C(n1362) );
  CKBD0 U1244 ( .CLK(n1362), .C(n1363) );
  CKBD0 U1245 ( .CLK(n1363), .C(n1364) );
  CKBD0 U1246 ( .CLK(n1364), .C(n1365) );
  CKBD0 U1247 ( .CLK(n1365), .C(n1366) );
  CKBD0 U1248 ( .CLK(n1366), .C(n1367) );
  CKBD0 U1249 ( .CLK(n1367), .C(n1368) );
  BUFFD0 U1250 ( .I(n1368), .Z(n1369) );
  CKBD0 U1251 ( .CLK(n1369), .C(n1370) );
  CKBD0 U1252 ( .CLK(n1370), .C(n1371) );
  CKBD0 U1253 ( .CLK(n1371), .C(n1372) );
  CKBD0 U1254 ( .CLK(n1372), .C(n1373) );
  CKBD0 U1255 ( .CLK(n1373), .C(n1374) );
  CKBD0 U1256 ( .CLK(n1374), .C(n1375) );
  CKBD0 U1257 ( .CLK(n1375), .C(n1376) );
  CKBD0 U1258 ( .CLK(n1376), .C(n1377) );
  CKBD0 U1259 ( .CLK(n1377), .C(n1378) );
  CKBD0 U1260 ( .CLK(n1378), .C(n1379) );
  BUFFD0 U1261 ( .I(n1379), .Z(n1380) );
  CKBD0 U1262 ( .CLK(n1380), .C(n1381) );
  CKBD0 U1263 ( .CLK(n1381), .C(n1382) );
  CKBD0 U1264 ( .CLK(n1382), .C(n1383) );
  CKBD0 U1265 ( .CLK(n1383), .C(n1384) );
  CKBD0 U1266 ( .CLK(n1384), .C(n1385) );
  CKBD0 U1267 ( .CLK(n1385), .C(n1386) );
  CKBD0 U1268 ( .CLK(n1386), .C(n1387) );
  CKBD0 U1269 ( .CLK(n1387), .C(n1388) );
  CKBD0 U1270 ( .CLK(n1388), .C(n1389) );
  CKBD0 U1271 ( .CLK(n1389), .C(n1390) );
  BUFFD0 U1272 ( .I(n1390), .Z(n1391) );
  CKBD0 U1273 ( .CLK(n1391), .C(n1392) );
  CKBD0 U1274 ( .CLK(n1392), .C(n1393) );
  CKBD0 U1275 ( .CLK(n1393), .C(n1394) );
  CKBD0 U1276 ( .CLK(n1394), .C(n1395) );
  CKBD0 U1277 ( .CLK(n1395), .C(n1396) );
  CKBD0 U1278 ( .CLK(n1396), .C(n1397) );
  CKBD0 U1279 ( .CLK(n1397), .C(n1398) );
  CKBD0 U1280 ( .CLK(n1398), .C(n1399) );
  CKBD0 U1281 ( .CLK(n1399), .C(n1400) );
  CKBD0 U1282 ( .CLK(n1400), .C(n1401) );
  BUFFD0 U1283 ( .I(n1401), .Z(n1402) );
  CKBD0 U1284 ( .CLK(n1402), .C(n1403) );
  CKBD0 U1285 ( .CLK(n1403), .C(n1404) );
  CKBD0 U1286 ( .CLK(n1404), .C(n1405) );
  CKBD0 U1287 ( .CLK(n1405), .C(n1406) );
  CKBD0 U1288 ( .CLK(n1406), .C(n1407) );
  CKBD0 U1289 ( .CLK(n1407), .C(n1408) );
  CKBD0 U1290 ( .CLK(n1408), .C(n1409) );
  CKBD0 U1291 ( .CLK(n1409), .C(n1410) );
  CKBD0 U1292 ( .CLK(n1410), .C(n1411) );
  CKBD0 U1293 ( .CLK(n1411), .C(n1412) );
  BUFFD0 U1294 ( .I(n1412), .Z(n1413) );
  CKBD0 U1295 ( .CLK(n1413), .C(n1414) );
  CKBD0 U1296 ( .CLK(n1414), .C(n1415) );
  CKBD0 U1297 ( .CLK(n1415), .C(n1416) );
  CKBD0 U1298 ( .CLK(n1416), .C(n1417) );
  CKBD0 U1299 ( .CLK(n1417), .C(n1418) );
  CKBD0 U1300 ( .CLK(n1418), .C(n1419) );
  CKBD0 U1301 ( .CLK(n1419), .C(n1420) );
  CKBD0 U1302 ( .CLK(n1420), .C(n1421) );
  CKBD0 U1303 ( .CLK(n1421), .C(n1422) );
  CKBD0 U1304 ( .CLK(n1422), .C(n1423) );
  BUFFD0 U1305 ( .I(n1423), .Z(n1424) );
  CKBD0 U1306 ( .CLK(n1424), .C(n1425) );
  CKBD0 U1307 ( .CLK(n1425), .C(n1426) );
  CKBD0 U1308 ( .CLK(n1426), .C(n1427) );
  CKBD0 U1309 ( .CLK(n1427), .C(n1428) );
  CKBD0 U1310 ( .CLK(n1428), .C(n1429) );
  CKBD0 U1311 ( .CLK(n1429), .C(n1430) );
  CKBD0 U1312 ( .CLK(n1430), .C(n1431) );
  CKBD0 U1313 ( .CLK(n1431), .C(n1432) );
  CKBD0 U1314 ( .CLK(n1432), .C(n1433) );
  BUFFD0 U1315 ( .I(n1433), .Z(n1434) );
  CKBD0 U1316 ( .CLK(n1434), .C(n1435) );
  CKBD0 U1317 ( .CLK(n1435), .C(n1436) );
  CKBD0 U1318 ( .CLK(n1436), .C(n1437) );
  CKBD0 U1319 ( .CLK(n1437), .C(n1438) );
  CKBD0 U1320 ( .CLK(n1438), .C(n1439) );
  CKBD0 U1321 ( .CLK(n1439), .C(n1440) );
  CKBD0 U1322 ( .CLK(n1440), .C(n1441) );
  CKBD0 U1323 ( .CLK(n1441), .C(n1442) );
  CKBD0 U1324 ( .CLK(n1442), .C(n1443) );
  CKBD0 U1325 ( .CLK(n1443), .C(n1444) );
  BUFFD0 U1326 ( .I(n1444), .Z(n1445) );
  CKBD0 U1327 ( .CLK(n1445), .C(n1446) );
  CKBD0 U1328 ( .CLK(n1446), .C(n1447) );
  CKBD0 U1329 ( .CLK(n1447), .C(n1448) );
  CKBD0 U1330 ( .CLK(n1448), .C(n1449) );
  CKBD0 U1331 ( .CLK(n1449), .C(n1450) );
  BUFFD0 U1332 ( .I(n8997), .Z(n1451) );
  CKBD0 U1333 ( .CLK(FrameSR[33]), .C(n1452) );
  CKBD0 U1334 ( .CLK(n1452), .C(n1453) );
  BUFFD0 U1335 ( .I(n1453), .Z(n1454) );
  CKBD0 U1336 ( .CLK(n1454), .C(n1455) );
  CKBD0 U1337 ( .CLK(n1455), .C(n1456) );
  CKBD0 U1338 ( .CLK(n1456), .C(n1457) );
  CKBD0 U1339 ( .CLK(n1457), .C(n1458) );
  CKBD0 U1340 ( .CLK(n1458), .C(n1459) );
  CKBD0 U1341 ( .CLK(n1459), .C(n1460) );
  CKBD0 U1342 ( .CLK(n1460), .C(n1461) );
  CKBD0 U1343 ( .CLK(n1461), .C(n1462) );
  CKBD0 U1344 ( .CLK(n1462), .C(n1463) );
  CKBD0 U1345 ( .CLK(n1463), .C(n1464) );
  BUFFD0 U1346 ( .I(n1464), .Z(n1465) );
  CKBD0 U1347 ( .CLK(n1465), .C(n1466) );
  CKBD0 U1348 ( .CLK(n1466), .C(n1467) );
  CKBD0 U1349 ( .CLK(n1467), .C(n1468) );
  CKBD0 U1350 ( .CLK(n1468), .C(n1469) );
  CKBD0 U1351 ( .CLK(n1469), .C(n1470) );
  CKBD0 U1352 ( .CLK(n1470), .C(n1471) );
  CKBD0 U1353 ( .CLK(n1471), .C(n1472) );
  CKBD0 U1354 ( .CLK(n1472), .C(n1473) );
  CKBD0 U1355 ( .CLK(n1473), .C(n1474) );
  BUFFD0 U1356 ( .I(n1474), .Z(n1475) );
  CKBD0 U1357 ( .CLK(n1475), .C(n1476) );
  CKBD0 U1358 ( .CLK(n1476), .C(n1477) );
  CKBD0 U1359 ( .CLK(n1477), .C(n1478) );
  CKBD0 U1360 ( .CLK(n1478), .C(n1479) );
  CKBD0 U1361 ( .CLK(n1479), .C(n1480) );
  CKBD0 U1362 ( .CLK(n1480), .C(n1481) );
  CKBD0 U1363 ( .CLK(n1481), .C(n1482) );
  CKBD0 U1364 ( .CLK(n1482), .C(n1483) );
  CKBD0 U1365 ( .CLK(n1483), .C(n1484) );
  CKBD0 U1366 ( .CLK(n1484), .C(n1485) );
  BUFFD0 U1367 ( .I(n1485), .Z(n1486) );
  CKBD0 U1368 ( .CLK(n1486), .C(n1487) );
  CKBD0 U1369 ( .CLK(n1487), .C(n1488) );
  CKBD0 U1370 ( .CLK(n1488), .C(n1489) );
  CKBD0 U1371 ( .CLK(n1489), .C(n1490) );
  CKBD0 U1372 ( .CLK(n1490), .C(n1491) );
  CKBD0 U1373 ( .CLK(n1491), .C(n1492) );
  CKBD0 U1374 ( .CLK(n1492), .C(n1493) );
  CKBD0 U1375 ( .CLK(n1493), .C(n1494) );
  CKBD0 U1376 ( .CLK(n1494), .C(n1495) );
  CKBD0 U1377 ( .CLK(n1495), .C(n1496) );
  BUFFD0 U1378 ( .I(n1496), .Z(n1497) );
  CKBD0 U1379 ( .CLK(n1497), .C(n1498) );
  CKBD0 U1380 ( .CLK(n1498), .C(n1499) );
  CKBD0 U1381 ( .CLK(n1499), .C(n1500) );
  CKBD0 U1382 ( .CLK(n1500), .C(n1501) );
  CKBD0 U1383 ( .CLK(n1501), .C(n1502) );
  CKBD0 U1384 ( .CLK(n1502), .C(n1503) );
  CKBD0 U1385 ( .CLK(n1503), .C(n1504) );
  CKBD0 U1386 ( .CLK(n1504), .C(n1505) );
  CKBD0 U1387 ( .CLK(n1505), .C(n1506) );
  CKBD0 U1388 ( .CLK(n1506), .C(n1507) );
  BUFFD0 U1389 ( .I(n1507), .Z(n1508) );
  CKBD0 U1390 ( .CLK(n1508), .C(n1509) );
  CKBD0 U1391 ( .CLK(n1509), .C(n1510) );
  CKBD0 U1392 ( .CLK(n1510), .C(n1511) );
  CKBD0 U1393 ( .CLK(n1511), .C(n1512) );
  CKBD0 U1394 ( .CLK(n1512), .C(n1513) );
  CKBD0 U1395 ( .CLK(n1513), .C(n1514) );
  CKBD0 U1396 ( .CLK(n1514), .C(n1515) );
  CKBD0 U1397 ( .CLK(n1515), .C(n1516) );
  CKBD0 U1398 ( .CLK(n1516), .C(n1517) );
  CKBD0 U1399 ( .CLK(n1517), .C(n1518) );
  BUFFD0 U1400 ( .I(n1518), .Z(n1519) );
  CKBD0 U1401 ( .CLK(n1519), .C(n1520) );
  CKBD0 U1402 ( .CLK(n1520), .C(n1521) );
  CKBD0 U1403 ( .CLK(n1521), .C(n1522) );
  CKBD0 U1404 ( .CLK(n1522), .C(n1523) );
  CKBD0 U1405 ( .CLK(n1523), .C(n1524) );
  CKBD0 U1406 ( .CLK(n1524), .C(n1525) );
  CKBD0 U1407 ( .CLK(n1525), .C(n1526) );
  CKBD0 U1408 ( .CLK(n1526), .C(n1527) );
  CKBD0 U1409 ( .CLK(n1527), .C(n1528) );
  CKBD0 U1410 ( .CLK(n1528), .C(n1529) );
  BUFFD0 U1411 ( .I(n1529), .Z(n1530) );
  CKBD0 U1412 ( .CLK(n1530), .C(n1531) );
  CKBD0 U1413 ( .CLK(n1531), .C(n1532) );
  CKBD0 U1414 ( .CLK(n1532), .C(n1533) );
  CKBD0 U1415 ( .CLK(n1533), .C(n1534) );
  CKBD0 U1416 ( .CLK(n1534), .C(n1535) );
  CKBD0 U1417 ( .CLK(n1535), .C(n1536) );
  CKBD0 U1418 ( .CLK(n1536), .C(n1537) );
  CKBD0 U1419 ( .CLK(n1537), .C(n1538) );
  CKBD0 U1420 ( .CLK(n1538), .C(n1539) );
  CKBD0 U1421 ( .CLK(n1539), .C(n1540) );
  BUFFD0 U1422 ( .I(n1540), .Z(n1541) );
  CKBD0 U1423 ( .CLK(n1541), .C(n1542) );
  CKBD0 U1424 ( .CLK(n1542), .C(n1543) );
  CKBD0 U1425 ( .CLK(n1543), .C(n1544) );
  CKBD0 U1426 ( .CLK(n1544), .C(n1545) );
  CKBD0 U1427 ( .CLK(n1545), .C(n1546) );
  BUFFD0 U1428 ( .I(n8996), .Z(n1547) );
  CKBD0 U1429 ( .CLK(FrameSR[48]), .C(n1548) );
  CKBD0 U1430 ( .CLK(n1548), .C(n1549) );
  BUFFD0 U1431 ( .I(n1549), .Z(n1550) );
  CKBD0 U1432 ( .CLK(n1550), .C(n1551) );
  CKBD0 U1433 ( .CLK(n1551), .C(n1552) );
  CKBD0 U1434 ( .CLK(n1552), .C(n1553) );
  CKBD0 U1435 ( .CLK(n1553), .C(n1554) );
  CKBD0 U1436 ( .CLK(n1554), .C(n1555) );
  CKBD0 U1437 ( .CLK(n1555), .C(n1556) );
  CKBD0 U1438 ( .CLK(n1556), .C(n1557) );
  CKBD0 U1439 ( .CLK(n1557), .C(n1558) );
  CKBD0 U1440 ( .CLK(n1558), .C(n1559) );
  CKBD0 U1441 ( .CLK(n1559), .C(n1560) );
  BUFFD0 U1442 ( .I(n1560), .Z(n1561) );
  CKBD0 U1443 ( .CLK(n1561), .C(n1562) );
  CKBD0 U1444 ( .CLK(n1562), .C(n1563) );
  CKBD0 U1445 ( .CLK(n1563), .C(n1564) );
  CKBD0 U1446 ( .CLK(n1564), .C(n1565) );
  CKBD0 U1447 ( .CLK(n1565), .C(n1566) );
  CKBD0 U1448 ( .CLK(n1566), .C(n1567) );
  CKBD0 U1449 ( .CLK(n1567), .C(n1568) );
  CKBD0 U1450 ( .CLK(n1568), .C(n1569) );
  CKBD0 U1451 ( .CLK(n1569), .C(n1570) );
  BUFFD0 U1452 ( .I(n1570), .Z(n1571) );
  CKBD0 U1453 ( .CLK(n1571), .C(n1572) );
  CKBD0 U1454 ( .CLK(n1572), .C(n1573) );
  CKBD0 U1455 ( .CLK(n1573), .C(n1574) );
  CKBD0 U1456 ( .CLK(n1574), .C(n1575) );
  CKBD0 U1457 ( .CLK(n1575), .C(n1576) );
  CKBD0 U1458 ( .CLK(n1576), .C(n1577) );
  CKBD0 U1459 ( .CLK(n1577), .C(n1578) );
  CKBD0 U1460 ( .CLK(n1578), .C(n1579) );
  CKBD0 U1461 ( .CLK(n1579), .C(n1580) );
  CKBD0 U1462 ( .CLK(n1580), .C(n1581) );
  BUFFD0 U1463 ( .I(n1581), .Z(n1582) );
  CKBD0 U1464 ( .CLK(n1582), .C(n1583) );
  CKBD0 U1465 ( .CLK(n1583), .C(n1584) );
  CKBD0 U1466 ( .CLK(n1584), .C(n1585) );
  CKBD0 U1467 ( .CLK(n1585), .C(n1586) );
  CKBD0 U1468 ( .CLK(n1586), .C(n1587) );
  CKBD0 U1469 ( .CLK(n1587), .C(n1588) );
  CKBD0 U1470 ( .CLK(n1588), .C(n1589) );
  CKBD0 U1471 ( .CLK(n1589), .C(n1590) );
  CKBD0 U1472 ( .CLK(n1590), .C(n1591) );
  CKBD0 U1473 ( .CLK(n1591), .C(n1592) );
  BUFFD0 U1474 ( .I(n1592), .Z(n1593) );
  CKBD0 U1475 ( .CLK(n1593), .C(n1594) );
  CKBD0 U1476 ( .CLK(n1594), .C(n1595) );
  CKBD0 U1477 ( .CLK(n1595), .C(n1596) );
  CKBD0 U1478 ( .CLK(n1596), .C(n1597) );
  CKBD0 U1479 ( .CLK(n1597), .C(n1598) );
  CKBD0 U1480 ( .CLK(n1598), .C(n1599) );
  CKBD0 U1481 ( .CLK(n1599), .C(n1600) );
  CKBD0 U1482 ( .CLK(n1600), .C(n1601) );
  CKBD0 U1483 ( .CLK(n1601), .C(n1602) );
  CKBD0 U1484 ( .CLK(n1602), .C(n1603) );
  BUFFD0 U1485 ( .I(n1603), .Z(n1604) );
  CKBD0 U1486 ( .CLK(n1604), .C(n1605) );
  CKBD0 U1487 ( .CLK(n1605), .C(n1606) );
  CKBD0 U1488 ( .CLK(n1606), .C(n1607) );
  CKBD0 U1489 ( .CLK(n1607), .C(n1608) );
  CKBD0 U1490 ( .CLK(n1608), .C(n1609) );
  CKBD0 U1491 ( .CLK(n1609), .C(n1610) );
  CKBD0 U1492 ( .CLK(n1610), .C(n1611) );
  CKBD0 U1493 ( .CLK(n1611), .C(n1612) );
  CKBD0 U1494 ( .CLK(n1612), .C(n1613) );
  CKBD0 U1495 ( .CLK(n1613), .C(n1614) );
  BUFFD0 U1496 ( .I(n1614), .Z(n1615) );
  CKBD0 U1497 ( .CLK(n1615), .C(n1616) );
  CKBD0 U1498 ( .CLK(n1616), .C(n1617) );
  CKBD0 U1499 ( .CLK(n1617), .C(n1618) );
  CKBD0 U1500 ( .CLK(n1618), .C(n1619) );
  CKBD0 U1501 ( .CLK(n1619), .C(n1620) );
  CKBD0 U1502 ( .CLK(n1620), .C(n1621) );
  CKBD0 U1503 ( .CLK(n1621), .C(n1622) );
  CKBD0 U1504 ( .CLK(n1622), .C(n1623) );
  CKBD0 U1505 ( .CLK(n1623), .C(n1624) );
  CKBD0 U1506 ( .CLK(n1624), .C(n1625) );
  BUFFD0 U1507 ( .I(n1625), .Z(n1626) );
  CKBD0 U1508 ( .CLK(n1626), .C(n1627) );
  CKBD0 U1509 ( .CLK(n1627), .C(n1628) );
  CKBD0 U1510 ( .CLK(n1628), .C(n1629) );
  CKBD0 U1511 ( .CLK(n1629), .C(n1630) );
  CKBD0 U1512 ( .CLK(n1630), .C(n1631) );
  CKBD0 U1513 ( .CLK(n1631), .C(n1632) );
  CKBD0 U1514 ( .CLK(n1632), .C(n1633) );
  CKBD0 U1515 ( .CLK(n1633), .C(n1634) );
  CKBD0 U1516 ( .CLK(n1634), .C(n1635) );
  CKBD0 U1517 ( .CLK(n1635), .C(n1636) );
  BUFFD0 U1518 ( .I(n1636), .Z(n1637) );
  CKBD0 U1519 ( .CLK(n1637), .C(n1638) );
  CKBD0 U1520 ( .CLK(n1638), .C(n1639) );
  CKBD0 U1521 ( .CLK(n1639), .C(n1640) );
  CKBD0 U1522 ( .CLK(n1640), .C(n1641) );
  CKBD0 U1523 ( .CLK(n1641), .C(n1642) );
  BUFFD0 U1524 ( .I(n9009), .Z(n1643) );
  CKBD0 U1525 ( .CLK(FrameSR[1]), .C(n1644) );
  CKBD0 U1526 ( .CLK(n1644), .C(n1645) );
  BUFFD0 U1527 ( .I(n9011), .Z(n1646) );
  CKBD0 U1528 ( .CLK(FrameSR[5]), .C(n1647) );
  CKBD0 U1529 ( .CLK(n1647), .C(n1648) );
  BUFFD0 U1530 ( .I(n1648), .Z(n1649) );
  BUFFD0 U1531 ( .I(n9008), .Z(n1650) );
  CKBD0 U1532 ( .CLK(FrameSR[17]), .C(n1651) );
  BUFFD0 U1533 ( .I(n1651), .Z(n1652) );
  CKBD0 U1534 ( .CLK(n1652), .C(n1653) );
  CKBD0 U1535 ( .CLK(n1653), .C(n1654) );
  CKBD0 U1536 ( .CLK(n1654), .C(n1655) );
  CKBD0 U1537 ( .CLK(n1655), .C(n1656) );
  CKBD0 U1538 ( .CLK(n1656), .C(n1657) );
  CKBD0 U1539 ( .CLK(n1657), .C(n1658) );
  CKBD0 U1540 ( .CLK(n1658), .C(n1659) );
  CKBD0 U1541 ( .CLK(n1659), .C(n1660) );
  CKBD0 U1542 ( .CLK(n1660), .C(n1661) );
  CKBD0 U1543 ( .CLK(n1661), .C(n1662) );
  BUFFD0 U1544 ( .I(n1662), .Z(n1663) );
  CKBD0 U1545 ( .CLK(n1663), .C(n1664) );
  CKBD0 U1546 ( .CLK(n1664), .C(n1665) );
  CKBD0 U1547 ( .CLK(n1665), .C(n1666) );
  CKBD0 U1548 ( .CLK(n1666), .C(n1667) );
  CKBD0 U1549 ( .CLK(n1667), .C(n1668) );
  CKBD0 U1550 ( .CLK(n1668), .C(n1669) );
  CKBD0 U1551 ( .CLK(n1669), .C(n1670) );
  CKBD0 U1552 ( .CLK(n1670), .C(n1671) );
  CKBD0 U1553 ( .CLK(n1671), .C(n1672) );
  CKBD0 U1554 ( .CLK(n1672), .C(n1673) );
  BUFFD0 U1555 ( .I(n1673), .Z(n1674) );
  CKBD0 U1556 ( .CLK(n1674), .C(n1675) );
  CKBD0 U1557 ( .CLK(n1675), .C(n1676) );
  CKBD0 U1558 ( .CLK(n1676), .C(n1677) );
  CKBD0 U1559 ( .CLK(n1677), .C(n1678) );
  CKBD0 U1560 ( .CLK(n1678), .C(n1679) );
  CKBD0 U1561 ( .CLK(n1679), .C(n1680) );
  CKBD0 U1562 ( .CLK(n1680), .C(n1681) );
  CKBD0 U1563 ( .CLK(n1681), .C(n1682) );
  CKBD0 U1564 ( .CLK(n1682), .C(n1683) );
  CKBD0 U1565 ( .CLK(n1683), .C(n1684) );
  BUFFD0 U1566 ( .I(n1684), .Z(n1685) );
  CKBD0 U1567 ( .CLK(n1685), .C(n1686) );
  CKBD0 U1568 ( .CLK(n1686), .C(n1687) );
  CKBD0 U1569 ( .CLK(n1687), .C(n1688) );
  CKBD0 U1570 ( .CLK(n1688), .C(n1689) );
  CKBD0 U1571 ( .CLK(n1689), .C(n1690) );
  CKBD0 U1572 ( .CLK(n1690), .C(n1691) );
  CKBD0 U1573 ( .CLK(n1691), .C(n1692) );
  CKBD0 U1574 ( .CLK(n1692), .C(n1693) );
  CKBD0 U1575 ( .CLK(n1693), .C(n1694) );
  CKBD0 U1576 ( .CLK(n1694), .C(n1695) );
  BUFFD0 U1577 ( .I(n1695), .Z(n1696) );
  CKBD0 U1578 ( .CLK(n1696), .C(n1697) );
  CKBD0 U1579 ( .CLK(n1697), .C(n1698) );
  CKBD0 U1580 ( .CLK(n1698), .C(n1699) );
  CKBD0 U1581 ( .CLK(n1699), .C(n1700) );
  CKBD0 U1582 ( .CLK(n1700), .C(n1701) );
  CKBD0 U1583 ( .CLK(n1701), .C(n1702) );
  CKBD0 U1584 ( .CLK(n1702), .C(n1703) );
  CKBD0 U1585 ( .CLK(n1703), .C(n1704) );
  CKBD0 U1586 ( .CLK(n1704), .C(n1705) );
  CKBD0 U1587 ( .CLK(n1705), .C(n1706) );
  BUFFD0 U1588 ( .I(n1706), .Z(n1707) );
  CKBD0 U1589 ( .CLK(n1707), .C(n1708) );
  CKBD0 U1590 ( .CLK(n1708), .C(n1709) );
  CKBD0 U1591 ( .CLK(n1709), .C(n1710) );
  CKBD0 U1592 ( .CLK(n1710), .C(n1711) );
  CKBD0 U1593 ( .CLK(n1711), .C(n1712) );
  CKBD0 U1594 ( .CLK(n1712), .C(n1713) );
  CKBD0 U1595 ( .CLK(n1713), .C(n1714) );
  CKBD0 U1596 ( .CLK(n1714), .C(n1715) );
  CKBD0 U1597 ( .CLK(n1715), .C(n1716) );
  BUFFD0 U1598 ( .I(n1716), .Z(n1717) );
  CKBD0 U1599 ( .CLK(n1717), .C(n1718) );
  CKBD0 U1600 ( .CLK(n1718), .C(n1719) );
  CKBD0 U1601 ( .CLK(n1719), .C(n1720) );
  CKBD0 U1602 ( .CLK(n1720), .C(n1721) );
  CKBD0 U1603 ( .CLK(n1721), .C(n1722) );
  CKBD0 U1604 ( .CLK(n1722), .C(n1723) );
  CKBD0 U1605 ( .CLK(n1723), .C(n1724) );
  CKBD0 U1606 ( .CLK(n1724), .C(n1725) );
  CKBD0 U1607 ( .CLK(n1725), .C(n1726) );
  CKBD0 U1608 ( .CLK(n1726), .C(n1727) );
  BUFFD0 U1609 ( .I(n1727), .Z(n1728) );
  CKBD0 U1610 ( .CLK(n1728), .C(n1729) );
  CKBD0 U1611 ( .CLK(n1729), .C(n1730) );
  CKBD0 U1612 ( .CLK(n1730), .C(n1731) );
  CKBD0 U1613 ( .CLK(n1731), .C(n1732) );
  CKBD0 U1614 ( .CLK(n1732), .C(n1733) );
  CKBD0 U1615 ( .CLK(n1733), .C(n1734) );
  CKBD0 U1616 ( .CLK(n1734), .C(n1735) );
  CKBD0 U1617 ( .CLK(n1735), .C(n1736) );
  CKBD0 U1618 ( .CLK(n1736), .C(n1737) );
  CKBD0 U1619 ( .CLK(n1737), .C(n1738) );
  BUFFD0 U1620 ( .I(n1738), .Z(n1739) );
  CKBD0 U1621 ( .CLK(n1739), .C(n1740) );
  CKBD0 U1622 ( .CLK(n1740), .C(n1741) );
  CKBD0 U1623 ( .CLK(n1741), .C(n1742) );
  CKBD0 U1624 ( .CLK(n1742), .C(n1743) );
  CKBD0 U1625 ( .CLK(n1743), .C(n1744) );
  CKBD0 U1626 ( .CLK(n1744), .C(n1745) );
  BUFFD0 U1627 ( .I(n8964), .Z(n1746) );
  CKBD0 U1628 ( .CLK(FrameSR[32]), .C(n1747) );
  BUFFD0 U1629 ( .I(n1747), .Z(n1748) );
  CKBD0 U1630 ( .CLK(n1748), .C(n1749) );
  CKBD0 U1631 ( .CLK(n1749), .C(n1750) );
  CKBD0 U1632 ( .CLK(n1750), .C(n1751) );
  CKBD0 U1633 ( .CLK(n1751), .C(n1752) );
  CKBD0 U1634 ( .CLK(n1752), .C(n1753) );
  CKBD0 U1635 ( .CLK(n1753), .C(n1754) );
  CKBD0 U1636 ( .CLK(n1754), .C(n1755) );
  CKBD0 U1637 ( .CLK(n1755), .C(n1756) );
  CKBD0 U1638 ( .CLK(n1756), .C(n1757) );
  BUFFD0 U1639 ( .I(n1757), .Z(n1758) );
  CKBD0 U1640 ( .CLK(n1758), .C(n1759) );
  CKBD0 U1641 ( .CLK(n1759), .C(n1760) );
  CKBD0 U1642 ( .CLK(n1760), .C(n1761) );
  CKBD0 U1643 ( .CLK(n1761), .C(n1762) );
  CKBD0 U1644 ( .CLK(n1762), .C(n1763) );
  CKBD0 U1645 ( .CLK(n1763), .C(n1764) );
  CKBD0 U1646 ( .CLK(n1764), .C(n1765) );
  CKBD0 U1647 ( .CLK(n1765), .C(n1766) );
  CKBD0 U1648 ( .CLK(n1766), .C(n1767) );
  CKBD0 U1649 ( .CLK(n1767), .C(n1768) );
  BUFFD0 U1650 ( .I(n1768), .Z(n1769) );
  CKBD0 U1651 ( .CLK(n1769), .C(n1770) );
  CKBD0 U1652 ( .CLK(n1770), .C(n1771) );
  CKBD0 U1653 ( .CLK(n1771), .C(n1772) );
  CKBD0 U1654 ( .CLK(n1772), .C(n1773) );
  CKBD0 U1655 ( .CLK(n1773), .C(n1774) );
  CKBD0 U1656 ( .CLK(n1774), .C(n1775) );
  CKBD0 U1657 ( .CLK(n1775), .C(n1776) );
  CKBD0 U1658 ( .CLK(n1776), .C(n1777) );
  CKBD0 U1659 ( .CLK(n1777), .C(n1778) );
  CKBD0 U1660 ( .CLK(n1778), .C(n1779) );
  BUFFD0 U1661 ( .I(n1779), .Z(n1780) );
  CKBD0 U1662 ( .CLK(n1780), .C(n1781) );
  CKBD0 U1663 ( .CLK(n1781), .C(n1782) );
  CKBD0 U1664 ( .CLK(n1782), .C(n1783) );
  CKBD0 U1665 ( .CLK(n1783), .C(n1784) );
  CKBD0 U1666 ( .CLK(n1784), .C(n1785) );
  CKBD0 U1667 ( .CLK(n1785), .C(n1786) );
  CKBD0 U1668 ( .CLK(n1786), .C(n1787) );
  CKBD0 U1669 ( .CLK(n1787), .C(n1788) );
  CKBD0 U1670 ( .CLK(n1788), .C(n1789) );
  CKBD0 U1671 ( .CLK(n1789), .C(n1790) );
  BUFFD0 U1672 ( .I(n1790), .Z(n1791) );
  CKBD0 U1673 ( .CLK(n1791), .C(n1792) );
  CKBD0 U1674 ( .CLK(n1792), .C(n1793) );
  CKBD0 U1675 ( .CLK(n1793), .C(n1794) );
  CKBD0 U1676 ( .CLK(n1794), .C(n1795) );
  CKBD0 U1677 ( .CLK(n1795), .C(n1796) );
  CKBD0 U1678 ( .CLK(n1796), .C(n1797) );
  CKBD0 U1679 ( .CLK(n1797), .C(n1798) );
  CKBD0 U1680 ( .CLK(n1798), .C(n1799) );
  CKBD0 U1681 ( .CLK(n1799), .C(n1800) );
  CKBD0 U1682 ( .CLK(n1800), .C(n1801) );
  BUFFD0 U1683 ( .I(n1801), .Z(n1802) );
  CKBD0 U1684 ( .CLK(n1802), .C(n1803) );
  CKBD0 U1685 ( .CLK(n1803), .C(n1804) );
  CKBD0 U1686 ( .CLK(n1804), .C(n1805) );
  CKBD0 U1687 ( .CLK(n1805), .C(n1806) );
  CKBD0 U1688 ( .CLK(n1806), .C(n1807) );
  CKBD0 U1689 ( .CLK(n1807), .C(n1808) );
  CKBD0 U1690 ( .CLK(n1808), .C(n1809) );
  CKBD0 U1691 ( .CLK(n1809), .C(n1810) );
  CKBD0 U1692 ( .CLK(n1810), .C(n1811) );
  CKBD0 U1693 ( .CLK(n1811), .C(n1812) );
  BUFFD0 U1694 ( .I(n1812), .Z(n1813) );
  CKBD0 U1695 ( .CLK(n1813), .C(n1814) );
  CKBD0 U1696 ( .CLK(n1814), .C(n1815) );
  CKBD0 U1697 ( .CLK(n1815), .C(n1816) );
  CKBD0 U1698 ( .CLK(n1816), .C(n1817) );
  CKBD0 U1699 ( .CLK(n1817), .C(n1818) );
  CKBD0 U1700 ( .CLK(n1818), .C(n1819) );
  CKBD0 U1701 ( .CLK(n1819), .C(n1820) );
  CKBD0 U1702 ( .CLK(n1820), .C(n1821) );
  CKBD0 U1703 ( .CLK(n1821), .C(n1822) );
  CKBD0 U1704 ( .CLK(n1822), .C(n1823) );
  BUFFD0 U1705 ( .I(n1823), .Z(n1824) );
  CKBD0 U1706 ( .CLK(n1824), .C(n1825) );
  CKBD0 U1707 ( .CLK(n1825), .C(n1826) );
  CKBD0 U1708 ( .CLK(n1826), .C(n1827) );
  CKBD0 U1709 ( .CLK(n1827), .C(n1828) );
  CKBD0 U1710 ( .CLK(n1828), .C(n1829) );
  CKBD0 U1711 ( .CLK(n1829), .C(n1830) );
  CKBD0 U1712 ( .CLK(n1830), .C(n1831) );
  CKBD0 U1713 ( .CLK(n1831), .C(n1832) );
  CKBD0 U1714 ( .CLK(n1832), .C(n1833) );
  BUFFD0 U1715 ( .I(n1833), .Z(n1834) );
  CKBD0 U1716 ( .CLK(n1834), .C(n1835) );
  CKBD0 U1717 ( .CLK(n1835), .C(n1836) );
  CKBD0 U1718 ( .CLK(n1836), .C(n1837) );
  CKBD0 U1719 ( .CLK(n1837), .C(n1838) );
  CKBD0 U1720 ( .CLK(n1838), .C(n1839) );
  CKBD0 U1721 ( .CLK(n1839), .C(n1840) );
  CKBD0 U1722 ( .CLK(n1840), .C(n1841) );
  CKBD0 U1723 ( .CLK(n1841), .C(n1842) );
  BUFFD0 U1724 ( .I(n3754), .Z(n1843) );
  CKBD0 U1725 ( .CLK(FrameSR[47]), .C(n1844) );
  BUFFD0 U1726 ( .I(n9006), .Z(n1845) );
  CKBD0 U1727 ( .CLK(FrameSR[0]), .C(n1846) );
  CKBD0 U1728 ( .CLK(n1846), .C(n1847) );
  BUFFD0 U1729 ( .I(n9013), .Z(n1848) );
  CKBD0 U1730 ( .CLK(FrameSR[2]), .C(n1849) );
  CKBD0 U1731 ( .CLK(n1849), .C(n1850) );
  BUFFD0 U1732 ( .I(n9010), .Z(n1851) );
  CKBD0 U1733 ( .CLK(FrameSR[4]), .C(n1852) );
  CKBD0 U1734 ( .CLK(n1852), .C(n1853) );
  BUFFD0 U1735 ( .I(n9014), .Z(n1854) );
  CKBD0 U1736 ( .CLK(FrameSR[6]), .C(n1855) );
  CKBD0 U1737 ( .CLK(n1855), .C(n1856) );
  BUFFD0 U1738 ( .I(n1856), .Z(n1857) );
  BUFFD0 U1739 ( .I(n8989), .Z(n1858) );
  CKBD0 U1740 ( .CLK(FrameSR[20]), .C(n1859) );
  CKBD0 U1741 ( .CLK(n1859), .C(n1860) );
  BUFFD0 U1742 ( .I(n1860), .Z(n1861) );
  CKBD0 U1743 ( .CLK(n1861), .C(n1862) );
  CKBD0 U1744 ( .CLK(n1862), .C(n1863) );
  CKBD0 U1745 ( .CLK(n1863), .C(n1864) );
  CKBD0 U1746 ( .CLK(n1864), .C(n1865) );
  CKBD0 U1747 ( .CLK(n1865), .C(n1866) );
  CKBD0 U1748 ( .CLK(n1866), .C(n1867) );
  CKBD0 U1749 ( .CLK(n1867), .C(n1868) );
  CKBD0 U1750 ( .CLK(n1868), .C(n1869) );
  CKBD0 U1751 ( .CLK(n1869), .C(n1870) );
  CKBD0 U1752 ( .CLK(n1870), .C(n1871) );
  BUFFD0 U1753 ( .I(n1871), .Z(n1872) );
  CKBD0 U1754 ( .CLK(n1872), .C(n1873) );
  CKBD0 U1755 ( .CLK(n1873), .C(n1874) );
  CKBD0 U1756 ( .CLK(n1874), .C(n1875) );
  CKBD0 U1757 ( .CLK(n1875), .C(n1876) );
  CKBD0 U1758 ( .CLK(n1876), .C(n1877) );
  CKBD0 U1759 ( .CLK(n1877), .C(n1878) );
  CKBD0 U1760 ( .CLK(n1878), .C(n1879) );
  CKBD0 U1761 ( .CLK(n1879), .C(n1880) );
  CKBD0 U1762 ( .CLK(n1880), .C(n1881) );
  BUFFD0 U1763 ( .I(n1881), .Z(n1882) );
  CKBD0 U1764 ( .CLK(n1882), .C(n1883) );
  CKBD0 U1765 ( .CLK(n1883), .C(n1884) );
  CKBD0 U1766 ( .CLK(n1884), .C(n1885) );
  CKBD0 U1767 ( .CLK(n1885), .C(n1886) );
  CKBD0 U1768 ( .CLK(n1886), .C(n1887) );
  CKBD0 U1769 ( .CLK(n1887), .C(n1888) );
  CKBD0 U1770 ( .CLK(n1888), .C(n1889) );
  CKBD0 U1771 ( .CLK(n1889), .C(n1890) );
  CKBD0 U1772 ( .CLK(n1890), .C(n1891) );
  CKBD0 U1773 ( .CLK(n1891), .C(n1892) );
  BUFFD0 U1774 ( .I(n1892), .Z(n1893) );
  CKBD0 U1775 ( .CLK(n1893), .C(n1894) );
  CKBD0 U1776 ( .CLK(n1894), .C(n1895) );
  CKBD0 U1777 ( .CLK(n1895), .C(n1896) );
  CKBD0 U1778 ( .CLK(n1896), .C(n1897) );
  CKBD0 U1779 ( .CLK(n1897), .C(n1898) );
  CKBD0 U1780 ( .CLK(n1898), .C(n1899) );
  CKBD0 U1781 ( .CLK(n1899), .C(n1900) );
  CKBD0 U1782 ( .CLK(n1900), .C(n1901) );
  CKBD0 U1783 ( .CLK(n1901), .C(n1902) );
  CKBD0 U1784 ( .CLK(n1902), .C(n1903) );
  BUFFD0 U1785 ( .I(n1903), .Z(n1904) );
  CKBD0 U1786 ( .CLK(n1904), .C(n1905) );
  CKBD0 U1787 ( .CLK(n1905), .C(n1906) );
  CKBD0 U1788 ( .CLK(n1906), .C(n1907) );
  CKBD0 U1789 ( .CLK(n1907), .C(n1908) );
  CKBD0 U1790 ( .CLK(n1908), .C(n1909) );
  CKBD0 U1791 ( .CLK(n1909), .C(n1910) );
  CKBD0 U1792 ( .CLK(n1910), .C(n1911) );
  CKBD0 U1793 ( .CLK(n1911), .C(n1912) );
  CKBD0 U1794 ( .CLK(n1912), .C(n1913) );
  CKBD0 U1795 ( .CLK(n1913), .C(n1914) );
  BUFFD0 U1796 ( .I(n1914), .Z(n1915) );
  CKBD0 U1797 ( .CLK(n1915), .C(n1916) );
  CKBD0 U1798 ( .CLK(n1916), .C(n1917) );
  CKBD0 U1799 ( .CLK(n1917), .C(n1918) );
  CKBD0 U1800 ( .CLK(n1918), .C(n1919) );
  CKBD0 U1801 ( .CLK(n1919), .C(n1920) );
  CKBD0 U1802 ( .CLK(n1920), .C(n1921) );
  CKBD0 U1803 ( .CLK(n1921), .C(n1922) );
  CKBD0 U1804 ( .CLK(n1922), .C(n1923) );
  CKBD0 U1805 ( .CLK(n1923), .C(n1924) );
  CKBD0 U1806 ( .CLK(n1924), .C(n1925) );
  BUFFD0 U1807 ( .I(n1925), .Z(n1926) );
  CKBD0 U1808 ( .CLK(n1926), .C(n1927) );
  CKBD0 U1809 ( .CLK(n1927), .C(n1928) );
  CKBD0 U1810 ( .CLK(n1928), .C(n1929) );
  CKBD0 U1811 ( .CLK(n1929), .C(n1930) );
  CKBD0 U1812 ( .CLK(n1930), .C(n1931) );
  CKBD0 U1813 ( .CLK(n1931), .C(n1932) );
  CKBD0 U1814 ( .CLK(n1932), .C(n1933) );
  CKBD0 U1815 ( .CLK(n1933), .C(n1934) );
  CKBD0 U1816 ( .CLK(n1934), .C(n1935) );
  CKBD0 U1817 ( .CLK(n1935), .C(n1936) );
  BUFFD0 U1818 ( .I(n1936), .Z(n1937) );
  CKBD0 U1819 ( .CLK(n1937), .C(n1938) );
  CKBD0 U1820 ( .CLK(n1938), .C(n1939) );
  CKBD0 U1821 ( .CLK(n1939), .C(n1940) );
  CKBD0 U1822 ( .CLK(n1940), .C(n1941) );
  CKBD0 U1823 ( .CLK(n1941), .C(n1942) );
  CKBD0 U1824 ( .CLK(n1942), .C(n1943) );
  CKBD0 U1825 ( .CLK(n1943), .C(n1944) );
  CKBD0 U1826 ( .CLK(n1944), .C(n1945) );
  CKBD0 U1827 ( .CLK(n1945), .C(n1946) );
  CKBD0 U1828 ( .CLK(n1946), .C(n1947) );
  BUFFD0 U1829 ( .I(n1947), .Z(n1948) );
  CKBD0 U1830 ( .CLK(n1948), .C(n1949) );
  CKBD0 U1831 ( .CLK(n1949), .C(n1950) );
  CKBD0 U1832 ( .CLK(n1950), .C(n1951) );
  CKBD0 U1833 ( .CLK(n1951), .C(n1952) );
  CKBD0 U1834 ( .CLK(n1952), .C(n1953) );
  BUFFD0 U1835 ( .I(n8990), .Z(n1954) );
  CKBD0 U1836 ( .CLK(FrameSR[34]), .C(n1955) );
  CKBD0 U1837 ( .CLK(n1955), .C(n1956) );
  BUFFD0 U1838 ( .I(n1956), .Z(n1957) );
  CKBD0 U1839 ( .CLK(n1957), .C(n1958) );
  CKBD0 U1840 ( .CLK(n1958), .C(n1959) );
  CKBD0 U1841 ( .CLK(n1959), .C(n1960) );
  CKBD0 U1842 ( .CLK(n1960), .C(n1961) );
  CKBD0 U1843 ( .CLK(n1961), .C(n1962) );
  CKBD0 U1844 ( .CLK(n1962), .C(n1963) );
  CKBD0 U1845 ( .CLK(n1963), .C(n1964) );
  CKBD0 U1846 ( .CLK(n1964), .C(n1965) );
  CKBD0 U1847 ( .CLK(n1965), .C(n1966) );
  CKBD0 U1848 ( .CLK(n1966), .C(n1967) );
  BUFFD0 U1849 ( .I(n1967), .Z(n1968) );
  CKBD0 U1850 ( .CLK(n1968), .C(n1969) );
  CKBD0 U1851 ( .CLK(n1969), .C(n1970) );
  CKBD0 U1852 ( .CLK(n1970), .C(n1971) );
  CKBD0 U1853 ( .CLK(n1971), .C(n1972) );
  CKBD0 U1854 ( .CLK(n1972), .C(n1973) );
  CKBD0 U1855 ( .CLK(n1973), .C(n1974) );
  CKBD0 U1856 ( .CLK(n1974), .C(n1975) );
  CKBD0 U1857 ( .CLK(n1975), .C(n1976) );
  CKBD0 U1858 ( .CLK(n1976), .C(n1977) );
  BUFFD0 U1859 ( .I(n1977), .Z(n1978) );
  CKBD0 U1860 ( .CLK(n1978), .C(n1979) );
  CKBD0 U1861 ( .CLK(n1979), .C(n1980) );
  CKBD0 U1862 ( .CLK(n1980), .C(n1981) );
  CKBD0 U1863 ( .CLK(n1981), .C(n1982) );
  CKBD0 U1864 ( .CLK(n1982), .C(n1983) );
  CKBD0 U1865 ( .CLK(n1983), .C(n1984) );
  CKBD0 U1866 ( .CLK(n1984), .C(n1985) );
  CKBD0 U1867 ( .CLK(n1985), .C(n1986) );
  CKBD0 U1868 ( .CLK(n1986), .C(n1987) );
  CKBD0 U1869 ( .CLK(n1987), .C(n1988) );
  BUFFD0 U1870 ( .I(n1988), .Z(n1989) );
  CKBD0 U1871 ( .CLK(n1989), .C(n1990) );
  CKBD0 U1872 ( .CLK(n1990), .C(n1991) );
  CKBD0 U1873 ( .CLK(n1991), .C(n1992) );
  CKBD0 U1874 ( .CLK(n1992), .C(n1993) );
  CKBD0 U1875 ( .CLK(n1993), .C(n1994) );
  CKBD0 U1876 ( .CLK(n1994), .C(n1995) );
  CKBD0 U1877 ( .CLK(n1995), .C(n1996) );
  CKBD0 U1878 ( .CLK(n1996), .C(n1997) );
  CKBD0 U1879 ( .CLK(n1997), .C(n1998) );
  CKBD0 U1880 ( .CLK(n1998), .C(n1999) );
  BUFFD0 U1881 ( .I(n1999), .Z(n2000) );
  CKBD0 U1882 ( .CLK(n2000), .C(n2001) );
  CKBD0 U1883 ( .CLK(n2001), .C(n2002) );
  CKBD0 U1884 ( .CLK(n2002), .C(n2003) );
  CKBD0 U1885 ( .CLK(n2003), .C(n2004) );
  CKBD0 U1886 ( .CLK(n2004), .C(n2005) );
  CKBD0 U1887 ( .CLK(n2005), .C(n2006) );
  CKBD0 U1888 ( .CLK(n2006), .C(n2007) );
  CKBD0 U1889 ( .CLK(n2007), .C(n2008) );
  CKBD0 U1890 ( .CLK(n2008), .C(n2009) );
  CKBD0 U1891 ( .CLK(n2009), .C(n2010) );
  BUFFD0 U1892 ( .I(n2010), .Z(n2011) );
  CKBD0 U1893 ( .CLK(n2011), .C(n2012) );
  CKBD0 U1894 ( .CLK(n2012), .C(n2013) );
  CKBD0 U1895 ( .CLK(n2013), .C(n2014) );
  CKBD0 U1896 ( .CLK(n2014), .C(n2015) );
  CKBD0 U1897 ( .CLK(n2015), .C(n2016) );
  CKBD0 U1898 ( .CLK(n2016), .C(n2017) );
  CKBD0 U1899 ( .CLK(n2017), .C(n2018) );
  CKBD0 U1900 ( .CLK(n2018), .C(n2019) );
  CKBD0 U1901 ( .CLK(n2019), .C(n2020) );
  CKBD0 U1902 ( .CLK(n2020), .C(n2021) );
  BUFFD0 U1903 ( .I(n2021), .Z(n2022) );
  CKBD0 U1904 ( .CLK(n2022), .C(n2023) );
  CKBD0 U1905 ( .CLK(n2023), .C(n2024) );
  CKBD0 U1906 ( .CLK(n2024), .C(n2025) );
  CKBD0 U1907 ( .CLK(n2025), .C(n2026) );
  CKBD0 U1908 ( .CLK(n2026), .C(n2027) );
  CKBD0 U1909 ( .CLK(n2027), .C(n2028) );
  CKBD0 U1910 ( .CLK(n2028), .C(n2029) );
  CKBD0 U1911 ( .CLK(n2029), .C(n2030) );
  CKBD0 U1912 ( .CLK(n2030), .C(n2031) );
  CKBD0 U1913 ( .CLK(n2031), .C(n2032) );
  BUFFD0 U1914 ( .I(n2032), .Z(n2033) );
  CKBD0 U1915 ( .CLK(n2033), .C(n2034) );
  CKBD0 U1916 ( .CLK(n2034), .C(n2035) );
  CKBD0 U1917 ( .CLK(n2035), .C(n2036) );
  CKBD0 U1918 ( .CLK(n2036), .C(n2037) );
  CKBD0 U1919 ( .CLK(n2037), .C(n2038) );
  CKBD0 U1920 ( .CLK(n2038), .C(n2039) );
  CKBD0 U1921 ( .CLK(n2039), .C(n2040) );
  CKBD0 U1922 ( .CLK(n2040), .C(n2041) );
  CKBD0 U1923 ( .CLK(n2041), .C(n2042) );
  CKBD0 U1924 ( .CLK(n2042), .C(n2043) );
  BUFFD0 U1925 ( .I(n2043), .Z(n2044) );
  CKBD0 U1926 ( .CLK(n2044), .C(n2045) );
  CKBD0 U1927 ( .CLK(n2045), .C(n2046) );
  CKBD0 U1928 ( .CLK(n2046), .C(n2047) );
  CKBD0 U1929 ( .CLK(n2047), .C(n2048) );
  CKBD0 U1930 ( .CLK(n2048), .C(n2049) );
  BUFFD0 U1931 ( .I(n8988), .Z(n2050) );
  CKBD0 U1932 ( .CLK(FrameSR[49]), .C(n2051) );
  CKBD0 U1933 ( .CLK(n2051), .C(n2052) );
  BUFFD0 U1934 ( .I(n2052), .Z(n2053) );
  CKBD0 U1935 ( .CLK(n2053), .C(n2054) );
  CKBD0 U1936 ( .CLK(n2054), .C(n2055) );
  CKBD0 U1937 ( .CLK(n2055), .C(n2056) );
  CKBD0 U1938 ( .CLK(n2056), .C(n2057) );
  CKBD0 U1939 ( .CLK(n2057), .C(n2058) );
  CKBD0 U1940 ( .CLK(n2058), .C(n2059) );
  CKBD0 U1941 ( .CLK(n2059), .C(n2060) );
  CKBD0 U1942 ( .CLK(n2060), .C(n2061) );
  CKBD0 U1943 ( .CLK(n2061), .C(n2062) );
  CKBD0 U1944 ( .CLK(n2062), .C(n2063) );
  BUFFD0 U1945 ( .I(n2063), .Z(n2064) );
  CKBD0 U1946 ( .CLK(n2064), .C(n2065) );
  CKBD0 U1947 ( .CLK(n2065), .C(n2066) );
  CKBD0 U1948 ( .CLK(n2066), .C(n2067) );
  CKBD0 U1949 ( .CLK(n2067), .C(n2068) );
  CKBD0 U1950 ( .CLK(n2068), .C(n2069) );
  CKBD0 U1951 ( .CLK(n2069), .C(n2070) );
  CKBD0 U1952 ( .CLK(n2070), .C(n2071) );
  CKBD0 U1953 ( .CLK(n2071), .C(n2072) );
  CKBD0 U1954 ( .CLK(n2072), .C(n2073) );
  BUFFD0 U1955 ( .I(n2073), .Z(n2074) );
  CKBD0 U1956 ( .CLK(n2074), .C(n2075) );
  CKBD0 U1957 ( .CLK(n2075), .C(n2076) );
  CKBD0 U1958 ( .CLK(n2076), .C(n2077) );
  CKBD0 U1959 ( .CLK(n2077), .C(n2078) );
  CKBD0 U1960 ( .CLK(n2078), .C(n2079) );
  CKBD0 U1961 ( .CLK(n2079), .C(n2080) );
  CKBD0 U1962 ( .CLK(n2080), .C(n2081) );
  CKBD0 U1963 ( .CLK(n2081), .C(n2082) );
  CKBD0 U1964 ( .CLK(n2082), .C(n2083) );
  CKBD0 U1965 ( .CLK(n2083), .C(n2084) );
  BUFFD0 U1966 ( .I(n2084), .Z(n2085) );
  CKBD0 U1967 ( .CLK(n2085), .C(n2086) );
  CKBD0 U1968 ( .CLK(n2086), .C(n2087) );
  CKBD0 U1969 ( .CLK(n2087), .C(n2088) );
  CKBD0 U1970 ( .CLK(n2088), .C(n2089) );
  CKBD0 U1971 ( .CLK(n2089), .C(n2090) );
  CKBD0 U1972 ( .CLK(n2090), .C(n2091) );
  CKBD0 U1973 ( .CLK(n2091), .C(n2092) );
  CKBD0 U1974 ( .CLK(n2092), .C(n2093) );
  CKBD0 U1975 ( .CLK(n2093), .C(n2094) );
  CKBD0 U1976 ( .CLK(n2094), .C(n2095) );
  BUFFD0 U1977 ( .I(n2095), .Z(n2096) );
  CKBD0 U1978 ( .CLK(n2096), .C(n2097) );
  CKBD0 U1979 ( .CLK(n2097), .C(n2098) );
  CKBD0 U1980 ( .CLK(n2098), .C(n2099) );
  CKBD0 U1981 ( .CLK(n2099), .C(n2100) );
  CKBD0 U1982 ( .CLK(n2100), .C(n2101) );
  CKBD0 U1983 ( .CLK(n2101), .C(n2102) );
  CKBD0 U1984 ( .CLK(n2102), .C(n2103) );
  CKBD0 U1985 ( .CLK(n2103), .C(n2104) );
  CKBD0 U1986 ( .CLK(n2104), .C(n2105) );
  CKBD0 U1987 ( .CLK(n2105), .C(n2106) );
  BUFFD0 U1988 ( .I(n2106), .Z(n2107) );
  CKBD0 U1989 ( .CLK(n2107), .C(n2108) );
  CKBD0 U1990 ( .CLK(n2108), .C(n2109) );
  CKBD0 U1991 ( .CLK(n2109), .C(n2110) );
  CKBD0 U1992 ( .CLK(n2110), .C(n2111) );
  CKBD0 U1993 ( .CLK(n2111), .C(n2112) );
  CKBD0 U1994 ( .CLK(n2112), .C(n2113) );
  CKBD0 U1995 ( .CLK(n2113), .C(n2114) );
  CKBD0 U1996 ( .CLK(n2114), .C(n2115) );
  CKBD0 U1997 ( .CLK(n2115), .C(n2116) );
  CKBD0 U1998 ( .CLK(n2116), .C(n2117) );
  BUFFD0 U1999 ( .I(n2117), .Z(n2118) );
  CKBD0 U2000 ( .CLK(n2118), .C(n2119) );
  CKBD0 U2001 ( .CLK(n2119), .C(n2120) );
  CKBD0 U2002 ( .CLK(n2120), .C(n2121) );
  CKBD0 U2003 ( .CLK(n2121), .C(n2122) );
  CKBD0 U2004 ( .CLK(n2122), .C(n2123) );
  CKBD0 U2005 ( .CLK(n2123), .C(n2124) );
  CKBD0 U2006 ( .CLK(n2124), .C(n2125) );
  CKBD0 U2007 ( .CLK(n2125), .C(n2126) );
  CKBD0 U2008 ( .CLK(n2126), .C(n2127) );
  CKBD0 U2009 ( .CLK(n2127), .C(n2128) );
  BUFFD0 U2010 ( .I(n2128), .Z(n2129) );
  CKBD0 U2011 ( .CLK(n2129), .C(n2130) );
  CKBD0 U2012 ( .CLK(n2130), .C(n2131) );
  CKBD0 U2013 ( .CLK(n2131), .C(n2132) );
  CKBD0 U2014 ( .CLK(n2132), .C(n2133) );
  CKBD0 U2015 ( .CLK(n2133), .C(n2134) );
  CKBD0 U2016 ( .CLK(n2134), .C(n2135) );
  CKBD0 U2017 ( .CLK(n2135), .C(n2136) );
  CKBD0 U2018 ( .CLK(n2136), .C(n2137) );
  CKBD0 U2019 ( .CLK(n2137), .C(n2138) );
  CKBD0 U2020 ( .CLK(n2138), .C(n2139) );
  BUFFD0 U2021 ( .I(n2139), .Z(n2140) );
  CKBD0 U2022 ( .CLK(n2140), .C(n2141) );
  CKBD0 U2023 ( .CLK(n2141), .C(n2142) );
  CKBD0 U2024 ( .CLK(n2142), .C(n2143) );
  CKBD0 U2025 ( .CLK(n2143), .C(n2144) );
  CKBD0 U2026 ( .CLK(n2144), .C(n2145) );
  BUFFD0 U2027 ( .I(n8991), .Z(n2146) );
  CKBD0 U2028 ( .CLK(FrameSR[50]), .C(n2147) );
  CKBD0 U2029 ( .CLK(n2147), .C(n2148) );
  BUFFD0 U2030 ( .I(n2148), .Z(n2149) );
  CKBD0 U2031 ( .CLK(n2149), .C(n2150) );
  CKBD0 U2032 ( .CLK(n2150), .C(n2151) );
  CKBD0 U2033 ( .CLK(n2151), .C(n2152) );
  CKBD0 U2034 ( .CLK(n2152), .C(n2153) );
  CKBD0 U2035 ( .CLK(n2153), .C(n2154) );
  CKBD0 U2036 ( .CLK(n2154), .C(n2155) );
  CKBD0 U2037 ( .CLK(n2155), .C(n2156) );
  CKBD0 U2038 ( .CLK(n2156), .C(n2157) );
  CKBD0 U2039 ( .CLK(n2157), .C(n2158) );
  CKBD0 U2040 ( .CLK(n2158), .C(n2159) );
  BUFFD0 U2041 ( .I(n2159), .Z(n2160) );
  CKBD0 U2042 ( .CLK(n2160), .C(n2161) );
  CKBD0 U2043 ( .CLK(n2161), .C(n2162) );
  CKBD0 U2044 ( .CLK(n2162), .C(n2163) );
  CKBD0 U2045 ( .CLK(n2163), .C(n2164) );
  CKBD0 U2046 ( .CLK(n2164), .C(n2165) );
  CKBD0 U2047 ( .CLK(n2165), .C(n2166) );
  CKBD0 U2048 ( .CLK(n2166), .C(n2167) );
  CKBD0 U2049 ( .CLK(n2167), .C(n2168) );
  CKBD0 U2050 ( .CLK(n2168), .C(n2169) );
  BUFFD0 U2051 ( .I(n2169), .Z(n2170) );
  CKBD0 U2052 ( .CLK(n2170), .C(n2171) );
  CKBD0 U2053 ( .CLK(n2171), .C(n2172) );
  CKBD0 U2054 ( .CLK(n2172), .C(n2173) );
  CKBD0 U2055 ( .CLK(n2173), .C(n2174) );
  CKBD0 U2056 ( .CLK(n2174), .C(n2175) );
  CKBD0 U2057 ( .CLK(n2175), .C(n2176) );
  CKBD0 U2058 ( .CLK(n2176), .C(n2177) );
  CKBD0 U2059 ( .CLK(n2177), .C(n2178) );
  CKBD0 U2060 ( .CLK(n2178), .C(n2179) );
  CKBD0 U2061 ( .CLK(n2179), .C(n2180) );
  BUFFD0 U2062 ( .I(n2180), .Z(n2181) );
  CKBD0 U2063 ( .CLK(n2181), .C(n2182) );
  CKBD0 U2064 ( .CLK(n2182), .C(n2183) );
  CKBD0 U2065 ( .CLK(n2183), .C(n2184) );
  CKBD0 U2066 ( .CLK(n2184), .C(n2185) );
  CKBD0 U2067 ( .CLK(n2185), .C(n2186) );
  CKBD0 U2068 ( .CLK(n2186), .C(n2187) );
  CKBD0 U2069 ( .CLK(n2187), .C(n2188) );
  CKBD0 U2070 ( .CLK(n2188), .C(n2189) );
  CKBD0 U2071 ( .CLK(n2189), .C(n2190) );
  CKBD0 U2072 ( .CLK(n2190), .C(n2191) );
  BUFFD0 U2073 ( .I(n2191), .Z(n2192) );
  CKBD0 U2074 ( .CLK(n2192), .C(n2193) );
  CKBD0 U2075 ( .CLK(n2193), .C(n2194) );
  CKBD0 U2076 ( .CLK(n2194), .C(n2195) );
  CKBD0 U2077 ( .CLK(n2195), .C(n2196) );
  CKBD0 U2078 ( .CLK(n2196), .C(n2197) );
  CKBD0 U2079 ( .CLK(n2197), .C(n2198) );
  CKBD0 U2080 ( .CLK(n2198), .C(n2199) );
  CKBD0 U2081 ( .CLK(n2199), .C(n2200) );
  CKBD0 U2082 ( .CLK(n2200), .C(n2201) );
  CKBD0 U2083 ( .CLK(n2201), .C(n2202) );
  BUFFD0 U2084 ( .I(n2202), .Z(n2203) );
  CKBD0 U2085 ( .CLK(n2203), .C(n2204) );
  CKBD0 U2086 ( .CLK(n2204), .C(n2205) );
  CKBD0 U2087 ( .CLK(n2205), .C(n2206) );
  CKBD0 U2088 ( .CLK(n2206), .C(n2207) );
  CKBD0 U2089 ( .CLK(n2207), .C(n2208) );
  CKBD0 U2090 ( .CLK(n2208), .C(n2209) );
  CKBD0 U2091 ( .CLK(n2209), .C(n2210) );
  CKBD0 U2092 ( .CLK(n2210), .C(n2211) );
  CKBD0 U2093 ( .CLK(n2211), .C(n2212) );
  CKBD0 U2094 ( .CLK(n2212), .C(n2213) );
  BUFFD0 U2095 ( .I(n2213), .Z(n2214) );
  CKBD0 U2096 ( .CLK(n2214), .C(n2215) );
  CKBD0 U2097 ( .CLK(n2215), .C(n2216) );
  CKBD0 U2098 ( .CLK(n2216), .C(n2217) );
  CKBD0 U2099 ( .CLK(n2217), .C(n2218) );
  CKBD0 U2100 ( .CLK(n2218), .C(n2219) );
  CKBD0 U2101 ( .CLK(n2219), .C(n2220) );
  CKBD0 U2102 ( .CLK(n2220), .C(n2221) );
  CKBD0 U2103 ( .CLK(n2221), .C(n2222) );
  CKBD0 U2104 ( .CLK(n2222), .C(n2223) );
  CKBD0 U2105 ( .CLK(n2223), .C(n2224) );
  BUFFD0 U2106 ( .I(n2224), .Z(n2225) );
  CKBD0 U2107 ( .CLK(n2225), .C(n2226) );
  CKBD0 U2108 ( .CLK(n2226), .C(n2227) );
  CKBD0 U2109 ( .CLK(n2227), .C(n2228) );
  CKBD0 U2110 ( .CLK(n2228), .C(n2229) );
  CKBD0 U2111 ( .CLK(n2229), .C(n2230) );
  CKBD0 U2112 ( .CLK(n2230), .C(n2231) );
  CKBD0 U2113 ( .CLK(n2231), .C(n2232) );
  CKBD0 U2114 ( .CLK(n2232), .C(n2233) );
  CKBD0 U2115 ( .CLK(n2233), .C(n2234) );
  CKBD0 U2116 ( .CLK(n2234), .C(n2235) );
  BUFFD0 U2117 ( .I(n2235), .Z(n2236) );
  CKBD0 U2118 ( .CLK(n2236), .C(n2237) );
  CKBD0 U2119 ( .CLK(n2237), .C(n2238) );
  CKBD0 U2120 ( .CLK(n2238), .C(n2239) );
  CKBD0 U2121 ( .CLK(n2239), .C(n2240) );
  CKBD0 U2122 ( .CLK(n2240), .C(n2241) );
  BUFFD0 U2123 ( .I(n8993), .Z(n2242) );
  CKBD0 U2124 ( .CLK(FrameSR[35]), .C(n2243) );
  CKBD0 U2125 ( .CLK(n2243), .C(n2244) );
  BUFFD0 U2126 ( .I(n2244), .Z(n2245) );
  CKBD0 U2127 ( .CLK(n2245), .C(n2246) );
  CKBD0 U2128 ( .CLK(n2246), .C(n2247) );
  CKBD0 U2129 ( .CLK(n2247), .C(n2248) );
  CKBD0 U2130 ( .CLK(n2248), .C(n2249) );
  CKBD0 U2131 ( .CLK(n2249), .C(n2250) );
  CKBD0 U2132 ( .CLK(n2250), .C(n2251) );
  CKBD0 U2133 ( .CLK(n2251), .C(n2252) );
  CKBD0 U2134 ( .CLK(n2252), .C(n2253) );
  CKBD0 U2135 ( .CLK(n2253), .C(n2254) );
  CKBD0 U2136 ( .CLK(n2254), .C(n2255) );
  BUFFD0 U2137 ( .I(n2255), .Z(n2256) );
  CKBD0 U2138 ( .CLK(n2256), .C(n2257) );
  CKBD0 U2139 ( .CLK(n2257), .C(n2258) );
  CKBD0 U2140 ( .CLK(n2258), .C(n2259) );
  CKBD0 U2141 ( .CLK(n2259), .C(n2260) );
  CKBD0 U2142 ( .CLK(n2260), .C(n2261) );
  CKBD0 U2143 ( .CLK(n2261), .C(n2262) );
  CKBD0 U2144 ( .CLK(n2262), .C(n2263) );
  CKBD0 U2145 ( .CLK(n2263), .C(n2264) );
  CKBD0 U2146 ( .CLK(n2264), .C(n2265) );
  BUFFD0 U2147 ( .I(n2265), .Z(n2266) );
  CKBD0 U2148 ( .CLK(n2266), .C(n2267) );
  CKBD0 U2149 ( .CLK(n2267), .C(n2268) );
  CKBD0 U2150 ( .CLK(n2268), .C(n2269) );
  CKBD0 U2151 ( .CLK(n2269), .C(n2270) );
  CKBD0 U2152 ( .CLK(n2270), .C(n2271) );
  CKBD0 U2153 ( .CLK(n2271), .C(n2272) );
  CKBD0 U2154 ( .CLK(n2272), .C(n2273) );
  CKBD0 U2155 ( .CLK(n2273), .C(n2274) );
  CKBD0 U2156 ( .CLK(n2274), .C(n2275) );
  CKBD0 U2157 ( .CLK(n2275), .C(n2276) );
  BUFFD0 U2158 ( .I(n2276), .Z(n2277) );
  CKBD0 U2159 ( .CLK(n2277), .C(n2278) );
  CKBD0 U2160 ( .CLK(n2278), .C(n2279) );
  CKBD0 U2161 ( .CLK(n2279), .C(n2280) );
  CKBD0 U2162 ( .CLK(n2280), .C(n2281) );
  CKBD0 U2163 ( .CLK(n2281), .C(n2282) );
  CKBD0 U2164 ( .CLK(n2282), .C(n2283) );
  CKBD0 U2165 ( .CLK(n2283), .C(n2284) );
  CKBD0 U2166 ( .CLK(n2284), .C(n2285) );
  CKBD0 U2167 ( .CLK(n2285), .C(n2286) );
  CKBD0 U2168 ( .CLK(n2286), .C(n2287) );
  BUFFD0 U2169 ( .I(n2287), .Z(n2288) );
  CKBD0 U2170 ( .CLK(n2288), .C(n2289) );
  CKBD0 U2171 ( .CLK(n2289), .C(n2290) );
  CKBD0 U2172 ( .CLK(n2290), .C(n2291) );
  CKBD0 U2173 ( .CLK(n2291), .C(n2292) );
  CKBD0 U2174 ( .CLK(n2292), .C(n2293) );
  CKBD0 U2175 ( .CLK(n2293), .C(n2294) );
  CKBD0 U2176 ( .CLK(n2294), .C(n2295) );
  CKBD0 U2177 ( .CLK(n2295), .C(n2296) );
  CKBD0 U2178 ( .CLK(n2296), .C(n2297) );
  CKBD0 U2179 ( .CLK(n2297), .C(n2298) );
  BUFFD0 U2180 ( .I(n2298), .Z(n2299) );
  CKBD0 U2181 ( .CLK(n2299), .C(n2300) );
  CKBD0 U2182 ( .CLK(n2300), .C(n2301) );
  CKBD0 U2183 ( .CLK(n2301), .C(n2302) );
  CKBD0 U2184 ( .CLK(n2302), .C(n2303) );
  CKBD0 U2185 ( .CLK(n2303), .C(n2304) );
  CKBD0 U2186 ( .CLK(n2304), .C(n2305) );
  CKBD0 U2187 ( .CLK(n2305), .C(n2306) );
  CKBD0 U2188 ( .CLK(n2306), .C(n2307) );
  CKBD0 U2189 ( .CLK(n2307), .C(n2308) );
  CKBD0 U2190 ( .CLK(n2308), .C(n2309) );
  BUFFD0 U2191 ( .I(n2309), .Z(n2310) );
  CKBD0 U2192 ( .CLK(n2310), .C(n2311) );
  CKBD0 U2193 ( .CLK(n2311), .C(n2312) );
  CKBD0 U2194 ( .CLK(n2312), .C(n2313) );
  CKBD0 U2195 ( .CLK(n2313), .C(n2314) );
  CKBD0 U2196 ( .CLK(n2314), .C(n2315) );
  CKBD0 U2197 ( .CLK(n2315), .C(n2316) );
  CKBD0 U2198 ( .CLK(n2316), .C(n2317) );
  CKBD0 U2199 ( .CLK(n2317), .C(n2318) );
  CKBD0 U2200 ( .CLK(n2318), .C(n2319) );
  CKBD0 U2201 ( .CLK(n2319), .C(n2320) );
  BUFFD0 U2202 ( .I(n2320), .Z(n2321) );
  CKBD0 U2203 ( .CLK(n2321), .C(n2322) );
  CKBD0 U2204 ( .CLK(n2322), .C(n2323) );
  CKBD0 U2205 ( .CLK(n2323), .C(n2324) );
  CKBD0 U2206 ( .CLK(n2324), .C(n2325) );
  CKBD0 U2207 ( .CLK(n2325), .C(n2326) );
  CKBD0 U2208 ( .CLK(n2326), .C(n2327) );
  CKBD0 U2209 ( .CLK(n2327), .C(n2328) );
  CKBD0 U2210 ( .CLK(n2328), .C(n2329) );
  CKBD0 U2211 ( .CLK(n2329), .C(n2330) );
  CKBD0 U2212 ( .CLK(n2330), .C(n2331) );
  BUFFD0 U2213 ( .I(n2331), .Z(n2332) );
  CKBD0 U2214 ( .CLK(n2332), .C(n2333) );
  CKBD0 U2215 ( .CLK(n2333), .C(n2334) );
  CKBD0 U2216 ( .CLK(n2334), .C(n2335) );
  CKBD0 U2217 ( .CLK(n2335), .C(n2336) );
  CKBD0 U2218 ( .CLK(n2336), .C(n2337) );
  BUFFD0 U2219 ( .I(n8980), .Z(n2338) );
  CKBD0 U2220 ( .CLK(FrameSR[51]), .C(n2339) );
  CKBD0 U2221 ( .CLK(n2339), .C(n2340) );
  CKBD0 U2222 ( .CLK(n2340), .C(n2341) );
  CKBD0 U2223 ( .CLK(n2341), .C(n2342) );
  CKBD0 U2224 ( .CLK(n2342), .C(n2343) );
  CKBD0 U2225 ( .CLK(n2343), .C(n2344) );
  CKBD0 U2226 ( .CLK(n2344), .C(n2345) );
  CKBD0 U2227 ( .CLK(n2345), .C(n2346) );
  CKBD0 U2228 ( .CLK(n2346), .C(n2347) );
  CKBD0 U2229 ( .CLK(n2347), .C(n2348) );
  BUFFD0 U2230 ( .I(n2348), .Z(n2349) );
  CKBD0 U2231 ( .CLK(n2349), .C(n2350) );
  CKBD0 U2232 ( .CLK(n2350), .C(n2351) );
  CKBD0 U2233 ( .CLK(n2351), .C(n2352) );
  CKBD0 U2234 ( .CLK(n2352), .C(n2353) );
  CKBD0 U2235 ( .CLK(n2353), .C(n2354) );
  CKBD0 U2236 ( .CLK(n2354), .C(n2355) );
  CKBD0 U2237 ( .CLK(n2355), .C(n2356) );
  CKBD0 U2238 ( .CLK(n2356), .C(n2357) );
  CKBD0 U2239 ( .CLK(n2357), .C(n2358) );
  BUFFD0 U2240 ( .I(n2358), .Z(n2359) );
  CKBD0 U2241 ( .CLK(n2359), .C(n2360) );
  CKBD0 U2242 ( .CLK(n2360), .C(n2361) );
  CKBD0 U2243 ( .CLK(n2361), .C(n2362) );
  CKBD0 U2244 ( .CLK(n2362), .C(n2363) );
  CKBD0 U2245 ( .CLK(n2363), .C(n2364) );
  CKBD0 U2246 ( .CLK(n2364), .C(n2365) );
  CKBD0 U2247 ( .CLK(n2365), .C(n2366) );
  CKBD0 U2248 ( .CLK(n2366), .C(n2367) );
  CKBD0 U2249 ( .CLK(n2367), .C(n2368) );
  CKBD0 U2250 ( .CLK(n2368), .C(n2369) );
  BUFFD0 U2251 ( .I(n2369), .Z(n2370) );
  CKBD0 U2252 ( .CLK(n2370), .C(n2371) );
  CKBD0 U2253 ( .CLK(n2371), .C(n2372) );
  CKBD0 U2254 ( .CLK(n2372), .C(n2373) );
  CKBD0 U2255 ( .CLK(n2373), .C(n2374) );
  CKBD0 U2256 ( .CLK(n2374), .C(n2375) );
  CKBD0 U2257 ( .CLK(n2375), .C(n2376) );
  CKBD0 U2258 ( .CLK(n2376), .C(n2377) );
  CKBD0 U2259 ( .CLK(n2377), .C(n2378) );
  CKBD0 U2260 ( .CLK(n2378), .C(n2379) );
  CKBD0 U2261 ( .CLK(n2379), .C(n2380) );
  BUFFD0 U2262 ( .I(n2380), .Z(n2381) );
  CKBD0 U2263 ( .CLK(n2381), .C(n2382) );
  CKBD0 U2264 ( .CLK(n2382), .C(n2383) );
  CKBD0 U2265 ( .CLK(n2383), .C(n2384) );
  CKBD0 U2266 ( .CLK(n2384), .C(n2385) );
  CKBD0 U2267 ( .CLK(n2385), .C(n2386) );
  CKBD0 U2268 ( .CLK(n2386), .C(n2387) );
  CKBD0 U2269 ( .CLK(n2387), .C(n2388) );
  CKBD0 U2270 ( .CLK(n2388), .C(n2389) );
  CKBD0 U2271 ( .CLK(n2389), .C(n2390) );
  CKBD0 U2272 ( .CLK(n2390), .C(n2391) );
  BUFFD0 U2273 ( .I(n2391), .Z(n2392) );
  CKBD0 U2274 ( .CLK(n2392), .C(n2393) );
  CKBD0 U2275 ( .CLK(n2393), .C(n2394) );
  CKBD0 U2276 ( .CLK(n2394), .C(n2395) );
  CKBD0 U2277 ( .CLK(n2395), .C(n2396) );
  CKBD0 U2278 ( .CLK(n2396), .C(n2397) );
  CKBD0 U2279 ( .CLK(n2397), .C(n2398) );
  CKBD0 U2280 ( .CLK(n2398), .C(n2399) );
  CKBD0 U2281 ( .CLK(n2399), .C(n2400) );
  CKBD0 U2282 ( .CLK(n2400), .C(n2401) );
  CKBD0 U2283 ( .CLK(n2401), .C(n2402) );
  BUFFD0 U2284 ( .I(n2402), .Z(n2403) );
  CKBD0 U2285 ( .CLK(n2403), .C(n2404) );
  CKBD0 U2286 ( .CLK(n2404), .C(n2405) );
  CKBD0 U2287 ( .CLK(n2405), .C(n2406) );
  CKBD0 U2288 ( .CLK(n2406), .C(n2407) );
  CKBD0 U2289 ( .CLK(n2407), .C(n2408) );
  CKBD0 U2290 ( .CLK(n2408), .C(n2409) );
  CKBD0 U2291 ( .CLK(n2409), .C(n2410) );
  CKBD0 U2292 ( .CLK(n2410), .C(n2411) );
  CKBD0 U2293 ( .CLK(n2411), .C(n2412) );
  CKBD0 U2294 ( .CLK(n2412), .C(n2413) );
  BUFFD0 U2295 ( .I(n2413), .Z(n2414) );
  CKBD0 U2296 ( .CLK(n2414), .C(n2415) );
  CKBD0 U2297 ( .CLK(n2415), .C(n2416) );
  CKBD0 U2298 ( .CLK(n2416), .C(n2417) );
  CKBD0 U2299 ( .CLK(n2417), .C(n2418) );
  CKBD0 U2300 ( .CLK(n2418), .C(n2419) );
  CKBD0 U2301 ( .CLK(n2419), .C(n2420) );
  CKBD0 U2302 ( .CLK(n2420), .C(n2421) );
  CKBD0 U2303 ( .CLK(n2421), .C(n2422) );
  CKBD0 U2304 ( .CLK(n2422), .C(n2423) );
  BUFFD0 U2305 ( .I(n2423), .Z(n2424) );
  CKBD0 U2306 ( .CLK(n2424), .C(n2425) );
  CKBD0 U2307 ( .CLK(n2425), .C(n2426) );
  CKBD0 U2308 ( .CLK(n2426), .C(n2427) );
  CKBD0 U2309 ( .CLK(n2427), .C(n2428) );
  CKBD0 U2310 ( .CLK(n2428), .C(n2429) );
  CKBD0 U2311 ( .CLK(n2429), .C(n2430) );
  CKBD0 U2312 ( .CLK(n2430), .C(n2431) );
  CKBD0 U2313 ( .CLK(n2431), .C(n2432) );
  CKBD0 U2314 ( .CLK(n2432), .C(n2433) );
  BUFFD0 U2315 ( .I(n9012), .Z(n2434) );
  CKBD0 U2316 ( .CLK(FrameSR[16]), .C(n2435) );
  BUFFD0 U2317 ( .I(n2435), .Z(n2436) );
  CKBD0 U2318 ( .CLK(n2436), .C(n2437) );
  CKBD0 U2319 ( .CLK(n2437), .C(n2438) );
  CKBD0 U2320 ( .CLK(n2438), .C(n2439) );
  CKBD0 U2321 ( .CLK(n2439), .C(n2440) );
  CKBD0 U2322 ( .CLK(n2440), .C(n2441) );
  CKBD0 U2323 ( .CLK(n2441), .C(n2442) );
  CKBD0 U2324 ( .CLK(n2442), .C(n2443) );
  CKBD0 U2325 ( .CLK(n2443), .C(n2444) );
  CKBD0 U2326 ( .CLK(n2444), .C(n2445) );
  CKBD0 U2327 ( .CLK(n2445), .C(n2446) );
  BUFFD0 U2328 ( .I(n2446), .Z(n2447) );
  CKBD0 U2329 ( .CLK(n2447), .C(n2448) );
  CKBD0 U2330 ( .CLK(n2448), .C(n2449) );
  CKBD0 U2331 ( .CLK(n2449), .C(n2450) );
  CKBD0 U2332 ( .CLK(n2450), .C(n2451) );
  CKBD0 U2333 ( .CLK(n2451), .C(n2452) );
  CKBD0 U2334 ( .CLK(n2452), .C(n2453) );
  CKBD0 U2335 ( .CLK(n2453), .C(n2454) );
  CKBD0 U2336 ( .CLK(n2454), .C(n2455) );
  CKBD0 U2337 ( .CLK(n2455), .C(n2456) );
  CKBD0 U2338 ( .CLK(n2456), .C(n2457) );
  BUFFD0 U2339 ( .I(n2457), .Z(n2458) );
  CKBD0 U2340 ( .CLK(n2458), .C(n2459) );
  CKBD0 U2341 ( .CLK(n2459), .C(n2460) );
  CKBD0 U2342 ( .CLK(n2460), .C(n2461) );
  CKBD0 U2343 ( .CLK(n2461), .C(n2462) );
  CKBD0 U2344 ( .CLK(n2462), .C(n2463) );
  CKBD0 U2345 ( .CLK(n2463), .C(n2464) );
  CKBD0 U2346 ( .CLK(n2464), .C(n2465) );
  CKBD0 U2347 ( .CLK(n2465), .C(n2466) );
  CKBD0 U2348 ( .CLK(n2466), .C(n2467) );
  CKBD0 U2349 ( .CLK(n2467), .C(n2468) );
  BUFFD0 U2350 ( .I(n2468), .Z(n2469) );
  CKBD0 U2351 ( .CLK(n2469), .C(n2470) );
  CKBD0 U2352 ( .CLK(n2470), .C(n2471) );
  CKBD0 U2353 ( .CLK(n2471), .C(n2472) );
  CKBD0 U2354 ( .CLK(n2472), .C(n2473) );
  CKBD0 U2355 ( .CLK(n2473), .C(n2474) );
  CKBD0 U2356 ( .CLK(n2474), .C(n2475) );
  CKBD0 U2357 ( .CLK(n2475), .C(n2476) );
  CKBD0 U2358 ( .CLK(n2476), .C(n2477) );
  CKBD0 U2359 ( .CLK(n2477), .C(n2478) );
  BUFFD0 U2360 ( .I(n2478), .Z(n2479) );
  CKBD0 U2361 ( .CLK(n2479), .C(n2480) );
  CKBD0 U2362 ( .CLK(n2480), .C(n2481) );
  CKBD0 U2363 ( .CLK(n2481), .C(n2482) );
  CKBD0 U2364 ( .CLK(n2482), .C(n2483) );
  CKBD0 U2365 ( .CLK(n2483), .C(n2484) );
  CKBD0 U2366 ( .CLK(n2484), .C(n2485) );
  CKBD0 U2367 ( .CLK(n2485), .C(n2486) );
  CKBD0 U2368 ( .CLK(n2486), .C(n2487) );
  CKBD0 U2369 ( .CLK(n2487), .C(n2488) );
  CKBD0 U2370 ( .CLK(n2488), .C(n2489) );
  BUFFD0 U2371 ( .I(n2489), .Z(n2490) );
  CKBD0 U2372 ( .CLK(n2490), .C(n2491) );
  CKBD0 U2373 ( .CLK(n2491), .C(n2492) );
  CKBD0 U2374 ( .CLK(n2492), .C(n2493) );
  CKBD0 U2375 ( .CLK(n2493), .C(n2494) );
  CKBD0 U2376 ( .CLK(n2494), .C(n2495) );
  CKBD0 U2377 ( .CLK(n2495), .C(n2496) );
  CKBD0 U2378 ( .CLK(n2496), .C(n2497) );
  CKBD0 U2379 ( .CLK(n2497), .C(n2498) );
  CKBD0 U2380 ( .CLK(n2498), .C(n2499) );
  CKBD0 U2381 ( .CLK(n2499), .C(n2500) );
  BUFFD0 U2382 ( .I(n2500), .Z(n2501) );
  CKBD0 U2383 ( .CLK(n2501), .C(n2502) );
  CKBD0 U2384 ( .CLK(n2502), .C(n2503) );
  CKBD0 U2385 ( .CLK(n2503), .C(n2504) );
  CKBD0 U2386 ( .CLK(n2504), .C(n2505) );
  CKBD0 U2387 ( .CLK(n2505), .C(n2506) );
  CKBD0 U2388 ( .CLK(n2506), .C(n2507) );
  CKBD0 U2389 ( .CLK(n2507), .C(n2508) );
  CKBD0 U2390 ( .CLK(n2508), .C(n2509) );
  CKBD0 U2391 ( .CLK(n2509), .C(n2510) );
  CKBD0 U2392 ( .CLK(n2510), .C(n2511) );
  BUFFD0 U2393 ( .I(n2511), .Z(n2512) );
  CKBD0 U2394 ( .CLK(n2512), .C(n2513) );
  CKBD0 U2395 ( .CLK(n2513), .C(n2514) );
  CKBD0 U2396 ( .CLK(n2514), .C(n2515) );
  CKBD0 U2397 ( .CLK(n2515), .C(n2516) );
  CKBD0 U2398 ( .CLK(n2516), .C(n2517) );
  CKBD0 U2399 ( .CLK(n2517), .C(n2518) );
  CKBD0 U2400 ( .CLK(n2518), .C(n2519) );
  CKBD0 U2401 ( .CLK(n2519), .C(n2520) );
  CKBD0 U2402 ( .CLK(n2520), .C(n2521) );
  CKBD0 U2403 ( .CLK(n2521), .C(n2522) );
  BUFFD0 U2404 ( .I(n2522), .Z(n2523) );
  CKBD0 U2405 ( .CLK(n2523), .C(n2524) );
  CKBD0 U2406 ( .CLK(n2524), .C(n2525) );
  CKBD0 U2407 ( .CLK(n2525), .C(n2526) );
  CKBD0 U2408 ( .CLK(n2526), .C(n2527) );
  CKBD0 U2409 ( .CLK(n2527), .C(n2528) );
  CKBD0 U2410 ( .CLK(n2528), .C(n2529) );
  BUFFD0 U2411 ( .I(n5932), .Z(n2530) );
  CKBD0 U2412 ( .CLK(FrameSR[15]), .C(n2531) );
  BUFFD0 U2413 ( .I(N42), .Z(n2532) );
  BUFFD0 U2414 ( .I(n2664), .Z(n2533) );
  CKBD0 U2415 ( .CLK(FrameSR[63]), .C(n2534) );
  CKBD0 U2416 ( .CLK(n2534), .C(n2535) );
  CKBD0 U2417 ( .CLK(n2535), .C(n2536) );
  CKBD0 U2418 ( .CLK(n2536), .C(n2537) );
  CKBD0 U2419 ( .CLK(n2537), .C(n2538) );
  CKBD0 U2420 ( .CLK(n2538), .C(n2539) );
  CKBD0 U2421 ( .CLK(n2539), .C(n2540) );
  CKBD0 U2422 ( .CLK(n2540), .C(n2541) );
  CKBD0 U2423 ( .CLK(n2541), .C(n2542) );
  CKBD0 U2424 ( .CLK(n2542), .C(n2543) );
  BUFFD0 U2425 ( .I(n2543), .Z(n2544) );
  CKBD0 U2426 ( .CLK(n2544), .C(n2545) );
  CKBD0 U2427 ( .CLK(n2545), .C(n2546) );
  CKBD0 U2428 ( .CLK(n2546), .C(n2547) );
  CKBD0 U2429 ( .CLK(n2547), .C(n2548) );
  CKBD0 U2430 ( .CLK(n2548), .C(n2549) );
  CKBD0 U2431 ( .CLK(n2549), .C(n2550) );
  CKBD0 U2432 ( .CLK(n2550), .C(n2551) );
  CKBD0 U2433 ( .CLK(n2551), .C(n2552) );
  CKBD0 U2434 ( .CLK(n2552), .C(n2553) );
  CKBD0 U2435 ( .CLK(n2553), .C(n2554) );
  BUFFD0 U2436 ( .I(n2554), .Z(n2555) );
  CKBD0 U2437 ( .CLK(n2555), .C(n2556) );
  CKBD0 U2438 ( .CLK(n2556), .C(n2557) );
  CKBD0 U2439 ( .CLK(n2557), .C(n2558) );
  CKBD0 U2440 ( .CLK(n2558), .C(n2559) );
  CKBD0 U2441 ( .CLK(n2559), .C(n2560) );
  CKBD0 U2442 ( .CLK(n2560), .C(n2561) );
  CKBD0 U2443 ( .CLK(n2561), .C(n2562) );
  CKBD0 U2444 ( .CLK(n2562), .C(n2563) );
  CKBD0 U2445 ( .CLK(n2563), .C(n2564) );
  CKBD0 U2446 ( .CLK(n2564), .C(n2565) );
  BUFFD0 U2447 ( .I(n2565), .Z(n2566) );
  CKBD0 U2448 ( .CLK(n2566), .C(n2567) );
  CKBD0 U2449 ( .CLK(n2567), .C(n2568) );
  CKBD0 U2450 ( .CLK(n2568), .C(n2569) );
  CKBD0 U2451 ( .CLK(n2569), .C(n2570) );
  CKBD0 U2452 ( .CLK(n2570), .C(n2571) );
  CKBD0 U2453 ( .CLK(n2571), .C(n2572) );
  CKBD0 U2454 ( .CLK(n2572), .C(n2573) );
  CKBD0 U2455 ( .CLK(n2573), .C(n2574) );
  CKBD0 U2456 ( .CLK(n2574), .C(n2575) );
  CKBD0 U2457 ( .CLK(n2575), .C(n2576) );
  BUFFD0 U2458 ( .I(n2576), .Z(n2577) );
  CKBD0 U2459 ( .CLK(n2577), .C(n2578) );
  CKBD0 U2460 ( .CLK(n2578), .C(n2579) );
  CKBD0 U2461 ( .CLK(n2579), .C(n2580) );
  CKBD0 U2462 ( .CLK(n2580), .C(n2581) );
  CKBD0 U2463 ( .CLK(n2581), .C(n2582) );
  CKBD0 U2464 ( .CLK(n2582), .C(n2583) );
  CKBD0 U2465 ( .CLK(n2583), .C(n2584) );
  CKBD0 U2466 ( .CLK(n2584), .C(n2585) );
  CKBD0 U2467 ( .CLK(n2585), .C(n2586) );
  CKBD0 U2468 ( .CLK(n2586), .C(n2587) );
  BUFFD0 U2469 ( .I(n2587), .Z(n2588) );
  CKBD0 U2470 ( .CLK(n2588), .C(n2589) );
  CKBD0 U2471 ( .CLK(n2589), .C(n2590) );
  CKBD0 U2472 ( .CLK(n2590), .C(n2591) );
  CKBD0 U2473 ( .CLK(n2591), .C(n2592) );
  CKBD0 U2474 ( .CLK(n2592), .C(n2593) );
  CKBD0 U2475 ( .CLK(n2593), .C(n2594) );
  CKBD0 U2476 ( .CLK(n2594), .C(n2595) );
  CKBD0 U2477 ( .CLK(n2595), .C(n2596) );
  CKBD0 U2478 ( .CLK(n2596), .C(n2597) );
  CKBD0 U2479 ( .CLK(n2597), .C(n2598) );
  BUFFD0 U2480 ( .I(n2598), .Z(n2599) );
  CKBD0 U2481 ( .CLK(n2599), .C(n2600) );
  CKBD0 U2482 ( .CLK(n2600), .C(n2601) );
  CKBD0 U2483 ( .CLK(n2601), .C(n2602) );
  CKBD0 U2484 ( .CLK(n2602), .C(n2603) );
  CKBD0 U2485 ( .CLK(n2603), .C(n2604) );
  CKBD0 U2486 ( .CLK(n2604), .C(n2605) );
  CKBD0 U2487 ( .CLK(n2605), .C(n2606) );
  CKBD0 U2488 ( .CLK(n2606), .C(n2607) );
  CKBD0 U2489 ( .CLK(n2607), .C(n2608) );
  BUFFD0 U2490 ( .I(n2608), .Z(n2609) );
  CKBD0 U2491 ( .CLK(n2609), .C(n2610) );
  CKBD0 U2492 ( .CLK(n2610), .C(n2611) );
  CKBD0 U2493 ( .CLK(n2611), .C(n2612) );
  CKBD0 U2494 ( .CLK(n2612), .C(n2613) );
  CKBD0 U2495 ( .CLK(n2613), .C(n2614) );
  CKBD0 U2496 ( .CLK(n2614), .C(n2615) );
  CKBD0 U2497 ( .CLK(n2615), .C(n2616) );
  CKBD0 U2498 ( .CLK(n2616), .C(n2617) );
  CKBD0 U2499 ( .CLK(n2617), .C(n2618) );
  CKBD0 U2500 ( .CLK(n2618), .C(n2619) );
  BUFFD0 U2501 ( .I(n2619), .Z(n2620) );
  CKBD0 U2502 ( .CLK(n2620), .C(n2621) );
  CKBD0 U2503 ( .CLK(n2621), .C(n2622) );
  CKBD0 U2504 ( .CLK(n2622), .C(n2623) );
  CKBD0 U2505 ( .CLK(n2623), .C(n2624) );
  CKBD0 U2506 ( .CLK(n2624), .C(n2625) );
  CKBD0 U2507 ( .CLK(n2625), .C(n2626) );
  CKBD0 U2508 ( .CLK(n2626), .C(n2627) );
  CKBD0 U2509 ( .CLK(n2627), .C(n2628) );
  CKBD0 U2510 ( .CLK(n2628), .C(n2629) );
  CKBD0 U2511 ( .CLK(n2629), .C(n2630) );
  BUFFD0 U2512 ( .I(n2630), .Z(n2631) );
  CKBD0 U2513 ( .CLK(n2631), .C(n2632) );
  CKBD0 U2514 ( .CLK(n2632), .C(n2633) );
  CKBD0 U2515 ( .CLK(n2633), .C(n2634) );
  CKBD0 U2516 ( .CLK(n2634), .C(n2635) );
  BUFFD0 U2517 ( .I(n2635), .Z(n2636) );
  CKBD0 U2518 ( .CLK(n2636), .C(n2637) );
  BUFFD0 U2519 ( .I(n2637), .Z(n2638) );
  CKBD0 U2520 ( .CLK(n2638), .C(n2639) );
  BUFFD0 U2521 ( .I(n2639), .Z(n2640) );
  CKBD0 U2522 ( .CLK(n2640), .C(n2641) );
  BUFFD0 U2523 ( .I(n2641), .Z(n2642) );
  CKBD0 U2524 ( .CLK(n2642), .C(n2643) );
  BUFFD0 U2525 ( .I(n2643), .Z(n2644) );
  CKBD0 U2526 ( .CLK(n2644), .C(n2645) );
  BUFFD0 U2527 ( .I(n2645), .Z(n2646) );
  CKBD0 U2528 ( .CLK(n2646), .C(n2647) );
  BUFFD0 U2529 ( .I(n2647), .Z(n2648) );
  CKBD0 U2530 ( .CLK(n2648), .C(n2649) );
  BUFFD0 U2531 ( .I(n2649), .Z(n2650) );
  CKBD0 U2532 ( .CLK(n2650), .C(n2651) );
  BUFFD0 U2533 ( .I(n2651), .Z(n2652) );
  CKBD0 U2534 ( .CLK(n2652), .C(n2653) );
  BUFFD0 U2535 ( .I(n2653), .Z(n2654) );
  CKBD0 U2536 ( .CLK(n2654), .C(n2655) );
  BUFFD0 U2537 ( .I(n2655), .Z(n2656) );
  CKBD0 U2538 ( .CLK(n2656), .C(n2657) );
  BUFFD0 U2539 ( .I(n2657), .Z(n2658) );
  CKBD0 U2540 ( .CLK(n2658), .C(n2659) );
  BUFFD0 U2541 ( .I(n2659), .Z(n2660) );
  CKBD0 U2542 ( .CLK(n2660), .C(n2661) );
  BUFFD0 U2543 ( .I(n2661), .Z(n2662) );
  CKBD0 U2544 ( .CLK(n2662), .C(n2663) );
  BUFFD0 U2545 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2546 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2547 ( .I(n164), .Z(n2666) );
  BUFFD0 U2548 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2549 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2550 ( .I(n163), .Z(n2669) );
  CKBD0 U2551 ( .CLK(n5), .C(n2670) );
  CKBD0 U2552 ( .CLK(n2670), .C(n2671) );
  CKBD0 U2553 ( .CLK(n2671), .C(n2672) );
  BUFFD0 U2554 ( .I(n2672), .Z(n2673) );
  CKBD0 U2555 ( .CLK(n2673), .C(n2674) );
  CKBD0 U2556 ( .CLK(n2674), .C(n2675) );
  CKBD0 U2557 ( .CLK(n2675), .C(n2676) );
  CKBD0 U2558 ( .CLK(n2676), .C(n2677) );
  CKBD0 U2559 ( .CLK(n2677), .C(n2678) );
  CKBD0 U2560 ( .CLK(n2678), .C(n2679) );
  CKBD0 U2561 ( .CLK(n2679), .C(n2680) );
  CKBD0 U2562 ( .CLK(n2680), .C(n2681) );
  CKBD0 U2563 ( .CLK(n2681), .C(n2682) );
  CKBD0 U2564 ( .CLK(n2682), .C(n2683) );
  BUFFD0 U2565 ( .I(n2683), .Z(n2684) );
  CKBD0 U2566 ( .CLK(n2684), .C(n2685) );
  CKBD0 U2567 ( .CLK(n2685), .C(n2686) );
  CKBD0 U2568 ( .CLK(n2686), .C(n2687) );
  CKBD0 U2569 ( .CLK(n2687), .C(n2688) );
  CKBD0 U2570 ( .CLK(n2688), .C(n2689) );
  CKBD0 U2571 ( .CLK(n2689), .C(n2690) );
  CKBD0 U2572 ( .CLK(n2690), .C(n2691) );
  CKBD0 U2573 ( .CLK(n2691), .C(n2692) );
  CKBD0 U2574 ( .CLK(n2692), .C(n2693) );
  BUFFD0 U2575 ( .I(n2693), .Z(n2694) );
  CKBD0 U2576 ( .CLK(n2694), .C(n2695) );
  CKBD0 U2577 ( .CLK(n2695), .C(n2696) );
  CKBD0 U2578 ( .CLK(n2696), .C(n2697) );
  CKBD0 U2579 ( .CLK(n2697), .C(n2698) );
  CKBD0 U2580 ( .CLK(n2698), .C(n2699) );
  CKBD0 U2581 ( .CLK(n2699), .C(n2700) );
  CKBD0 U2582 ( .CLK(n2700), .C(n2701) );
  CKBD0 U2583 ( .CLK(n2701), .C(n2702) );
  CKBD0 U2584 ( .CLK(n2702), .C(n2703) );
  CKBD0 U2585 ( .CLK(n2703), .C(n2704) );
  BUFFD0 U2586 ( .I(n2704), .Z(n2705) );
  CKBD0 U2587 ( .CLK(n2705), .C(n2706) );
  CKBD0 U2588 ( .CLK(n2706), .C(n2707) );
  CKBD0 U2589 ( .CLK(n2707), .C(n2708) );
  CKBD0 U2590 ( .CLK(n2708), .C(n2709) );
  CKBD0 U2591 ( .CLK(n2709), .C(n2710) );
  CKBD0 U2592 ( .CLK(n2710), .C(n2711) );
  CKBD0 U2593 ( .CLK(n2711), .C(n2712) );
  CKBD0 U2594 ( .CLK(n2712), .C(n2713) );
  CKBD0 U2595 ( .CLK(n2713), .C(n2714) );
  CKBD0 U2596 ( .CLK(n2714), .C(n2715) );
  BUFFD0 U2597 ( .I(n2715), .Z(n2716) );
  CKBD0 U2598 ( .CLK(n2716), .C(n2717) );
  CKBD0 U2599 ( .CLK(n2717), .C(n2718) );
  CKBD0 U2600 ( .CLK(n2718), .C(n2719) );
  CKBD0 U2601 ( .CLK(n2719), .C(n2720) );
  CKBD0 U2602 ( .CLK(n2720), .C(n2721) );
  CKBD0 U2603 ( .CLK(n2721), .C(n2722) );
  CKBD0 U2604 ( .CLK(n2722), .C(n2723) );
  CKBD0 U2605 ( .CLK(n2723), .C(n2724) );
  CKBD0 U2606 ( .CLK(n2724), .C(n2725) );
  CKBD0 U2607 ( .CLK(n2725), .C(n2726) );
  BUFFD0 U2608 ( .I(n2726), .Z(n2727) );
  CKBD0 U2609 ( .CLK(n2727), .C(n2728) );
  CKBD0 U2610 ( .CLK(n2728), .C(n2729) );
  CKBD0 U2611 ( .CLK(n2729), .C(n2730) );
  CKBD0 U2612 ( .CLK(n2730), .C(n2731) );
  CKBD0 U2613 ( .CLK(n2731), .C(n2732) );
  CKBD0 U2614 ( .CLK(n2732), .C(n2733) );
  CKBD0 U2615 ( .CLK(n2733), .C(n2734) );
  CKBD0 U2616 ( .CLK(n2734), .C(n2735) );
  CKBD0 U2617 ( .CLK(n2735), .C(n2736) );
  CKBD0 U2618 ( .CLK(n2736), .C(n2737) );
  BUFFD0 U2619 ( .I(n2737), .Z(n2738) );
  CKBD0 U2620 ( .CLK(n2738), .C(n2739) );
  CKBD0 U2621 ( .CLK(n2739), .C(n2740) );
  CKBD0 U2622 ( .CLK(n2740), .C(n2741) );
  CKBD0 U2623 ( .CLK(n2741), .C(n2742) );
  CKBD0 U2624 ( .CLK(n2742), .C(n2743) );
  CKBD0 U2625 ( .CLK(n2743), .C(n2744) );
  CKBD0 U2626 ( .CLK(n2744), .C(n2745) );
  CKBD0 U2627 ( .CLK(n2745), .C(n2746) );
  CKBD0 U2628 ( .CLK(n2746), .C(n2747) );
  CKBD0 U2629 ( .CLK(n2747), .C(n2748) );
  BUFFD0 U2630 ( .I(n2748), .Z(n2749) );
  CKBD0 U2631 ( .CLK(n2749), .C(n2750) );
  CKBD0 U2632 ( .CLK(n2750), .C(n2751) );
  CKBD0 U2633 ( .CLK(n2751), .C(n2752) );
  CKBD0 U2634 ( .CLK(n2752), .C(n2753) );
  CKBD0 U2635 ( .CLK(n2753), .C(n2754) );
  CKBD0 U2636 ( .CLK(n2754), .C(n2755) );
  CKBD0 U2637 ( .CLK(n2755), .C(n2756) );
  CKBD0 U2638 ( .CLK(n2756), .C(n2757) );
  CKBD0 U2639 ( .CLK(n2757), .C(n2758) );
  BUFFD0 U2640 ( .I(n2758), .Z(n2759) );
  CKBD0 U2641 ( .CLK(n2759), .C(n2760) );
  CKBD0 U2642 ( .CLK(n2760), .C(n2761) );
  CKBD0 U2643 ( .CLK(n2761), .C(n2762) );
  CKBD0 U2644 ( .CLK(n2762), .C(n2763) );
  CKBD0 U2645 ( .CLK(n2763), .C(n2764) );
  CKBD0 U2646 ( .CLK(n2764), .C(n2765) );
  CKBD0 U2647 ( .CLK(n2765), .C(n2766) );
  CKBD0 U2648 ( .CLK(n2766), .C(n2767) );
  CKBD0 U2649 ( .CLK(n2767), .C(n2768) );
  CKBD0 U2650 ( .CLK(n2768), .C(n2769) );
  BUFFD0 U2651 ( .I(n2769), .Z(n2770) );
  CKBD0 U2652 ( .CLK(n2770), .C(n2771) );
  CKBD0 U2653 ( .CLK(n2771), .C(n2772) );
  CKBD0 U2654 ( .CLK(n2772), .C(n2773) );
  CKBD0 U2655 ( .CLK(n2773), .C(n2774) );
  CKBD0 U2656 ( .CLK(n2774), .C(n2775) );
  CKBD0 U2657 ( .CLK(n2775), .C(n2776) );
  CKBD0 U2658 ( .CLK(n2776), .C(n2777) );
  CKBD0 U2659 ( .CLK(n2777), .C(n2778) );
  CKBD0 U2660 ( .CLK(n2778), .C(n2779) );
  CKBD0 U2661 ( .CLK(n2779), .C(n2780) );
  BUFFD0 U2662 ( .I(n2780), .Z(n2781) );
  CKBD0 U2663 ( .CLK(n2781), .C(n2782) );
  CKBD0 U2664 ( .CLK(n2782), .C(n2783) );
  CKBD0 U2665 ( .CLK(n2783), .C(n2784) );
  CKBD0 U2666 ( .CLK(n2784), .C(n2785) );
  CKBD0 U2667 ( .CLK(n2785), .C(n2786) );
  CKBD0 U2668 ( .CLK(n2786), .C(n2787) );
  BUFFD0 U2669 ( .I(n2787), .Z(n2788) );
  CKBD0 U2670 ( .CLK(n2788), .C(n2789) );
  BUFFD0 U2671 ( .I(n2789), .Z(n2790) );
  CKBD0 U2672 ( .CLK(n2790), .C(n2791) );
  BUFFD0 U2673 ( .I(n2791), .Z(n2792) );
  CKBD0 U2674 ( .CLK(n2792), .C(n2793) );
  BUFFD0 U2675 ( .I(n2793), .Z(n2794) );
  CKBD0 U2676 ( .CLK(n2794), .C(n2795) );
  BUFFD0 U2677 ( .I(n2795), .Z(n2796) );
  CKBD0 U2678 ( .CLK(n2796), .C(n2797) );
  BUFFD0 U2679 ( .I(n2797), .Z(n2798) );
  CKBD0 U2680 ( .CLK(n2798), .C(n2799) );
  BUFFD0 U2681 ( .I(n2799), .Z(n2800) );
  CKBD0 U2682 ( .CLK(n2800), .C(n2801) );
  BUFFD0 U2683 ( .I(n2801), .Z(n2802) );
  BUFFD0 U2684 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2685 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2686 ( .I(n162), .Z(n2805) );
  CKBD0 U2687 ( .CLK(n1352), .C(n2806) );
  CKBD0 U2688 ( .CLK(n2806), .C(n2807) );
  CKBD0 U2689 ( .CLK(n2807), .C(n2808) );
  BUFFD0 U2690 ( .I(n2808), .Z(n2809) );
  CKBD0 U2691 ( .CLK(n2809), .C(n2810) );
  CKBD0 U2692 ( .CLK(n2810), .C(n2811) );
  CKBD0 U2693 ( .CLK(n2811), .C(n2812) );
  CKBD0 U2694 ( .CLK(n2812), .C(n2813) );
  CKBD0 U2695 ( .CLK(n2813), .C(n2814) );
  CKBD0 U2696 ( .CLK(n2814), .C(n2815) );
  CKBD0 U2697 ( .CLK(n2815), .C(n2816) );
  CKBD0 U2698 ( .CLK(n2816), .C(n2817) );
  CKBD0 U2699 ( .CLK(n2817), .C(n2818) );
  CKBD0 U2700 ( .CLK(n2818), .C(n2819) );
  BUFFD0 U2701 ( .I(n2819), .Z(n2820) );
  CKBD0 U2702 ( .CLK(n2820), .C(n2821) );
  CKBD0 U2703 ( .CLK(n2821), .C(n2822) );
  CKBD0 U2704 ( .CLK(n2822), .C(n2823) );
  CKBD0 U2705 ( .CLK(n2823), .C(n2824) );
  CKBD0 U2706 ( .CLK(n2824), .C(n2825) );
  CKBD0 U2707 ( .CLK(n2825), .C(n2826) );
  CKBD0 U2708 ( .CLK(n2826), .C(n2827) );
  CKBD0 U2709 ( .CLK(n2827), .C(n2828) );
  CKBD0 U2710 ( .CLK(n2828), .C(n2829) );
  BUFFD0 U2711 ( .I(n2829), .Z(n2830) );
  CKBD0 U2712 ( .CLK(n2830), .C(n2831) );
  CKBD0 U2713 ( .CLK(n2831), .C(n2832) );
  CKBD0 U2714 ( .CLK(n2832), .C(n2833) );
  CKBD0 U2715 ( .CLK(n2833), .C(n2834) );
  CKBD0 U2716 ( .CLK(n2834), .C(n2835) );
  CKBD0 U2717 ( .CLK(n2835), .C(n2836) );
  CKBD0 U2718 ( .CLK(n2836), .C(n2837) );
  CKBD0 U2719 ( .CLK(n2837), .C(n2838) );
  CKBD0 U2720 ( .CLK(n2838), .C(n2839) );
  CKBD0 U2721 ( .CLK(n2839), .C(n2840) );
  BUFFD0 U2722 ( .I(n2840), .Z(n2841) );
  CKBD0 U2723 ( .CLK(n2841), .C(n2842) );
  CKBD0 U2724 ( .CLK(n2842), .C(n2843) );
  CKBD0 U2725 ( .CLK(n2843), .C(n2844) );
  CKBD0 U2726 ( .CLK(n2844), .C(n2845) );
  CKBD0 U2727 ( .CLK(n2845), .C(n2846) );
  CKBD0 U2728 ( .CLK(n2846), .C(n2847) );
  CKBD0 U2729 ( .CLK(n2847), .C(n2848) );
  CKBD0 U2730 ( .CLK(n2848), .C(n2849) );
  CKBD0 U2731 ( .CLK(n2849), .C(n2850) );
  CKBD0 U2732 ( .CLK(n2850), .C(n2851) );
  BUFFD0 U2733 ( .I(n2851), .Z(n2852) );
  CKBD0 U2734 ( .CLK(n2852), .C(n2853) );
  CKBD0 U2735 ( .CLK(n2853), .C(n2854) );
  CKBD0 U2736 ( .CLK(n2854), .C(n2855) );
  CKBD0 U2737 ( .CLK(n2855), .C(n2856) );
  CKBD0 U2738 ( .CLK(n2856), .C(n2857) );
  CKBD0 U2739 ( .CLK(n2857), .C(n2858) );
  CKBD0 U2740 ( .CLK(n2858), .C(n2859) );
  CKBD0 U2741 ( .CLK(n2859), .C(n2860) );
  CKBD0 U2742 ( .CLK(n2860), .C(n2861) );
  CKBD0 U2743 ( .CLK(n2861), .C(n2862) );
  BUFFD0 U2744 ( .I(n2862), .Z(n2863) );
  CKBD0 U2745 ( .CLK(n2863), .C(n2864) );
  CKBD0 U2746 ( .CLK(n2864), .C(n2865) );
  CKBD0 U2747 ( .CLK(n2865), .C(n2866) );
  CKBD0 U2748 ( .CLK(n2866), .C(n2867) );
  CKBD0 U2749 ( .CLK(n2867), .C(n2868) );
  CKBD0 U2750 ( .CLK(n2868), .C(n2869) );
  CKBD0 U2751 ( .CLK(n2869), .C(n2870) );
  CKBD0 U2752 ( .CLK(n2870), .C(n2871) );
  CKBD0 U2753 ( .CLK(n2871), .C(n2872) );
  CKBD0 U2754 ( .CLK(n2872), .C(n2873) );
  BUFFD0 U2755 ( .I(n2873), .Z(n2874) );
  CKBD0 U2756 ( .CLK(n2874), .C(n2875) );
  CKBD0 U2757 ( .CLK(n2875), .C(n2876) );
  CKBD0 U2758 ( .CLK(n2876), .C(n2877) );
  CKBD0 U2759 ( .CLK(n2877), .C(n2878) );
  CKBD0 U2760 ( .CLK(n2878), .C(n2879) );
  CKBD0 U2761 ( .CLK(n2879), .C(n2880) );
  CKBD0 U2762 ( .CLK(n2880), .C(n2881) );
  CKBD0 U2763 ( .CLK(n2881), .C(n2882) );
  CKBD0 U2764 ( .CLK(n2882), .C(n2883) );
  CKBD0 U2765 ( .CLK(n2883), .C(n2884) );
  BUFFD0 U2766 ( .I(n2884), .Z(n2885) );
  CKBD0 U2767 ( .CLK(n2885), .C(n2886) );
  CKBD0 U2768 ( .CLK(n2886), .C(n2887) );
  CKBD0 U2769 ( .CLK(n2887), .C(n2888) );
  CKBD0 U2770 ( .CLK(n2888), .C(n2889) );
  CKBD0 U2771 ( .CLK(n2889), .C(n2890) );
  CKBD0 U2772 ( .CLK(n2890), .C(n2891) );
  CKBD0 U2773 ( .CLK(n2891), .C(n2892) );
  CKBD0 U2774 ( .CLK(n2892), .C(n2893) );
  CKBD0 U2775 ( .CLK(n2893), .C(n2894) );
  BUFFD0 U2776 ( .I(n2894), .Z(n2895) );
  CKBD0 U2777 ( .CLK(n2895), .C(n2896) );
  CKBD0 U2778 ( .CLK(n2896), .C(n2897) );
  CKBD0 U2779 ( .CLK(n2897), .C(n2898) );
  CKBD0 U2780 ( .CLK(n2898), .C(n2899) );
  CKBD0 U2781 ( .CLK(n2899), .C(n2900) );
  CKBD0 U2782 ( .CLK(n2900), .C(n2901) );
  CKBD0 U2783 ( .CLK(n2901), .C(n2902) );
  CKBD0 U2784 ( .CLK(n2902), .C(n2903) );
  CKBD0 U2785 ( .CLK(n2903), .C(n2904) );
  CKBD0 U2786 ( .CLK(n2904), .C(n2905) );
  BUFFD0 U2787 ( .I(n2905), .Z(n2906) );
  CKBD0 U2788 ( .CLK(n2906), .C(n2907) );
  CKBD0 U2789 ( .CLK(n2907), .C(n2908) );
  CKBD0 U2790 ( .CLK(n2908), .C(n2909) );
  CKBD0 U2791 ( .CLK(n2909), .C(n2910) );
  CKBD0 U2792 ( .CLK(n2910), .C(n2911) );
  CKBD0 U2793 ( .CLK(n2911), .C(n2912) );
  CKBD0 U2794 ( .CLK(n2912), .C(n2913) );
  CKBD0 U2795 ( .CLK(n2913), .C(n2914) );
  CKBD0 U2796 ( .CLK(n2914), .C(n2915) );
  CKBD0 U2797 ( .CLK(n2915), .C(n2916) );
  BUFFD0 U2798 ( .I(n2916), .Z(n2917) );
  CKBD0 U2799 ( .CLK(n2917), .C(n2918) );
  CKBD0 U2800 ( .CLK(n2918), .C(n2919) );
  CKBD0 U2801 ( .CLK(n2919), .C(n2920) );
  CKBD0 U2802 ( .CLK(n2920), .C(n2921) );
  CKBD0 U2803 ( .CLK(n2921), .C(n2922) );
  CKBD0 U2804 ( .CLK(n2922), .C(n2923) );
  BUFFD0 U2805 ( .I(n2923), .Z(n2924) );
  CKBD0 U2806 ( .CLK(n2924), .C(n2925) );
  BUFFD0 U2807 ( .I(n2925), .Z(n2926) );
  CKBD0 U2808 ( .CLK(n2926), .C(n2927) );
  BUFFD0 U2809 ( .I(n2927), .Z(n2928) );
  CKBD0 U2810 ( .CLK(n2928), .C(n2929) );
  BUFFD0 U2811 ( .I(n2929), .Z(n2930) );
  CKBD0 U2812 ( .CLK(n2930), .C(n2931) );
  BUFFD0 U2813 ( .I(n2931), .Z(n2932) );
  CKBD0 U2814 ( .CLK(n2932), .C(n2933) );
  BUFFD0 U2815 ( .I(n2933), .Z(n2934) );
  CKBD0 U2816 ( .CLK(n2934), .C(n2935) );
  BUFFD0 U2817 ( .I(n2935), .Z(n2936) );
  CKBD0 U2818 ( .CLK(n2936), .C(n2937) );
  BUFFD0 U2819 ( .I(n2937), .Z(n2938) );
  BUFFD0 U2820 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2821 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2822 ( .I(n161), .Z(n2941) );
  CKBD0 U2823 ( .CLK(n1350), .C(n2942) );
  CKBD0 U2824 ( .CLK(n2942), .C(n2943) );
  CKBD0 U2825 ( .CLK(n2943), .C(n2944) );
  BUFFD0 U2826 ( .I(n2944), .Z(n2945) );
  CKBD0 U2827 ( .CLK(n2945), .C(n2946) );
  CKBD0 U2828 ( .CLK(n2946), .C(n2947) );
  CKBD0 U2829 ( .CLK(n2947), .C(n2948) );
  CKBD0 U2830 ( .CLK(n2948), .C(n2949) );
  CKBD0 U2831 ( .CLK(n2949), .C(n2950) );
  CKBD0 U2832 ( .CLK(n2950), .C(n2951) );
  CKBD0 U2833 ( .CLK(n2951), .C(n2952) );
  CKBD0 U2834 ( .CLK(n2952), .C(n2953) );
  CKBD0 U2835 ( .CLK(n2953), .C(n2954) );
  CKBD0 U2836 ( .CLK(n2954), .C(n2955) );
  BUFFD0 U2837 ( .I(n2955), .Z(n2956) );
  CKBD0 U2838 ( .CLK(n2956), .C(n2957) );
  CKBD0 U2839 ( .CLK(n2957), .C(n2958) );
  CKBD0 U2840 ( .CLK(n2958), .C(n2959) );
  CKBD0 U2841 ( .CLK(n2959), .C(n2960) );
  CKBD0 U2842 ( .CLK(n2960), .C(n2961) );
  CKBD0 U2843 ( .CLK(n2961), .C(n2962) );
  CKBD0 U2844 ( .CLK(n2962), .C(n2963) );
  CKBD0 U2845 ( .CLK(n2963), .C(n2964) );
  CKBD0 U2846 ( .CLK(n2964), .C(n2965) );
  BUFFD0 U2847 ( .I(n2965), .Z(n2966) );
  CKBD0 U2848 ( .CLK(n2966), .C(n2967) );
  CKBD0 U2849 ( .CLK(n2967), .C(n2968) );
  CKBD0 U2850 ( .CLK(n2968), .C(n2969) );
  CKBD0 U2851 ( .CLK(n2969), .C(n2970) );
  CKBD0 U2852 ( .CLK(n2970), .C(n2971) );
  CKBD0 U2853 ( .CLK(n2971), .C(n2972) );
  CKBD0 U2854 ( .CLK(n2972), .C(n2973) );
  CKBD0 U2855 ( .CLK(n2973), .C(n2974) );
  CKBD0 U2856 ( .CLK(n2974), .C(n2975) );
  CKBD0 U2857 ( .CLK(n2975), .C(n2976) );
  BUFFD0 U2858 ( .I(n2976), .Z(n2977) );
  CKBD0 U2859 ( .CLK(n2977), .C(n2978) );
  CKBD0 U2860 ( .CLK(n2978), .C(n2979) );
  CKBD0 U2861 ( .CLK(n2979), .C(n2980) );
  CKBD0 U2862 ( .CLK(n2980), .C(n2981) );
  CKBD0 U2863 ( .CLK(n2981), .C(n2982) );
  CKBD0 U2864 ( .CLK(n2982), .C(n2983) );
  CKBD0 U2865 ( .CLK(n2983), .C(n2984) );
  CKBD0 U2866 ( .CLK(n2984), .C(n2985) );
  CKBD0 U2867 ( .CLK(n2985), .C(n2986) );
  CKBD0 U2868 ( .CLK(n2986), .C(n2987) );
  BUFFD0 U2869 ( .I(n2987), .Z(n2988) );
  CKBD0 U2870 ( .CLK(n2988), .C(n2989) );
  CKBD0 U2871 ( .CLK(n2989), .C(n2990) );
  CKBD0 U2872 ( .CLK(n2990), .C(n2991) );
  CKBD0 U2873 ( .CLK(n2991), .C(n2992) );
  CKBD0 U2874 ( .CLK(n2992), .C(n2993) );
  CKBD0 U2875 ( .CLK(n2993), .C(n2994) );
  CKBD0 U2876 ( .CLK(n2994), .C(n2995) );
  CKBD0 U2877 ( .CLK(n2995), .C(n2996) );
  CKBD0 U2878 ( .CLK(n2996), .C(n2997) );
  CKBD0 U2879 ( .CLK(n2997), .C(n2998) );
  BUFFD0 U2880 ( .I(n2998), .Z(n2999) );
  CKBD0 U2881 ( .CLK(n2999), .C(n3000) );
  CKBD0 U2882 ( .CLK(n3000), .C(n3001) );
  CKBD0 U2883 ( .CLK(n3001), .C(n3002) );
  CKBD0 U2884 ( .CLK(n3002), .C(n3003) );
  CKBD0 U2885 ( .CLK(n3003), .C(n3004) );
  CKBD0 U2886 ( .CLK(n3004), .C(n3005) );
  CKBD0 U2887 ( .CLK(n3005), .C(n3006) );
  CKBD0 U2888 ( .CLK(n3006), .C(n3007) );
  CKBD0 U2889 ( .CLK(n3007), .C(n3008) );
  CKBD0 U2890 ( .CLK(n3008), .C(n3009) );
  BUFFD0 U2891 ( .I(n3009), .Z(n3010) );
  CKBD0 U2892 ( .CLK(n3010), .C(n3011) );
  CKBD0 U2893 ( .CLK(n3011), .C(n3012) );
  CKBD0 U2894 ( .CLK(n3012), .C(n3013) );
  CKBD0 U2895 ( .CLK(n3013), .C(n3014) );
  CKBD0 U2896 ( .CLK(n3014), .C(n3015) );
  CKBD0 U2897 ( .CLK(n3015), .C(n3016) );
  CKBD0 U2898 ( .CLK(n3016), .C(n3017) );
  CKBD0 U2899 ( .CLK(n3017), .C(n3018) );
  CKBD0 U2900 ( .CLK(n3018), .C(n3019) );
  CKBD0 U2901 ( .CLK(n3019), .C(n3020) );
  BUFFD0 U2902 ( .I(n3020), .Z(n3021) );
  CKBD0 U2903 ( .CLK(n3021), .C(n3022) );
  CKBD0 U2904 ( .CLK(n3022), .C(n3023) );
  CKBD0 U2905 ( .CLK(n3023), .C(n3024) );
  CKBD0 U2906 ( .CLK(n3024), .C(n3025) );
  CKBD0 U2907 ( .CLK(n3025), .C(n3026) );
  CKBD0 U2908 ( .CLK(n3026), .C(n3027) );
  CKBD0 U2909 ( .CLK(n3027), .C(n3028) );
  CKBD0 U2910 ( .CLK(n3028), .C(n3029) );
  CKBD0 U2911 ( .CLK(n3029), .C(n3030) );
  BUFFD0 U2912 ( .I(n3030), .Z(n3031) );
  CKBD0 U2913 ( .CLK(n3031), .C(n3032) );
  CKBD0 U2914 ( .CLK(n3032), .C(n3033) );
  CKBD0 U2915 ( .CLK(n3033), .C(n3034) );
  CKBD0 U2916 ( .CLK(n3034), .C(n3035) );
  CKBD0 U2917 ( .CLK(n3035), .C(n3036) );
  CKBD0 U2918 ( .CLK(n3036), .C(n3037) );
  CKBD0 U2919 ( .CLK(n3037), .C(n3038) );
  CKBD0 U2920 ( .CLK(n3038), .C(n3039) );
  CKBD0 U2921 ( .CLK(n3039), .C(n3040) );
  CKBD0 U2922 ( .CLK(n3040), .C(n3041) );
  BUFFD0 U2923 ( .I(n3041), .Z(n3042) );
  CKBD0 U2924 ( .CLK(n3042), .C(n3043) );
  CKBD0 U2925 ( .CLK(n3043), .C(n3044) );
  CKBD0 U2926 ( .CLK(n3044), .C(n3045) );
  CKBD0 U2927 ( .CLK(n3045), .C(n3046) );
  CKBD0 U2928 ( .CLK(n3046), .C(n3047) );
  CKBD0 U2929 ( .CLK(n3047), .C(n3048) );
  CKBD0 U2930 ( .CLK(n3048), .C(n3049) );
  CKBD0 U2931 ( .CLK(n3049), .C(n3050) );
  CKBD0 U2932 ( .CLK(n3050), .C(n3051) );
  CKBD0 U2933 ( .CLK(n3051), .C(n3052) );
  BUFFD0 U2934 ( .I(n3052), .Z(n3053) );
  CKBD0 U2935 ( .CLK(n3053), .C(n3054) );
  CKBD0 U2936 ( .CLK(n3054), .C(n3055) );
  CKBD0 U2937 ( .CLK(n3055), .C(n3056) );
  CKBD0 U2938 ( .CLK(n3056), .C(n3057) );
  CKBD0 U2939 ( .CLK(n3057), .C(n3058) );
  CKBD0 U2940 ( .CLK(n3058), .C(n3059) );
  BUFFD0 U2941 ( .I(n3059), .Z(n3060) );
  CKBD0 U2942 ( .CLK(n3060), .C(n3061) );
  BUFFD0 U2943 ( .I(n3061), .Z(n3062) );
  CKBD0 U2944 ( .CLK(n3062), .C(n3063) );
  BUFFD0 U2945 ( .I(n3063), .Z(n3064) );
  CKBD0 U2946 ( .CLK(n3064), .C(n3065) );
  BUFFD0 U2947 ( .I(n3065), .Z(n3066) );
  CKBD0 U2948 ( .CLK(n3066), .C(n3067) );
  BUFFD0 U2949 ( .I(n3067), .Z(n3068) );
  CKBD0 U2950 ( .CLK(n3068), .C(n3069) );
  BUFFD0 U2951 ( .I(n3069), .Z(n3070) );
  CKBD0 U2952 ( .CLK(n3070), .C(n3071) );
  BUFFD0 U2953 ( .I(n3071), .Z(n3072) );
  CKBD0 U2954 ( .CLK(n3072), .C(n3073) );
  BUFFD0 U2955 ( .I(n3073), .Z(n3074) );
  BUFFD0 U2956 ( .I(n3076), .Z(n3075) );
  BUFFD0 U2957 ( .I(n3077), .Z(n3076) );
  BUFFD0 U2958 ( .I(n160), .Z(n3077) );
  CKBD0 U2959 ( .CLK(n1348), .C(n3078) );
  CKBD0 U2960 ( .CLK(n3078), .C(n3079) );
  CKBD0 U2961 ( .CLK(n3079), .C(n3080) );
  BUFFD0 U2962 ( .I(n3080), .Z(n3081) );
  CKBD0 U2963 ( .CLK(n3081), .C(n3082) );
  CKBD0 U2964 ( .CLK(n3082), .C(n3083) );
  CKBD0 U2965 ( .CLK(n3083), .C(n3084) );
  CKBD0 U2966 ( .CLK(n3084), .C(n3085) );
  CKBD0 U2967 ( .CLK(n3085), .C(n3086) );
  CKBD0 U2968 ( .CLK(n3086), .C(n3087) );
  CKBD0 U2969 ( .CLK(n3087), .C(n3088) );
  CKBD0 U2970 ( .CLK(n3088), .C(n3089) );
  CKBD0 U2971 ( .CLK(n3089), .C(n3090) );
  CKBD0 U2972 ( .CLK(n3090), .C(n3091) );
  BUFFD0 U2973 ( .I(n3091), .Z(n3092) );
  CKBD0 U2974 ( .CLK(n3092), .C(n3093) );
  CKBD0 U2975 ( .CLK(n3093), .C(n3094) );
  CKBD0 U2976 ( .CLK(n3094), .C(n3095) );
  CKBD0 U2977 ( .CLK(n3095), .C(n3096) );
  CKBD0 U2978 ( .CLK(n3096), .C(n3097) );
  CKBD0 U2979 ( .CLK(n3097), .C(n3098) );
  CKBD0 U2980 ( .CLK(n3098), .C(n3099) );
  CKBD0 U2981 ( .CLK(n3099), .C(n3100) );
  CKBD0 U2982 ( .CLK(n3100), .C(n3101) );
  BUFFD0 U2983 ( .I(n3101), .Z(n3102) );
  CKBD0 U2984 ( .CLK(n3102), .C(n3103) );
  CKBD0 U2985 ( .CLK(n3103), .C(n3104) );
  CKBD0 U2986 ( .CLK(n3104), .C(n3105) );
  CKBD0 U2987 ( .CLK(n3105), .C(n3106) );
  CKBD0 U2988 ( .CLK(n3106), .C(n3107) );
  CKBD0 U2989 ( .CLK(n3107), .C(n3108) );
  CKBD0 U2990 ( .CLK(n3108), .C(n3109) );
  CKBD0 U2991 ( .CLK(n3109), .C(n3110) );
  CKBD0 U2992 ( .CLK(n3110), .C(n3111) );
  CKBD0 U2993 ( .CLK(n3111), .C(n3112) );
  BUFFD0 U2994 ( .I(n3112), .Z(n3113) );
  CKBD0 U2995 ( .CLK(n3113), .C(n3114) );
  CKBD0 U2996 ( .CLK(n3114), .C(n3115) );
  CKBD0 U2997 ( .CLK(n3115), .C(n3116) );
  CKBD0 U2998 ( .CLK(n3116), .C(n3117) );
  CKBD0 U2999 ( .CLK(n3117), .C(n3118) );
  CKBD0 U3000 ( .CLK(n3118), .C(n3119) );
  CKBD0 U3001 ( .CLK(n3119), .C(n3120) );
  CKBD0 U3002 ( .CLK(n3120), .C(n3121) );
  CKBD0 U3003 ( .CLK(n3121), .C(n3122) );
  CKBD0 U3004 ( .CLK(n3122), .C(n3123) );
  BUFFD0 U3005 ( .I(n3123), .Z(n3124) );
  CKBD0 U3006 ( .CLK(n3124), .C(n3125) );
  CKBD0 U3007 ( .CLK(n3125), .C(n3126) );
  CKBD0 U3008 ( .CLK(n3126), .C(n3127) );
  CKBD0 U3009 ( .CLK(n3127), .C(n3128) );
  CKBD0 U3010 ( .CLK(n3128), .C(n3129) );
  CKBD0 U3011 ( .CLK(n3129), .C(n3130) );
  CKBD0 U3012 ( .CLK(n3130), .C(n3131) );
  CKBD0 U3013 ( .CLK(n3131), .C(n3132) );
  CKBD0 U3014 ( .CLK(n3132), .C(n3133) );
  CKBD0 U3015 ( .CLK(n3133), .C(n3134) );
  BUFFD0 U3016 ( .I(n3134), .Z(n3135) );
  CKBD0 U3017 ( .CLK(n3135), .C(n3136) );
  CKBD0 U3018 ( .CLK(n3136), .C(n3137) );
  CKBD0 U3019 ( .CLK(n3137), .C(n3138) );
  CKBD0 U3020 ( .CLK(n3138), .C(n3139) );
  CKBD0 U3021 ( .CLK(n3139), .C(n3140) );
  CKBD0 U3022 ( .CLK(n3140), .C(n3141) );
  CKBD0 U3023 ( .CLK(n3141), .C(n3142) );
  CKBD0 U3024 ( .CLK(n3142), .C(n3143) );
  CKBD0 U3025 ( .CLK(n3143), .C(n3144) );
  CKBD0 U3026 ( .CLK(n3144), .C(n3145) );
  BUFFD0 U3027 ( .I(n3145), .Z(n3146) );
  CKBD0 U3028 ( .CLK(n3146), .C(n3147) );
  CKBD0 U3029 ( .CLK(n3147), .C(n3148) );
  CKBD0 U3030 ( .CLK(n3148), .C(n3149) );
  CKBD0 U3031 ( .CLK(n3149), .C(n3150) );
  CKBD0 U3032 ( .CLK(n3150), .C(n3151) );
  CKBD0 U3033 ( .CLK(n3151), .C(n3152) );
  CKBD0 U3034 ( .CLK(n3152), .C(n3153) );
  CKBD0 U3035 ( .CLK(n3153), .C(n3154) );
  CKBD0 U3036 ( .CLK(n3154), .C(n3155) );
  CKBD0 U3037 ( .CLK(n3155), .C(n3156) );
  BUFFD0 U3038 ( .I(n3156), .Z(n3157) );
  CKBD0 U3039 ( .CLK(n3157), .C(n3158) );
  CKBD0 U3040 ( .CLK(n3158), .C(n3159) );
  CKBD0 U3041 ( .CLK(n3159), .C(n3160) );
  CKBD0 U3042 ( .CLK(n3160), .C(n3161) );
  CKBD0 U3043 ( .CLK(n3161), .C(n3162) );
  CKBD0 U3044 ( .CLK(n3162), .C(n3163) );
  CKBD0 U3045 ( .CLK(n3163), .C(n3164) );
  CKBD0 U3046 ( .CLK(n3164), .C(n3165) );
  CKBD0 U3047 ( .CLK(n3165), .C(n3166) );
  BUFFD0 U3048 ( .I(n3166), .Z(n3167) );
  CKBD0 U3049 ( .CLK(n3167), .C(n3168) );
  CKBD0 U3050 ( .CLK(n3168), .C(n3169) );
  CKBD0 U3051 ( .CLK(n3169), .C(n3170) );
  CKBD0 U3052 ( .CLK(n3170), .C(n3171) );
  CKBD0 U3053 ( .CLK(n3171), .C(n3172) );
  CKBD0 U3054 ( .CLK(n3172), .C(n3173) );
  CKBD0 U3055 ( .CLK(n3173), .C(n3174) );
  CKBD0 U3056 ( .CLK(n3174), .C(n3175) );
  CKBD0 U3057 ( .CLK(n3175), .C(n3176) );
  CKBD0 U3058 ( .CLK(n3176), .C(n3177) );
  BUFFD0 U3059 ( .I(n3177), .Z(n3178) );
  CKBD0 U3060 ( .CLK(n3178), .C(n3179) );
  CKBD0 U3061 ( .CLK(n3179), .C(n3180) );
  CKBD0 U3062 ( .CLK(n3180), .C(n3181) );
  CKBD0 U3063 ( .CLK(n3181), .C(n3182) );
  CKBD0 U3064 ( .CLK(n3182), .C(n3183) );
  CKBD0 U3065 ( .CLK(n3183), .C(n3184) );
  CKBD0 U3066 ( .CLK(n3184), .C(n3185) );
  CKBD0 U3067 ( .CLK(n3185), .C(n3186) );
  CKBD0 U3068 ( .CLK(n3186), .C(n3187) );
  CKBD0 U3069 ( .CLK(n3187), .C(n3188) );
  BUFFD0 U3070 ( .I(n3188), .Z(n3189) );
  CKBD0 U3071 ( .CLK(n3189), .C(n3190) );
  CKBD0 U3072 ( .CLK(n3190), .C(n3191) );
  CKBD0 U3073 ( .CLK(n3191), .C(n3192) );
  CKBD0 U3074 ( .CLK(n3192), .C(n3193) );
  CKBD0 U3075 ( .CLK(n3193), .C(n3194) );
  CKBD0 U3076 ( .CLK(n3194), .C(n3195) );
  BUFFD0 U3077 ( .I(n3195), .Z(n3196) );
  CKBD0 U3078 ( .CLK(n3196), .C(n3197) );
  BUFFD0 U3079 ( .I(n3197), .Z(n3198) );
  CKBD0 U3080 ( .CLK(n3198), .C(n3199) );
  BUFFD0 U3081 ( .I(n3199), .Z(n3200) );
  CKBD0 U3082 ( .CLK(n3200), .C(n3201) );
  BUFFD0 U3083 ( .I(n3201), .Z(n3202) );
  CKBD0 U3084 ( .CLK(n3202), .C(n3203) );
  BUFFD0 U3085 ( .I(n3203), .Z(n3204) );
  CKBD0 U3086 ( .CLK(n3204), .C(n3205) );
  BUFFD0 U3087 ( .I(n3205), .Z(n3206) );
  CKBD0 U3088 ( .CLK(n3206), .C(n3207) );
  BUFFD0 U3089 ( .I(n3207), .Z(n3208) );
  CKBD0 U3090 ( .CLK(n3208), .C(n3209) );
  BUFFD0 U3091 ( .I(n3209), .Z(n3210) );
  BUFFD0 U3092 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3093 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3094 ( .I(n159), .Z(n3213) );
  CKBD0 U3095 ( .CLK(n1346), .C(n3214) );
  CKBD0 U3096 ( .CLK(n3214), .C(n3215) );
  CKBD0 U3097 ( .CLK(n3215), .C(n3216) );
  BUFFD0 U3098 ( .I(n3216), .Z(n3217) );
  CKBD0 U3099 ( .CLK(n3217), .C(n3218) );
  CKBD0 U3100 ( .CLK(n3218), .C(n3219) );
  CKBD0 U3101 ( .CLK(n3219), .C(n3220) );
  CKBD0 U3102 ( .CLK(n3220), .C(n3221) );
  CKBD0 U3103 ( .CLK(n3221), .C(n3222) );
  CKBD0 U3104 ( .CLK(n3222), .C(n3223) );
  CKBD0 U3105 ( .CLK(n3223), .C(n3224) );
  CKBD0 U3106 ( .CLK(n3224), .C(n3225) );
  CKBD0 U3107 ( .CLK(n3225), .C(n3226) );
  CKBD0 U3108 ( .CLK(n3226), .C(n3227) );
  BUFFD0 U3109 ( .I(n3227), .Z(n3228) );
  CKBD0 U3110 ( .CLK(n3228), .C(n3229) );
  CKBD0 U3111 ( .CLK(n3229), .C(n3230) );
  CKBD0 U3112 ( .CLK(n3230), .C(n3231) );
  CKBD0 U3113 ( .CLK(n3231), .C(n3232) );
  CKBD0 U3114 ( .CLK(n3232), .C(n3233) );
  CKBD0 U3115 ( .CLK(n3233), .C(n3234) );
  CKBD0 U3116 ( .CLK(n3234), .C(n3235) );
  CKBD0 U3117 ( .CLK(n3235), .C(n3236) );
  CKBD0 U3118 ( .CLK(n3236), .C(n3237) );
  BUFFD0 U3119 ( .I(n3237), .Z(n3238) );
  CKBD0 U3120 ( .CLK(n3238), .C(n3239) );
  CKBD0 U3121 ( .CLK(n3239), .C(n3240) );
  CKBD0 U3122 ( .CLK(n3240), .C(n3241) );
  CKBD0 U3123 ( .CLK(n3241), .C(n3242) );
  CKBD0 U3124 ( .CLK(n3242), .C(n3243) );
  CKBD0 U3125 ( .CLK(n3243), .C(n3244) );
  CKBD0 U3126 ( .CLK(n3244), .C(n3245) );
  CKBD0 U3127 ( .CLK(n3245), .C(n3246) );
  CKBD0 U3128 ( .CLK(n3246), .C(n3247) );
  CKBD0 U3129 ( .CLK(n3247), .C(n3248) );
  BUFFD0 U3130 ( .I(n3248), .Z(n3249) );
  CKBD0 U3131 ( .CLK(n3249), .C(n3250) );
  CKBD0 U3132 ( .CLK(n3250), .C(n3251) );
  CKBD0 U3133 ( .CLK(n3251), .C(n3252) );
  CKBD0 U3134 ( .CLK(n3252), .C(n3253) );
  CKBD0 U3135 ( .CLK(n3253), .C(n3254) );
  CKBD0 U3136 ( .CLK(n3254), .C(n3255) );
  CKBD0 U3137 ( .CLK(n3255), .C(n3256) );
  CKBD0 U3138 ( .CLK(n3256), .C(n3257) );
  CKBD0 U3139 ( .CLK(n3257), .C(n3258) );
  CKBD0 U3140 ( .CLK(n3258), .C(n3259) );
  BUFFD0 U3141 ( .I(n3259), .Z(n3260) );
  CKBD0 U3142 ( .CLK(n3260), .C(n3261) );
  CKBD0 U3143 ( .CLK(n3261), .C(n3262) );
  CKBD0 U3144 ( .CLK(n3262), .C(n3263) );
  CKBD0 U3145 ( .CLK(n3263), .C(n3264) );
  CKBD0 U3146 ( .CLK(n3264), .C(n3265) );
  CKBD0 U3147 ( .CLK(n3265), .C(n3266) );
  CKBD0 U3148 ( .CLK(n3266), .C(n3267) );
  CKBD0 U3149 ( .CLK(n3267), .C(n3268) );
  CKBD0 U3150 ( .CLK(n3268), .C(n3269) );
  CKBD0 U3151 ( .CLK(n3269), .C(n3270) );
  BUFFD0 U3152 ( .I(n3270), .Z(n3271) );
  CKBD0 U3153 ( .CLK(n3271), .C(n3272) );
  CKBD0 U3154 ( .CLK(n3272), .C(n3273) );
  CKBD0 U3155 ( .CLK(n3273), .C(n3274) );
  CKBD0 U3156 ( .CLK(n3274), .C(n3275) );
  CKBD0 U3157 ( .CLK(n3275), .C(n3276) );
  CKBD0 U3158 ( .CLK(n3276), .C(n3277) );
  CKBD0 U3159 ( .CLK(n3277), .C(n3278) );
  CKBD0 U3160 ( .CLK(n3278), .C(n3279) );
  CKBD0 U3161 ( .CLK(n3279), .C(n3280) );
  CKBD0 U3162 ( .CLK(n3280), .C(n3281) );
  BUFFD0 U3163 ( .I(n3281), .Z(n3282) );
  CKBD0 U3164 ( .CLK(n3282), .C(n3283) );
  CKBD0 U3165 ( .CLK(n3283), .C(n3284) );
  CKBD0 U3166 ( .CLK(n3284), .C(n3285) );
  CKBD0 U3167 ( .CLK(n3285), .C(n3286) );
  CKBD0 U3168 ( .CLK(n3286), .C(n3287) );
  CKBD0 U3169 ( .CLK(n3287), .C(n3288) );
  CKBD0 U3170 ( .CLK(n3288), .C(n3289) );
  CKBD0 U3171 ( .CLK(n3289), .C(n3290) );
  CKBD0 U3172 ( .CLK(n3290), .C(n3291) );
  CKBD0 U3173 ( .CLK(n3291), .C(n3292) );
  BUFFD0 U3174 ( .I(n3292), .Z(n3293) );
  CKBD0 U3175 ( .CLK(n3293), .C(n3294) );
  CKBD0 U3176 ( .CLK(n3294), .C(n3295) );
  CKBD0 U3177 ( .CLK(n3295), .C(n3296) );
  CKBD0 U3178 ( .CLK(n3296), .C(n3297) );
  CKBD0 U3179 ( .CLK(n3297), .C(n3298) );
  CKBD0 U3180 ( .CLK(n3298), .C(n3299) );
  CKBD0 U3181 ( .CLK(n3299), .C(n3300) );
  CKBD0 U3182 ( .CLK(n3300), .C(n3301) );
  CKBD0 U3183 ( .CLK(n3301), .C(n3302) );
  BUFFD0 U3184 ( .I(n3302), .Z(n3303) );
  CKBD0 U3185 ( .CLK(n3303), .C(n3304) );
  CKBD0 U3186 ( .CLK(n3304), .C(n3305) );
  CKBD0 U3187 ( .CLK(n3305), .C(n3306) );
  CKBD0 U3188 ( .CLK(n3306), .C(n3307) );
  CKBD0 U3189 ( .CLK(n3307), .C(n3308) );
  CKBD0 U3190 ( .CLK(n3308), .C(n3309) );
  CKBD0 U3191 ( .CLK(n3309), .C(n3310) );
  CKBD0 U3192 ( .CLK(n3310), .C(n3311) );
  CKBD0 U3193 ( .CLK(n3311), .C(n3312) );
  CKBD0 U3194 ( .CLK(n3312), .C(n3313) );
  BUFFD0 U3195 ( .I(n3313), .Z(n3314) );
  CKBD0 U3196 ( .CLK(n3314), .C(n3315) );
  CKBD0 U3197 ( .CLK(n3315), .C(n3316) );
  CKBD0 U3198 ( .CLK(n3316), .C(n3317) );
  CKBD0 U3199 ( .CLK(n3317), .C(n3318) );
  CKBD0 U3200 ( .CLK(n3318), .C(n3319) );
  CKBD0 U3201 ( .CLK(n3319), .C(n3320) );
  CKBD0 U3202 ( .CLK(n3320), .C(n3321) );
  CKBD0 U3203 ( .CLK(n3321), .C(n3322) );
  CKBD0 U3204 ( .CLK(n3322), .C(n3323) );
  CKBD0 U3205 ( .CLK(n3323), .C(n3324) );
  BUFFD0 U3206 ( .I(n3324), .Z(n3325) );
  CKBD0 U3207 ( .CLK(n3325), .C(n3326) );
  CKBD0 U3208 ( .CLK(n3326), .C(n3327) );
  CKBD0 U3209 ( .CLK(n3327), .C(n3328) );
  CKBD0 U3210 ( .CLK(n3328), .C(n3329) );
  CKBD0 U3211 ( .CLK(n3329), .C(n3330) );
  CKBD0 U3212 ( .CLK(n3330), .C(n3331) );
  BUFFD0 U3213 ( .I(n3331), .Z(n3332) );
  CKBD0 U3214 ( .CLK(n3332), .C(n3333) );
  BUFFD0 U3215 ( .I(n3333), .Z(n3334) );
  CKBD0 U3216 ( .CLK(n3334), .C(n3335) );
  BUFFD0 U3217 ( .I(n3335), .Z(n3336) );
  CKBD0 U3218 ( .CLK(n3336), .C(n3337) );
  BUFFD0 U3219 ( .I(n3337), .Z(n3338) );
  CKBD0 U3220 ( .CLK(n3338), .C(n3339) );
  BUFFD0 U3221 ( .I(n3339), .Z(n3340) );
  CKBD0 U3222 ( .CLK(n3340), .C(n3341) );
  BUFFD0 U3223 ( .I(n3341), .Z(n3342) );
  CKBD0 U3224 ( .CLK(n3342), .C(n3343) );
  BUFFD0 U3225 ( .I(n3343), .Z(n3344) );
  CKBD0 U3226 ( .CLK(n3344), .C(n3345) );
  BUFFD0 U3227 ( .I(n3345), .Z(n3346) );
  BUFFD0 U3228 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3229 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3230 ( .I(n158), .Z(n3349) );
  CKBD0 U3231 ( .CLK(n1344), .C(n3350) );
  CKBD0 U3232 ( .CLK(n3350), .C(n3351) );
  CKBD0 U3233 ( .CLK(n3351), .C(n3352) );
  BUFFD0 U3234 ( .I(n3352), .Z(n3353) );
  CKBD0 U3235 ( .CLK(n3353), .C(n3354) );
  CKBD0 U3236 ( .CLK(n3354), .C(n3355) );
  CKBD0 U3237 ( .CLK(n3355), .C(n3356) );
  CKBD0 U3238 ( .CLK(n3356), .C(n3357) );
  CKBD0 U3239 ( .CLK(n3357), .C(n3358) );
  CKBD0 U3240 ( .CLK(n3358), .C(n3359) );
  CKBD0 U3241 ( .CLK(n3359), .C(n3360) );
  CKBD0 U3242 ( .CLK(n3360), .C(n3361) );
  CKBD0 U3243 ( .CLK(n3361), .C(n3362) );
  CKBD0 U3244 ( .CLK(n3362), .C(n3363) );
  BUFFD0 U3245 ( .I(n3363), .Z(n3364) );
  CKBD0 U3246 ( .CLK(n3364), .C(n3365) );
  CKBD0 U3247 ( .CLK(n3365), .C(n3366) );
  CKBD0 U3248 ( .CLK(n3366), .C(n3367) );
  CKBD0 U3249 ( .CLK(n3367), .C(n3368) );
  CKBD0 U3250 ( .CLK(n3368), .C(n3369) );
  CKBD0 U3251 ( .CLK(n3369), .C(n3370) );
  CKBD0 U3252 ( .CLK(n3370), .C(n3371) );
  CKBD0 U3253 ( .CLK(n3371), .C(n3372) );
  CKBD0 U3254 ( .CLK(n3372), .C(n3373) );
  BUFFD0 U3255 ( .I(n3373), .Z(n3374) );
  CKBD0 U3256 ( .CLK(n3374), .C(n3375) );
  CKBD0 U3257 ( .CLK(n3375), .C(n3376) );
  CKBD0 U3258 ( .CLK(n3376), .C(n3377) );
  CKBD0 U3259 ( .CLK(n3377), .C(n3378) );
  CKBD0 U3260 ( .CLK(n3378), .C(n3379) );
  CKBD0 U3261 ( .CLK(n3379), .C(n3380) );
  CKBD0 U3262 ( .CLK(n3380), .C(n3381) );
  CKBD0 U3263 ( .CLK(n3381), .C(n3382) );
  CKBD0 U3264 ( .CLK(n3382), .C(n3383) );
  CKBD0 U3265 ( .CLK(n3383), .C(n3384) );
  BUFFD0 U3266 ( .I(n3384), .Z(n3385) );
  CKBD0 U3267 ( .CLK(n3385), .C(n3386) );
  CKBD0 U3268 ( .CLK(n3386), .C(n3387) );
  CKBD0 U3269 ( .CLK(n3387), .C(n3388) );
  CKBD0 U3270 ( .CLK(n3388), .C(n3389) );
  CKBD0 U3271 ( .CLK(n3389), .C(n3390) );
  CKBD0 U3272 ( .CLK(n3390), .C(n3391) );
  CKBD0 U3273 ( .CLK(n3391), .C(n3392) );
  CKBD0 U3274 ( .CLK(n3392), .C(n3393) );
  CKBD0 U3275 ( .CLK(n3393), .C(n3394) );
  CKBD0 U3276 ( .CLK(n3394), .C(n3395) );
  BUFFD0 U3277 ( .I(n3395), .Z(n3396) );
  CKBD0 U3278 ( .CLK(n3396), .C(n3397) );
  CKBD0 U3279 ( .CLK(n3397), .C(n3398) );
  CKBD0 U3280 ( .CLK(n3398), .C(n3399) );
  CKBD0 U3281 ( .CLK(n3399), .C(n3400) );
  CKBD0 U3282 ( .CLK(n3400), .C(n3401) );
  CKBD0 U3283 ( .CLK(n3401), .C(n3402) );
  CKBD0 U3284 ( .CLK(n3402), .C(n3403) );
  CKBD0 U3285 ( .CLK(n3403), .C(n3404) );
  CKBD0 U3286 ( .CLK(n3404), .C(n3405) );
  CKBD0 U3287 ( .CLK(n3405), .C(n3406) );
  BUFFD0 U3288 ( .I(n3406), .Z(n3407) );
  CKBD0 U3289 ( .CLK(n3407), .C(n3408) );
  CKBD0 U3290 ( .CLK(n3408), .C(n3409) );
  CKBD0 U3291 ( .CLK(n3409), .C(n3410) );
  CKBD0 U3292 ( .CLK(n3410), .C(n3411) );
  CKBD0 U3293 ( .CLK(n3411), .C(n3412) );
  CKBD0 U3294 ( .CLK(n3412), .C(n3413) );
  CKBD0 U3295 ( .CLK(n3413), .C(n3414) );
  CKBD0 U3296 ( .CLK(n3414), .C(n3415) );
  CKBD0 U3297 ( .CLK(n3415), .C(n3416) );
  CKBD0 U3298 ( .CLK(n3416), .C(n3417) );
  BUFFD0 U3299 ( .I(n3417), .Z(n3418) );
  CKBD0 U3300 ( .CLK(n3418), .C(n3419) );
  CKBD0 U3301 ( .CLK(n3419), .C(n3420) );
  CKBD0 U3302 ( .CLK(n3420), .C(n3421) );
  CKBD0 U3303 ( .CLK(n3421), .C(n3422) );
  CKBD0 U3304 ( .CLK(n3422), .C(n3423) );
  CKBD0 U3305 ( .CLK(n3423), .C(n3424) );
  CKBD0 U3306 ( .CLK(n3424), .C(n3425) );
  CKBD0 U3307 ( .CLK(n3425), .C(n3426) );
  CKBD0 U3308 ( .CLK(n3426), .C(n3427) );
  CKBD0 U3309 ( .CLK(n3427), .C(n3428) );
  BUFFD0 U3310 ( .I(n3428), .Z(n3429) );
  CKBD0 U3311 ( .CLK(n3429), .C(n3430) );
  CKBD0 U3312 ( .CLK(n3430), .C(n3431) );
  CKBD0 U3313 ( .CLK(n3431), .C(n3432) );
  CKBD0 U3314 ( .CLK(n3432), .C(n3433) );
  CKBD0 U3315 ( .CLK(n3433), .C(n3434) );
  CKBD0 U3316 ( .CLK(n3434), .C(n3435) );
  CKBD0 U3317 ( .CLK(n3435), .C(n3436) );
  CKBD0 U3318 ( .CLK(n3436), .C(n3437) );
  CKBD0 U3319 ( .CLK(n3437), .C(n3438) );
  BUFFD0 U3320 ( .I(n3438), .Z(n3439) );
  CKBD0 U3321 ( .CLK(n3439), .C(n3440) );
  CKBD0 U3322 ( .CLK(n3440), .C(n3441) );
  CKBD0 U3323 ( .CLK(n3441), .C(n3442) );
  CKBD0 U3324 ( .CLK(n3442), .C(n3443) );
  CKBD0 U3325 ( .CLK(n3443), .C(n3444) );
  CKBD0 U3326 ( .CLK(n3444), .C(n3445) );
  CKBD0 U3327 ( .CLK(n3445), .C(n3446) );
  CKBD0 U3328 ( .CLK(n3446), .C(n3447) );
  CKBD0 U3329 ( .CLK(n3447), .C(n3448) );
  CKBD0 U3330 ( .CLK(n3448), .C(n3449) );
  BUFFD0 U3331 ( .I(n3449), .Z(n3450) );
  CKBD0 U3332 ( .CLK(n3450), .C(n3451) );
  CKBD0 U3333 ( .CLK(n3451), .C(n3452) );
  CKBD0 U3334 ( .CLK(n3452), .C(n3453) );
  CKBD0 U3335 ( .CLK(n3453), .C(n3454) );
  CKBD0 U3336 ( .CLK(n3454), .C(n3455) );
  CKBD0 U3337 ( .CLK(n3455), .C(n3456) );
  CKBD0 U3338 ( .CLK(n3456), .C(n3457) );
  CKBD0 U3339 ( .CLK(n3457), .C(n3458) );
  CKBD0 U3340 ( .CLK(n3458), .C(n3459) );
  CKBD0 U3341 ( .CLK(n3459), .C(n3460) );
  BUFFD0 U3342 ( .I(n3460), .Z(n3461) );
  CKBD0 U3343 ( .CLK(n3461), .C(n3462) );
  CKBD0 U3344 ( .CLK(n3462), .C(n3463) );
  CKBD0 U3345 ( .CLK(n3463), .C(n3464) );
  CKBD0 U3346 ( .CLK(n3464), .C(n3465) );
  CKBD0 U3347 ( .CLK(n3465), .C(n3466) );
  CKBD0 U3348 ( .CLK(n3466), .C(n3467) );
  BUFFD0 U3349 ( .I(n3467), .Z(n3468) );
  CKBD0 U3350 ( .CLK(n3468), .C(n3469) );
  BUFFD0 U3351 ( .I(n3469), .Z(n3470) );
  CKBD0 U3352 ( .CLK(n3470), .C(n3471) );
  BUFFD0 U3353 ( .I(n3471), .Z(n3472) );
  CKBD0 U3354 ( .CLK(n3472), .C(n3473) );
  BUFFD0 U3355 ( .I(n3473), .Z(n3474) );
  CKBD0 U3356 ( .CLK(n3474), .C(n3475) );
  BUFFD0 U3357 ( .I(n3475), .Z(n3476) );
  CKBD0 U3358 ( .CLK(n3476), .C(n3477) );
  BUFFD0 U3359 ( .I(n3477), .Z(n3478) );
  CKBD0 U3360 ( .CLK(n3478), .C(n3479) );
  BUFFD0 U3361 ( .I(n3479), .Z(n3480) );
  CKBD0 U3362 ( .CLK(n3480), .C(n3481) );
  BUFFD0 U3363 ( .I(n3481), .Z(n3482) );
  BUFFD0 U3364 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3365 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3366 ( .I(n157), .Z(n3485) );
  CKBD0 U3367 ( .CLK(n1342), .C(n3486) );
  CKBD0 U3368 ( .CLK(n3486), .C(n3487) );
  CKBD0 U3369 ( .CLK(n3487), .C(n3488) );
  BUFFD0 U3370 ( .I(n3488), .Z(n3489) );
  CKBD0 U3371 ( .CLK(n3489), .C(n3490) );
  CKBD0 U3372 ( .CLK(n3490), .C(n3491) );
  CKBD0 U3373 ( .CLK(n3491), .C(n3492) );
  CKBD0 U3374 ( .CLK(n3492), .C(n3493) );
  CKBD0 U3375 ( .CLK(n3493), .C(n3494) );
  CKBD0 U3376 ( .CLK(n3494), .C(n3495) );
  CKBD0 U3377 ( .CLK(n3495), .C(n3496) );
  CKBD0 U3378 ( .CLK(n3496), .C(n3497) );
  CKBD0 U3379 ( .CLK(n3497), .C(n3498) );
  CKBD0 U3380 ( .CLK(n3498), .C(n3499) );
  BUFFD0 U3381 ( .I(n3499), .Z(n3500) );
  CKBD0 U3382 ( .CLK(n3500), .C(n3501) );
  CKBD0 U3383 ( .CLK(n3501), .C(n3502) );
  CKBD0 U3384 ( .CLK(n3502), .C(n3503) );
  CKBD0 U3385 ( .CLK(n3503), .C(n3504) );
  CKBD0 U3386 ( .CLK(n3504), .C(n3505) );
  CKBD0 U3387 ( .CLK(n3505), .C(n3506) );
  CKBD0 U3388 ( .CLK(n3506), .C(n3507) );
  CKBD0 U3389 ( .CLK(n3507), .C(n3508) );
  CKBD0 U3390 ( .CLK(n3508), .C(n3509) );
  BUFFD0 U3391 ( .I(n3509), .Z(n3510) );
  CKBD0 U3392 ( .CLK(n3510), .C(n3511) );
  CKBD0 U3393 ( .CLK(n3511), .C(n3512) );
  CKBD0 U3394 ( .CLK(n3512), .C(n3513) );
  CKBD0 U3395 ( .CLK(n3513), .C(n3514) );
  CKBD0 U3396 ( .CLK(n3514), .C(n3515) );
  CKBD0 U3397 ( .CLK(n3515), .C(n3516) );
  CKBD0 U3398 ( .CLK(n3516), .C(n3517) );
  CKBD0 U3399 ( .CLK(n3517), .C(n3518) );
  CKBD0 U3400 ( .CLK(n3518), .C(n3519) );
  CKBD0 U3401 ( .CLK(n3519), .C(n3520) );
  BUFFD0 U3402 ( .I(n3520), .Z(n3521) );
  CKBD0 U3403 ( .CLK(n3521), .C(n3522) );
  CKBD0 U3404 ( .CLK(n3522), .C(n3523) );
  CKBD0 U3405 ( .CLK(n3523), .C(n3524) );
  CKBD0 U3406 ( .CLK(n3524), .C(n3525) );
  CKBD0 U3407 ( .CLK(n3525), .C(n3526) );
  CKBD0 U3408 ( .CLK(n3526), .C(n3527) );
  CKBD0 U3409 ( .CLK(n3527), .C(n3528) );
  CKBD0 U3410 ( .CLK(n3528), .C(n3529) );
  CKBD0 U3411 ( .CLK(n3529), .C(n3530) );
  CKBD0 U3412 ( .CLK(n3530), .C(n3531) );
  BUFFD0 U3413 ( .I(n3531), .Z(n3532) );
  CKBD0 U3414 ( .CLK(n3532), .C(n3533) );
  CKBD0 U3415 ( .CLK(n3533), .C(n3534) );
  CKBD0 U3416 ( .CLK(n3534), .C(n3535) );
  CKBD0 U3417 ( .CLK(n3535), .C(n3536) );
  CKBD0 U3418 ( .CLK(n3536), .C(n3537) );
  CKBD0 U3419 ( .CLK(n3537), .C(n3538) );
  CKBD0 U3420 ( .CLK(n3538), .C(n3539) );
  CKBD0 U3421 ( .CLK(n3539), .C(n3540) );
  CKBD0 U3422 ( .CLK(n3540), .C(n3541) );
  CKBD0 U3423 ( .CLK(n3541), .C(n3542) );
  BUFFD0 U3424 ( .I(n3542), .Z(n3543) );
  CKBD0 U3425 ( .CLK(n3543), .C(n3544) );
  CKBD0 U3426 ( .CLK(n3544), .C(n3545) );
  CKBD0 U3427 ( .CLK(n3545), .C(n3546) );
  CKBD0 U3428 ( .CLK(n3546), .C(n3547) );
  CKBD0 U3429 ( .CLK(n3547), .C(n3548) );
  CKBD0 U3430 ( .CLK(n3548), .C(n3549) );
  CKBD0 U3431 ( .CLK(n3549), .C(n3550) );
  CKBD0 U3432 ( .CLK(n3550), .C(n3551) );
  CKBD0 U3433 ( .CLK(n3551), .C(n3552) );
  CKBD0 U3434 ( .CLK(n3552), .C(n3553) );
  BUFFD0 U3435 ( .I(n3553), .Z(n3554) );
  CKBD0 U3436 ( .CLK(n3554), .C(n3555) );
  CKBD0 U3437 ( .CLK(n3555), .C(n3556) );
  CKBD0 U3438 ( .CLK(n3556), .C(n3557) );
  CKBD0 U3439 ( .CLK(n3557), .C(n3558) );
  CKBD0 U3440 ( .CLK(n3558), .C(n3559) );
  CKBD0 U3441 ( .CLK(n3559), .C(n3560) );
  CKBD0 U3442 ( .CLK(n3560), .C(n3561) );
  CKBD0 U3443 ( .CLK(n3561), .C(n3562) );
  CKBD0 U3444 ( .CLK(n3562), .C(n3563) );
  CKBD0 U3445 ( .CLK(n3563), .C(n3564) );
  BUFFD0 U3446 ( .I(n3564), .Z(n3565) );
  CKBD0 U3447 ( .CLK(n3565), .C(n3566) );
  CKBD0 U3448 ( .CLK(n3566), .C(n3567) );
  CKBD0 U3449 ( .CLK(n3567), .C(n3568) );
  CKBD0 U3450 ( .CLK(n3568), .C(n3569) );
  CKBD0 U3451 ( .CLK(n3569), .C(n3570) );
  CKBD0 U3452 ( .CLK(n3570), .C(n3571) );
  CKBD0 U3453 ( .CLK(n3571), .C(n3572) );
  CKBD0 U3454 ( .CLK(n3572), .C(n3573) );
  CKBD0 U3455 ( .CLK(n3573), .C(n3574) );
  BUFFD0 U3456 ( .I(n3574), .Z(n3575) );
  CKBD0 U3457 ( .CLK(n3575), .C(n3576) );
  CKBD0 U3458 ( .CLK(n3576), .C(n3577) );
  CKBD0 U3459 ( .CLK(n3577), .C(n3578) );
  CKBD0 U3460 ( .CLK(n3578), .C(n3579) );
  CKBD0 U3461 ( .CLK(n3579), .C(n3580) );
  CKBD0 U3462 ( .CLK(n3580), .C(n3581) );
  CKBD0 U3463 ( .CLK(n3581), .C(n3582) );
  CKBD0 U3464 ( .CLK(n3582), .C(n3583) );
  CKBD0 U3465 ( .CLK(n3583), .C(n3584) );
  CKBD0 U3466 ( .CLK(n3584), .C(n3585) );
  BUFFD0 U3467 ( .I(n3585), .Z(n3586) );
  CKBD0 U3468 ( .CLK(n3586), .C(n3587) );
  CKBD0 U3469 ( .CLK(n3587), .C(n3588) );
  CKBD0 U3470 ( .CLK(n3588), .C(n3589) );
  CKBD0 U3471 ( .CLK(n3589), .C(n3590) );
  CKBD0 U3472 ( .CLK(n3590), .C(n3591) );
  CKBD0 U3473 ( .CLK(n3591), .C(n3592) );
  CKBD0 U3474 ( .CLK(n3592), .C(n3593) );
  CKBD0 U3475 ( .CLK(n3593), .C(n3594) );
  CKBD0 U3476 ( .CLK(n3594), .C(n3595) );
  CKBD0 U3477 ( .CLK(n3595), .C(n3596) );
  BUFFD0 U3478 ( .I(n3596), .Z(n3597) );
  CKBD0 U3479 ( .CLK(n3597), .C(n3598) );
  CKBD0 U3480 ( .CLK(n3598), .C(n3599) );
  CKBD0 U3481 ( .CLK(n3599), .C(n3600) );
  CKBD0 U3482 ( .CLK(n3600), .C(n3601) );
  CKBD0 U3483 ( .CLK(n3601), .C(n3602) );
  CKBD0 U3484 ( .CLK(n3602), .C(n3603) );
  BUFFD0 U3485 ( .I(n3603), .Z(n3604) );
  CKBD0 U3486 ( .CLK(n3604), .C(n3605) );
  BUFFD0 U3487 ( .I(n3605), .Z(n3606) );
  CKBD0 U3488 ( .CLK(n3606), .C(n3607) );
  BUFFD0 U3489 ( .I(n3607), .Z(n3608) );
  CKBD0 U3490 ( .CLK(n3608), .C(n3609) );
  BUFFD0 U3491 ( .I(n3609), .Z(n3610) );
  CKBD0 U3492 ( .CLK(n3610), .C(n3611) );
  BUFFD0 U3493 ( .I(n3611), .Z(n3612) );
  CKBD0 U3494 ( .CLK(n3612), .C(n3613) );
  BUFFD0 U3495 ( .I(n3613), .Z(n3614) );
  CKBD0 U3496 ( .CLK(n3614), .C(n3615) );
  BUFFD0 U3497 ( .I(n3615), .Z(n3616) );
  CKBD0 U3498 ( .CLK(n3616), .C(n3617) );
  BUFFD0 U3499 ( .I(n3617), .Z(n3618) );
  BUFFD0 U3500 ( .I(n3620), .Z(n3619) );
  BUFFD0 U3501 ( .I(n3621), .Z(n3620) );
  BUFFD0 U3502 ( .I(n156), .Z(n3621) );
  CKBD0 U3503 ( .CLK(n1844), .C(n3622) );
  CKBD0 U3504 ( .CLK(n3622), .C(n3623) );
  CKBD0 U3505 ( .CLK(n3623), .C(n3624) );
  BUFFD0 U3506 ( .I(n3624), .Z(n3625) );
  CKBD0 U3507 ( .CLK(n3625), .C(n3626) );
  CKBD0 U3508 ( .CLK(n3626), .C(n3627) );
  CKBD0 U3509 ( .CLK(n3627), .C(n3628) );
  CKBD0 U3510 ( .CLK(n3628), .C(n3629) );
  CKBD0 U3511 ( .CLK(n3629), .C(n3630) );
  CKBD0 U3512 ( .CLK(n3630), .C(n3631) );
  CKBD0 U3513 ( .CLK(n3631), .C(n3632) );
  CKBD0 U3514 ( .CLK(n3632), .C(n3633) );
  CKBD0 U3515 ( .CLK(n3633), .C(n3634) );
  CKBD0 U3516 ( .CLK(n3634), .C(n3635) );
  BUFFD0 U3517 ( .I(n3635), .Z(n3636) );
  CKBD0 U3518 ( .CLK(n3636), .C(n3637) );
  CKBD0 U3519 ( .CLK(n3637), .C(n3638) );
  CKBD0 U3520 ( .CLK(n3638), .C(n3639) );
  CKBD0 U3521 ( .CLK(n3639), .C(n3640) );
  CKBD0 U3522 ( .CLK(n3640), .C(n3641) );
  CKBD0 U3523 ( .CLK(n3641), .C(n3642) );
  CKBD0 U3524 ( .CLK(n3642), .C(n3643) );
  CKBD0 U3525 ( .CLK(n3643), .C(n3644) );
  CKBD0 U3526 ( .CLK(n3644), .C(n3645) );
  BUFFD0 U3527 ( .I(n3645), .Z(n3646) );
  CKBD0 U3528 ( .CLK(n3646), .C(n3647) );
  CKBD0 U3529 ( .CLK(n3647), .C(n3648) );
  CKBD0 U3530 ( .CLK(n3648), .C(n3649) );
  CKBD0 U3531 ( .CLK(n3649), .C(n3650) );
  CKBD0 U3532 ( .CLK(n3650), .C(n3651) );
  CKBD0 U3533 ( .CLK(n3651), .C(n3652) );
  CKBD0 U3534 ( .CLK(n3652), .C(n3653) );
  CKBD0 U3535 ( .CLK(n3653), .C(n3654) );
  CKBD0 U3536 ( .CLK(n3654), .C(n3655) );
  CKBD0 U3537 ( .CLK(n3655), .C(n3656) );
  BUFFD0 U3538 ( .I(n3656), .Z(n3657) );
  CKBD0 U3539 ( .CLK(n3657), .C(n3658) );
  CKBD0 U3540 ( .CLK(n3658), .C(n3659) );
  CKBD0 U3541 ( .CLK(n3659), .C(n3660) );
  CKBD0 U3542 ( .CLK(n3660), .C(n3661) );
  CKBD0 U3543 ( .CLK(n3661), .C(n3662) );
  CKBD0 U3544 ( .CLK(n3662), .C(n3663) );
  CKBD0 U3545 ( .CLK(n3663), .C(n3664) );
  CKBD0 U3546 ( .CLK(n3664), .C(n3665) );
  CKBD0 U3547 ( .CLK(n3665), .C(n3666) );
  CKBD0 U3548 ( .CLK(n3666), .C(n3667) );
  BUFFD0 U3549 ( .I(n3667), .Z(n3668) );
  CKBD0 U3550 ( .CLK(n3668), .C(n3669) );
  CKBD0 U3551 ( .CLK(n3669), .C(n3670) );
  CKBD0 U3552 ( .CLK(n3670), .C(n3671) );
  CKBD0 U3553 ( .CLK(n3671), .C(n3672) );
  CKBD0 U3554 ( .CLK(n3672), .C(n3673) );
  CKBD0 U3555 ( .CLK(n3673), .C(n3674) );
  CKBD0 U3556 ( .CLK(n3674), .C(n3675) );
  CKBD0 U3557 ( .CLK(n3675), .C(n3676) );
  CKBD0 U3558 ( .CLK(n3676), .C(n3677) );
  CKBD0 U3559 ( .CLK(n3677), .C(n3678) );
  BUFFD0 U3560 ( .I(n3678), .Z(n3679) );
  CKBD0 U3561 ( .CLK(n3679), .C(n3680) );
  CKBD0 U3562 ( .CLK(n3680), .C(n3681) );
  CKBD0 U3563 ( .CLK(n3681), .C(n3682) );
  CKBD0 U3564 ( .CLK(n3682), .C(n3683) );
  CKBD0 U3565 ( .CLK(n3683), .C(n3684) );
  CKBD0 U3566 ( .CLK(n3684), .C(n3685) );
  CKBD0 U3567 ( .CLK(n3685), .C(n3686) );
  CKBD0 U3568 ( .CLK(n3686), .C(n3687) );
  CKBD0 U3569 ( .CLK(n3687), .C(n3688) );
  CKBD0 U3570 ( .CLK(n3688), .C(n3689) );
  BUFFD0 U3571 ( .I(n3689), .Z(n3690) );
  CKBD0 U3572 ( .CLK(n3690), .C(n3691) );
  CKBD0 U3573 ( .CLK(n3691), .C(n3692) );
  CKBD0 U3574 ( .CLK(n3692), .C(n3693) );
  CKBD0 U3575 ( .CLK(n3693), .C(n3694) );
  CKBD0 U3576 ( .CLK(n3694), .C(n3695) );
  CKBD0 U3577 ( .CLK(n3695), .C(n3696) );
  CKBD0 U3578 ( .CLK(n3696), .C(n3697) );
  CKBD0 U3579 ( .CLK(n3697), .C(n3698) );
  CKBD0 U3580 ( .CLK(n3698), .C(n3699) );
  CKBD0 U3581 ( .CLK(n3699), .C(n3700) );
  BUFFD0 U3582 ( .I(n3700), .Z(n3701) );
  CKBD0 U3583 ( .CLK(n3701), .C(n3702) );
  CKBD0 U3584 ( .CLK(n3702), .C(n3703) );
  CKBD0 U3585 ( .CLK(n3703), .C(n3704) );
  CKBD0 U3586 ( .CLK(n3704), .C(n3705) );
  CKBD0 U3587 ( .CLK(n3705), .C(n3706) );
  CKBD0 U3588 ( .CLK(n3706), .C(n3707) );
  CKBD0 U3589 ( .CLK(n3707), .C(n3708) );
  CKBD0 U3590 ( .CLK(n3708), .C(n3709) );
  CKBD0 U3591 ( .CLK(n3709), .C(n3710) );
  BUFFD0 U3592 ( .I(n3710), .Z(n3711) );
  CKBD0 U3593 ( .CLK(n3711), .C(n3712) );
  CKBD0 U3594 ( .CLK(n3712), .C(n3713) );
  CKBD0 U3595 ( .CLK(n3713), .C(n3714) );
  CKBD0 U3596 ( .CLK(n3714), .C(n3715) );
  CKBD0 U3597 ( .CLK(n3715), .C(n3716) );
  CKBD0 U3598 ( .CLK(n3716), .C(n3717) );
  CKBD0 U3599 ( .CLK(n3717), .C(n3718) );
  CKBD0 U3600 ( .CLK(n3718), .C(n3719) );
  CKBD0 U3601 ( .CLK(n3719), .C(n3720) );
  CKBD0 U3602 ( .CLK(n3720), .C(n3721) );
  BUFFD0 U3603 ( .I(n3721), .Z(n3722) );
  CKBD0 U3604 ( .CLK(n3722), .C(n3723) );
  CKBD0 U3605 ( .CLK(n3723), .C(n3724) );
  CKBD0 U3606 ( .CLK(n3724), .C(n3725) );
  CKBD0 U3607 ( .CLK(n3725), .C(n3726) );
  CKBD0 U3608 ( .CLK(n3726), .C(n3727) );
  CKBD0 U3609 ( .CLK(n3727), .C(n3728) );
  CKBD0 U3610 ( .CLK(n3728), .C(n3729) );
  CKBD0 U3611 ( .CLK(n3729), .C(n3730) );
  CKBD0 U3612 ( .CLK(n3730), .C(n3731) );
  CKBD0 U3613 ( .CLK(n3731), .C(n3732) );
  BUFFD0 U3614 ( .I(n3732), .Z(n3733) );
  CKBD0 U3615 ( .CLK(n3733), .C(n3734) );
  CKBD0 U3616 ( .CLK(n3734), .C(n3735) );
  CKBD0 U3617 ( .CLK(n3735), .C(n3736) );
  CKBD0 U3618 ( .CLK(n3736), .C(n3737) );
  CKBD0 U3619 ( .CLK(n3737), .C(n3738) );
  CKBD0 U3620 ( .CLK(n3738), .C(n3739) );
  BUFFD0 U3621 ( .I(n3739), .Z(n3740) );
  CKBD0 U3622 ( .CLK(n3740), .C(n3741) );
  BUFFD0 U3623 ( .I(n3741), .Z(n3742) );
  CKBD0 U3624 ( .CLK(n3742), .C(n3743) );
  BUFFD0 U3625 ( .I(n3743), .Z(n3744) );
  CKBD0 U3626 ( .CLK(n3744), .C(n3745) );
  BUFFD0 U3627 ( .I(n3745), .Z(n3746) );
  CKBD0 U3628 ( .CLK(n3746), .C(n3747) );
  BUFFD0 U3629 ( .I(n3747), .Z(n3748) );
  CKBD0 U3630 ( .CLK(n3748), .C(n3749) );
  BUFFD0 U3631 ( .I(n3749), .Z(n3750) );
  CKBD0 U3632 ( .CLK(n3750), .C(n3751) );
  BUFFD0 U3633 ( .I(n3751), .Z(n3752) );
  CKBD0 U3634 ( .CLK(n3752), .C(n3753) );
  BUFFD0 U3635 ( .I(n3753), .Z(n3754) );
  BUFFD0 U3636 ( .I(n3756), .Z(n3755) );
  BUFFD0 U3637 ( .I(n3757), .Z(n3756) );
  BUFFD0 U3638 ( .I(n155), .Z(n3757) );
  CKBD0 U3639 ( .CLK(n1243), .C(n3758) );
  CKBD0 U3640 ( .CLK(n3758), .C(n3759) );
  CKBD0 U3641 ( .CLK(n3759), .C(n3760) );
  BUFFD0 U3642 ( .I(n3760), .Z(n3761) );
  CKBD0 U3643 ( .CLK(n3761), .C(n3762) );
  CKBD0 U3644 ( .CLK(n3762), .C(n3763) );
  CKBD0 U3645 ( .CLK(n3763), .C(n3764) );
  CKBD0 U3646 ( .CLK(n3764), .C(n3765) );
  CKBD0 U3647 ( .CLK(n3765), .C(n3766) );
  CKBD0 U3648 ( .CLK(n3766), .C(n3767) );
  CKBD0 U3649 ( .CLK(n3767), .C(n3768) );
  CKBD0 U3650 ( .CLK(n3768), .C(n3769) );
  CKBD0 U3651 ( .CLK(n3769), .C(n3770) );
  CKBD0 U3652 ( .CLK(n3770), .C(n3771) );
  BUFFD0 U3653 ( .I(n3771), .Z(n3772) );
  CKBD0 U3654 ( .CLK(n3772), .C(n3773) );
  CKBD0 U3655 ( .CLK(n3773), .C(n3774) );
  CKBD0 U3656 ( .CLK(n3774), .C(n3775) );
  CKBD0 U3657 ( .CLK(n3775), .C(n3776) );
  CKBD0 U3658 ( .CLK(n3776), .C(n3777) );
  CKBD0 U3659 ( .CLK(n3777), .C(n3778) );
  CKBD0 U3660 ( .CLK(n3778), .C(n3779) );
  CKBD0 U3661 ( .CLK(n3779), .C(n3780) );
  CKBD0 U3662 ( .CLK(n3780), .C(n3781) );
  BUFFD0 U3663 ( .I(n3781), .Z(n3782) );
  CKBD0 U3664 ( .CLK(n3782), .C(n3783) );
  CKBD0 U3665 ( .CLK(n3783), .C(n3784) );
  CKBD0 U3666 ( .CLK(n3784), .C(n3785) );
  CKBD0 U3667 ( .CLK(n3785), .C(n3786) );
  CKBD0 U3668 ( .CLK(n3786), .C(n3787) );
  CKBD0 U3669 ( .CLK(n3787), .C(n3788) );
  CKBD0 U3670 ( .CLK(n3788), .C(n3789) );
  CKBD0 U3671 ( .CLK(n3789), .C(n3790) );
  CKBD0 U3672 ( .CLK(n3790), .C(n3791) );
  CKBD0 U3673 ( .CLK(n3791), .C(n3792) );
  BUFFD0 U3674 ( .I(n3792), .Z(n3793) );
  CKBD0 U3675 ( .CLK(n3793), .C(n3794) );
  CKBD0 U3676 ( .CLK(n3794), .C(n3795) );
  CKBD0 U3677 ( .CLK(n3795), .C(n3796) );
  CKBD0 U3678 ( .CLK(n3796), .C(n3797) );
  CKBD0 U3679 ( .CLK(n3797), .C(n3798) );
  CKBD0 U3680 ( .CLK(n3798), .C(n3799) );
  CKBD0 U3681 ( .CLK(n3799), .C(n3800) );
  CKBD0 U3682 ( .CLK(n3800), .C(n3801) );
  CKBD0 U3683 ( .CLK(n3801), .C(n3802) );
  CKBD0 U3684 ( .CLK(n3802), .C(n3803) );
  BUFFD0 U3685 ( .I(n3803), .Z(n3804) );
  CKBD0 U3686 ( .CLK(n3804), .C(n3805) );
  CKBD0 U3687 ( .CLK(n3805), .C(n3806) );
  CKBD0 U3688 ( .CLK(n3806), .C(n3807) );
  CKBD0 U3689 ( .CLK(n3807), .C(n3808) );
  CKBD0 U3690 ( .CLK(n3808), .C(n3809) );
  CKBD0 U3691 ( .CLK(n3809), .C(n3810) );
  CKBD0 U3692 ( .CLK(n3810), .C(n3811) );
  CKBD0 U3693 ( .CLK(n3811), .C(n3812) );
  CKBD0 U3694 ( .CLK(n3812), .C(n3813) );
  CKBD0 U3695 ( .CLK(n3813), .C(n3814) );
  BUFFD0 U3696 ( .I(n3814), .Z(n3815) );
  CKBD0 U3697 ( .CLK(n3815), .C(n3816) );
  CKBD0 U3698 ( .CLK(n3816), .C(n3817) );
  CKBD0 U3699 ( .CLK(n3817), .C(n3818) );
  CKBD0 U3700 ( .CLK(n3818), .C(n3819) );
  CKBD0 U3701 ( .CLK(n3819), .C(n3820) );
  CKBD0 U3702 ( .CLK(n3820), .C(n3821) );
  CKBD0 U3703 ( .CLK(n3821), .C(n3822) );
  CKBD0 U3704 ( .CLK(n3822), .C(n3823) );
  CKBD0 U3705 ( .CLK(n3823), .C(n3824) );
  CKBD0 U3706 ( .CLK(n3824), .C(n3825) );
  BUFFD0 U3707 ( .I(n3825), .Z(n3826) );
  CKBD0 U3708 ( .CLK(n3826), .C(n3827) );
  CKBD0 U3709 ( .CLK(n3827), .C(n3828) );
  CKBD0 U3710 ( .CLK(n3828), .C(n3829) );
  CKBD0 U3711 ( .CLK(n3829), .C(n3830) );
  CKBD0 U3712 ( .CLK(n3830), .C(n3831) );
  CKBD0 U3713 ( .CLK(n3831), .C(n3832) );
  CKBD0 U3714 ( .CLK(n3832), .C(n3833) );
  CKBD0 U3715 ( .CLK(n3833), .C(n3834) );
  CKBD0 U3716 ( .CLK(n3834), .C(n3835) );
  CKBD0 U3717 ( .CLK(n3835), .C(n3836) );
  BUFFD0 U3718 ( .I(n3836), .Z(n3837) );
  CKBD0 U3719 ( .CLK(n3837), .C(n3838) );
  CKBD0 U3720 ( .CLK(n3838), .C(n3839) );
  CKBD0 U3721 ( .CLK(n3839), .C(n3840) );
  CKBD0 U3722 ( .CLK(n3840), .C(n3841) );
  CKBD0 U3723 ( .CLK(n3841), .C(n3842) );
  CKBD0 U3724 ( .CLK(n3842), .C(n3843) );
  CKBD0 U3725 ( .CLK(n3843), .C(n3844) );
  CKBD0 U3726 ( .CLK(n3844), .C(n3845) );
  CKBD0 U3727 ( .CLK(n3845), .C(n3846) );
  BUFFD0 U3728 ( .I(n3846), .Z(n3847) );
  CKBD0 U3729 ( .CLK(n3847), .C(n3848) );
  CKBD0 U3730 ( .CLK(n3848), .C(n3849) );
  CKBD0 U3731 ( .CLK(n3849), .C(n3850) );
  CKBD0 U3732 ( .CLK(n3850), .C(n3851) );
  CKBD0 U3733 ( .CLK(n3851), .C(n3852) );
  CKBD0 U3734 ( .CLK(n3852), .C(n3853) );
  CKBD0 U3735 ( .CLK(n3853), .C(n3854) );
  CKBD0 U3736 ( .CLK(n3854), .C(n3855) );
  CKBD0 U3737 ( .CLK(n3855), .C(n3856) );
  CKBD0 U3738 ( .CLK(n3856), .C(n3857) );
  BUFFD0 U3739 ( .I(n3857), .Z(n3858) );
  CKBD0 U3740 ( .CLK(n3858), .C(n3859) );
  CKBD0 U3741 ( .CLK(n3859), .C(n3860) );
  CKBD0 U3742 ( .CLK(n3860), .C(n3861) );
  CKBD0 U3743 ( .CLK(n3861), .C(n3862) );
  CKBD0 U3744 ( .CLK(n3862), .C(n3863) );
  CKBD0 U3745 ( .CLK(n3863), .C(n3864) );
  CKBD0 U3746 ( .CLK(n3864), .C(n3865) );
  CKBD0 U3747 ( .CLK(n3865), .C(n3866) );
  CKBD0 U3748 ( .CLK(n3866), .C(n3867) );
  CKBD0 U3749 ( .CLK(n3867), .C(n3868) );
  BUFFD0 U3750 ( .I(n3868), .Z(n3869) );
  CKBD0 U3751 ( .CLK(n3869), .C(n3870) );
  CKBD0 U3752 ( .CLK(n3870), .C(n3871) );
  CKBD0 U3753 ( .CLK(n3871), .C(n3872) );
  CKBD0 U3754 ( .CLK(n3872), .C(n3873) );
  CKBD0 U3755 ( .CLK(n3873), .C(n3874) );
  CKBD0 U3756 ( .CLK(n3874), .C(n3875) );
  BUFFD0 U3757 ( .I(n3875), .Z(n3876) );
  CKBD0 U3758 ( .CLK(n3876), .C(n3877) );
  BUFFD0 U3759 ( .I(n3877), .Z(n3878) );
  CKBD0 U3760 ( .CLK(n3878), .C(n3879) );
  BUFFD0 U3761 ( .I(n3879), .Z(n3880) );
  CKBD0 U3762 ( .CLK(n3880), .C(n3881) );
  BUFFD0 U3763 ( .I(n3881), .Z(n3882) );
  CKBD0 U3764 ( .CLK(n3882), .C(n3883) );
  BUFFD0 U3765 ( .I(n3883), .Z(n3884) );
  CKBD0 U3766 ( .CLK(n3884), .C(n3885) );
  BUFFD0 U3767 ( .I(n3885), .Z(n3886) );
  CKBD0 U3768 ( .CLK(n3886), .C(n3887) );
  BUFFD0 U3769 ( .I(n3887), .Z(n3888) );
  CKBD0 U3770 ( .CLK(n3888), .C(n3889) );
  BUFFD0 U3771 ( .I(n3889), .Z(n3890) );
  BUFFD0 U3772 ( .I(n3892), .Z(n3891) );
  BUFFD0 U3773 ( .I(n3893), .Z(n3892) );
  BUFFD0 U3774 ( .I(n154), .Z(n3893) );
  CKBD0 U3775 ( .CLK(n1241), .C(n3894) );
  CKBD0 U3776 ( .CLK(n3894), .C(n3895) );
  CKBD0 U3777 ( .CLK(n3895), .C(n3896) );
  BUFFD0 U3778 ( .I(n3896), .Z(n3897) );
  CKBD0 U3779 ( .CLK(n3897), .C(n3898) );
  CKBD0 U3780 ( .CLK(n3898), .C(n3899) );
  CKBD0 U3781 ( .CLK(n3899), .C(n3900) );
  CKBD0 U3782 ( .CLK(n3900), .C(n3901) );
  CKBD0 U3783 ( .CLK(n3901), .C(n3902) );
  CKBD0 U3784 ( .CLK(n3902), .C(n3903) );
  CKBD0 U3785 ( .CLK(n3903), .C(n3904) );
  CKBD0 U3786 ( .CLK(n3904), .C(n3905) );
  CKBD0 U3787 ( .CLK(n3905), .C(n3906) );
  CKBD0 U3788 ( .CLK(n3906), .C(n3907) );
  BUFFD0 U3789 ( .I(n3907), .Z(n3908) );
  CKBD0 U3790 ( .CLK(n3908), .C(n3909) );
  CKBD0 U3791 ( .CLK(n3909), .C(n3910) );
  CKBD0 U3792 ( .CLK(n3910), .C(n3911) );
  CKBD0 U3793 ( .CLK(n3911), .C(n3912) );
  CKBD0 U3794 ( .CLK(n3912), .C(n3913) );
  CKBD0 U3795 ( .CLK(n3913), .C(n3914) );
  CKBD0 U3796 ( .CLK(n3914), .C(n3915) );
  CKBD0 U3797 ( .CLK(n3915), .C(n3916) );
  CKBD0 U3798 ( .CLK(n3916), .C(n3917) );
  BUFFD0 U3799 ( .I(n3917), .Z(n3918) );
  CKBD0 U3800 ( .CLK(n3918), .C(n3919) );
  CKBD0 U3801 ( .CLK(n3919), .C(n3920) );
  CKBD0 U3802 ( .CLK(n3920), .C(n3921) );
  CKBD0 U3803 ( .CLK(n3921), .C(n3922) );
  CKBD0 U3804 ( .CLK(n3922), .C(n3923) );
  CKBD0 U3805 ( .CLK(n3923), .C(n3924) );
  CKBD0 U3806 ( .CLK(n3924), .C(n3925) );
  CKBD0 U3807 ( .CLK(n3925), .C(n3926) );
  CKBD0 U3808 ( .CLK(n3926), .C(n3927) );
  CKBD0 U3809 ( .CLK(n3927), .C(n3928) );
  BUFFD0 U3810 ( .I(n3928), .Z(n3929) );
  CKBD0 U3811 ( .CLK(n3929), .C(n3930) );
  CKBD0 U3812 ( .CLK(n3930), .C(n3931) );
  CKBD0 U3813 ( .CLK(n3931), .C(n3932) );
  CKBD0 U3814 ( .CLK(n3932), .C(n3933) );
  CKBD0 U3815 ( .CLK(n3933), .C(n3934) );
  CKBD0 U3816 ( .CLK(n3934), .C(n3935) );
  CKBD0 U3817 ( .CLK(n3935), .C(n3936) );
  CKBD0 U3818 ( .CLK(n3936), .C(n3937) );
  CKBD0 U3819 ( .CLK(n3937), .C(n3938) );
  CKBD0 U3820 ( .CLK(n3938), .C(n3939) );
  BUFFD0 U3821 ( .I(n3939), .Z(n3940) );
  CKBD0 U3822 ( .CLK(n3940), .C(n3941) );
  CKBD0 U3823 ( .CLK(n3941), .C(n3942) );
  CKBD0 U3824 ( .CLK(n3942), .C(n3943) );
  CKBD0 U3825 ( .CLK(n3943), .C(n3944) );
  CKBD0 U3826 ( .CLK(n3944), .C(n3945) );
  CKBD0 U3827 ( .CLK(n3945), .C(n3946) );
  CKBD0 U3828 ( .CLK(n3946), .C(n3947) );
  CKBD0 U3829 ( .CLK(n3947), .C(n3948) );
  CKBD0 U3830 ( .CLK(n3948), .C(n3949) );
  CKBD0 U3831 ( .CLK(n3949), .C(n3950) );
  BUFFD0 U3832 ( .I(n3950), .Z(n3951) );
  CKBD0 U3833 ( .CLK(n3951), .C(n3952) );
  CKBD0 U3834 ( .CLK(n3952), .C(n3953) );
  CKBD0 U3835 ( .CLK(n3953), .C(n3954) );
  CKBD0 U3836 ( .CLK(n3954), .C(n3955) );
  CKBD0 U3837 ( .CLK(n3955), .C(n3956) );
  CKBD0 U3838 ( .CLK(n3956), .C(n3957) );
  CKBD0 U3839 ( .CLK(n3957), .C(n3958) );
  CKBD0 U3840 ( .CLK(n3958), .C(n3959) );
  CKBD0 U3841 ( .CLK(n3959), .C(n3960) );
  CKBD0 U3842 ( .CLK(n3960), .C(n3961) );
  BUFFD0 U3843 ( .I(n3961), .Z(n3962) );
  CKBD0 U3844 ( .CLK(n3962), .C(n3963) );
  CKBD0 U3845 ( .CLK(n3963), .C(n3964) );
  CKBD0 U3846 ( .CLK(n3964), .C(n3965) );
  CKBD0 U3847 ( .CLK(n3965), .C(n3966) );
  CKBD0 U3848 ( .CLK(n3966), .C(n3967) );
  CKBD0 U3849 ( .CLK(n3967), .C(n3968) );
  CKBD0 U3850 ( .CLK(n3968), .C(n3969) );
  CKBD0 U3851 ( .CLK(n3969), .C(n3970) );
  CKBD0 U3852 ( .CLK(n3970), .C(n3971) );
  CKBD0 U3853 ( .CLK(n3971), .C(n3972) );
  BUFFD0 U3854 ( .I(n3972), .Z(n3973) );
  CKBD0 U3855 ( .CLK(n3973), .C(n3974) );
  CKBD0 U3856 ( .CLK(n3974), .C(n3975) );
  CKBD0 U3857 ( .CLK(n3975), .C(n3976) );
  CKBD0 U3858 ( .CLK(n3976), .C(n3977) );
  CKBD0 U3859 ( .CLK(n3977), .C(n3978) );
  CKBD0 U3860 ( .CLK(n3978), .C(n3979) );
  CKBD0 U3861 ( .CLK(n3979), .C(n3980) );
  CKBD0 U3862 ( .CLK(n3980), .C(n3981) );
  CKBD0 U3863 ( .CLK(n3981), .C(n3982) );
  BUFFD0 U3864 ( .I(n3982), .Z(n3983) );
  CKBD0 U3865 ( .CLK(n3983), .C(n3984) );
  CKBD0 U3866 ( .CLK(n3984), .C(n3985) );
  CKBD0 U3867 ( .CLK(n3985), .C(n3986) );
  CKBD0 U3868 ( .CLK(n3986), .C(n3987) );
  CKBD0 U3869 ( .CLK(n3987), .C(n3988) );
  CKBD0 U3870 ( .CLK(n3988), .C(n3989) );
  CKBD0 U3871 ( .CLK(n3989), .C(n3990) );
  CKBD0 U3872 ( .CLK(n3990), .C(n3991) );
  CKBD0 U3873 ( .CLK(n3991), .C(n3992) );
  CKBD0 U3874 ( .CLK(n3992), .C(n3993) );
  BUFFD0 U3875 ( .I(n3993), .Z(n3994) );
  CKBD0 U3876 ( .CLK(n3994), .C(n3995) );
  CKBD0 U3877 ( .CLK(n3995), .C(n3996) );
  CKBD0 U3878 ( .CLK(n3996), .C(n3997) );
  CKBD0 U3879 ( .CLK(n3997), .C(n3998) );
  CKBD0 U3880 ( .CLK(n3998), .C(n3999) );
  CKBD0 U3881 ( .CLK(n3999), .C(n4000) );
  CKBD0 U3882 ( .CLK(n4000), .C(n4001) );
  CKBD0 U3883 ( .CLK(n4001), .C(n4002) );
  CKBD0 U3884 ( .CLK(n4002), .C(n4003) );
  CKBD0 U3885 ( .CLK(n4003), .C(n4004) );
  BUFFD0 U3886 ( .I(n4004), .Z(n4005) );
  CKBD0 U3887 ( .CLK(n4005), .C(n4006) );
  CKBD0 U3888 ( .CLK(n4006), .C(n4007) );
  CKBD0 U3889 ( .CLK(n4007), .C(n4008) );
  CKBD0 U3890 ( .CLK(n4008), .C(n4009) );
  CKBD0 U3891 ( .CLK(n4009), .C(n4010) );
  CKBD0 U3892 ( .CLK(n4010), .C(n4011) );
  BUFFD0 U3893 ( .I(n4011), .Z(n4012) );
  CKBD0 U3894 ( .CLK(n4012), .C(n4013) );
  BUFFD0 U3895 ( .I(n4013), .Z(n4014) );
  CKBD0 U3896 ( .CLK(n4014), .C(n4015) );
  BUFFD0 U3897 ( .I(n4015), .Z(n4016) );
  CKBD0 U3898 ( .CLK(n4016), .C(n4017) );
  BUFFD0 U3899 ( .I(n4017), .Z(n4018) );
  CKBD0 U3900 ( .CLK(n4018), .C(n4019) );
  BUFFD0 U3901 ( .I(n4019), .Z(n4020) );
  CKBD0 U3902 ( .CLK(n4020), .C(n4021) );
  BUFFD0 U3903 ( .I(n4021), .Z(n4022) );
  CKBD0 U3904 ( .CLK(n4022), .C(n4023) );
  BUFFD0 U3905 ( .I(n4023), .Z(n4024) );
  CKBD0 U3906 ( .CLK(n4024), .C(n4025) );
  BUFFD0 U3907 ( .I(n4025), .Z(n4026) );
  BUFFD0 U3908 ( .I(n4028), .Z(n4027) );
  BUFFD0 U3909 ( .I(n4029), .Z(n4028) );
  BUFFD0 U3910 ( .I(n153), .Z(n4029) );
  CKBD0 U3911 ( .CLK(n1239), .C(n4030) );
  CKBD0 U3912 ( .CLK(n4030), .C(n4031) );
  CKBD0 U3913 ( .CLK(n4031), .C(n4032) );
  BUFFD0 U3914 ( .I(n4032), .Z(n4033) );
  CKBD0 U3915 ( .CLK(n4033), .C(n4034) );
  CKBD0 U3916 ( .CLK(n4034), .C(n4035) );
  CKBD0 U3917 ( .CLK(n4035), .C(n4036) );
  CKBD0 U3918 ( .CLK(n4036), .C(n4037) );
  CKBD0 U3919 ( .CLK(n4037), .C(n4038) );
  CKBD0 U3920 ( .CLK(n4038), .C(n4039) );
  CKBD0 U3921 ( .CLK(n4039), .C(n4040) );
  CKBD0 U3922 ( .CLK(n4040), .C(n4041) );
  CKBD0 U3923 ( .CLK(n4041), .C(n4042) );
  CKBD0 U3924 ( .CLK(n4042), .C(n4043) );
  BUFFD0 U3925 ( .I(n4043), .Z(n4044) );
  CKBD0 U3926 ( .CLK(n4044), .C(n4045) );
  CKBD0 U3927 ( .CLK(n4045), .C(n4046) );
  CKBD0 U3928 ( .CLK(n4046), .C(n4047) );
  CKBD0 U3929 ( .CLK(n4047), .C(n4048) );
  CKBD0 U3930 ( .CLK(n4048), .C(n4049) );
  CKBD0 U3931 ( .CLK(n4049), .C(n4050) );
  CKBD0 U3932 ( .CLK(n4050), .C(n4051) );
  CKBD0 U3933 ( .CLK(n4051), .C(n4052) );
  CKBD0 U3934 ( .CLK(n4052), .C(n4053) );
  BUFFD0 U3935 ( .I(n4053), .Z(n4054) );
  CKBD0 U3936 ( .CLK(n4054), .C(n4055) );
  CKBD0 U3937 ( .CLK(n4055), .C(n4056) );
  CKBD0 U3938 ( .CLK(n4056), .C(n4057) );
  CKBD0 U3939 ( .CLK(n4057), .C(n4058) );
  CKBD0 U3940 ( .CLK(n4058), .C(n4059) );
  CKBD0 U3941 ( .CLK(n4059), .C(n4060) );
  CKBD0 U3942 ( .CLK(n4060), .C(n4061) );
  CKBD0 U3943 ( .CLK(n4061), .C(n4062) );
  CKBD0 U3944 ( .CLK(n4062), .C(n4063) );
  CKBD0 U3945 ( .CLK(n4063), .C(n4064) );
  BUFFD0 U3946 ( .I(n4064), .Z(n4065) );
  CKBD0 U3947 ( .CLK(n4065), .C(n4066) );
  CKBD0 U3948 ( .CLK(n4066), .C(n4067) );
  CKBD0 U3949 ( .CLK(n4067), .C(n4068) );
  CKBD0 U3950 ( .CLK(n4068), .C(n4069) );
  CKBD0 U3951 ( .CLK(n4069), .C(n4070) );
  CKBD0 U3952 ( .CLK(n4070), .C(n4071) );
  CKBD0 U3953 ( .CLK(n4071), .C(n4072) );
  CKBD0 U3954 ( .CLK(n4072), .C(n4073) );
  CKBD0 U3955 ( .CLK(n4073), .C(n4074) );
  CKBD0 U3956 ( .CLK(n4074), .C(n4075) );
  BUFFD0 U3957 ( .I(n4075), .Z(n4076) );
  CKBD0 U3958 ( .CLK(n4076), .C(n4077) );
  CKBD0 U3959 ( .CLK(n4077), .C(n4078) );
  CKBD0 U3960 ( .CLK(n4078), .C(n4079) );
  CKBD0 U3961 ( .CLK(n4079), .C(n4080) );
  CKBD0 U3962 ( .CLK(n4080), .C(n4081) );
  CKBD0 U3963 ( .CLK(n4081), .C(n4082) );
  CKBD0 U3964 ( .CLK(n4082), .C(n4083) );
  CKBD0 U3965 ( .CLK(n4083), .C(n4084) );
  CKBD0 U3966 ( .CLK(n4084), .C(n4085) );
  CKBD0 U3967 ( .CLK(n4085), .C(n4086) );
  BUFFD0 U3968 ( .I(n4086), .Z(n4087) );
  CKBD0 U3969 ( .CLK(n4087), .C(n4088) );
  CKBD0 U3970 ( .CLK(n4088), .C(n4089) );
  CKBD0 U3971 ( .CLK(n4089), .C(n4090) );
  CKBD0 U3972 ( .CLK(n4090), .C(n4091) );
  CKBD0 U3973 ( .CLK(n4091), .C(n4092) );
  CKBD0 U3974 ( .CLK(n4092), .C(n4093) );
  CKBD0 U3975 ( .CLK(n4093), .C(n4094) );
  CKBD0 U3976 ( .CLK(n4094), .C(n4095) );
  CKBD0 U3977 ( .CLK(n4095), .C(n4096) );
  CKBD0 U3978 ( .CLK(n4096), .C(n4097) );
  BUFFD0 U3979 ( .I(n4097), .Z(n4098) );
  CKBD0 U3980 ( .CLK(n4098), .C(n4099) );
  CKBD0 U3981 ( .CLK(n4099), .C(n4100) );
  CKBD0 U3982 ( .CLK(n4100), .C(n4101) );
  CKBD0 U3983 ( .CLK(n4101), .C(n4102) );
  CKBD0 U3984 ( .CLK(n4102), .C(n4103) );
  CKBD0 U3985 ( .CLK(n4103), .C(n4104) );
  CKBD0 U3986 ( .CLK(n4104), .C(n4105) );
  CKBD0 U3987 ( .CLK(n4105), .C(n4106) );
  CKBD0 U3988 ( .CLK(n4106), .C(n4107) );
  CKBD0 U3989 ( .CLK(n4107), .C(n4108) );
  BUFFD0 U3990 ( .I(n4108), .Z(n4109) );
  CKBD0 U3991 ( .CLK(n4109), .C(n4110) );
  CKBD0 U3992 ( .CLK(n4110), .C(n4111) );
  CKBD0 U3993 ( .CLK(n4111), .C(n4112) );
  CKBD0 U3994 ( .CLK(n4112), .C(n4113) );
  CKBD0 U3995 ( .CLK(n4113), .C(n4114) );
  CKBD0 U3996 ( .CLK(n4114), .C(n4115) );
  CKBD0 U3997 ( .CLK(n4115), .C(n4116) );
  CKBD0 U3998 ( .CLK(n4116), .C(n4117) );
  CKBD0 U3999 ( .CLK(n4117), .C(n4118) );
  BUFFD0 U4000 ( .I(n4118), .Z(n4119) );
  CKBD0 U4001 ( .CLK(n4119), .C(n4120) );
  CKBD0 U4002 ( .CLK(n4120), .C(n4121) );
  CKBD0 U4003 ( .CLK(n4121), .C(n4122) );
  CKBD0 U4004 ( .CLK(n4122), .C(n4123) );
  CKBD0 U4005 ( .CLK(n4123), .C(n4124) );
  CKBD0 U4006 ( .CLK(n4124), .C(n4125) );
  CKBD0 U4007 ( .CLK(n4125), .C(n4126) );
  CKBD0 U4008 ( .CLK(n4126), .C(n4127) );
  CKBD0 U4009 ( .CLK(n4127), .C(n4128) );
  CKBD0 U4010 ( .CLK(n4128), .C(n4129) );
  BUFFD0 U4011 ( .I(n4129), .Z(n4130) );
  CKBD0 U4012 ( .CLK(n4130), .C(n4131) );
  CKBD0 U4013 ( .CLK(n4131), .C(n4132) );
  CKBD0 U4014 ( .CLK(n4132), .C(n4133) );
  CKBD0 U4015 ( .CLK(n4133), .C(n4134) );
  CKBD0 U4016 ( .CLK(n4134), .C(n4135) );
  CKBD0 U4017 ( .CLK(n4135), .C(n4136) );
  CKBD0 U4018 ( .CLK(n4136), .C(n4137) );
  CKBD0 U4019 ( .CLK(n4137), .C(n4138) );
  CKBD0 U4020 ( .CLK(n4138), .C(n4139) );
  CKBD0 U4021 ( .CLK(n4139), .C(n4140) );
  BUFFD0 U4022 ( .I(n4140), .Z(n4141) );
  CKBD0 U4023 ( .CLK(n4141), .C(n4142) );
  CKBD0 U4024 ( .CLK(n4142), .C(n4143) );
  CKBD0 U4025 ( .CLK(n4143), .C(n4144) );
  CKBD0 U4026 ( .CLK(n4144), .C(n4145) );
  CKBD0 U4027 ( .CLK(n4145), .C(n4146) );
  CKBD0 U4028 ( .CLK(n4146), .C(n4147) );
  BUFFD0 U4029 ( .I(n4147), .Z(n4148) );
  CKBD0 U4030 ( .CLK(n4148), .C(n4149) );
  BUFFD0 U4031 ( .I(n4149), .Z(n4150) );
  CKBD0 U4032 ( .CLK(n4150), .C(n4151) );
  BUFFD0 U4033 ( .I(n4151), .Z(n4152) );
  CKBD0 U4034 ( .CLK(n4152), .C(n4153) );
  BUFFD0 U4035 ( .I(n4153), .Z(n4154) );
  CKBD0 U4036 ( .CLK(n4154), .C(n4155) );
  BUFFD0 U4037 ( .I(n4155), .Z(n4156) );
  CKBD0 U4038 ( .CLK(n4156), .C(n4157) );
  BUFFD0 U4039 ( .I(n4157), .Z(n4158) );
  CKBD0 U4040 ( .CLK(n4158), .C(n4159) );
  BUFFD0 U4041 ( .I(n4159), .Z(n4160) );
  CKBD0 U4042 ( .CLK(n4160), .C(n4161) );
  BUFFD0 U4043 ( .I(n4161), .Z(n4162) );
  BUFFD0 U4044 ( .I(n4164), .Z(n4163) );
  BUFFD0 U4045 ( .I(n4165), .Z(n4164) );
  BUFFD0 U4046 ( .I(n152), .Z(n4165) );
  CKBD0 U4047 ( .CLK(n1237), .C(n4166) );
  CKBD0 U4048 ( .CLK(n4166), .C(n4167) );
  CKBD0 U4049 ( .CLK(n4167), .C(n4168) );
  BUFFD0 U4050 ( .I(n4168), .Z(n4169) );
  CKBD0 U4051 ( .CLK(n4169), .C(n4170) );
  CKBD0 U4052 ( .CLK(n4170), .C(n4171) );
  CKBD0 U4053 ( .CLK(n4171), .C(n4172) );
  CKBD0 U4054 ( .CLK(n4172), .C(n4173) );
  CKBD0 U4055 ( .CLK(n4173), .C(n4174) );
  CKBD0 U4056 ( .CLK(n4174), .C(n4175) );
  CKBD0 U4057 ( .CLK(n4175), .C(n4176) );
  CKBD0 U4058 ( .CLK(n4176), .C(n4177) );
  CKBD0 U4059 ( .CLK(n4177), .C(n4178) );
  CKBD0 U4060 ( .CLK(n4178), .C(n4179) );
  BUFFD0 U4061 ( .I(n4179), .Z(n4180) );
  CKBD0 U4062 ( .CLK(n4180), .C(n4181) );
  CKBD0 U4063 ( .CLK(n4181), .C(n4182) );
  CKBD0 U4064 ( .CLK(n4182), .C(n4183) );
  CKBD0 U4065 ( .CLK(n4183), .C(n4184) );
  CKBD0 U4066 ( .CLK(n4184), .C(n4185) );
  CKBD0 U4067 ( .CLK(n4185), .C(n4186) );
  CKBD0 U4068 ( .CLK(n4186), .C(n4187) );
  CKBD0 U4069 ( .CLK(n4187), .C(n4188) );
  CKBD0 U4070 ( .CLK(n4188), .C(n4189) );
  BUFFD0 U4071 ( .I(n4189), .Z(n4190) );
  CKBD0 U4072 ( .CLK(n4190), .C(n4191) );
  CKBD0 U4073 ( .CLK(n4191), .C(n4192) );
  CKBD0 U4074 ( .CLK(n4192), .C(n4193) );
  CKBD0 U4075 ( .CLK(n4193), .C(n4194) );
  CKBD0 U4076 ( .CLK(n4194), .C(n4195) );
  CKBD0 U4077 ( .CLK(n4195), .C(n4196) );
  CKBD0 U4078 ( .CLK(n4196), .C(n4197) );
  CKBD0 U4079 ( .CLK(n4197), .C(n4198) );
  CKBD0 U4080 ( .CLK(n4198), .C(n4199) );
  CKBD0 U4081 ( .CLK(n4199), .C(n4200) );
  BUFFD0 U4082 ( .I(n4200), .Z(n4201) );
  CKBD0 U4083 ( .CLK(n4201), .C(n4202) );
  CKBD0 U4084 ( .CLK(n4202), .C(n4203) );
  CKBD0 U4085 ( .CLK(n4203), .C(n4204) );
  CKBD0 U4086 ( .CLK(n4204), .C(n4205) );
  CKBD0 U4087 ( .CLK(n4205), .C(n4206) );
  CKBD0 U4088 ( .CLK(n4206), .C(n4207) );
  CKBD0 U4089 ( .CLK(n4207), .C(n4208) );
  CKBD0 U4090 ( .CLK(n4208), .C(n4209) );
  CKBD0 U4091 ( .CLK(n4209), .C(n4210) );
  CKBD0 U4092 ( .CLK(n4210), .C(n4211) );
  BUFFD0 U4093 ( .I(n4211), .Z(n4212) );
  CKBD0 U4094 ( .CLK(n4212), .C(n4213) );
  CKBD0 U4095 ( .CLK(n4213), .C(n4214) );
  CKBD0 U4096 ( .CLK(n4214), .C(n4215) );
  CKBD0 U4097 ( .CLK(n4215), .C(n4216) );
  CKBD0 U4098 ( .CLK(n4216), .C(n4217) );
  CKBD0 U4099 ( .CLK(n4217), .C(n4218) );
  CKBD0 U4100 ( .CLK(n4218), .C(n4219) );
  CKBD0 U4101 ( .CLK(n4219), .C(n4220) );
  CKBD0 U4102 ( .CLK(n4220), .C(n4221) );
  CKBD0 U4103 ( .CLK(n4221), .C(n4222) );
  BUFFD0 U4104 ( .I(n4222), .Z(n4223) );
  CKBD0 U4105 ( .CLK(n4223), .C(n4224) );
  CKBD0 U4106 ( .CLK(n4224), .C(n4225) );
  CKBD0 U4107 ( .CLK(n4225), .C(n4226) );
  CKBD0 U4108 ( .CLK(n4226), .C(n4227) );
  CKBD0 U4109 ( .CLK(n4227), .C(n4228) );
  CKBD0 U4110 ( .CLK(n4228), .C(n4229) );
  CKBD0 U4111 ( .CLK(n4229), .C(n4230) );
  CKBD0 U4112 ( .CLK(n4230), .C(n4231) );
  CKBD0 U4113 ( .CLK(n4231), .C(n4232) );
  CKBD0 U4114 ( .CLK(n4232), .C(n4233) );
  BUFFD0 U4115 ( .I(n4233), .Z(n4234) );
  CKBD0 U4116 ( .CLK(n4234), .C(n4235) );
  CKBD0 U4117 ( .CLK(n4235), .C(n4236) );
  CKBD0 U4118 ( .CLK(n4236), .C(n4237) );
  CKBD0 U4119 ( .CLK(n4237), .C(n4238) );
  CKBD0 U4120 ( .CLK(n4238), .C(n4239) );
  CKBD0 U4121 ( .CLK(n4239), .C(n4240) );
  CKBD0 U4122 ( .CLK(n4240), .C(n4241) );
  CKBD0 U4123 ( .CLK(n4241), .C(n4242) );
  CKBD0 U4124 ( .CLK(n4242), .C(n4243) );
  CKBD0 U4125 ( .CLK(n4243), .C(n4244) );
  BUFFD0 U4126 ( .I(n4244), .Z(n4245) );
  CKBD0 U4127 ( .CLK(n4245), .C(n4246) );
  CKBD0 U4128 ( .CLK(n4246), .C(n4247) );
  CKBD0 U4129 ( .CLK(n4247), .C(n4248) );
  CKBD0 U4130 ( .CLK(n4248), .C(n4249) );
  CKBD0 U4131 ( .CLK(n4249), .C(n4250) );
  CKBD0 U4132 ( .CLK(n4250), .C(n4251) );
  CKBD0 U4133 ( .CLK(n4251), .C(n4252) );
  CKBD0 U4134 ( .CLK(n4252), .C(n4253) );
  CKBD0 U4135 ( .CLK(n4253), .C(n4254) );
  BUFFD0 U4136 ( .I(n4254), .Z(n4255) );
  CKBD0 U4137 ( .CLK(n4255), .C(n4256) );
  CKBD0 U4138 ( .CLK(n4256), .C(n4257) );
  CKBD0 U4139 ( .CLK(n4257), .C(n4258) );
  CKBD0 U4140 ( .CLK(n4258), .C(n4259) );
  CKBD0 U4141 ( .CLK(n4259), .C(n4260) );
  CKBD0 U4142 ( .CLK(n4260), .C(n4261) );
  CKBD0 U4143 ( .CLK(n4261), .C(n4262) );
  CKBD0 U4144 ( .CLK(n4262), .C(n4263) );
  CKBD0 U4145 ( .CLK(n4263), .C(n4264) );
  CKBD0 U4146 ( .CLK(n4264), .C(n4265) );
  BUFFD0 U4147 ( .I(n4265), .Z(n4266) );
  CKBD0 U4148 ( .CLK(n4266), .C(n4267) );
  CKBD0 U4149 ( .CLK(n4267), .C(n4268) );
  CKBD0 U4150 ( .CLK(n4268), .C(n4269) );
  CKBD0 U4151 ( .CLK(n4269), .C(n4270) );
  CKBD0 U4152 ( .CLK(n4270), .C(n4271) );
  CKBD0 U4153 ( .CLK(n4271), .C(n4272) );
  CKBD0 U4154 ( .CLK(n4272), .C(n4273) );
  CKBD0 U4155 ( .CLK(n4273), .C(n4274) );
  CKBD0 U4156 ( .CLK(n4274), .C(n4275) );
  CKBD0 U4157 ( .CLK(n4275), .C(n4276) );
  BUFFD0 U4158 ( .I(n4276), .Z(n4277) );
  CKBD0 U4159 ( .CLK(n4277), .C(n4278) );
  CKBD0 U4160 ( .CLK(n4278), .C(n4279) );
  CKBD0 U4161 ( .CLK(n4279), .C(n4280) );
  CKBD0 U4162 ( .CLK(n4280), .C(n4281) );
  CKBD0 U4163 ( .CLK(n4281), .C(n4282) );
  CKBD0 U4164 ( .CLK(n4282), .C(n4283) );
  BUFFD0 U4165 ( .I(n4283), .Z(n4284) );
  CKBD0 U4166 ( .CLK(n4284), .C(n4285) );
  BUFFD0 U4167 ( .I(n4285), .Z(n4286) );
  CKBD0 U4168 ( .CLK(n4286), .C(n4287) );
  BUFFD0 U4169 ( .I(n4287), .Z(n4288) );
  CKBD0 U4170 ( .CLK(n4288), .C(n4289) );
  BUFFD0 U4171 ( .I(n4289), .Z(n4290) );
  CKBD0 U4172 ( .CLK(n4290), .C(n4291) );
  BUFFD0 U4173 ( .I(n4291), .Z(n4292) );
  CKBD0 U4174 ( .CLK(n4292), .C(n4293) );
  BUFFD0 U4175 ( .I(n4293), .Z(n4294) );
  CKBD0 U4176 ( .CLK(n4294), .C(n4295) );
  BUFFD0 U4177 ( .I(n4295), .Z(n4296) );
  CKBD0 U4178 ( .CLK(n4296), .C(n4297) );
  BUFFD0 U4179 ( .I(n4297), .Z(n4298) );
  BUFFD0 U4180 ( .I(n4300), .Z(n4299) );
  BUFFD0 U4181 ( .I(n4301), .Z(n4300) );
  BUFFD0 U4182 ( .I(n151), .Z(n4301) );
  CKBD0 U4183 ( .CLK(n1235), .C(n4302) );
  CKBD0 U4184 ( .CLK(n4302), .C(n4303) );
  CKBD0 U4185 ( .CLK(n4303), .C(n4304) );
  BUFFD0 U4186 ( .I(n4304), .Z(n4305) );
  CKBD0 U4187 ( .CLK(n4305), .C(n4306) );
  CKBD0 U4188 ( .CLK(n4306), .C(n4307) );
  CKBD0 U4189 ( .CLK(n4307), .C(n4308) );
  CKBD0 U4190 ( .CLK(n4308), .C(n4309) );
  CKBD0 U4191 ( .CLK(n4309), .C(n4310) );
  CKBD0 U4192 ( .CLK(n4310), .C(n4311) );
  CKBD0 U4193 ( .CLK(n4311), .C(n4312) );
  CKBD0 U4194 ( .CLK(n4312), .C(n4313) );
  CKBD0 U4195 ( .CLK(n4313), .C(n4314) );
  CKBD0 U4196 ( .CLK(n4314), .C(n4315) );
  BUFFD0 U4197 ( .I(n4315), .Z(n4316) );
  CKBD0 U4198 ( .CLK(n4316), .C(n4317) );
  CKBD0 U4199 ( .CLK(n4317), .C(n4318) );
  CKBD0 U4200 ( .CLK(n4318), .C(n4319) );
  CKBD0 U4201 ( .CLK(n4319), .C(n4320) );
  CKBD0 U4202 ( .CLK(n4320), .C(n4321) );
  CKBD0 U4203 ( .CLK(n4321), .C(n4322) );
  CKBD0 U4204 ( .CLK(n4322), .C(n4323) );
  CKBD0 U4205 ( .CLK(n4323), .C(n4324) );
  CKBD0 U4206 ( .CLK(n4324), .C(n4325) );
  BUFFD0 U4207 ( .I(n4325), .Z(n4326) );
  CKBD0 U4208 ( .CLK(n4326), .C(n4327) );
  CKBD0 U4209 ( .CLK(n4327), .C(n4328) );
  CKBD0 U4210 ( .CLK(n4328), .C(n4329) );
  CKBD0 U4211 ( .CLK(n4329), .C(n4330) );
  CKBD0 U4212 ( .CLK(n4330), .C(n4331) );
  CKBD0 U4213 ( .CLK(n4331), .C(n4332) );
  CKBD0 U4214 ( .CLK(n4332), .C(n4333) );
  CKBD0 U4215 ( .CLK(n4333), .C(n4334) );
  CKBD0 U4216 ( .CLK(n4334), .C(n4335) );
  CKBD0 U4217 ( .CLK(n4335), .C(n4336) );
  BUFFD0 U4218 ( .I(n4336), .Z(n4337) );
  CKBD0 U4219 ( .CLK(n4337), .C(n4338) );
  CKBD0 U4220 ( .CLK(n4338), .C(n4339) );
  CKBD0 U4221 ( .CLK(n4339), .C(n4340) );
  CKBD0 U4222 ( .CLK(n4340), .C(n4341) );
  CKBD0 U4223 ( .CLK(n4341), .C(n4342) );
  CKBD0 U4224 ( .CLK(n4342), .C(n4343) );
  CKBD0 U4225 ( .CLK(n4343), .C(n4344) );
  CKBD0 U4226 ( .CLK(n4344), .C(n4345) );
  CKBD0 U4227 ( .CLK(n4345), .C(n4346) );
  CKBD0 U4228 ( .CLK(n4346), .C(n4347) );
  BUFFD0 U4229 ( .I(n4347), .Z(n4348) );
  CKBD0 U4230 ( .CLK(n4348), .C(n4349) );
  CKBD0 U4231 ( .CLK(n4349), .C(n4350) );
  CKBD0 U4232 ( .CLK(n4350), .C(n4351) );
  CKBD0 U4233 ( .CLK(n4351), .C(n4352) );
  CKBD0 U4234 ( .CLK(n4352), .C(n4353) );
  CKBD0 U4235 ( .CLK(n4353), .C(n4354) );
  CKBD0 U4236 ( .CLK(n4354), .C(n4355) );
  CKBD0 U4237 ( .CLK(n4355), .C(n4356) );
  CKBD0 U4238 ( .CLK(n4356), .C(n4357) );
  CKBD0 U4239 ( .CLK(n4357), .C(n4358) );
  BUFFD0 U4240 ( .I(n4358), .Z(n4359) );
  CKBD0 U4241 ( .CLK(n4359), .C(n4360) );
  CKBD0 U4242 ( .CLK(n4360), .C(n4361) );
  CKBD0 U4243 ( .CLK(n4361), .C(n4362) );
  CKBD0 U4244 ( .CLK(n4362), .C(n4363) );
  CKBD0 U4245 ( .CLK(n4363), .C(n4364) );
  CKBD0 U4246 ( .CLK(n4364), .C(n4365) );
  CKBD0 U4247 ( .CLK(n4365), .C(n4366) );
  CKBD0 U4248 ( .CLK(n4366), .C(n4367) );
  CKBD0 U4249 ( .CLK(n4367), .C(n4368) );
  CKBD0 U4250 ( .CLK(n4368), .C(n4369) );
  BUFFD0 U4251 ( .I(n4369), .Z(n4370) );
  CKBD0 U4252 ( .CLK(n4370), .C(n4371) );
  CKBD0 U4253 ( .CLK(n4371), .C(n4372) );
  CKBD0 U4254 ( .CLK(n4372), .C(n4373) );
  CKBD0 U4255 ( .CLK(n4373), .C(n4374) );
  CKBD0 U4256 ( .CLK(n4374), .C(n4375) );
  CKBD0 U4257 ( .CLK(n4375), .C(n4376) );
  CKBD0 U4258 ( .CLK(n4376), .C(n4377) );
  CKBD0 U4259 ( .CLK(n4377), .C(n4378) );
  CKBD0 U4260 ( .CLK(n4378), .C(n4379) );
  CKBD0 U4261 ( .CLK(n4379), .C(n4380) );
  BUFFD0 U4262 ( .I(n4380), .Z(n4381) );
  CKBD0 U4263 ( .CLK(n4381), .C(n4382) );
  CKBD0 U4264 ( .CLK(n4382), .C(n4383) );
  CKBD0 U4265 ( .CLK(n4383), .C(n4384) );
  CKBD0 U4266 ( .CLK(n4384), .C(n4385) );
  CKBD0 U4267 ( .CLK(n4385), .C(n4386) );
  CKBD0 U4268 ( .CLK(n4386), .C(n4387) );
  CKBD0 U4269 ( .CLK(n4387), .C(n4388) );
  CKBD0 U4270 ( .CLK(n4388), .C(n4389) );
  CKBD0 U4271 ( .CLK(n4389), .C(n4390) );
  BUFFD0 U4272 ( .I(n4390), .Z(n4391) );
  CKBD0 U4273 ( .CLK(n4391), .C(n4392) );
  CKBD0 U4274 ( .CLK(n4392), .C(n4393) );
  CKBD0 U4275 ( .CLK(n4393), .C(n4394) );
  CKBD0 U4276 ( .CLK(n4394), .C(n4395) );
  CKBD0 U4277 ( .CLK(n4395), .C(n4396) );
  CKBD0 U4278 ( .CLK(n4396), .C(n4397) );
  CKBD0 U4279 ( .CLK(n4397), .C(n4398) );
  CKBD0 U4280 ( .CLK(n4398), .C(n4399) );
  CKBD0 U4281 ( .CLK(n4399), .C(n4400) );
  CKBD0 U4282 ( .CLK(n4400), .C(n4401) );
  BUFFD0 U4283 ( .I(n4401), .Z(n4402) );
  CKBD0 U4284 ( .CLK(n4402), .C(n4403) );
  CKBD0 U4285 ( .CLK(n4403), .C(n4404) );
  CKBD0 U4286 ( .CLK(n4404), .C(n4405) );
  CKBD0 U4287 ( .CLK(n4405), .C(n4406) );
  CKBD0 U4288 ( .CLK(n4406), .C(n4407) );
  CKBD0 U4289 ( .CLK(n4407), .C(n4408) );
  CKBD0 U4290 ( .CLK(n4408), .C(n4409) );
  CKBD0 U4291 ( .CLK(n4409), .C(n4410) );
  CKBD0 U4292 ( .CLK(n4410), .C(n4411) );
  CKBD0 U4293 ( .CLK(n4411), .C(n4412) );
  BUFFD0 U4294 ( .I(n4412), .Z(n4413) );
  CKBD0 U4295 ( .CLK(n4413), .C(n4414) );
  CKBD0 U4296 ( .CLK(n4414), .C(n4415) );
  CKBD0 U4297 ( .CLK(n4415), .C(n4416) );
  CKBD0 U4298 ( .CLK(n4416), .C(n4417) );
  CKBD0 U4299 ( .CLK(n4417), .C(n4418) );
  CKBD0 U4300 ( .CLK(n4418), .C(n4419) );
  BUFFD0 U4301 ( .I(n4419), .Z(n4420) );
  CKBD0 U4302 ( .CLK(n4420), .C(n4421) );
  BUFFD0 U4303 ( .I(n4421), .Z(n4422) );
  CKBD0 U4304 ( .CLK(n4422), .C(n4423) );
  BUFFD0 U4305 ( .I(n4423), .Z(n4424) );
  CKBD0 U4306 ( .CLK(n4424), .C(n4425) );
  BUFFD0 U4307 ( .I(n4425), .Z(n4426) );
  CKBD0 U4308 ( .CLK(n4426), .C(n4427) );
  BUFFD0 U4309 ( .I(n4427), .Z(n4428) );
  CKBD0 U4310 ( .CLK(n4428), .C(n4429) );
  BUFFD0 U4311 ( .I(n4429), .Z(n4430) );
  CKBD0 U4312 ( .CLK(n4430), .C(n4431) );
  BUFFD0 U4313 ( .I(n4431), .Z(n4432) );
  CKBD0 U4314 ( .CLK(n4432), .C(n4433) );
  BUFFD0 U4315 ( .I(n4433), .Z(n4434) );
  BUFFD0 U4316 ( .I(n4436), .Z(n4435) );
  BUFFD0 U4317 ( .I(n4437), .Z(n4436) );
  BUFFD0 U4318 ( .I(n150), .Z(n4437) );
  CKBD0 U4319 ( .CLK(n1233), .C(n4438) );
  CKBD0 U4320 ( .CLK(n4438), .C(n4439) );
  CKBD0 U4321 ( .CLK(n4439), .C(n4440) );
  BUFFD0 U4322 ( .I(n4440), .Z(n4441) );
  CKBD0 U4323 ( .CLK(n4441), .C(n4442) );
  CKBD0 U4324 ( .CLK(n4442), .C(n4443) );
  CKBD0 U4325 ( .CLK(n4443), .C(n4444) );
  CKBD0 U4326 ( .CLK(n4444), .C(n4445) );
  CKBD0 U4327 ( .CLK(n4445), .C(n4446) );
  CKBD0 U4328 ( .CLK(n4446), .C(n4447) );
  CKBD0 U4329 ( .CLK(n4447), .C(n4448) );
  CKBD0 U4330 ( .CLK(n4448), .C(n4449) );
  CKBD0 U4331 ( .CLK(n4449), .C(n4450) );
  CKBD0 U4332 ( .CLK(n4450), .C(n4451) );
  BUFFD0 U4333 ( .I(n4451), .Z(n4452) );
  CKBD0 U4334 ( .CLK(n4452), .C(n4453) );
  CKBD0 U4335 ( .CLK(n4453), .C(n4454) );
  CKBD0 U4336 ( .CLK(n4454), .C(n4455) );
  CKBD0 U4337 ( .CLK(n4455), .C(n4456) );
  CKBD0 U4338 ( .CLK(n4456), .C(n4457) );
  CKBD0 U4339 ( .CLK(n4457), .C(n4458) );
  CKBD0 U4340 ( .CLK(n4458), .C(n4459) );
  CKBD0 U4341 ( .CLK(n4459), .C(n4460) );
  CKBD0 U4342 ( .CLK(n4460), .C(n4461) );
  BUFFD0 U4343 ( .I(n4461), .Z(n4462) );
  CKBD0 U4344 ( .CLK(n4462), .C(n4463) );
  CKBD0 U4345 ( .CLK(n4463), .C(n4464) );
  CKBD0 U4346 ( .CLK(n4464), .C(n4465) );
  CKBD0 U4347 ( .CLK(n4465), .C(n4466) );
  CKBD0 U4348 ( .CLK(n4466), .C(n4467) );
  CKBD0 U4349 ( .CLK(n4467), .C(n4468) );
  CKBD0 U4350 ( .CLK(n4468), .C(n4469) );
  CKBD0 U4351 ( .CLK(n4469), .C(n4470) );
  CKBD0 U4352 ( .CLK(n4470), .C(n4471) );
  CKBD0 U4353 ( .CLK(n4471), .C(n4472) );
  BUFFD0 U4354 ( .I(n4472), .Z(n4473) );
  CKBD0 U4355 ( .CLK(n4473), .C(n4474) );
  CKBD0 U4356 ( .CLK(n4474), .C(n4475) );
  CKBD0 U4357 ( .CLK(n4475), .C(n4476) );
  CKBD0 U4358 ( .CLK(n4476), .C(n4477) );
  CKBD0 U4359 ( .CLK(n4477), .C(n4478) );
  CKBD0 U4360 ( .CLK(n4478), .C(n4479) );
  CKBD0 U4361 ( .CLK(n4479), .C(n4480) );
  CKBD0 U4362 ( .CLK(n4480), .C(n4481) );
  CKBD0 U4363 ( .CLK(n4481), .C(n4482) );
  CKBD0 U4364 ( .CLK(n4482), .C(n4483) );
  BUFFD0 U4365 ( .I(n4483), .Z(n4484) );
  CKBD0 U4366 ( .CLK(n4484), .C(n4485) );
  CKBD0 U4367 ( .CLK(n4485), .C(n4486) );
  CKBD0 U4368 ( .CLK(n4486), .C(n4487) );
  CKBD0 U4369 ( .CLK(n4487), .C(n4488) );
  CKBD0 U4370 ( .CLK(n4488), .C(n4489) );
  CKBD0 U4371 ( .CLK(n4489), .C(n4490) );
  CKBD0 U4372 ( .CLK(n4490), .C(n4491) );
  CKBD0 U4373 ( .CLK(n4491), .C(n4492) );
  CKBD0 U4374 ( .CLK(n4492), .C(n4493) );
  CKBD0 U4375 ( .CLK(n4493), .C(n4494) );
  BUFFD0 U4376 ( .I(n4494), .Z(n4495) );
  CKBD0 U4377 ( .CLK(n4495), .C(n4496) );
  CKBD0 U4378 ( .CLK(n4496), .C(n4497) );
  CKBD0 U4379 ( .CLK(n4497), .C(n4498) );
  CKBD0 U4380 ( .CLK(n4498), .C(n4499) );
  CKBD0 U4381 ( .CLK(n4499), .C(n4500) );
  CKBD0 U4382 ( .CLK(n4500), .C(n4501) );
  CKBD0 U4383 ( .CLK(n4501), .C(n4502) );
  CKBD0 U4384 ( .CLK(n4502), .C(n4503) );
  CKBD0 U4385 ( .CLK(n4503), .C(n4504) );
  CKBD0 U4386 ( .CLK(n4504), .C(n4505) );
  BUFFD0 U4387 ( .I(n4505), .Z(n4506) );
  CKBD0 U4388 ( .CLK(n4506), .C(n4507) );
  CKBD0 U4389 ( .CLK(n4507), .C(n4508) );
  CKBD0 U4390 ( .CLK(n4508), .C(n4509) );
  CKBD0 U4391 ( .CLK(n4509), .C(n4510) );
  CKBD0 U4392 ( .CLK(n4510), .C(n4511) );
  CKBD0 U4393 ( .CLK(n4511), .C(n4512) );
  CKBD0 U4394 ( .CLK(n4512), .C(n4513) );
  CKBD0 U4395 ( .CLK(n4513), .C(n4514) );
  CKBD0 U4396 ( .CLK(n4514), .C(n4515) );
  CKBD0 U4397 ( .CLK(n4515), .C(n4516) );
  BUFFD0 U4398 ( .I(n4516), .Z(n4517) );
  CKBD0 U4399 ( .CLK(n4517), .C(n4518) );
  CKBD0 U4400 ( .CLK(n4518), .C(n4519) );
  CKBD0 U4401 ( .CLK(n4519), .C(n4520) );
  CKBD0 U4402 ( .CLK(n4520), .C(n4521) );
  CKBD0 U4403 ( .CLK(n4521), .C(n4522) );
  CKBD0 U4404 ( .CLK(n4522), .C(n4523) );
  CKBD0 U4405 ( .CLK(n4523), .C(n4524) );
  CKBD0 U4406 ( .CLK(n4524), .C(n4525) );
  CKBD0 U4407 ( .CLK(n4525), .C(n4526) );
  BUFFD0 U4408 ( .I(n4526), .Z(n4527) );
  CKBD0 U4409 ( .CLK(n4527), .C(n4528) );
  CKBD0 U4410 ( .CLK(n4528), .C(n4529) );
  CKBD0 U4411 ( .CLK(n4529), .C(n4530) );
  CKBD0 U4412 ( .CLK(n4530), .C(n4531) );
  CKBD0 U4413 ( .CLK(n4531), .C(n4532) );
  CKBD0 U4414 ( .CLK(n4532), .C(n4533) );
  CKBD0 U4415 ( .CLK(n4533), .C(n4534) );
  CKBD0 U4416 ( .CLK(n4534), .C(n4535) );
  CKBD0 U4417 ( .CLK(n4535), .C(n4536) );
  CKBD0 U4418 ( .CLK(n4536), .C(n4537) );
  BUFFD0 U4419 ( .I(n4537), .Z(n4538) );
  CKBD0 U4420 ( .CLK(n4538), .C(n4539) );
  CKBD0 U4421 ( .CLK(n4539), .C(n4540) );
  CKBD0 U4422 ( .CLK(n4540), .C(n4541) );
  CKBD0 U4423 ( .CLK(n4541), .C(n4542) );
  CKBD0 U4424 ( .CLK(n4542), .C(n4543) );
  CKBD0 U4425 ( .CLK(n4543), .C(n4544) );
  CKBD0 U4426 ( .CLK(n4544), .C(n4545) );
  CKBD0 U4427 ( .CLK(n4545), .C(n4546) );
  CKBD0 U4428 ( .CLK(n4546), .C(n4547) );
  CKBD0 U4429 ( .CLK(n4547), .C(n4548) );
  BUFFD0 U4430 ( .I(n4548), .Z(n4549) );
  CKBD0 U4431 ( .CLK(n4549), .C(n4550) );
  CKBD0 U4432 ( .CLK(n4550), .C(n4551) );
  CKBD0 U4433 ( .CLK(n4551), .C(n4552) );
  CKBD0 U4434 ( .CLK(n4552), .C(n4553) );
  CKBD0 U4435 ( .CLK(n4553), .C(n4554) );
  CKBD0 U4436 ( .CLK(n4554), .C(n4555) );
  BUFFD0 U4437 ( .I(n4555), .Z(n4556) );
  CKBD0 U4438 ( .CLK(n4556), .C(n4557) );
  BUFFD0 U4439 ( .I(n4557), .Z(n4558) );
  CKBD0 U4440 ( .CLK(n4558), .C(n4559) );
  BUFFD0 U4441 ( .I(n4559), .Z(n4560) );
  CKBD0 U4442 ( .CLK(n4560), .C(n4561) );
  BUFFD0 U4443 ( .I(n4561), .Z(n4562) );
  CKBD0 U4444 ( .CLK(n4562), .C(n4563) );
  BUFFD0 U4445 ( .I(n4563), .Z(n4564) );
  CKBD0 U4446 ( .CLK(n4564), .C(n4565) );
  BUFFD0 U4447 ( .I(n4565), .Z(n4566) );
  CKBD0 U4448 ( .CLK(n4566), .C(n4567) );
  BUFFD0 U4449 ( .I(n4567), .Z(n4568) );
  CKBD0 U4450 ( .CLK(n4568), .C(n4569) );
  BUFFD0 U4451 ( .I(n4569), .Z(n4570) );
  BUFFD0 U4452 ( .I(n4572), .Z(n4571) );
  BUFFD0 U4453 ( .I(n4573), .Z(n4572) );
  BUFFD0 U4454 ( .I(n149), .Z(n4573) );
  CKBD0 U4455 ( .CLK(n1231), .C(n4574) );
  CKBD0 U4456 ( .CLK(n4574), .C(n4575) );
  CKBD0 U4457 ( .CLK(n4575), .C(n4576) );
  BUFFD0 U4458 ( .I(n4576), .Z(n4577) );
  CKBD0 U4459 ( .CLK(n4577), .C(n4578) );
  CKBD0 U4460 ( .CLK(n4578), .C(n4579) );
  CKBD0 U4461 ( .CLK(n4579), .C(n4580) );
  CKBD0 U4462 ( .CLK(n4580), .C(n4581) );
  CKBD0 U4463 ( .CLK(n4581), .C(n4582) );
  CKBD0 U4464 ( .CLK(n4582), .C(n4583) );
  CKBD0 U4465 ( .CLK(n4583), .C(n4584) );
  CKBD0 U4466 ( .CLK(n4584), .C(n4585) );
  CKBD0 U4467 ( .CLK(n4585), .C(n4586) );
  CKBD0 U4468 ( .CLK(n4586), .C(n4587) );
  BUFFD0 U4469 ( .I(n4587), .Z(n4588) );
  CKBD0 U4470 ( .CLK(n4588), .C(n4589) );
  CKBD0 U4471 ( .CLK(n4589), .C(n4590) );
  CKBD0 U4472 ( .CLK(n4590), .C(n4591) );
  CKBD0 U4473 ( .CLK(n4591), .C(n4592) );
  CKBD0 U4474 ( .CLK(n4592), .C(n4593) );
  CKBD0 U4475 ( .CLK(n4593), .C(n4594) );
  CKBD0 U4476 ( .CLK(n4594), .C(n4595) );
  CKBD0 U4477 ( .CLK(n4595), .C(n4596) );
  CKBD0 U4478 ( .CLK(n4596), .C(n4597) );
  BUFFD0 U4479 ( .I(n4597), .Z(n4598) );
  CKBD0 U4480 ( .CLK(n4598), .C(n4599) );
  CKBD0 U4481 ( .CLK(n4599), .C(n4600) );
  CKBD0 U4482 ( .CLK(n4600), .C(n4601) );
  CKBD0 U4483 ( .CLK(n4601), .C(n4602) );
  CKBD0 U4484 ( .CLK(n4602), .C(n4603) );
  CKBD0 U4485 ( .CLK(n4603), .C(n4604) );
  CKBD0 U4486 ( .CLK(n4604), .C(n4605) );
  CKBD0 U4487 ( .CLK(n4605), .C(n4606) );
  CKBD0 U4488 ( .CLK(n4606), .C(n4607) );
  CKBD0 U4489 ( .CLK(n4607), .C(n4608) );
  BUFFD0 U4490 ( .I(n4608), .Z(n4609) );
  CKBD0 U4491 ( .CLK(n4609), .C(n4610) );
  CKBD0 U4492 ( .CLK(n4610), .C(n4611) );
  CKBD0 U4493 ( .CLK(n4611), .C(n4612) );
  CKBD0 U4494 ( .CLK(n4612), .C(n4613) );
  CKBD0 U4495 ( .CLK(n4613), .C(n4614) );
  CKBD0 U4496 ( .CLK(n4614), .C(n4615) );
  CKBD0 U4497 ( .CLK(n4615), .C(n4616) );
  CKBD0 U4498 ( .CLK(n4616), .C(n4617) );
  CKBD0 U4499 ( .CLK(n4617), .C(n4618) );
  CKBD0 U4500 ( .CLK(n4618), .C(n4619) );
  BUFFD0 U4501 ( .I(n4619), .Z(n4620) );
  CKBD0 U4502 ( .CLK(n4620), .C(n4621) );
  CKBD0 U4503 ( .CLK(n4621), .C(n4622) );
  CKBD0 U4504 ( .CLK(n4622), .C(n4623) );
  CKBD0 U4505 ( .CLK(n4623), .C(n4624) );
  CKBD0 U4506 ( .CLK(n4624), .C(n4625) );
  CKBD0 U4507 ( .CLK(n4625), .C(n4626) );
  CKBD0 U4508 ( .CLK(n4626), .C(n4627) );
  CKBD0 U4509 ( .CLK(n4627), .C(n4628) );
  CKBD0 U4510 ( .CLK(n4628), .C(n4629) );
  CKBD0 U4511 ( .CLK(n4629), .C(n4630) );
  BUFFD0 U4512 ( .I(n4630), .Z(n4631) );
  CKBD0 U4513 ( .CLK(n4631), .C(n4632) );
  CKBD0 U4514 ( .CLK(n4632), .C(n4633) );
  CKBD0 U4515 ( .CLK(n4633), .C(n4634) );
  CKBD0 U4516 ( .CLK(n4634), .C(n4635) );
  CKBD0 U4517 ( .CLK(n4635), .C(n4636) );
  CKBD0 U4518 ( .CLK(n4636), .C(n4637) );
  CKBD0 U4519 ( .CLK(n4637), .C(n4638) );
  CKBD0 U4520 ( .CLK(n4638), .C(n4639) );
  CKBD0 U4521 ( .CLK(n4639), .C(n4640) );
  CKBD0 U4522 ( .CLK(n4640), .C(n4641) );
  BUFFD0 U4523 ( .I(n4641), .Z(n4642) );
  CKBD0 U4524 ( .CLK(n4642), .C(n4643) );
  CKBD0 U4525 ( .CLK(n4643), .C(n4644) );
  CKBD0 U4526 ( .CLK(n4644), .C(n4645) );
  CKBD0 U4527 ( .CLK(n4645), .C(n4646) );
  CKBD0 U4528 ( .CLK(n4646), .C(n4647) );
  CKBD0 U4529 ( .CLK(n4647), .C(n4648) );
  CKBD0 U4530 ( .CLK(n4648), .C(n4649) );
  CKBD0 U4531 ( .CLK(n4649), .C(n4650) );
  CKBD0 U4532 ( .CLK(n4650), .C(n4651) );
  CKBD0 U4533 ( .CLK(n4651), .C(n4652) );
  BUFFD0 U4534 ( .I(n4652), .Z(n4653) );
  CKBD0 U4535 ( .CLK(n4653), .C(n4654) );
  CKBD0 U4536 ( .CLK(n4654), .C(n4655) );
  CKBD0 U4537 ( .CLK(n4655), .C(n4656) );
  CKBD0 U4538 ( .CLK(n4656), .C(n4657) );
  CKBD0 U4539 ( .CLK(n4657), .C(n4658) );
  CKBD0 U4540 ( .CLK(n4658), .C(n4659) );
  CKBD0 U4541 ( .CLK(n4659), .C(n4660) );
  CKBD0 U4542 ( .CLK(n4660), .C(n4661) );
  CKBD0 U4543 ( .CLK(n4661), .C(n4662) );
  BUFFD0 U4544 ( .I(n4662), .Z(n4663) );
  CKBD0 U4545 ( .CLK(n4663), .C(n4664) );
  CKBD0 U4546 ( .CLK(n4664), .C(n4665) );
  CKBD0 U4547 ( .CLK(n4665), .C(n4666) );
  CKBD0 U4548 ( .CLK(n4666), .C(n4667) );
  CKBD0 U4549 ( .CLK(n4667), .C(n4668) );
  CKBD0 U4550 ( .CLK(n4668), .C(n4669) );
  CKBD0 U4551 ( .CLK(n4669), .C(n4670) );
  CKBD0 U4552 ( .CLK(n4670), .C(n4671) );
  CKBD0 U4553 ( .CLK(n4671), .C(n4672) );
  CKBD0 U4554 ( .CLK(n4672), .C(n4673) );
  BUFFD0 U4555 ( .I(n4673), .Z(n4674) );
  CKBD0 U4556 ( .CLK(n4674), .C(n4675) );
  CKBD0 U4557 ( .CLK(n4675), .C(n4676) );
  CKBD0 U4558 ( .CLK(n4676), .C(n4677) );
  CKBD0 U4559 ( .CLK(n4677), .C(n4678) );
  CKBD0 U4560 ( .CLK(n4678), .C(n4679) );
  CKBD0 U4561 ( .CLK(n4679), .C(n4680) );
  CKBD0 U4562 ( .CLK(n4680), .C(n4681) );
  CKBD0 U4563 ( .CLK(n4681), .C(n4682) );
  CKBD0 U4564 ( .CLK(n4682), .C(n4683) );
  CKBD0 U4565 ( .CLK(n4683), .C(n4684) );
  BUFFD0 U4566 ( .I(n4684), .Z(n4685) );
  CKBD0 U4567 ( .CLK(n4685), .C(n4686) );
  CKBD0 U4568 ( .CLK(n4686), .C(n4687) );
  CKBD0 U4569 ( .CLK(n4687), .C(n4688) );
  CKBD0 U4570 ( .CLK(n4688), .C(n4689) );
  CKBD0 U4571 ( .CLK(n4689), .C(n4690) );
  CKBD0 U4572 ( .CLK(n4690), .C(n4691) );
  BUFFD0 U4573 ( .I(n4691), .Z(n4692) );
  CKBD0 U4574 ( .CLK(n4692), .C(n4693) );
  BUFFD0 U4575 ( .I(n4693), .Z(n4694) );
  CKBD0 U4576 ( .CLK(n4694), .C(n4695) );
  BUFFD0 U4577 ( .I(n4695), .Z(n4696) );
  CKBD0 U4578 ( .CLK(n4696), .C(n4697) );
  BUFFD0 U4579 ( .I(n4697), .Z(n4698) );
  CKBD0 U4580 ( .CLK(n4698), .C(n4699) );
  BUFFD0 U4581 ( .I(n4699), .Z(n4700) );
  CKBD0 U4582 ( .CLK(n4700), .C(n4701) );
  BUFFD0 U4583 ( .I(n4701), .Z(n4702) );
  CKBD0 U4584 ( .CLK(n4702), .C(n4703) );
  BUFFD0 U4585 ( .I(n4703), .Z(n4704) );
  CKBD0 U4586 ( .CLK(n4704), .C(n4705) );
  BUFFD0 U4587 ( .I(n4705), .Z(n4706) );
  BUFFD0 U4588 ( .I(n4708), .Z(n4707) );
  BUFFD0 U4589 ( .I(n4709), .Z(n4708) );
  BUFFD0 U4590 ( .I(n148), .Z(n4709) );
  CKBD0 U4591 ( .CLK(n714), .C(n4710) );
  CKBD0 U4592 ( .CLK(n4710), .C(n4711) );
  CKBD0 U4593 ( .CLK(n4711), .C(n4712) );
  BUFFD0 U4594 ( .I(n4712), .Z(n4713) );
  CKBD0 U4595 ( .CLK(n4713), .C(n4714) );
  CKBD0 U4596 ( .CLK(n4714), .C(n4715) );
  CKBD0 U4597 ( .CLK(n4715), .C(n4716) );
  CKBD0 U4598 ( .CLK(n4716), .C(n4717) );
  CKBD0 U4599 ( .CLK(n4717), .C(n4718) );
  CKBD0 U4600 ( .CLK(n4718), .C(n4719) );
  CKBD0 U4601 ( .CLK(n4719), .C(n4720) );
  CKBD0 U4602 ( .CLK(n4720), .C(n4721) );
  CKBD0 U4603 ( .CLK(n4721), .C(n4722) );
  CKBD0 U4604 ( .CLK(n4722), .C(n4723) );
  BUFFD0 U4605 ( .I(n4723), .Z(n4724) );
  CKBD0 U4606 ( .CLK(n4724), .C(n4725) );
  CKBD0 U4607 ( .CLK(n4725), .C(n4726) );
  CKBD0 U4608 ( .CLK(n4726), .C(n4727) );
  CKBD0 U4609 ( .CLK(n4727), .C(n4728) );
  CKBD0 U4610 ( .CLK(n4728), .C(n4729) );
  CKBD0 U4611 ( .CLK(n4729), .C(n4730) );
  CKBD0 U4612 ( .CLK(n4730), .C(n4731) );
  CKBD0 U4613 ( .CLK(n4731), .C(n4732) );
  CKBD0 U4614 ( .CLK(n4732), .C(n4733) );
  BUFFD0 U4615 ( .I(n4733), .Z(n4734) );
  CKBD0 U4616 ( .CLK(n4734), .C(n4735) );
  CKBD0 U4617 ( .CLK(n4735), .C(n4736) );
  CKBD0 U4618 ( .CLK(n4736), .C(n4737) );
  CKBD0 U4619 ( .CLK(n4737), .C(n4738) );
  CKBD0 U4620 ( .CLK(n4738), .C(n4739) );
  CKBD0 U4621 ( .CLK(n4739), .C(n4740) );
  CKBD0 U4622 ( .CLK(n4740), .C(n4741) );
  CKBD0 U4623 ( .CLK(n4741), .C(n4742) );
  CKBD0 U4624 ( .CLK(n4742), .C(n4743) );
  CKBD0 U4625 ( .CLK(n4743), .C(n4744) );
  BUFFD0 U4626 ( .I(n4744), .Z(n4745) );
  CKBD0 U4627 ( .CLK(n4745), .C(n4746) );
  CKBD0 U4628 ( .CLK(n4746), .C(n4747) );
  CKBD0 U4629 ( .CLK(n4747), .C(n4748) );
  CKBD0 U4630 ( .CLK(n4748), .C(n4749) );
  CKBD0 U4631 ( .CLK(n4749), .C(n4750) );
  CKBD0 U4632 ( .CLK(n4750), .C(n4751) );
  CKBD0 U4633 ( .CLK(n4751), .C(n4752) );
  CKBD0 U4634 ( .CLK(n4752), .C(n4753) );
  CKBD0 U4635 ( .CLK(n4753), .C(n4754) );
  CKBD0 U4636 ( .CLK(n4754), .C(n4755) );
  BUFFD0 U4637 ( .I(n4755), .Z(n4756) );
  CKBD0 U4638 ( .CLK(n4756), .C(n4757) );
  CKBD0 U4639 ( .CLK(n4757), .C(n4758) );
  CKBD0 U4640 ( .CLK(n4758), .C(n4759) );
  CKBD0 U4641 ( .CLK(n4759), .C(n4760) );
  CKBD0 U4642 ( .CLK(n4760), .C(n4761) );
  CKBD0 U4643 ( .CLK(n4761), .C(n4762) );
  CKBD0 U4644 ( .CLK(n4762), .C(n4763) );
  CKBD0 U4645 ( .CLK(n4763), .C(n4764) );
  CKBD0 U4646 ( .CLK(n4764), .C(n4765) );
  CKBD0 U4647 ( .CLK(n4765), .C(n4766) );
  BUFFD0 U4648 ( .I(n4766), .Z(n4767) );
  CKBD0 U4649 ( .CLK(n4767), .C(n4768) );
  CKBD0 U4650 ( .CLK(n4768), .C(n4769) );
  CKBD0 U4651 ( .CLK(n4769), .C(n4770) );
  CKBD0 U4652 ( .CLK(n4770), .C(n4771) );
  CKBD0 U4653 ( .CLK(n4771), .C(n4772) );
  CKBD0 U4654 ( .CLK(n4772), .C(n4773) );
  CKBD0 U4655 ( .CLK(n4773), .C(n4774) );
  CKBD0 U4656 ( .CLK(n4774), .C(n4775) );
  CKBD0 U4657 ( .CLK(n4775), .C(n4776) );
  CKBD0 U4658 ( .CLK(n4776), .C(n4777) );
  BUFFD0 U4659 ( .I(n4777), .Z(n4778) );
  CKBD0 U4660 ( .CLK(n4778), .C(n4779) );
  CKBD0 U4661 ( .CLK(n4779), .C(n4780) );
  CKBD0 U4662 ( .CLK(n4780), .C(n4781) );
  CKBD0 U4663 ( .CLK(n4781), .C(n4782) );
  CKBD0 U4664 ( .CLK(n4782), .C(n4783) );
  CKBD0 U4665 ( .CLK(n4783), .C(n4784) );
  CKBD0 U4666 ( .CLK(n4784), .C(n4785) );
  CKBD0 U4667 ( .CLK(n4785), .C(n4786) );
  CKBD0 U4668 ( .CLK(n4786), .C(n4787) );
  CKBD0 U4669 ( .CLK(n4787), .C(n4788) );
  BUFFD0 U4670 ( .I(n4788), .Z(n4789) );
  CKBD0 U4671 ( .CLK(n4789), .C(n4790) );
  CKBD0 U4672 ( .CLK(n4790), .C(n4791) );
  CKBD0 U4673 ( .CLK(n4791), .C(n4792) );
  CKBD0 U4674 ( .CLK(n4792), .C(n4793) );
  CKBD0 U4675 ( .CLK(n4793), .C(n4794) );
  CKBD0 U4676 ( .CLK(n4794), .C(n4795) );
  CKBD0 U4677 ( .CLK(n4795), .C(n4796) );
  CKBD0 U4678 ( .CLK(n4796), .C(n4797) );
  CKBD0 U4679 ( .CLK(n4797), .C(n4798) );
  BUFFD0 U4680 ( .I(n4798), .Z(n4799) );
  CKBD0 U4681 ( .CLK(n4799), .C(n4800) );
  CKBD0 U4682 ( .CLK(n4800), .C(n4801) );
  CKBD0 U4683 ( .CLK(n4801), .C(n4802) );
  CKBD0 U4684 ( .CLK(n4802), .C(n4803) );
  CKBD0 U4685 ( .CLK(n4803), .C(n4804) );
  CKBD0 U4686 ( .CLK(n4804), .C(n4805) );
  CKBD0 U4687 ( .CLK(n4805), .C(n4806) );
  CKBD0 U4688 ( .CLK(n4806), .C(n4807) );
  CKBD0 U4689 ( .CLK(n4807), .C(n4808) );
  CKBD0 U4690 ( .CLK(n4808), .C(n4809) );
  BUFFD0 U4691 ( .I(n4809), .Z(n4810) );
  CKBD0 U4692 ( .CLK(n4810), .C(n4811) );
  CKBD0 U4693 ( .CLK(n4811), .C(n4812) );
  CKBD0 U4694 ( .CLK(n4812), .C(n4813) );
  CKBD0 U4695 ( .CLK(n4813), .C(n4814) );
  CKBD0 U4696 ( .CLK(n4814), .C(n4815) );
  CKBD0 U4697 ( .CLK(n4815), .C(n4816) );
  CKBD0 U4698 ( .CLK(n4816), .C(n4817) );
  CKBD0 U4699 ( .CLK(n4817), .C(n4818) );
  CKBD0 U4700 ( .CLK(n4818), .C(n4819) );
  CKBD0 U4701 ( .CLK(n4819), .C(n4820) );
  BUFFD0 U4702 ( .I(n4820), .Z(n4821) );
  CKBD0 U4703 ( .CLK(n4821), .C(n4822) );
  CKBD0 U4704 ( .CLK(n4822), .C(n4823) );
  CKBD0 U4705 ( .CLK(n4823), .C(n4824) );
  CKBD0 U4706 ( .CLK(n4824), .C(n4825) );
  CKBD0 U4707 ( .CLK(n4825), .C(n4826) );
  CKBD0 U4708 ( .CLK(n4826), .C(n4827) );
  BUFFD0 U4709 ( .I(n4827), .Z(n4828) );
  CKBD0 U4710 ( .CLK(n4828), .C(n4829) );
  BUFFD0 U4711 ( .I(n4829), .Z(n4830) );
  CKBD0 U4712 ( .CLK(n4830), .C(n4831) );
  BUFFD0 U4713 ( .I(n4831), .Z(n4832) );
  CKBD0 U4714 ( .CLK(n4832), .C(n4833) );
  BUFFD0 U4715 ( .I(n4833), .Z(n4834) );
  CKBD0 U4716 ( .CLK(n4834), .C(n4835) );
  BUFFD0 U4717 ( .I(n4835), .Z(n4836) );
  CKBD0 U4718 ( .CLK(n4836), .C(n4837) );
  BUFFD0 U4719 ( .I(n4837), .Z(n4838) );
  CKBD0 U4720 ( .CLK(n4838), .C(n4839) );
  BUFFD0 U4721 ( .I(n4839), .Z(n4840) );
  CKBD0 U4722 ( .CLK(n4840), .C(n4841) );
  BUFFD0 U4723 ( .I(n4841), .Z(n4842) );
  BUFFD0 U4724 ( .I(n4844), .Z(n4843) );
  BUFFD0 U4725 ( .I(n4845), .Z(n4844) );
  BUFFD0 U4726 ( .I(n147), .Z(n4845) );
  CKBD0 U4727 ( .CLK(n1132), .C(n4846) );
  CKBD0 U4728 ( .CLK(n4846), .C(n4847) );
  CKBD0 U4729 ( .CLK(n4847), .C(n4848) );
  BUFFD0 U4730 ( .I(n4848), .Z(n4849) );
  CKBD0 U4731 ( .CLK(n4849), .C(n4850) );
  CKBD0 U4732 ( .CLK(n4850), .C(n4851) );
  CKBD0 U4733 ( .CLK(n4851), .C(n4852) );
  CKBD0 U4734 ( .CLK(n4852), .C(n4853) );
  CKBD0 U4735 ( .CLK(n4853), .C(n4854) );
  CKBD0 U4736 ( .CLK(n4854), .C(n4855) );
  CKBD0 U4737 ( .CLK(n4855), .C(n4856) );
  CKBD0 U4738 ( .CLK(n4856), .C(n4857) );
  CKBD0 U4739 ( .CLK(n4857), .C(n4858) );
  CKBD0 U4740 ( .CLK(n4858), .C(n4859) );
  BUFFD0 U4741 ( .I(n4859), .Z(n4860) );
  CKBD0 U4742 ( .CLK(n4860), .C(n4861) );
  CKBD0 U4743 ( .CLK(n4861), .C(n4862) );
  CKBD0 U4744 ( .CLK(n4862), .C(n4863) );
  CKBD0 U4745 ( .CLK(n4863), .C(n4864) );
  CKBD0 U4746 ( .CLK(n4864), .C(n4865) );
  CKBD0 U4747 ( .CLK(n4865), .C(n4866) );
  CKBD0 U4748 ( .CLK(n4866), .C(n4867) );
  CKBD0 U4749 ( .CLK(n4867), .C(n4868) );
  CKBD0 U4750 ( .CLK(n4868), .C(n4869) );
  BUFFD0 U4751 ( .I(n4869), .Z(n4870) );
  CKBD0 U4752 ( .CLK(n4870), .C(n4871) );
  CKBD0 U4753 ( .CLK(n4871), .C(n4872) );
  CKBD0 U4754 ( .CLK(n4872), .C(n4873) );
  CKBD0 U4755 ( .CLK(n4873), .C(n4874) );
  CKBD0 U4756 ( .CLK(n4874), .C(n4875) );
  CKBD0 U4757 ( .CLK(n4875), .C(n4876) );
  CKBD0 U4758 ( .CLK(n4876), .C(n4877) );
  CKBD0 U4759 ( .CLK(n4877), .C(n4878) );
  CKBD0 U4760 ( .CLK(n4878), .C(n4879) );
  CKBD0 U4761 ( .CLK(n4879), .C(n4880) );
  BUFFD0 U4762 ( .I(n4880), .Z(n4881) );
  CKBD0 U4763 ( .CLK(n4881), .C(n4882) );
  CKBD0 U4764 ( .CLK(n4882), .C(n4883) );
  CKBD0 U4765 ( .CLK(n4883), .C(n4884) );
  CKBD0 U4766 ( .CLK(n4884), .C(n4885) );
  CKBD0 U4767 ( .CLK(n4885), .C(n4886) );
  CKBD0 U4768 ( .CLK(n4886), .C(n4887) );
  CKBD0 U4769 ( .CLK(n4887), .C(n4888) );
  CKBD0 U4770 ( .CLK(n4888), .C(n4889) );
  CKBD0 U4771 ( .CLK(n4889), .C(n4890) );
  CKBD0 U4772 ( .CLK(n4890), .C(n4891) );
  BUFFD0 U4773 ( .I(n4891), .Z(n4892) );
  CKBD0 U4774 ( .CLK(n4892), .C(n4893) );
  CKBD0 U4775 ( .CLK(n4893), .C(n4894) );
  CKBD0 U4776 ( .CLK(n4894), .C(n4895) );
  CKBD0 U4777 ( .CLK(n4895), .C(n4896) );
  CKBD0 U4778 ( .CLK(n4896), .C(n4897) );
  CKBD0 U4779 ( .CLK(n4897), .C(n4898) );
  CKBD0 U4780 ( .CLK(n4898), .C(n4899) );
  CKBD0 U4781 ( .CLK(n4899), .C(n4900) );
  CKBD0 U4782 ( .CLK(n4900), .C(n4901) );
  CKBD0 U4783 ( .CLK(n4901), .C(n4902) );
  BUFFD0 U4784 ( .I(n4902), .Z(n4903) );
  CKBD0 U4785 ( .CLK(n4903), .C(n4904) );
  CKBD0 U4786 ( .CLK(n4904), .C(n4905) );
  CKBD0 U4787 ( .CLK(n4905), .C(n4906) );
  CKBD0 U4788 ( .CLK(n4906), .C(n4907) );
  CKBD0 U4789 ( .CLK(n4907), .C(n4908) );
  CKBD0 U4790 ( .CLK(n4908), .C(n4909) );
  CKBD0 U4791 ( .CLK(n4909), .C(n4910) );
  CKBD0 U4792 ( .CLK(n4910), .C(n4911) );
  CKBD0 U4793 ( .CLK(n4911), .C(n4912) );
  CKBD0 U4794 ( .CLK(n4912), .C(n4913) );
  BUFFD0 U4795 ( .I(n4913), .Z(n4914) );
  CKBD0 U4796 ( .CLK(n4914), .C(n4915) );
  CKBD0 U4797 ( .CLK(n4915), .C(n4916) );
  CKBD0 U4798 ( .CLK(n4916), .C(n4917) );
  CKBD0 U4799 ( .CLK(n4917), .C(n4918) );
  CKBD0 U4800 ( .CLK(n4918), .C(n4919) );
  CKBD0 U4801 ( .CLK(n4919), .C(n4920) );
  CKBD0 U4802 ( .CLK(n4920), .C(n4921) );
  CKBD0 U4803 ( .CLK(n4921), .C(n4922) );
  CKBD0 U4804 ( .CLK(n4922), .C(n4923) );
  CKBD0 U4805 ( .CLK(n4923), .C(n4924) );
  BUFFD0 U4806 ( .I(n4924), .Z(n4925) );
  CKBD0 U4807 ( .CLK(n4925), .C(n4926) );
  CKBD0 U4808 ( .CLK(n4926), .C(n4927) );
  CKBD0 U4809 ( .CLK(n4927), .C(n4928) );
  CKBD0 U4810 ( .CLK(n4928), .C(n4929) );
  CKBD0 U4811 ( .CLK(n4929), .C(n4930) );
  CKBD0 U4812 ( .CLK(n4930), .C(n4931) );
  CKBD0 U4813 ( .CLK(n4931), .C(n4932) );
  CKBD0 U4814 ( .CLK(n4932), .C(n4933) );
  CKBD0 U4815 ( .CLK(n4933), .C(n4934) );
  BUFFD0 U4816 ( .I(n4934), .Z(n4935) );
  CKBD0 U4817 ( .CLK(n4935), .C(n4936) );
  CKBD0 U4818 ( .CLK(n4936), .C(n4937) );
  CKBD0 U4819 ( .CLK(n4937), .C(n4938) );
  CKBD0 U4820 ( .CLK(n4938), .C(n4939) );
  CKBD0 U4821 ( .CLK(n4939), .C(n4940) );
  CKBD0 U4822 ( .CLK(n4940), .C(n4941) );
  CKBD0 U4823 ( .CLK(n4941), .C(n4942) );
  CKBD0 U4824 ( .CLK(n4942), .C(n4943) );
  CKBD0 U4825 ( .CLK(n4943), .C(n4944) );
  CKBD0 U4826 ( .CLK(n4944), .C(n4945) );
  BUFFD0 U4827 ( .I(n4945), .Z(n4946) );
  CKBD0 U4828 ( .CLK(n4946), .C(n4947) );
  CKBD0 U4829 ( .CLK(n4947), .C(n4948) );
  CKBD0 U4830 ( .CLK(n4948), .C(n4949) );
  CKBD0 U4831 ( .CLK(n4949), .C(n4950) );
  CKBD0 U4832 ( .CLK(n4950), .C(n4951) );
  CKBD0 U4833 ( .CLK(n4951), .C(n4952) );
  CKBD0 U4834 ( .CLK(n4952), .C(n4953) );
  CKBD0 U4835 ( .CLK(n4953), .C(n4954) );
  CKBD0 U4836 ( .CLK(n4954), .C(n4955) );
  CKBD0 U4837 ( .CLK(n4955), .C(n4956) );
  BUFFD0 U4838 ( .I(n4956), .Z(n4957) );
  CKBD0 U4839 ( .CLK(n4957), .C(n4958) );
  CKBD0 U4840 ( .CLK(n4958), .C(n4959) );
  CKBD0 U4841 ( .CLK(n4959), .C(n4960) );
  CKBD0 U4842 ( .CLK(n4960), .C(n4961) );
  CKBD0 U4843 ( .CLK(n4961), .C(n4962) );
  CKBD0 U4844 ( .CLK(n4962), .C(n4963) );
  BUFFD0 U4845 ( .I(n4963), .Z(n4964) );
  CKBD0 U4846 ( .CLK(n4964), .C(n4965) );
  BUFFD0 U4847 ( .I(n4965), .Z(n4966) );
  CKBD0 U4848 ( .CLK(n4966), .C(n4967) );
  BUFFD0 U4849 ( .I(n4967), .Z(n4968) );
  CKBD0 U4850 ( .CLK(n4968), .C(n4969) );
  BUFFD0 U4851 ( .I(n4969), .Z(n4970) );
  CKBD0 U4852 ( .CLK(n4970), .C(n4971) );
  BUFFD0 U4853 ( .I(n4971), .Z(n4972) );
  CKBD0 U4854 ( .CLK(n4972), .C(n4973) );
  BUFFD0 U4855 ( .I(n4973), .Z(n4974) );
  CKBD0 U4856 ( .CLK(n4974), .C(n4975) );
  BUFFD0 U4857 ( .I(n4975), .Z(n4976) );
  CKBD0 U4858 ( .CLK(n4976), .C(n4977) );
  BUFFD0 U4859 ( .I(n4977), .Z(n4978) );
  BUFFD0 U4860 ( .I(n4980), .Z(n4979) );
  BUFFD0 U4861 ( .I(n4981), .Z(n4980) );
  BUFFD0 U4862 ( .I(n146), .Z(n4981) );
  CKBD0 U4863 ( .CLK(n1130), .C(n4982) );
  CKBD0 U4864 ( .CLK(n4982), .C(n4983) );
  CKBD0 U4865 ( .CLK(n4983), .C(n4984) );
  BUFFD0 U4866 ( .I(n4984), .Z(n4985) );
  CKBD0 U4867 ( .CLK(n4985), .C(n4986) );
  CKBD0 U4868 ( .CLK(n4986), .C(n4987) );
  CKBD0 U4869 ( .CLK(n4987), .C(n4988) );
  CKBD0 U4870 ( .CLK(n4988), .C(n4989) );
  CKBD0 U4871 ( .CLK(n4989), .C(n4990) );
  CKBD0 U4872 ( .CLK(n4990), .C(n4991) );
  CKBD0 U4873 ( .CLK(n4991), .C(n4992) );
  CKBD0 U4874 ( .CLK(n4992), .C(n4993) );
  CKBD0 U4875 ( .CLK(n4993), .C(n4994) );
  CKBD0 U4876 ( .CLK(n4994), .C(n4995) );
  BUFFD0 U4877 ( .I(n4995), .Z(n4996) );
  CKBD0 U4878 ( .CLK(n4996), .C(n4997) );
  CKBD0 U4879 ( .CLK(n4997), .C(n4998) );
  CKBD0 U4880 ( .CLK(n4998), .C(n4999) );
  CKBD0 U4881 ( .CLK(n4999), .C(n5000) );
  CKBD0 U4882 ( .CLK(n5000), .C(n5001) );
  CKBD0 U4883 ( .CLK(n5001), .C(n5002) );
  CKBD0 U4884 ( .CLK(n5002), .C(n5003) );
  CKBD0 U4885 ( .CLK(n5003), .C(n5004) );
  CKBD0 U4886 ( .CLK(n5004), .C(n5005) );
  BUFFD0 U4887 ( .I(n5005), .Z(n5006) );
  CKBD0 U4888 ( .CLK(n5006), .C(n5007) );
  CKBD0 U4889 ( .CLK(n5007), .C(n5008) );
  CKBD0 U4890 ( .CLK(n5008), .C(n5009) );
  CKBD0 U4891 ( .CLK(n5009), .C(n5010) );
  CKBD0 U4892 ( .CLK(n5010), .C(n5011) );
  CKBD0 U4893 ( .CLK(n5011), .C(n5012) );
  CKBD0 U4894 ( .CLK(n5012), .C(n5013) );
  CKBD0 U4895 ( .CLK(n5013), .C(n5014) );
  CKBD0 U4896 ( .CLK(n5014), .C(n5015) );
  CKBD0 U4897 ( .CLK(n5015), .C(n5016) );
  BUFFD0 U4898 ( .I(n5016), .Z(n5017) );
  CKBD0 U4899 ( .CLK(n5017), .C(n5018) );
  CKBD0 U4900 ( .CLK(n5018), .C(n5019) );
  CKBD0 U4901 ( .CLK(n5019), .C(n5020) );
  CKBD0 U4902 ( .CLK(n5020), .C(n5021) );
  CKBD0 U4903 ( .CLK(n5021), .C(n5022) );
  CKBD0 U4904 ( .CLK(n5022), .C(n5023) );
  CKBD0 U4905 ( .CLK(n5023), .C(n5024) );
  CKBD0 U4906 ( .CLK(n5024), .C(n5025) );
  CKBD0 U4907 ( .CLK(n5025), .C(n5026) );
  CKBD0 U4908 ( .CLK(n5026), .C(n5027) );
  BUFFD0 U4909 ( .I(n5027), .Z(n5028) );
  CKBD0 U4910 ( .CLK(n5028), .C(n5029) );
  CKBD0 U4911 ( .CLK(n5029), .C(n5030) );
  CKBD0 U4912 ( .CLK(n5030), .C(n5031) );
  CKBD0 U4913 ( .CLK(n5031), .C(n5032) );
  CKBD0 U4914 ( .CLK(n5032), .C(n5033) );
  CKBD0 U4915 ( .CLK(n5033), .C(n5034) );
  CKBD0 U4916 ( .CLK(n5034), .C(n5035) );
  CKBD0 U4917 ( .CLK(n5035), .C(n5036) );
  CKBD0 U4918 ( .CLK(n5036), .C(n5037) );
  CKBD0 U4919 ( .CLK(n5037), .C(n5038) );
  BUFFD0 U4920 ( .I(n5038), .Z(n5039) );
  CKBD0 U4921 ( .CLK(n5039), .C(n5040) );
  CKBD0 U4922 ( .CLK(n5040), .C(n5041) );
  CKBD0 U4923 ( .CLK(n5041), .C(n5042) );
  CKBD0 U4924 ( .CLK(n5042), .C(n5043) );
  CKBD0 U4925 ( .CLK(n5043), .C(n5044) );
  CKBD0 U4926 ( .CLK(n5044), .C(n5045) );
  CKBD0 U4927 ( .CLK(n5045), .C(n5046) );
  CKBD0 U4928 ( .CLK(n5046), .C(n5047) );
  CKBD0 U4929 ( .CLK(n5047), .C(n5048) );
  CKBD0 U4930 ( .CLK(n5048), .C(n5049) );
  BUFFD0 U4931 ( .I(n5049), .Z(n5050) );
  CKBD0 U4932 ( .CLK(n5050), .C(n5051) );
  CKBD0 U4933 ( .CLK(n5051), .C(n5052) );
  CKBD0 U4934 ( .CLK(n5052), .C(n5053) );
  CKBD0 U4935 ( .CLK(n5053), .C(n5054) );
  CKBD0 U4936 ( .CLK(n5054), .C(n5055) );
  CKBD0 U4937 ( .CLK(n5055), .C(n5056) );
  CKBD0 U4938 ( .CLK(n5056), .C(n5057) );
  CKBD0 U4939 ( .CLK(n5057), .C(n5058) );
  CKBD0 U4940 ( .CLK(n5058), .C(n5059) );
  CKBD0 U4941 ( .CLK(n5059), .C(n5060) );
  BUFFD0 U4942 ( .I(n5060), .Z(n5061) );
  CKBD0 U4943 ( .CLK(n5061), .C(n5062) );
  CKBD0 U4944 ( .CLK(n5062), .C(n5063) );
  CKBD0 U4945 ( .CLK(n5063), .C(n5064) );
  CKBD0 U4946 ( .CLK(n5064), .C(n5065) );
  CKBD0 U4947 ( .CLK(n5065), .C(n5066) );
  CKBD0 U4948 ( .CLK(n5066), .C(n5067) );
  CKBD0 U4949 ( .CLK(n5067), .C(n5068) );
  CKBD0 U4950 ( .CLK(n5068), .C(n5069) );
  CKBD0 U4951 ( .CLK(n5069), .C(n5070) );
  BUFFD0 U4952 ( .I(n5070), .Z(n5071) );
  CKBD0 U4953 ( .CLK(n5071), .C(n5072) );
  CKBD0 U4954 ( .CLK(n5072), .C(n5073) );
  CKBD0 U4955 ( .CLK(n5073), .C(n5074) );
  CKBD0 U4956 ( .CLK(n5074), .C(n5075) );
  CKBD0 U4957 ( .CLK(n5075), .C(n5076) );
  CKBD0 U4958 ( .CLK(n5076), .C(n5077) );
  CKBD0 U4959 ( .CLK(n5077), .C(n5078) );
  CKBD0 U4960 ( .CLK(n5078), .C(n5079) );
  CKBD0 U4961 ( .CLK(n5079), .C(n5080) );
  CKBD0 U4962 ( .CLK(n5080), .C(n5081) );
  BUFFD0 U4963 ( .I(n5081), .Z(n5082) );
  CKBD0 U4964 ( .CLK(n5082), .C(n5083) );
  CKBD0 U4965 ( .CLK(n5083), .C(n5084) );
  CKBD0 U4966 ( .CLK(n5084), .C(n5085) );
  CKBD0 U4967 ( .CLK(n5085), .C(n5086) );
  CKBD0 U4968 ( .CLK(n5086), .C(n5087) );
  CKBD0 U4969 ( .CLK(n5087), .C(n5088) );
  CKBD0 U4970 ( .CLK(n5088), .C(n5089) );
  CKBD0 U4971 ( .CLK(n5089), .C(n5090) );
  CKBD0 U4972 ( .CLK(n5090), .C(n5091) );
  CKBD0 U4973 ( .CLK(n5091), .C(n5092) );
  BUFFD0 U4974 ( .I(n5092), .Z(n5093) );
  CKBD0 U4975 ( .CLK(n5093), .C(n5094) );
  CKBD0 U4976 ( .CLK(n5094), .C(n5095) );
  CKBD0 U4977 ( .CLK(n5095), .C(n5096) );
  CKBD0 U4978 ( .CLK(n5096), .C(n5097) );
  CKBD0 U4979 ( .CLK(n5097), .C(n5098) );
  CKBD0 U4980 ( .CLK(n5098), .C(n5099) );
  BUFFD0 U4981 ( .I(n5099), .Z(n5100) );
  CKBD0 U4982 ( .CLK(n5100), .C(n5101) );
  BUFFD0 U4983 ( .I(n5101), .Z(n5102) );
  CKBD0 U4984 ( .CLK(n5102), .C(n5103) );
  BUFFD0 U4985 ( .I(n5103), .Z(n5104) );
  CKBD0 U4986 ( .CLK(n5104), .C(n5105) );
  BUFFD0 U4987 ( .I(n5105), .Z(n5106) );
  CKBD0 U4988 ( .CLK(n5106), .C(n5107) );
  BUFFD0 U4989 ( .I(n5107), .Z(n5108) );
  CKBD0 U4990 ( .CLK(n5108), .C(n5109) );
  BUFFD0 U4991 ( .I(n5109), .Z(n5110) );
  CKBD0 U4992 ( .CLK(n5110), .C(n5111) );
  BUFFD0 U4993 ( .I(n5111), .Z(n5112) );
  CKBD0 U4994 ( .CLK(n5112), .C(n5113) );
  BUFFD0 U4995 ( .I(n5113), .Z(n5114) );
  BUFFD0 U4996 ( .I(n5116), .Z(n5115) );
  BUFFD0 U4997 ( .I(n5117), .Z(n5116) );
  BUFFD0 U4998 ( .I(n145), .Z(n5117) );
  CKBD0 U4999 ( .CLK(n1128), .C(n5118) );
  CKBD0 U5000 ( .CLK(n5118), .C(n5119) );
  CKBD0 U5001 ( .CLK(n5119), .C(n5120) );
  BUFFD0 U5002 ( .I(n5120), .Z(n5121) );
  CKBD0 U5003 ( .CLK(n5121), .C(n5122) );
  CKBD0 U5004 ( .CLK(n5122), .C(n5123) );
  CKBD0 U5005 ( .CLK(n5123), .C(n5124) );
  CKBD0 U5006 ( .CLK(n5124), .C(n5125) );
  CKBD0 U5007 ( .CLK(n5125), .C(n5126) );
  CKBD0 U5008 ( .CLK(n5126), .C(n5127) );
  CKBD0 U5009 ( .CLK(n5127), .C(n5128) );
  CKBD0 U5010 ( .CLK(n5128), .C(n5129) );
  CKBD0 U5011 ( .CLK(n5129), .C(n5130) );
  BUFFD0 U5012 ( .I(n5130), .Z(n5131) );
  CKBD0 U5013 ( .CLK(n5131), .C(n5132) );
  CKBD0 U5014 ( .CLK(n5132), .C(n5133) );
  CKBD0 U5015 ( .CLK(n5133), .C(n5134) );
  CKBD0 U5016 ( .CLK(n5134), .C(n5135) );
  CKBD0 U5017 ( .CLK(n5135), .C(n5136) );
  CKBD0 U5018 ( .CLK(n5136), .C(n5137) );
  CKBD0 U5019 ( .CLK(n5137), .C(n5138) );
  CKBD0 U5020 ( .CLK(n5138), .C(n5139) );
  CKBD0 U5021 ( .CLK(n5139), .C(n5140) );
  CKBD0 U5022 ( .CLK(n5140), .C(n5141) );
  BUFFD0 U5023 ( .I(n5141), .Z(n5142) );
  CKBD0 U5024 ( .CLK(n5142), .C(n5143) );
  CKBD0 U5025 ( .CLK(n5143), .C(n5144) );
  CKBD0 U5026 ( .CLK(n5144), .C(n5145) );
  CKBD0 U5027 ( .CLK(n5145), .C(n5146) );
  CKBD0 U5028 ( .CLK(n5146), .C(n5147) );
  CKBD0 U5029 ( .CLK(n5147), .C(n5148) );
  CKBD0 U5030 ( .CLK(n5148), .C(n5149) );
  CKBD0 U5031 ( .CLK(n5149), .C(n5150) );
  CKBD0 U5032 ( .CLK(n5150), .C(n5151) );
  CKBD0 U5033 ( .CLK(n5151), .C(n5152) );
  BUFFD0 U5034 ( .I(n5152), .Z(n5153) );
  CKBD0 U5035 ( .CLK(n5153), .C(n5154) );
  CKBD0 U5036 ( .CLK(n5154), .C(n5155) );
  CKBD0 U5037 ( .CLK(n5155), .C(n5156) );
  CKBD0 U5038 ( .CLK(n5156), .C(n5157) );
  CKBD0 U5039 ( .CLK(n5157), .C(n5158) );
  CKBD0 U5040 ( .CLK(n5158), .C(n5159) );
  CKBD0 U5041 ( .CLK(n5159), .C(n5160) );
  CKBD0 U5042 ( .CLK(n5160), .C(n5161) );
  CKBD0 U5043 ( .CLK(n5161), .C(n5162) );
  CKBD0 U5044 ( .CLK(n5162), .C(n5163) );
  BUFFD0 U5045 ( .I(n5163), .Z(n5164) );
  CKBD0 U5046 ( .CLK(n5164), .C(n5165) );
  CKBD0 U5047 ( .CLK(n5165), .C(n5166) );
  CKBD0 U5048 ( .CLK(n5166), .C(n5167) );
  CKBD0 U5049 ( .CLK(n5167), .C(n5168) );
  CKBD0 U5050 ( .CLK(n5168), .C(n5169) );
  CKBD0 U5051 ( .CLK(n5169), .C(n5170) );
  CKBD0 U5052 ( .CLK(n5170), .C(n5171) );
  CKBD0 U5053 ( .CLK(n5171), .C(n5172) );
  CKBD0 U5054 ( .CLK(n5172), .C(n5173) );
  CKBD0 U5055 ( .CLK(n5173), .C(n5174) );
  BUFFD0 U5056 ( .I(n5174), .Z(n5175) );
  CKBD0 U5057 ( .CLK(n5175), .C(n5176) );
  CKBD0 U5058 ( .CLK(n5176), .C(n5177) );
  CKBD0 U5059 ( .CLK(n5177), .C(n5178) );
  CKBD0 U5060 ( .CLK(n5178), .C(n5179) );
  CKBD0 U5061 ( .CLK(n5179), .C(n5180) );
  CKBD0 U5062 ( .CLK(n5180), .C(n5181) );
  CKBD0 U5063 ( .CLK(n5181), .C(n5182) );
  CKBD0 U5064 ( .CLK(n5182), .C(n5183) );
  CKBD0 U5065 ( .CLK(n5183), .C(n5184) );
  CKBD0 U5066 ( .CLK(n5184), .C(n5185) );
  BUFFD0 U5067 ( .I(n5185), .Z(n5186) );
  CKBD0 U5068 ( .CLK(n5186), .C(n5187) );
  CKBD0 U5069 ( .CLK(n5187), .C(n5188) );
  CKBD0 U5070 ( .CLK(n5188), .C(n5189) );
  CKBD0 U5071 ( .CLK(n5189), .C(n5190) );
  CKBD0 U5072 ( .CLK(n5190), .C(n5191) );
  CKBD0 U5073 ( .CLK(n5191), .C(n5192) );
  CKBD0 U5074 ( .CLK(n5192), .C(n5193) );
  CKBD0 U5075 ( .CLK(n5193), .C(n5194) );
  CKBD0 U5076 ( .CLK(n5194), .C(n5195) );
  CKBD0 U5077 ( .CLK(n5195), .C(n5196) );
  BUFFD0 U5078 ( .I(n5196), .Z(n5197) );
  CKBD0 U5079 ( .CLK(n5197), .C(n5198) );
  CKBD0 U5080 ( .CLK(n5198), .C(n5199) );
  CKBD0 U5081 ( .CLK(n5199), .C(n5200) );
  CKBD0 U5082 ( .CLK(n5200), .C(n5201) );
  CKBD0 U5083 ( .CLK(n5201), .C(n5202) );
  CKBD0 U5084 ( .CLK(n5202), .C(n5203) );
  CKBD0 U5085 ( .CLK(n5203), .C(n5204) );
  CKBD0 U5086 ( .CLK(n5204), .C(n5205) );
  CKBD0 U5087 ( .CLK(n5205), .C(n5206) );
  BUFFD0 U5088 ( .I(n5206), .Z(n5207) );
  CKBD0 U5089 ( .CLK(n5207), .C(n5208) );
  CKBD0 U5090 ( .CLK(n5208), .C(n5209) );
  CKBD0 U5091 ( .CLK(n5209), .C(n5210) );
  CKBD0 U5092 ( .CLK(n5210), .C(n5211) );
  CKBD0 U5093 ( .CLK(n5211), .C(n5212) );
  CKBD0 U5094 ( .CLK(n5212), .C(n5213) );
  CKBD0 U5095 ( .CLK(n5213), .C(n5214) );
  CKBD0 U5096 ( .CLK(n5214), .C(n5215) );
  CKBD0 U5097 ( .CLK(n5215), .C(n5216) );
  CKBD0 U5098 ( .CLK(n5216), .C(n5217) );
  BUFFD0 U5099 ( .I(n5217), .Z(n5218) );
  CKBD0 U5100 ( .CLK(n5218), .C(n5219) );
  CKBD0 U5101 ( .CLK(n5219), .C(n5220) );
  CKBD0 U5102 ( .CLK(n5220), .C(n5221) );
  CKBD0 U5103 ( .CLK(n5221), .C(n5222) );
  CKBD0 U5104 ( .CLK(n5222), .C(n5223) );
  CKBD0 U5105 ( .CLK(n5223), .C(n5224) );
  CKBD0 U5106 ( .CLK(n5224), .C(n5225) );
  CKBD0 U5107 ( .CLK(n5225), .C(n5226) );
  CKBD0 U5108 ( .CLK(n5226), .C(n5227) );
  CKBD0 U5109 ( .CLK(n5227), .C(n5228) );
  BUFFD0 U5110 ( .I(n5228), .Z(n5229) );
  CKBD0 U5111 ( .CLK(n5229), .C(n5230) );
  CKBD0 U5112 ( .CLK(n5230), .C(n5231) );
  CKBD0 U5113 ( .CLK(n5231), .C(n5232) );
  CKBD0 U5114 ( .CLK(n5232), .C(n5233) );
  CKBD0 U5115 ( .CLK(n5233), .C(n5234) );
  CKBD0 U5116 ( .CLK(n5234), .C(n5235) );
  BUFFD0 U5117 ( .I(n5235), .Z(n5236) );
  CKBD0 U5118 ( .CLK(n5236), .C(n5237) );
  BUFFD0 U5119 ( .I(n5237), .Z(n5238) );
  CKBD0 U5120 ( .CLK(n5238), .C(n5239) );
  BUFFD0 U5121 ( .I(n5239), .Z(n5240) );
  CKBD0 U5122 ( .CLK(n5240), .C(n5241) );
  BUFFD0 U5123 ( .I(n5241), .Z(n5242) );
  CKBD0 U5124 ( .CLK(n5242), .C(n5243) );
  BUFFD0 U5125 ( .I(n5243), .Z(n5244) );
  CKBD0 U5126 ( .CLK(n5244), .C(n5245) );
  BUFFD0 U5127 ( .I(n5245), .Z(n5246) );
  CKBD0 U5128 ( .CLK(n5246), .C(n5247) );
  BUFFD0 U5129 ( .I(n5247), .Z(n5248) );
  CKBD0 U5130 ( .CLK(n5248), .C(n5249) );
  BUFFD0 U5131 ( .I(n5249), .Z(n5250) );
  BUFFD0 U5132 ( .I(n5252), .Z(n5251) );
  BUFFD0 U5133 ( .I(n5253), .Z(n5252) );
  BUFFD0 U5134 ( .I(n144), .Z(n5253) );
  CKBD0 U5135 ( .CLK(n1126), .C(n5254) );
  CKBD0 U5136 ( .CLK(n5254), .C(n5255) );
  CKBD0 U5137 ( .CLK(n5255), .C(n5256) );
  BUFFD0 U5138 ( .I(n5256), .Z(n5257) );
  CKBD0 U5139 ( .CLK(n5257), .C(n5258) );
  CKBD0 U5140 ( .CLK(n5258), .C(n5259) );
  CKBD0 U5141 ( .CLK(n5259), .C(n5260) );
  CKBD0 U5142 ( .CLK(n5260), .C(n5261) );
  CKBD0 U5143 ( .CLK(n5261), .C(n5262) );
  CKBD0 U5144 ( .CLK(n5262), .C(n5263) );
  CKBD0 U5145 ( .CLK(n5263), .C(n5264) );
  CKBD0 U5146 ( .CLK(n5264), .C(n5265) );
  CKBD0 U5147 ( .CLK(n5265), .C(n5266) );
  BUFFD0 U5148 ( .I(n5266), .Z(n5267) );
  CKBD0 U5149 ( .CLK(n5267), .C(n5268) );
  CKBD0 U5150 ( .CLK(n5268), .C(n5269) );
  CKBD0 U5151 ( .CLK(n5269), .C(n5270) );
  CKBD0 U5152 ( .CLK(n5270), .C(n5271) );
  CKBD0 U5153 ( .CLK(n5271), .C(n5272) );
  CKBD0 U5154 ( .CLK(n5272), .C(n5273) );
  CKBD0 U5155 ( .CLK(n5273), .C(n5274) );
  CKBD0 U5156 ( .CLK(n5274), .C(n5275) );
  CKBD0 U5157 ( .CLK(n5275), .C(n5276) );
  CKBD0 U5158 ( .CLK(n5276), .C(n5277) );
  BUFFD0 U5159 ( .I(n5277), .Z(n5278) );
  CKBD0 U5160 ( .CLK(n5278), .C(n5279) );
  CKBD0 U5161 ( .CLK(n5279), .C(n5280) );
  CKBD0 U5162 ( .CLK(n5280), .C(n5281) );
  CKBD0 U5163 ( .CLK(n5281), .C(n5282) );
  CKBD0 U5164 ( .CLK(n5282), .C(n5283) );
  CKBD0 U5165 ( .CLK(n5283), .C(n5284) );
  CKBD0 U5166 ( .CLK(n5284), .C(n5285) );
  CKBD0 U5167 ( .CLK(n5285), .C(n5286) );
  CKBD0 U5168 ( .CLK(n5286), .C(n5287) );
  CKBD0 U5169 ( .CLK(n5287), .C(n5288) );
  BUFFD0 U5170 ( .I(n5288), .Z(n5289) );
  CKBD0 U5171 ( .CLK(n5289), .C(n5290) );
  CKBD0 U5172 ( .CLK(n5290), .C(n5291) );
  CKBD0 U5173 ( .CLK(n5291), .C(n5292) );
  CKBD0 U5174 ( .CLK(n5292), .C(n5293) );
  CKBD0 U5175 ( .CLK(n5293), .C(n5294) );
  CKBD0 U5176 ( .CLK(n5294), .C(n5295) );
  CKBD0 U5177 ( .CLK(n5295), .C(n5296) );
  CKBD0 U5178 ( .CLK(n5296), .C(n5297) );
  CKBD0 U5179 ( .CLK(n5297), .C(n5298) );
  CKBD0 U5180 ( .CLK(n5298), .C(n5299) );
  BUFFD0 U5181 ( .I(n5299), .Z(n5300) );
  CKBD0 U5182 ( .CLK(n5300), .C(n5301) );
  CKBD0 U5183 ( .CLK(n5301), .C(n5302) );
  CKBD0 U5184 ( .CLK(n5302), .C(n5303) );
  CKBD0 U5185 ( .CLK(n5303), .C(n5304) );
  CKBD0 U5186 ( .CLK(n5304), .C(n5305) );
  CKBD0 U5187 ( .CLK(n5305), .C(n5306) );
  CKBD0 U5188 ( .CLK(n5306), .C(n5307) );
  CKBD0 U5189 ( .CLK(n5307), .C(n5308) );
  CKBD0 U5190 ( .CLK(n5308), .C(n5309) );
  CKBD0 U5191 ( .CLK(n5309), .C(n5310) );
  BUFFD0 U5192 ( .I(n5310), .Z(n5311) );
  CKBD0 U5193 ( .CLK(n5311), .C(n5312) );
  CKBD0 U5194 ( .CLK(n5312), .C(n5313) );
  CKBD0 U5195 ( .CLK(n5313), .C(n5314) );
  CKBD0 U5196 ( .CLK(n5314), .C(n5315) );
  CKBD0 U5197 ( .CLK(n5315), .C(n5316) );
  CKBD0 U5198 ( .CLK(n5316), .C(n5317) );
  CKBD0 U5199 ( .CLK(n5317), .C(n5318) );
  CKBD0 U5200 ( .CLK(n5318), .C(n5319) );
  CKBD0 U5201 ( .CLK(n5319), .C(n5320) );
  CKBD0 U5202 ( .CLK(n5320), .C(n5321) );
  BUFFD0 U5203 ( .I(n5321), .Z(n5322) );
  CKBD0 U5204 ( .CLK(n5322), .C(n5323) );
  CKBD0 U5205 ( .CLK(n5323), .C(n5324) );
  CKBD0 U5206 ( .CLK(n5324), .C(n5325) );
  CKBD0 U5207 ( .CLK(n5325), .C(n5326) );
  CKBD0 U5208 ( .CLK(n5326), .C(n5327) );
  CKBD0 U5209 ( .CLK(n5327), .C(n5328) );
  CKBD0 U5210 ( .CLK(n5328), .C(n5329) );
  CKBD0 U5211 ( .CLK(n5329), .C(n5330) );
  CKBD0 U5212 ( .CLK(n5330), .C(n5331) );
  CKBD0 U5213 ( .CLK(n5331), .C(n5332) );
  BUFFD0 U5214 ( .I(n5332), .Z(n5333) );
  CKBD0 U5215 ( .CLK(n5333), .C(n5334) );
  CKBD0 U5216 ( .CLK(n5334), .C(n5335) );
  CKBD0 U5217 ( .CLK(n5335), .C(n5336) );
  CKBD0 U5218 ( .CLK(n5336), .C(n5337) );
  CKBD0 U5219 ( .CLK(n5337), .C(n5338) );
  CKBD0 U5220 ( .CLK(n5338), .C(n5339) );
  CKBD0 U5221 ( .CLK(n5339), .C(n5340) );
  CKBD0 U5222 ( .CLK(n5340), .C(n5341) );
  CKBD0 U5223 ( .CLK(n5341), .C(n5342) );
  BUFFD0 U5224 ( .I(n5342), .Z(n5343) );
  CKBD0 U5225 ( .CLK(n5343), .C(n5344) );
  CKBD0 U5226 ( .CLK(n5344), .C(n5345) );
  CKBD0 U5227 ( .CLK(n5345), .C(n5346) );
  CKBD0 U5228 ( .CLK(n5346), .C(n5347) );
  CKBD0 U5229 ( .CLK(n5347), .C(n5348) );
  CKBD0 U5230 ( .CLK(n5348), .C(n5349) );
  CKBD0 U5231 ( .CLK(n5349), .C(n5350) );
  CKBD0 U5232 ( .CLK(n5350), .C(n5351) );
  CKBD0 U5233 ( .CLK(n5351), .C(n5352) );
  CKBD0 U5234 ( .CLK(n5352), .C(n5353) );
  BUFFD0 U5235 ( .I(n5353), .Z(n5354) );
  CKBD0 U5236 ( .CLK(n5354), .C(n5355) );
  CKBD0 U5237 ( .CLK(n5355), .C(n5356) );
  CKBD0 U5238 ( .CLK(n5356), .C(n5357) );
  CKBD0 U5239 ( .CLK(n5357), .C(n5358) );
  CKBD0 U5240 ( .CLK(n5358), .C(n5359) );
  CKBD0 U5241 ( .CLK(n5359), .C(n5360) );
  CKBD0 U5242 ( .CLK(n5360), .C(n5361) );
  CKBD0 U5243 ( .CLK(n5361), .C(n5362) );
  CKBD0 U5244 ( .CLK(n5362), .C(n5363) );
  CKBD0 U5245 ( .CLK(n5363), .C(n5364) );
  BUFFD0 U5246 ( .I(n5364), .Z(n5365) );
  CKBD0 U5247 ( .CLK(n5365), .C(n5366) );
  CKBD0 U5248 ( .CLK(n5366), .C(n5367) );
  CKBD0 U5249 ( .CLK(n5367), .C(n5368) );
  CKBD0 U5250 ( .CLK(n5368), .C(n5369) );
  CKBD0 U5251 ( .CLK(n5369), .C(n5370) );
  CKBD0 U5252 ( .CLK(n5370), .C(n5371) );
  BUFFD0 U5253 ( .I(n5371), .Z(n5372) );
  CKBD0 U5254 ( .CLK(n5372), .C(n5373) );
  BUFFD0 U5255 ( .I(n5373), .Z(n5374) );
  CKBD0 U5256 ( .CLK(n5374), .C(n5375) );
  BUFFD0 U5257 ( .I(n5375), .Z(n5376) );
  CKBD0 U5258 ( .CLK(n5376), .C(n5377) );
  BUFFD0 U5259 ( .I(n5377), .Z(n5378) );
  CKBD0 U5260 ( .CLK(n5378), .C(n5379) );
  BUFFD0 U5261 ( .I(n5379), .Z(n5380) );
  CKBD0 U5262 ( .CLK(n5380), .C(n5381) );
  BUFFD0 U5263 ( .I(n5381), .Z(n5382) );
  CKBD0 U5264 ( .CLK(n5382), .C(n5383) );
  BUFFD0 U5265 ( .I(n5383), .Z(n5384) );
  CKBD0 U5266 ( .CLK(n5384), .C(n5385) );
  BUFFD0 U5267 ( .I(n5385), .Z(n5386) );
  BUFFD0 U5268 ( .I(n5388), .Z(n5387) );
  BUFFD0 U5269 ( .I(n5389), .Z(n5388) );
  BUFFD0 U5270 ( .I(n143), .Z(n5389) );
  CKBD0 U5271 ( .CLK(n1124), .C(n5390) );
  CKBD0 U5272 ( .CLK(n5390), .C(n5391) );
  CKBD0 U5273 ( .CLK(n5391), .C(n5392) );
  BUFFD0 U5274 ( .I(n5392), .Z(n5393) );
  CKBD0 U5275 ( .CLK(n5393), .C(n5394) );
  CKBD0 U5276 ( .CLK(n5394), .C(n5395) );
  CKBD0 U5277 ( .CLK(n5395), .C(n5396) );
  CKBD0 U5278 ( .CLK(n5396), .C(n5397) );
  CKBD0 U5279 ( .CLK(n5397), .C(n5398) );
  CKBD0 U5280 ( .CLK(n5398), .C(n5399) );
  CKBD0 U5281 ( .CLK(n5399), .C(n5400) );
  CKBD0 U5282 ( .CLK(n5400), .C(n5401) );
  CKBD0 U5283 ( .CLK(n5401), .C(n5402) );
  CKBD0 U5284 ( .CLK(n5402), .C(n5403) );
  BUFFD0 U5285 ( .I(n5403), .Z(n5404) );
  CKBD0 U5286 ( .CLK(n5404), .C(n5405) );
  CKBD0 U5287 ( .CLK(n5405), .C(n5406) );
  CKBD0 U5288 ( .CLK(n5406), .C(n5407) );
  CKBD0 U5289 ( .CLK(n5407), .C(n5408) );
  CKBD0 U5290 ( .CLK(n5408), .C(n5409) );
  CKBD0 U5291 ( .CLK(n5409), .C(n5410) );
  CKBD0 U5292 ( .CLK(n5410), .C(n5411) );
  CKBD0 U5293 ( .CLK(n5411), .C(n5412) );
  CKBD0 U5294 ( .CLK(n5412), .C(n5413) );
  BUFFD0 U5295 ( .I(n5413), .Z(n5414) );
  CKBD0 U5296 ( .CLK(n5414), .C(n5415) );
  CKBD0 U5297 ( .CLK(n5415), .C(n5416) );
  CKBD0 U5298 ( .CLK(n5416), .C(n5417) );
  CKBD0 U5299 ( .CLK(n5417), .C(n5418) );
  CKBD0 U5300 ( .CLK(n5418), .C(n5419) );
  CKBD0 U5301 ( .CLK(n5419), .C(n5420) );
  CKBD0 U5302 ( .CLK(n5420), .C(n5421) );
  CKBD0 U5303 ( .CLK(n5421), .C(n5422) );
  CKBD0 U5304 ( .CLK(n5422), .C(n5423) );
  CKBD0 U5305 ( .CLK(n5423), .C(n5424) );
  BUFFD0 U5306 ( .I(n5424), .Z(n5425) );
  CKBD0 U5307 ( .CLK(n5425), .C(n5426) );
  CKBD0 U5308 ( .CLK(n5426), .C(n5427) );
  CKBD0 U5309 ( .CLK(n5427), .C(n5428) );
  CKBD0 U5310 ( .CLK(n5428), .C(n5429) );
  CKBD0 U5311 ( .CLK(n5429), .C(n5430) );
  CKBD0 U5312 ( .CLK(n5430), .C(n5431) );
  CKBD0 U5313 ( .CLK(n5431), .C(n5432) );
  CKBD0 U5314 ( .CLK(n5432), .C(n5433) );
  CKBD0 U5315 ( .CLK(n5433), .C(n5434) );
  CKBD0 U5316 ( .CLK(n5434), .C(n5435) );
  BUFFD0 U5317 ( .I(n5435), .Z(n5436) );
  CKBD0 U5318 ( .CLK(n5436), .C(n5437) );
  CKBD0 U5319 ( .CLK(n5437), .C(n5438) );
  CKBD0 U5320 ( .CLK(n5438), .C(n5439) );
  CKBD0 U5321 ( .CLK(n5439), .C(n5440) );
  CKBD0 U5322 ( .CLK(n5440), .C(n5441) );
  CKBD0 U5323 ( .CLK(n5441), .C(n5442) );
  CKBD0 U5324 ( .CLK(n5442), .C(n5443) );
  CKBD0 U5325 ( .CLK(n5443), .C(n5444) );
  CKBD0 U5326 ( .CLK(n5444), .C(n5445) );
  CKBD0 U5327 ( .CLK(n5445), .C(n5446) );
  BUFFD0 U5328 ( .I(n5446), .Z(n5447) );
  CKBD0 U5329 ( .CLK(n5447), .C(n5448) );
  CKBD0 U5330 ( .CLK(n5448), .C(n5449) );
  CKBD0 U5331 ( .CLK(n5449), .C(n5450) );
  CKBD0 U5332 ( .CLK(n5450), .C(n5451) );
  CKBD0 U5333 ( .CLK(n5451), .C(n5452) );
  CKBD0 U5334 ( .CLK(n5452), .C(n5453) );
  CKBD0 U5335 ( .CLK(n5453), .C(n5454) );
  CKBD0 U5336 ( .CLK(n5454), .C(n5455) );
  CKBD0 U5337 ( .CLK(n5455), .C(n5456) );
  CKBD0 U5338 ( .CLK(n5456), .C(n5457) );
  BUFFD0 U5339 ( .I(n5457), .Z(n5458) );
  CKBD0 U5340 ( .CLK(n5458), .C(n5459) );
  CKBD0 U5341 ( .CLK(n5459), .C(n5460) );
  CKBD0 U5342 ( .CLK(n5460), .C(n5461) );
  CKBD0 U5343 ( .CLK(n5461), .C(n5462) );
  CKBD0 U5344 ( .CLK(n5462), .C(n5463) );
  CKBD0 U5345 ( .CLK(n5463), .C(n5464) );
  CKBD0 U5346 ( .CLK(n5464), .C(n5465) );
  CKBD0 U5347 ( .CLK(n5465), .C(n5466) );
  CKBD0 U5348 ( .CLK(n5466), .C(n5467) );
  CKBD0 U5349 ( .CLK(n5467), .C(n5468) );
  BUFFD0 U5350 ( .I(n5468), .Z(n5469) );
  CKBD0 U5351 ( .CLK(n5469), .C(n5470) );
  CKBD0 U5352 ( .CLK(n5470), .C(n5471) );
  CKBD0 U5353 ( .CLK(n5471), .C(n5472) );
  CKBD0 U5354 ( .CLK(n5472), .C(n5473) );
  CKBD0 U5355 ( .CLK(n5473), .C(n5474) );
  CKBD0 U5356 ( .CLK(n5474), .C(n5475) );
  CKBD0 U5357 ( .CLK(n5475), .C(n5476) );
  CKBD0 U5358 ( .CLK(n5476), .C(n5477) );
  CKBD0 U5359 ( .CLK(n5477), .C(n5478) );
  BUFFD0 U5360 ( .I(n5478), .Z(n5479) );
  CKBD0 U5361 ( .CLK(n5479), .C(n5480) );
  CKBD0 U5362 ( .CLK(n5480), .C(n5481) );
  CKBD0 U5363 ( .CLK(n5481), .C(n5482) );
  CKBD0 U5364 ( .CLK(n5482), .C(n5483) );
  CKBD0 U5365 ( .CLK(n5483), .C(n5484) );
  CKBD0 U5366 ( .CLK(n5484), .C(n5485) );
  CKBD0 U5367 ( .CLK(n5485), .C(n5486) );
  CKBD0 U5368 ( .CLK(n5486), .C(n5487) );
  CKBD0 U5369 ( .CLK(n5487), .C(n5488) );
  CKBD0 U5370 ( .CLK(n5488), .C(n5489) );
  BUFFD0 U5371 ( .I(n5489), .Z(n5490) );
  CKBD0 U5372 ( .CLK(n5490), .C(n5491) );
  CKBD0 U5373 ( .CLK(n5491), .C(n5492) );
  CKBD0 U5374 ( .CLK(n5492), .C(n5493) );
  CKBD0 U5375 ( .CLK(n5493), .C(n5494) );
  CKBD0 U5376 ( .CLK(n5494), .C(n5495) );
  CKBD0 U5377 ( .CLK(n5495), .C(n5496) );
  CKBD0 U5378 ( .CLK(n5496), .C(n5497) );
  CKBD0 U5379 ( .CLK(n5497), .C(n5498) );
  CKBD0 U5380 ( .CLK(n5498), .C(n5499) );
  CKBD0 U5381 ( .CLK(n5499), .C(n5500) );
  BUFFD0 U5382 ( .I(n5500), .Z(n5501) );
  CKBD0 U5383 ( .CLK(n5501), .C(n5502) );
  CKBD0 U5384 ( .CLK(n5502), .C(n5503) );
  CKBD0 U5385 ( .CLK(n5503), .C(n5504) );
  CKBD0 U5386 ( .CLK(n5504), .C(n5505) );
  CKBD0 U5387 ( .CLK(n5505), .C(n5506) );
  CKBD0 U5388 ( .CLK(n5506), .C(n5507) );
  BUFFD0 U5389 ( .I(n5507), .Z(n5508) );
  CKBD0 U5390 ( .CLK(n5508), .C(n5509) );
  BUFFD0 U5391 ( .I(n5509), .Z(n5510) );
  CKBD0 U5392 ( .CLK(n5510), .C(n5511) );
  BUFFD0 U5393 ( .I(n5511), .Z(n5512) );
  CKBD0 U5394 ( .CLK(n5512), .C(n5513) );
  BUFFD0 U5395 ( .I(n5513), .Z(n5514) );
  CKBD0 U5396 ( .CLK(n5514), .C(n5515) );
  BUFFD0 U5397 ( .I(n5515), .Z(n5516) );
  CKBD0 U5398 ( .CLK(n5516), .C(n5517) );
  BUFFD0 U5399 ( .I(n5517), .Z(n5518) );
  CKBD0 U5400 ( .CLK(n5518), .C(n5519) );
  BUFFD0 U5401 ( .I(n5519), .Z(n5520) );
  CKBD0 U5402 ( .CLK(n5520), .C(n5521) );
  BUFFD0 U5403 ( .I(n5521), .Z(n5522) );
  BUFFD0 U5404 ( .I(Decoder[9]), .Z(n5523) );
  BUFFD0 U5405 ( .I(n5525), .Z(n5524) );
  BUFFD0 U5406 ( .I(n5526), .Z(n5525) );
  BUFFD0 U5407 ( .I(n142), .Z(n5526) );
  CKBD0 U5408 ( .CLK(n1122), .C(n5527) );
  CKBD0 U5409 ( .CLK(n5527), .C(n5528) );
  CKBD0 U5410 ( .CLK(n5528), .C(n5529) );
  BUFFD0 U5411 ( .I(n5529), .Z(n5530) );
  CKBD0 U5412 ( .CLK(n5530), .C(n5531) );
  CKBD0 U5413 ( .CLK(n5531), .C(n5532) );
  CKBD0 U5414 ( .CLK(n5532), .C(n5533) );
  CKBD0 U5415 ( .CLK(n5533), .C(n5534) );
  CKBD0 U5416 ( .CLK(n5534), .C(n5535) );
  CKBD0 U5417 ( .CLK(n5535), .C(n5536) );
  CKBD0 U5418 ( .CLK(n5536), .C(n5537) );
  CKBD0 U5419 ( .CLK(n5537), .C(n5538) );
  CKBD0 U5420 ( .CLK(n5538), .C(n5539) );
  CKBD0 U5421 ( .CLK(n5539), .C(n5540) );
  BUFFD0 U5422 ( .I(n5540), .Z(n5541) );
  CKBD0 U5423 ( .CLK(n5541), .C(n5542) );
  CKBD0 U5424 ( .CLK(n5542), .C(n5543) );
  CKBD0 U5425 ( .CLK(n5543), .C(n5544) );
  CKBD0 U5426 ( .CLK(n5544), .C(n5545) );
  CKBD0 U5427 ( .CLK(n5545), .C(n5546) );
  CKBD0 U5428 ( .CLK(n5546), .C(n5547) );
  CKBD0 U5429 ( .CLK(n5547), .C(n5548) );
  CKBD0 U5430 ( .CLK(n5548), .C(n5549) );
  CKBD0 U5431 ( .CLK(n5549), .C(n5550) );
  BUFFD0 U5432 ( .I(n5550), .Z(n5551) );
  CKBD0 U5433 ( .CLK(n5551), .C(n5552) );
  CKBD0 U5434 ( .CLK(n5552), .C(n5553) );
  CKBD0 U5435 ( .CLK(n5553), .C(n5554) );
  CKBD0 U5436 ( .CLK(n5554), .C(n5555) );
  CKBD0 U5437 ( .CLK(n5555), .C(n5556) );
  CKBD0 U5438 ( .CLK(n5556), .C(n5557) );
  CKBD0 U5439 ( .CLK(n5557), .C(n5558) );
  CKBD0 U5440 ( .CLK(n5558), .C(n5559) );
  CKBD0 U5441 ( .CLK(n5559), .C(n5560) );
  CKBD0 U5442 ( .CLK(n5560), .C(n5561) );
  BUFFD0 U5443 ( .I(n5561), .Z(n5562) );
  CKBD0 U5444 ( .CLK(n5562), .C(n5563) );
  CKBD0 U5445 ( .CLK(n5563), .C(n5564) );
  CKBD0 U5446 ( .CLK(n5564), .C(n5565) );
  CKBD0 U5447 ( .CLK(n5565), .C(n5566) );
  CKBD0 U5448 ( .CLK(n5566), .C(n5567) );
  CKBD0 U5449 ( .CLK(n5567), .C(n5568) );
  CKBD0 U5450 ( .CLK(n5568), .C(n5569) );
  CKBD0 U5451 ( .CLK(n5569), .C(n5570) );
  CKBD0 U5452 ( .CLK(n5570), .C(n5571) );
  CKBD0 U5453 ( .CLK(n5571), .C(n5572) );
  BUFFD0 U5454 ( .I(n5572), .Z(n5573) );
  CKBD0 U5455 ( .CLK(n5573), .C(n5574) );
  CKBD0 U5456 ( .CLK(n5574), .C(n5575) );
  CKBD0 U5457 ( .CLK(n5575), .C(n5576) );
  CKBD0 U5458 ( .CLK(n5576), .C(n5577) );
  CKBD0 U5459 ( .CLK(n5577), .C(n5578) );
  CKBD0 U5460 ( .CLK(n5578), .C(n5579) );
  CKBD0 U5461 ( .CLK(n5579), .C(n5580) );
  CKBD0 U5462 ( .CLK(n5580), .C(n5581) );
  CKBD0 U5463 ( .CLK(n5581), .C(n5582) );
  CKBD0 U5464 ( .CLK(n5582), .C(n5583) );
  BUFFD0 U5465 ( .I(n5583), .Z(n5584) );
  CKBD0 U5466 ( .CLK(n5584), .C(n5585) );
  CKBD0 U5467 ( .CLK(n5585), .C(n5586) );
  CKBD0 U5468 ( .CLK(n5586), .C(n5587) );
  CKBD0 U5469 ( .CLK(n5587), .C(n5588) );
  CKBD0 U5470 ( .CLK(n5588), .C(n5589) );
  CKBD0 U5471 ( .CLK(n5589), .C(n5590) );
  CKBD0 U5472 ( .CLK(n5590), .C(n5591) );
  CKBD0 U5473 ( .CLK(n5591), .C(n5592) );
  CKBD0 U5474 ( .CLK(n5592), .C(n5593) );
  CKBD0 U5475 ( .CLK(n5593), .C(n5594) );
  BUFFD0 U5476 ( .I(n5594), .Z(n5595) );
  CKBD0 U5477 ( .CLK(n5595), .C(n5596) );
  CKBD0 U5478 ( .CLK(n5596), .C(n5597) );
  CKBD0 U5479 ( .CLK(n5597), .C(n5598) );
  CKBD0 U5480 ( .CLK(n5598), .C(n5599) );
  CKBD0 U5481 ( .CLK(n5599), .C(n5600) );
  CKBD0 U5482 ( .CLK(n5600), .C(n5601) );
  CKBD0 U5483 ( .CLK(n5601), .C(n5602) );
  CKBD0 U5484 ( .CLK(n5602), .C(n5603) );
  CKBD0 U5485 ( .CLK(n5603), .C(n5604) );
  CKBD0 U5486 ( .CLK(n5604), .C(n5605) );
  BUFFD0 U5487 ( .I(n5605), .Z(n5606) );
  CKBD0 U5488 ( .CLK(n5606), .C(n5607) );
  CKBD0 U5489 ( .CLK(n5607), .C(n5608) );
  CKBD0 U5490 ( .CLK(n5608), .C(n5609) );
  CKBD0 U5491 ( .CLK(n5609), .C(n5610) );
  CKBD0 U5492 ( .CLK(n5610), .C(n5611) );
  CKBD0 U5493 ( .CLK(n5611), .C(n5612) );
  CKBD0 U5494 ( .CLK(n5612), .C(n5613) );
  CKBD0 U5495 ( .CLK(n5613), .C(n5614) );
  CKBD0 U5496 ( .CLK(n5614), .C(n5615) );
  CKBD0 U5497 ( .CLK(n5615), .C(n5616) );
  BUFFD0 U5498 ( .I(n5616), .Z(n5617) );
  CKBD0 U5499 ( .CLK(n5617), .C(n5618) );
  CKBD0 U5500 ( .CLK(n5618), .C(n5619) );
  CKBD0 U5501 ( .CLK(n5619), .C(n5620) );
  CKBD0 U5502 ( .CLK(n5620), .C(n5621) );
  CKBD0 U5503 ( .CLK(n5621), .C(n5622) );
  CKBD0 U5504 ( .CLK(n5622), .C(n5623) );
  CKBD0 U5505 ( .CLK(n5623), .C(n5624) );
  CKBD0 U5506 ( .CLK(n5624), .C(n5625) );
  CKBD0 U5507 ( .CLK(n5625), .C(n5626) );
  BUFFD0 U5508 ( .I(n5626), .Z(n5627) );
  CKBD0 U5509 ( .CLK(n5627), .C(n5628) );
  CKBD0 U5510 ( .CLK(n5628), .C(n5629) );
  CKBD0 U5511 ( .CLK(n5629), .C(n5630) );
  CKBD0 U5512 ( .CLK(n5630), .C(n5631) );
  CKBD0 U5513 ( .CLK(n5631), .C(n5632) );
  CKBD0 U5514 ( .CLK(n5632), .C(n5633) );
  CKBD0 U5515 ( .CLK(n5633), .C(n5634) );
  CKBD0 U5516 ( .CLK(n5634), .C(n5635) );
  CKBD0 U5517 ( .CLK(n5635), .C(n5636) );
  CKBD0 U5518 ( .CLK(n5636), .C(n5637) );
  BUFFD0 U5519 ( .I(n5637), .Z(n5638) );
  CKBD0 U5520 ( .CLK(n5638), .C(n5639) );
  CKBD0 U5521 ( .CLK(n5639), .C(n5640) );
  CKBD0 U5522 ( .CLK(n5640), .C(n5641) );
  CKBD0 U5523 ( .CLK(n5641), .C(n5642) );
  CKBD0 U5524 ( .CLK(n5642), .C(n5643) );
  CKBD0 U5525 ( .CLK(n5643), .C(n5644) );
  BUFFD0 U5526 ( .I(n5644), .Z(n5645) );
  CKBD0 U5527 ( .CLK(n5645), .C(n5646) );
  BUFFD0 U5528 ( .I(n5646), .Z(n5647) );
  CKBD0 U5529 ( .CLK(n5647), .C(n5648) );
  BUFFD0 U5530 ( .I(n5648), .Z(n5649) );
  CKBD0 U5531 ( .CLK(n5649), .C(n5650) );
  BUFFD0 U5532 ( .I(n5650), .Z(n5651) );
  CKBD0 U5533 ( .CLK(n5651), .C(n5652) );
  BUFFD0 U5534 ( .I(n5652), .Z(n5653) );
  CKBD0 U5535 ( .CLK(n5653), .C(n5654) );
  BUFFD0 U5536 ( .I(n5654), .Z(n5655) );
  CKBD0 U5537 ( .CLK(n5655), .C(n5656) );
  BUFFD0 U5538 ( .I(n5656), .Z(n5657) );
  CKBD0 U5539 ( .CLK(n5657), .C(n5658) );
  BUFFD0 U5540 ( .I(n5658), .Z(n5659) );
  BUFFD0 U5541 ( .I(Decoder[8]), .Z(n5660) );
  BUFFD0 U5542 ( .I(n5662), .Z(n5661) );
  BUFFD0 U5543 ( .I(n5663), .Z(n5662) );
  BUFFD0 U5544 ( .I(n141), .Z(n5663) );
  CKBD0 U5545 ( .CLK(n1120), .C(n5664) );
  CKBD0 U5546 ( .CLK(n5664), .C(n5665) );
  CKBD0 U5547 ( .CLK(n5665), .C(n5666) );
  BUFFD0 U5548 ( .I(n5666), .Z(n5667) );
  CKBD0 U5549 ( .CLK(n5667), .C(n5668) );
  CKBD0 U5550 ( .CLK(n5668), .C(n5669) );
  CKBD0 U5551 ( .CLK(n5669), .C(n5670) );
  CKBD0 U5552 ( .CLK(n5670), .C(n5671) );
  CKBD0 U5553 ( .CLK(n5671), .C(n5672) );
  CKBD0 U5554 ( .CLK(n5672), .C(n5673) );
  CKBD0 U5555 ( .CLK(n5673), .C(n5674) );
  CKBD0 U5556 ( .CLK(n5674), .C(n5675) );
  CKBD0 U5557 ( .CLK(n5675), .C(n5676) );
  CKBD0 U5558 ( .CLK(n5676), .C(n5677) );
  BUFFD0 U5559 ( .I(n5677), .Z(n5678) );
  CKBD0 U5560 ( .CLK(n5678), .C(n5679) );
  CKBD0 U5561 ( .CLK(n5679), .C(n5680) );
  CKBD0 U5562 ( .CLK(n5680), .C(n5681) );
  CKBD0 U5563 ( .CLK(n5681), .C(n5682) );
  CKBD0 U5564 ( .CLK(n5682), .C(n5683) );
  CKBD0 U5565 ( .CLK(n5683), .C(n5684) );
  CKBD0 U5566 ( .CLK(n5684), .C(n5685) );
  CKBD0 U5567 ( .CLK(n5685), .C(n5686) );
  CKBD0 U5568 ( .CLK(n5686), .C(n5687) );
  BUFFD0 U5569 ( .I(n5687), .Z(n5688) );
  CKBD0 U5570 ( .CLK(n5688), .C(n5689) );
  CKBD0 U5571 ( .CLK(n5689), .C(n5690) );
  CKBD0 U5572 ( .CLK(n5690), .C(n5691) );
  CKBD0 U5573 ( .CLK(n5691), .C(n5692) );
  CKBD0 U5574 ( .CLK(n5692), .C(n5693) );
  CKBD0 U5575 ( .CLK(n5693), .C(n5694) );
  CKBD0 U5576 ( .CLK(n5694), .C(n5695) );
  CKBD0 U5577 ( .CLK(n5695), .C(n5696) );
  CKBD0 U5578 ( .CLK(n5696), .C(n5697) );
  CKBD0 U5579 ( .CLK(n5697), .C(n5698) );
  BUFFD0 U5580 ( .I(n5698), .Z(n5699) );
  CKBD0 U5581 ( .CLK(n5699), .C(n5700) );
  CKBD0 U5582 ( .CLK(n5700), .C(n5701) );
  CKBD0 U5583 ( .CLK(n5701), .C(n5702) );
  CKBD0 U5584 ( .CLK(n5702), .C(n5703) );
  CKBD0 U5585 ( .CLK(n5703), .C(n5704) );
  CKBD0 U5586 ( .CLK(n5704), .C(n5705) );
  CKBD0 U5587 ( .CLK(n5705), .C(n5706) );
  CKBD0 U5588 ( .CLK(n5706), .C(n5707) );
  CKBD0 U5589 ( .CLK(n5707), .C(n5708) );
  CKBD0 U5590 ( .CLK(n5708), .C(n5709) );
  BUFFD0 U5591 ( .I(n5709), .Z(n5710) );
  CKBD0 U5592 ( .CLK(n5710), .C(n5711) );
  CKBD0 U5593 ( .CLK(n5711), .C(n5712) );
  CKBD0 U5594 ( .CLK(n5712), .C(n5713) );
  CKBD0 U5595 ( .CLK(n5713), .C(n5714) );
  CKBD0 U5596 ( .CLK(n5714), .C(n5715) );
  CKBD0 U5597 ( .CLK(n5715), .C(n5716) );
  CKBD0 U5598 ( .CLK(n5716), .C(n5717) );
  CKBD0 U5599 ( .CLK(n5717), .C(n5718) );
  CKBD0 U5600 ( .CLK(n5718), .C(n5719) );
  CKBD0 U5601 ( .CLK(n5719), .C(n5720) );
  BUFFD0 U5602 ( .I(n5720), .Z(n5721) );
  CKBD0 U5603 ( .CLK(n5721), .C(n5722) );
  CKBD0 U5604 ( .CLK(n5722), .C(n5723) );
  CKBD0 U5605 ( .CLK(n5723), .C(n5724) );
  CKBD0 U5606 ( .CLK(n5724), .C(n5725) );
  CKBD0 U5607 ( .CLK(n5725), .C(n5726) );
  CKBD0 U5608 ( .CLK(n5726), .C(n5727) );
  CKBD0 U5609 ( .CLK(n5727), .C(n5728) );
  CKBD0 U5610 ( .CLK(n5728), .C(n5729) );
  CKBD0 U5611 ( .CLK(n5729), .C(n5730) );
  CKBD0 U5612 ( .CLK(n5730), .C(n5731) );
  BUFFD0 U5613 ( .I(n5731), .Z(n5732) );
  CKBD0 U5614 ( .CLK(n5732), .C(n5733) );
  CKBD0 U5615 ( .CLK(n5733), .C(n5734) );
  CKBD0 U5616 ( .CLK(n5734), .C(n5735) );
  CKBD0 U5617 ( .CLK(n5735), .C(n5736) );
  CKBD0 U5618 ( .CLK(n5736), .C(n5737) );
  CKBD0 U5619 ( .CLK(n5737), .C(n5738) );
  CKBD0 U5620 ( .CLK(n5738), .C(n5739) );
  CKBD0 U5621 ( .CLK(n5739), .C(n5740) );
  CKBD0 U5622 ( .CLK(n5740), .C(n5741) );
  CKBD0 U5623 ( .CLK(n5741), .C(n5742) );
  BUFFD0 U5624 ( .I(n5742), .Z(n5743) );
  CKBD0 U5625 ( .CLK(n5743), .C(n5744) );
  CKBD0 U5626 ( .CLK(n5744), .C(n5745) );
  CKBD0 U5627 ( .CLK(n5745), .C(n5746) );
  CKBD0 U5628 ( .CLK(n5746), .C(n5747) );
  CKBD0 U5629 ( .CLK(n5747), .C(n5748) );
  CKBD0 U5630 ( .CLK(n5748), .C(n5749) );
  CKBD0 U5631 ( .CLK(n5749), .C(n5750) );
  CKBD0 U5632 ( .CLK(n5750), .C(n5751) );
  CKBD0 U5633 ( .CLK(n5751), .C(n5752) );
  CKBD0 U5634 ( .CLK(n5752), .C(n5753) );
  BUFFD0 U5635 ( .I(n5753), .Z(n5754) );
  CKBD0 U5636 ( .CLK(n5754), .C(n5755) );
  CKBD0 U5637 ( .CLK(n5755), .C(n5756) );
  CKBD0 U5638 ( .CLK(n5756), .C(n5757) );
  CKBD0 U5639 ( .CLK(n5757), .C(n5758) );
  CKBD0 U5640 ( .CLK(n5758), .C(n5759) );
  CKBD0 U5641 ( .CLK(n5759), .C(n5760) );
  CKBD0 U5642 ( .CLK(n5760), .C(n5761) );
  CKBD0 U5643 ( .CLK(n5761), .C(n5762) );
  CKBD0 U5644 ( .CLK(n5762), .C(n5763) );
  BUFFD0 U5645 ( .I(n5763), .Z(n5764) );
  CKBD0 U5646 ( .CLK(n5764), .C(n5765) );
  CKBD0 U5647 ( .CLK(n5765), .C(n5766) );
  CKBD0 U5648 ( .CLK(n5766), .C(n5767) );
  CKBD0 U5649 ( .CLK(n5767), .C(n5768) );
  CKBD0 U5650 ( .CLK(n5768), .C(n5769) );
  CKBD0 U5651 ( .CLK(n5769), .C(n5770) );
  CKBD0 U5652 ( .CLK(n5770), .C(n5771) );
  CKBD0 U5653 ( .CLK(n5771), .C(n5772) );
  CKBD0 U5654 ( .CLK(n5772), .C(n5773) );
  CKBD0 U5655 ( .CLK(n5773), .C(n5774) );
  BUFFD0 U5656 ( .I(n5774), .Z(n5775) );
  CKBD0 U5657 ( .CLK(n5775), .C(n5776) );
  CKBD0 U5658 ( .CLK(n5776), .C(n5777) );
  CKBD0 U5659 ( .CLK(n5777), .C(n5778) );
  CKBD0 U5660 ( .CLK(n5778), .C(n5779) );
  CKBD0 U5661 ( .CLK(n5779), .C(n5780) );
  CKBD0 U5662 ( .CLK(n5780), .C(n5781) );
  BUFFD0 U5663 ( .I(n5781), .Z(n5782) );
  CKBD0 U5664 ( .CLK(n5782), .C(n5783) );
  BUFFD0 U5665 ( .I(n5783), .Z(n5784) );
  CKBD0 U5666 ( .CLK(n5784), .C(n5785) );
  BUFFD0 U5667 ( .I(n5785), .Z(n5786) );
  CKBD0 U5668 ( .CLK(n5786), .C(n5787) );
  BUFFD0 U5669 ( .I(n5787), .Z(n5788) );
  CKBD0 U5670 ( .CLK(n5788), .C(n5789) );
  BUFFD0 U5671 ( .I(n5789), .Z(n5790) );
  CKBD0 U5672 ( .CLK(n5790), .C(n5791) );
  BUFFD0 U5673 ( .I(n5791), .Z(n5792) );
  CKBD0 U5674 ( .CLK(n5792), .C(n5793) );
  BUFFD0 U5675 ( .I(n5793), .Z(n5794) );
  CKBD0 U5676 ( .CLK(n5794), .C(n5795) );
  BUFFD0 U5677 ( .I(n5795), .Z(n5796) );
  BUFFD0 U5678 ( .I(n5798), .Z(n5797) );
  BUFFD0 U5679 ( .I(n5799), .Z(n5798) );
  BUFFD0 U5680 ( .I(n140), .Z(n5799) );
  CKBD0 U5681 ( .CLK(n2531), .C(n5800) );
  CKBD0 U5682 ( .CLK(n5800), .C(n5801) );
  CKBD0 U5683 ( .CLK(n5801), .C(n5802) );
  BUFFD0 U5684 ( .I(n5802), .Z(n5803) );
  CKBD0 U5685 ( .CLK(n5803), .C(n5804) );
  CKBD0 U5686 ( .CLK(n5804), .C(n5805) );
  CKBD0 U5687 ( .CLK(n5805), .C(n5806) );
  CKBD0 U5688 ( .CLK(n5806), .C(n5807) );
  CKBD0 U5689 ( .CLK(n5807), .C(n5808) );
  CKBD0 U5690 ( .CLK(n5808), .C(n5809) );
  CKBD0 U5691 ( .CLK(n5809), .C(n5810) );
  CKBD0 U5692 ( .CLK(n5810), .C(n5811) );
  CKBD0 U5693 ( .CLK(n5811), .C(n5812) );
  CKBD0 U5694 ( .CLK(n5812), .C(n5813) );
  BUFFD0 U5695 ( .I(n5813), .Z(n5814) );
  CKBD0 U5696 ( .CLK(n5814), .C(n5815) );
  CKBD0 U5697 ( .CLK(n5815), .C(n5816) );
  CKBD0 U5698 ( .CLK(n5816), .C(n5817) );
  CKBD0 U5699 ( .CLK(n5817), .C(n5818) );
  CKBD0 U5700 ( .CLK(n5818), .C(n5819) );
  CKBD0 U5701 ( .CLK(n5819), .C(n5820) );
  CKBD0 U5702 ( .CLK(n5820), .C(n5821) );
  CKBD0 U5703 ( .CLK(n5821), .C(n5822) );
  CKBD0 U5704 ( .CLK(n5822), .C(n5823) );
  BUFFD0 U5705 ( .I(n5823), .Z(n5824) );
  CKBD0 U5706 ( .CLK(n5824), .C(n5825) );
  CKBD0 U5707 ( .CLK(n5825), .C(n5826) );
  CKBD0 U5708 ( .CLK(n5826), .C(n5827) );
  CKBD0 U5709 ( .CLK(n5827), .C(n5828) );
  CKBD0 U5710 ( .CLK(n5828), .C(n5829) );
  CKBD0 U5711 ( .CLK(n5829), .C(n5830) );
  CKBD0 U5712 ( .CLK(n5830), .C(n5831) );
  CKBD0 U5713 ( .CLK(n5831), .C(n5832) );
  CKBD0 U5714 ( .CLK(n5832), .C(n5833) );
  CKBD0 U5715 ( .CLK(n5833), .C(n5834) );
  BUFFD0 U5716 ( .I(n5834), .Z(n5835) );
  CKBD0 U5717 ( .CLK(n5835), .C(n5836) );
  CKBD0 U5718 ( .CLK(n5836), .C(n5837) );
  CKBD0 U5719 ( .CLK(n5837), .C(n5838) );
  CKBD0 U5720 ( .CLK(n5838), .C(n5839) );
  CKBD0 U5721 ( .CLK(n5839), .C(n5840) );
  CKBD0 U5722 ( .CLK(n5840), .C(n5841) );
  CKBD0 U5723 ( .CLK(n5841), .C(n5842) );
  CKBD0 U5724 ( .CLK(n5842), .C(n5843) );
  CKBD0 U5725 ( .CLK(n5843), .C(n5844) );
  CKBD0 U5726 ( .CLK(n5844), .C(n5845) );
  BUFFD0 U5727 ( .I(n5845), .Z(n5846) );
  CKBD0 U5728 ( .CLK(n5846), .C(n5847) );
  CKBD0 U5729 ( .CLK(n5847), .C(n5848) );
  CKBD0 U5730 ( .CLK(n5848), .C(n5849) );
  CKBD0 U5731 ( .CLK(n5849), .C(n5850) );
  CKBD0 U5732 ( .CLK(n5850), .C(n5851) );
  CKBD0 U5733 ( .CLK(n5851), .C(n5852) );
  CKBD0 U5734 ( .CLK(n5852), .C(n5853) );
  CKBD0 U5735 ( .CLK(n5853), .C(n5854) );
  CKBD0 U5736 ( .CLK(n5854), .C(n5855) );
  CKBD0 U5737 ( .CLK(n5855), .C(n5856) );
  BUFFD0 U5738 ( .I(n5856), .Z(n5857) );
  CKBD0 U5739 ( .CLK(n5857), .C(n5858) );
  CKBD0 U5740 ( .CLK(n5858), .C(n5859) );
  CKBD0 U5741 ( .CLK(n5859), .C(n5860) );
  CKBD0 U5742 ( .CLK(n5860), .C(n5861) );
  CKBD0 U5743 ( .CLK(n5861), .C(n5862) );
  CKBD0 U5744 ( .CLK(n5862), .C(n5863) );
  CKBD0 U5745 ( .CLK(n5863), .C(n5864) );
  CKBD0 U5746 ( .CLK(n5864), .C(n5865) );
  CKBD0 U5747 ( .CLK(n5865), .C(n5866) );
  CKBD0 U5748 ( .CLK(n5866), .C(n5867) );
  BUFFD0 U5749 ( .I(n5867), .Z(n5868) );
  CKBD0 U5750 ( .CLK(n5868), .C(n5869) );
  CKBD0 U5751 ( .CLK(n5869), .C(n5870) );
  CKBD0 U5752 ( .CLK(n5870), .C(n5871) );
  CKBD0 U5753 ( .CLK(n5871), .C(n5872) );
  CKBD0 U5754 ( .CLK(n5872), .C(n5873) );
  CKBD0 U5755 ( .CLK(n5873), .C(n5874) );
  CKBD0 U5756 ( .CLK(n5874), .C(n5875) );
  CKBD0 U5757 ( .CLK(n5875), .C(n5876) );
  CKBD0 U5758 ( .CLK(n5876), .C(n5877) );
  CKBD0 U5759 ( .CLK(n5877), .C(n5878) );
  BUFFD0 U5760 ( .I(n5878), .Z(n5879) );
  CKBD0 U5761 ( .CLK(n5879), .C(n5880) );
  CKBD0 U5762 ( .CLK(n5880), .C(n5881) );
  CKBD0 U5763 ( .CLK(n5881), .C(n5882) );
  CKBD0 U5764 ( .CLK(n5882), .C(n5883) );
  CKBD0 U5765 ( .CLK(n5883), .C(n5884) );
  CKBD0 U5766 ( .CLK(n5884), .C(n5885) );
  CKBD0 U5767 ( .CLK(n5885), .C(n5886) );
  CKBD0 U5768 ( .CLK(n5886), .C(n5887) );
  CKBD0 U5769 ( .CLK(n5887), .C(n5888) );
  BUFFD0 U5770 ( .I(n5888), .Z(n5889) );
  CKBD0 U5771 ( .CLK(n5889), .C(n5890) );
  CKBD0 U5772 ( .CLK(n5890), .C(n5891) );
  CKBD0 U5773 ( .CLK(n5891), .C(n5892) );
  CKBD0 U5774 ( .CLK(n5892), .C(n5893) );
  CKBD0 U5775 ( .CLK(n5893), .C(n5894) );
  CKBD0 U5776 ( .CLK(n5894), .C(n5895) );
  CKBD0 U5777 ( .CLK(n5895), .C(n5896) );
  CKBD0 U5778 ( .CLK(n5896), .C(n5897) );
  CKBD0 U5779 ( .CLK(n5897), .C(n5898) );
  CKBD0 U5780 ( .CLK(n5898), .C(n5899) );
  BUFFD0 U5781 ( .I(n5899), .Z(n5900) );
  CKBD0 U5782 ( .CLK(n5900), .C(n5901) );
  CKBD0 U5783 ( .CLK(n5901), .C(n5902) );
  CKBD0 U5784 ( .CLK(n5902), .C(n5903) );
  CKBD0 U5785 ( .CLK(n5903), .C(n5904) );
  CKBD0 U5786 ( .CLK(n5904), .C(n5905) );
  CKBD0 U5787 ( .CLK(n5905), .C(n5906) );
  CKBD0 U5788 ( .CLK(n5906), .C(n5907) );
  CKBD0 U5789 ( .CLK(n5907), .C(n5908) );
  CKBD0 U5790 ( .CLK(n5908), .C(n5909) );
  CKBD0 U5791 ( .CLK(n5909), .C(n5910) );
  BUFFD0 U5792 ( .I(n5910), .Z(n5911) );
  CKBD0 U5793 ( .CLK(n5911), .C(n5912) );
  CKBD0 U5794 ( .CLK(n5912), .C(n5913) );
  CKBD0 U5795 ( .CLK(n5913), .C(n5914) );
  CKBD0 U5796 ( .CLK(n5914), .C(n5915) );
  CKBD0 U5797 ( .CLK(n5915), .C(n5916) );
  CKBD0 U5798 ( .CLK(n5916), .C(n5917) );
  BUFFD0 U5799 ( .I(n5917), .Z(n5918) );
  CKBD0 U5800 ( .CLK(n5918), .C(n5919) );
  BUFFD0 U5801 ( .I(n5919), .Z(n5920) );
  CKBD0 U5802 ( .CLK(n5920), .C(n5921) );
  BUFFD0 U5803 ( .I(n5921), .Z(n5922) );
  CKBD0 U5804 ( .CLK(n5922), .C(n5923) );
  BUFFD0 U5805 ( .I(n5923), .Z(n5924) );
  CKBD0 U5806 ( .CLK(n5924), .C(n5925) );
  BUFFD0 U5807 ( .I(n5925), .Z(n5926) );
  CKBD0 U5808 ( .CLK(n5926), .C(n5927) );
  BUFFD0 U5809 ( .I(n5927), .Z(n5928) );
  CKBD0 U5810 ( .CLK(n5928), .C(n5929) );
  BUFFD0 U5811 ( .I(n5929), .Z(n5930) );
  CKBD0 U5812 ( .CLK(n5930), .C(n5931) );
  BUFFD0 U5813 ( .I(n5931), .Z(n5932) );
  BUFFD0 U5814 ( .I(Decoder[6]), .Z(n5933) );
  BUFFD0 U5815 ( .I(n5935), .Z(n5934) );
  BUFFD0 U5816 ( .I(n5936), .Z(n5935) );
  BUFFD0 U5817 ( .I(n139), .Z(n5936) );
  CKBD0 U5818 ( .CLK(n925), .C(n5937) );
  CKBD0 U5819 ( .CLK(n5937), .C(n5938) );
  CKBD0 U5820 ( .CLK(n5938), .C(n5939) );
  BUFFD0 U5821 ( .I(n5939), .Z(n5940) );
  CKBD0 U5822 ( .CLK(n5940), .C(n5941) );
  CKBD0 U5823 ( .CLK(n5941), .C(n5942) );
  CKBD0 U5824 ( .CLK(n5942), .C(n5943) );
  CKBD0 U5825 ( .CLK(n5943), .C(n5944) );
  CKBD0 U5826 ( .CLK(n5944), .C(n5945) );
  CKBD0 U5827 ( .CLK(n5945), .C(n5946) );
  CKBD0 U5828 ( .CLK(n5946), .C(n5947) );
  CKBD0 U5829 ( .CLK(n5947), .C(n5948) );
  CKBD0 U5830 ( .CLK(n5948), .C(n5949) );
  BUFFD0 U5831 ( .I(n5949), .Z(n5950) );
  CKBD0 U5832 ( .CLK(n5950), .C(n5951) );
  CKBD0 U5833 ( .CLK(n5951), .C(n5952) );
  CKBD0 U5834 ( .CLK(n5952), .C(n5953) );
  CKBD0 U5835 ( .CLK(n5953), .C(n5954) );
  CKBD0 U5836 ( .CLK(n5954), .C(n5955) );
  CKBD0 U5837 ( .CLK(n5955), .C(n5956) );
  CKBD0 U5838 ( .CLK(n5956), .C(n5957) );
  CKBD0 U5839 ( .CLK(n5957), .C(n5958) );
  CKBD0 U5840 ( .CLK(n5958), .C(n5959) );
  CKBD0 U5841 ( .CLK(n5959), .C(n5960) );
  BUFFD0 U5842 ( .I(n5960), .Z(n5961) );
  CKBD0 U5843 ( .CLK(n5961), .C(n5962) );
  CKBD0 U5844 ( .CLK(n5962), .C(n5963) );
  CKBD0 U5845 ( .CLK(n5963), .C(n5964) );
  CKBD0 U5846 ( .CLK(n5964), .C(n5965) );
  CKBD0 U5847 ( .CLK(n5965), .C(n5966) );
  CKBD0 U5848 ( .CLK(n5966), .C(n5967) );
  CKBD0 U5849 ( .CLK(n5967), .C(n5968) );
  CKBD0 U5850 ( .CLK(n5968), .C(n5969) );
  CKBD0 U5851 ( .CLK(n5969), .C(n5970) );
  CKBD0 U5852 ( .CLK(n5970), .C(n5971) );
  BUFFD0 U5853 ( .I(n5971), .Z(n5972) );
  CKBD0 U5854 ( .CLK(n5972), .C(n5973) );
  CKBD0 U5855 ( .CLK(n5973), .C(n5974) );
  CKBD0 U5856 ( .CLK(n5974), .C(n5975) );
  CKBD0 U5857 ( .CLK(n5975), .C(n5976) );
  CKBD0 U5858 ( .CLK(n5976), .C(n5977) );
  CKBD0 U5859 ( .CLK(n5977), .C(n5978) );
  CKBD0 U5860 ( .CLK(n5978), .C(n5979) );
  CKBD0 U5861 ( .CLK(n5979), .C(n5980) );
  CKBD0 U5862 ( .CLK(n5980), .C(n5981) );
  CKBD0 U5863 ( .CLK(n5981), .C(n5982) );
  BUFFD0 U5864 ( .I(n5982), .Z(n5983) );
  CKBD0 U5865 ( .CLK(n5983), .C(n5984) );
  CKBD0 U5866 ( .CLK(n5984), .C(n5985) );
  CKBD0 U5867 ( .CLK(n5985), .C(n5986) );
  CKBD0 U5868 ( .CLK(n5986), .C(n5987) );
  CKBD0 U5869 ( .CLK(n5987), .C(n5988) );
  CKBD0 U5870 ( .CLK(n5988), .C(n5989) );
  CKBD0 U5871 ( .CLK(n5989), .C(n5990) );
  CKBD0 U5872 ( .CLK(n5990), .C(n5991) );
  CKBD0 U5873 ( .CLK(n5991), .C(n5992) );
  CKBD0 U5874 ( .CLK(n5992), .C(n5993) );
  BUFFD0 U5875 ( .I(n5993), .Z(n5994) );
  CKBD0 U5876 ( .CLK(n5994), .C(n5995) );
  CKBD0 U5877 ( .CLK(n5995), .C(n5996) );
  CKBD0 U5878 ( .CLK(n5996), .C(n5997) );
  CKBD0 U5879 ( .CLK(n5997), .C(n5998) );
  CKBD0 U5880 ( .CLK(n5998), .C(n5999) );
  CKBD0 U5881 ( .CLK(n5999), .C(n6000) );
  CKBD0 U5882 ( .CLK(n6000), .C(n6001) );
  CKBD0 U5883 ( .CLK(n6001), .C(n6002) );
  CKBD0 U5884 ( .CLK(n6002), .C(n6003) );
  CKBD0 U5885 ( .CLK(n6003), .C(n6004) );
  BUFFD0 U5886 ( .I(n6004), .Z(n6005) );
  CKBD0 U5887 ( .CLK(n6005), .C(n6006) );
  CKBD0 U5888 ( .CLK(n6006), .C(n6007) );
  CKBD0 U5889 ( .CLK(n6007), .C(n6008) );
  CKBD0 U5890 ( .CLK(n6008), .C(n6009) );
  CKBD0 U5891 ( .CLK(n6009), .C(n6010) );
  CKBD0 U5892 ( .CLK(n6010), .C(n6011) );
  CKBD0 U5893 ( .CLK(n6011), .C(n6012) );
  CKBD0 U5894 ( .CLK(n6012), .C(n6013) );
  CKBD0 U5895 ( .CLK(n6013), .C(n6014) );
  CKBD0 U5896 ( .CLK(n6014), .C(n6015) );
  BUFFD0 U5897 ( .I(n6015), .Z(n6016) );
  CKBD0 U5898 ( .CLK(n6016), .C(n6017) );
  CKBD0 U5899 ( .CLK(n6017), .C(n6018) );
  CKBD0 U5900 ( .CLK(n6018), .C(n6019) );
  CKBD0 U5901 ( .CLK(n6019), .C(n6020) );
  CKBD0 U5902 ( .CLK(n6020), .C(n6021) );
  CKBD0 U5903 ( .CLK(n6021), .C(n6022) );
  CKBD0 U5904 ( .CLK(n6022), .C(n6023) );
  CKBD0 U5905 ( .CLK(n6023), .C(n6024) );
  CKBD0 U5906 ( .CLK(n6024), .C(n6025) );
  BUFFD0 U5907 ( .I(n6025), .Z(n6026) );
  CKBD0 U5908 ( .CLK(n6026), .C(n6027) );
  CKBD0 U5909 ( .CLK(n6027), .C(n6028) );
  CKBD0 U5910 ( .CLK(n6028), .C(n6029) );
  CKBD0 U5911 ( .CLK(n6029), .C(n6030) );
  CKBD0 U5912 ( .CLK(n6030), .C(n6031) );
  CKBD0 U5913 ( .CLK(n6031), .C(n6032) );
  CKBD0 U5914 ( .CLK(n6032), .C(n6033) );
  CKBD0 U5915 ( .CLK(n6033), .C(n6034) );
  CKBD0 U5916 ( .CLK(n6034), .C(n6035) );
  CKBD0 U5917 ( .CLK(n6035), .C(n6036) );
  BUFFD0 U5918 ( .I(n6036), .Z(n6037) );
  CKBD0 U5919 ( .CLK(n6037), .C(n6038) );
  CKBD0 U5920 ( .CLK(n6038), .C(n6039) );
  CKBD0 U5921 ( .CLK(n6039), .C(n6040) );
  CKBD0 U5922 ( .CLK(n6040), .C(n6041) );
  CKBD0 U5923 ( .CLK(n6041), .C(n6042) );
  CKBD0 U5924 ( .CLK(n6042), .C(n6043) );
  CKBD0 U5925 ( .CLK(n6043), .C(n6044) );
  CKBD0 U5926 ( .CLK(n6044), .C(n6045) );
  CKBD0 U5927 ( .CLK(n6045), .C(n6046) );
  CKBD0 U5928 ( .CLK(n6046), .C(n6047) );
  BUFFD0 U5929 ( .I(n6047), .Z(n6048) );
  CKBD0 U5930 ( .CLK(n6048), .C(n6049) );
  CKBD0 U5931 ( .CLK(n6049), .C(n6050) );
  CKBD0 U5932 ( .CLK(n6050), .C(n6051) );
  CKBD0 U5933 ( .CLK(n6051), .C(n6052) );
  CKBD0 U5934 ( .CLK(n6052), .C(n6053) );
  CKBD0 U5935 ( .CLK(n6053), .C(n6054) );
  BUFFD0 U5936 ( .I(n6054), .Z(n6055) );
  CKBD0 U5937 ( .CLK(n6055), .C(n6056) );
  BUFFD0 U5938 ( .I(n6056), .Z(n6057) );
  CKBD0 U5939 ( .CLK(n6057), .C(n6058) );
  BUFFD0 U5940 ( .I(n6058), .Z(n6059) );
  CKBD0 U5941 ( .CLK(n6059), .C(n6060) );
  BUFFD0 U5942 ( .I(n6060), .Z(n6061) );
  CKBD0 U5943 ( .CLK(n6061), .C(n6062) );
  BUFFD0 U5944 ( .I(n6062), .Z(n6063) );
  CKBD0 U5945 ( .CLK(n6063), .C(n6064) );
  BUFFD0 U5946 ( .I(n6064), .Z(n6065) );
  CKBD0 U5947 ( .CLK(n6065), .C(n6066) );
  BUFFD0 U5948 ( .I(n6066), .Z(n6067) );
  CKBD0 U5949 ( .CLK(n6067), .C(n6068) );
  BUFFD0 U5950 ( .I(n6068), .Z(n6069) );
  BUFFD0 U5951 ( .I(n138), .Z(n6070) );
  BUFFD0 U5952 ( .I(n6072), .Z(n6071) );
  BUFFD0 U5953 ( .I(n6073), .Z(n6072) );
  BUFFD0 U5954 ( .I(Decoder[5]), .Z(n6073) );
  CKBD0 U5955 ( .CLK(n923), .C(n6074) );
  CKBD0 U5956 ( .CLK(n6074), .C(n6075) );
  CKBD0 U5957 ( .CLK(n6075), .C(n6076) );
  BUFFD0 U5958 ( .I(n6076), .Z(n6077) );
  CKBD0 U5959 ( .CLK(n6077), .C(n6078) );
  CKBD0 U5960 ( .CLK(n6078), .C(n6079) );
  CKBD0 U5961 ( .CLK(n6079), .C(n6080) );
  CKBD0 U5962 ( .CLK(n6080), .C(n6081) );
  CKBD0 U5963 ( .CLK(n6081), .C(n6082) );
  CKBD0 U5964 ( .CLK(n6082), .C(n6083) );
  CKBD0 U5965 ( .CLK(n6083), .C(n6084) );
  CKBD0 U5966 ( .CLK(n6084), .C(n6085) );
  CKBD0 U5967 ( .CLK(n6085), .C(n6086) );
  CKBD0 U5968 ( .CLK(n6086), .C(n6087) );
  BUFFD0 U5969 ( .I(n6087), .Z(n6088) );
  CKBD0 U5970 ( .CLK(n6088), .C(n6089) );
  CKBD0 U5971 ( .CLK(n6089), .C(n6090) );
  CKBD0 U5972 ( .CLK(n6090), .C(n6091) );
  CKBD0 U5973 ( .CLK(n6091), .C(n6092) );
  CKBD0 U5974 ( .CLK(n6092), .C(n6093) );
  CKBD0 U5975 ( .CLK(n6093), .C(n6094) );
  CKBD0 U5976 ( .CLK(n6094), .C(n6095) );
  CKBD0 U5977 ( .CLK(n6095), .C(n6096) );
  CKBD0 U5978 ( .CLK(n6096), .C(n6097) );
  BUFFD0 U5979 ( .I(n6097), .Z(n6098) );
  CKBD0 U5980 ( .CLK(n6098), .C(n6099) );
  CKBD0 U5981 ( .CLK(n6099), .C(n6100) );
  CKBD0 U5982 ( .CLK(n6100), .C(n6101) );
  CKBD0 U5983 ( .CLK(n6101), .C(n6102) );
  CKBD0 U5984 ( .CLK(n6102), .C(n6103) );
  CKBD0 U5985 ( .CLK(n6103), .C(n6104) );
  CKBD0 U5986 ( .CLK(n6104), .C(n6105) );
  CKBD0 U5987 ( .CLK(n6105), .C(n6106) );
  CKBD0 U5988 ( .CLK(n6106), .C(n6107) );
  CKBD0 U5989 ( .CLK(n6107), .C(n6108) );
  BUFFD0 U5990 ( .I(n6108), .Z(n6109) );
  CKBD0 U5991 ( .CLK(n6109), .C(n6110) );
  CKBD0 U5992 ( .CLK(n6110), .C(n6111) );
  CKBD0 U5993 ( .CLK(n6111), .C(n6112) );
  CKBD0 U5994 ( .CLK(n6112), .C(n6113) );
  CKBD0 U5995 ( .CLK(n6113), .C(n6114) );
  CKBD0 U5996 ( .CLK(n6114), .C(n6115) );
  CKBD0 U5997 ( .CLK(n6115), .C(n6116) );
  CKBD0 U5998 ( .CLK(n6116), .C(n6117) );
  CKBD0 U5999 ( .CLK(n6117), .C(n6118) );
  CKBD0 U6000 ( .CLK(n6118), .C(n6119) );
  BUFFD0 U6001 ( .I(n6119), .Z(n6120) );
  CKBD0 U6002 ( .CLK(n6120), .C(n6121) );
  CKBD0 U6003 ( .CLK(n6121), .C(n6122) );
  CKBD0 U6004 ( .CLK(n6122), .C(n6123) );
  CKBD0 U6005 ( .CLK(n6123), .C(n6124) );
  CKBD0 U6006 ( .CLK(n6124), .C(n6125) );
  CKBD0 U6007 ( .CLK(n6125), .C(n6126) );
  CKBD0 U6008 ( .CLK(n6126), .C(n6127) );
  CKBD0 U6009 ( .CLK(n6127), .C(n6128) );
  CKBD0 U6010 ( .CLK(n6128), .C(n6129) );
  CKBD0 U6011 ( .CLK(n6129), .C(n6130) );
  BUFFD0 U6012 ( .I(n6130), .Z(n6131) );
  CKBD0 U6013 ( .CLK(n6131), .C(n6132) );
  CKBD0 U6014 ( .CLK(n6132), .C(n6133) );
  CKBD0 U6015 ( .CLK(n6133), .C(n6134) );
  CKBD0 U6016 ( .CLK(n6134), .C(n6135) );
  CKBD0 U6017 ( .CLK(n6135), .C(n6136) );
  CKBD0 U6018 ( .CLK(n6136), .C(n6137) );
  CKBD0 U6019 ( .CLK(n6137), .C(n6138) );
  CKBD0 U6020 ( .CLK(n6138), .C(n6139) );
  CKBD0 U6021 ( .CLK(n6139), .C(n6140) );
  CKBD0 U6022 ( .CLK(n6140), .C(n6141) );
  BUFFD0 U6023 ( .I(n6141), .Z(n6142) );
  CKBD0 U6024 ( .CLK(n6142), .C(n6143) );
  CKBD0 U6025 ( .CLK(n6143), .C(n6144) );
  CKBD0 U6026 ( .CLK(n6144), .C(n6145) );
  CKBD0 U6027 ( .CLK(n6145), .C(n6146) );
  CKBD0 U6028 ( .CLK(n6146), .C(n6147) );
  CKBD0 U6029 ( .CLK(n6147), .C(n6148) );
  CKBD0 U6030 ( .CLK(n6148), .C(n6149) );
  CKBD0 U6031 ( .CLK(n6149), .C(n6150) );
  CKBD0 U6032 ( .CLK(n6150), .C(n6151) );
  CKBD0 U6033 ( .CLK(n6151), .C(n6152) );
  BUFFD0 U6034 ( .I(n6152), .Z(n6153) );
  CKBD0 U6035 ( .CLK(n6153), .C(n6154) );
  CKBD0 U6036 ( .CLK(n6154), .C(n6155) );
  CKBD0 U6037 ( .CLK(n6155), .C(n6156) );
  CKBD0 U6038 ( .CLK(n6156), .C(n6157) );
  CKBD0 U6039 ( .CLK(n6157), .C(n6158) );
  CKBD0 U6040 ( .CLK(n6158), .C(n6159) );
  CKBD0 U6041 ( .CLK(n6159), .C(n6160) );
  CKBD0 U6042 ( .CLK(n6160), .C(n6161) );
  CKBD0 U6043 ( .CLK(n6161), .C(n6162) );
  BUFFD0 U6044 ( .I(n6162), .Z(n6163) );
  CKBD0 U6045 ( .CLK(n6163), .C(n6164) );
  CKBD0 U6046 ( .CLK(n6164), .C(n6165) );
  CKBD0 U6047 ( .CLK(n6165), .C(n6166) );
  CKBD0 U6048 ( .CLK(n6166), .C(n6167) );
  CKBD0 U6049 ( .CLK(n6167), .C(n6168) );
  CKBD0 U6050 ( .CLK(n6168), .C(n6169) );
  CKBD0 U6051 ( .CLK(n6169), .C(n6170) );
  CKBD0 U6052 ( .CLK(n6170), .C(n6171) );
  CKBD0 U6053 ( .CLK(n6171), .C(n6172) );
  CKBD0 U6054 ( .CLK(n6172), .C(n6173) );
  BUFFD0 U6055 ( .I(n6173), .Z(n6174) );
  CKBD0 U6056 ( .CLK(n6174), .C(n6175) );
  CKBD0 U6057 ( .CLK(n6175), .C(n6176) );
  CKBD0 U6058 ( .CLK(n6176), .C(n6177) );
  CKBD0 U6059 ( .CLK(n6177), .C(n6178) );
  CKBD0 U6060 ( .CLK(n6178), .C(n6179) );
  CKBD0 U6061 ( .CLK(n6179), .C(n6180) );
  CKBD0 U6062 ( .CLK(n6180), .C(n6181) );
  CKBD0 U6063 ( .CLK(n6181), .C(n6182) );
  CKBD0 U6064 ( .CLK(n6182), .C(n6183) );
  CKBD0 U6065 ( .CLK(n6183), .C(n6184) );
  BUFFD0 U6066 ( .I(n6184), .Z(n6185) );
  CKBD0 U6067 ( .CLK(n6185), .C(n6186) );
  CKBD0 U6068 ( .CLK(n6186), .C(n6187) );
  CKBD0 U6069 ( .CLK(n6187), .C(n6188) );
  CKBD0 U6070 ( .CLK(n6188), .C(n6189) );
  CKBD0 U6071 ( .CLK(n6189), .C(n6190) );
  CKBD0 U6072 ( .CLK(n6190), .C(n6191) );
  BUFFD0 U6073 ( .I(n6191), .Z(n6192) );
  CKBD0 U6074 ( .CLK(n6192), .C(n6193) );
  BUFFD0 U6075 ( .I(n6193), .Z(n6194) );
  CKBD0 U6076 ( .CLK(n6194), .C(n6195) );
  BUFFD0 U6077 ( .I(n6195), .Z(n6196) );
  CKBD0 U6078 ( .CLK(n6196), .C(n6197) );
  BUFFD0 U6079 ( .I(n6197), .Z(n6198) );
  CKBD0 U6080 ( .CLK(n6198), .C(n6199) );
  BUFFD0 U6081 ( .I(n6199), .Z(n6200) );
  CKBD0 U6082 ( .CLK(n6200), .C(n6201) );
  BUFFD0 U6083 ( .I(n6201), .Z(n6202) );
  CKBD0 U6084 ( .CLK(n6202), .C(n6203) );
  BUFFD0 U6085 ( .I(n6203), .Z(n6204) );
  CKBD0 U6086 ( .CLK(n6204), .C(n6205) );
  BUFFD0 U6087 ( .I(n6205), .Z(n6206) );
  BUFFD0 U6088 ( .I(n137), .Z(n6207) );
  BUFFD0 U6089 ( .I(n6209), .Z(n6208) );
  BUFFD0 U6090 ( .I(n6210), .Z(n6209) );
  BUFFD0 U6091 ( .I(Decoder[4]), .Z(n6210) );
  CKBD0 U6092 ( .CLK(n921), .C(n6211) );
  CKBD0 U6093 ( .CLK(n6211), .C(n6212) );
  CKBD0 U6094 ( .CLK(n6212), .C(n6213) );
  BUFFD0 U6095 ( .I(n6213), .Z(n6214) );
  CKBD0 U6096 ( .CLK(n6214), .C(n6215) );
  CKBD0 U6097 ( .CLK(n6215), .C(n6216) );
  CKBD0 U6098 ( .CLK(n6216), .C(n6217) );
  CKBD0 U6099 ( .CLK(n6217), .C(n6218) );
  CKBD0 U6100 ( .CLK(n6218), .C(n6219) );
  CKBD0 U6101 ( .CLK(n6219), .C(n6220) );
  CKBD0 U6102 ( .CLK(n6220), .C(n6221) );
  CKBD0 U6103 ( .CLK(n6221), .C(n6222) );
  CKBD0 U6104 ( .CLK(n6222), .C(n6223) );
  CKBD0 U6105 ( .CLK(n6223), .C(n6224) );
  BUFFD0 U6106 ( .I(n6224), .Z(n6225) );
  CKBD0 U6107 ( .CLK(n6225), .C(n6226) );
  CKBD0 U6108 ( .CLK(n6226), .C(n6227) );
  CKBD0 U6109 ( .CLK(n6227), .C(n6228) );
  CKBD0 U6110 ( .CLK(n6228), .C(n6229) );
  CKBD0 U6111 ( .CLK(n6229), .C(n6230) );
  CKBD0 U6112 ( .CLK(n6230), .C(n6231) );
  CKBD0 U6113 ( .CLK(n6231), .C(n6232) );
  CKBD0 U6114 ( .CLK(n6232), .C(n6233) );
  CKBD0 U6115 ( .CLK(n6233), .C(n6234) );
  BUFFD0 U6116 ( .I(n6234), .Z(n6235) );
  CKBD0 U6117 ( .CLK(n6235), .C(n6236) );
  CKBD0 U6118 ( .CLK(n6236), .C(n6237) );
  CKBD0 U6119 ( .CLK(n6237), .C(n6238) );
  CKBD0 U6120 ( .CLK(n6238), .C(n6239) );
  CKBD0 U6121 ( .CLK(n6239), .C(n6240) );
  CKBD0 U6122 ( .CLK(n6240), .C(n6241) );
  CKBD0 U6123 ( .CLK(n6241), .C(n6242) );
  CKBD0 U6124 ( .CLK(n6242), .C(n6243) );
  CKBD0 U6125 ( .CLK(n6243), .C(n6244) );
  CKBD0 U6126 ( .CLK(n6244), .C(n6245) );
  BUFFD0 U6127 ( .I(n6245), .Z(n6246) );
  CKBD0 U6128 ( .CLK(n6246), .C(n6247) );
  CKBD0 U6129 ( .CLK(n6247), .C(n6248) );
  CKBD0 U6130 ( .CLK(n6248), .C(n6249) );
  CKBD0 U6131 ( .CLK(n6249), .C(n6250) );
  CKBD0 U6132 ( .CLK(n6250), .C(n6251) );
  CKBD0 U6133 ( .CLK(n6251), .C(n6252) );
  CKBD0 U6134 ( .CLK(n6252), .C(n6253) );
  CKBD0 U6135 ( .CLK(n6253), .C(n6254) );
  CKBD0 U6136 ( .CLK(n6254), .C(n6255) );
  CKBD0 U6137 ( .CLK(n6255), .C(n6256) );
  BUFFD0 U6138 ( .I(n6256), .Z(n6257) );
  CKBD0 U6139 ( .CLK(n6257), .C(n6258) );
  CKBD0 U6140 ( .CLK(n6258), .C(n6259) );
  CKBD0 U6141 ( .CLK(n6259), .C(n6260) );
  CKBD0 U6142 ( .CLK(n6260), .C(n6261) );
  CKBD0 U6143 ( .CLK(n6261), .C(n6262) );
  CKBD0 U6144 ( .CLK(n6262), .C(n6263) );
  CKBD0 U6145 ( .CLK(n6263), .C(n6264) );
  CKBD0 U6146 ( .CLK(n6264), .C(n6265) );
  CKBD0 U6147 ( .CLK(n6265), .C(n6266) );
  CKBD0 U6148 ( .CLK(n6266), .C(n6267) );
  BUFFD0 U6149 ( .I(n6267), .Z(n6268) );
  CKBD0 U6150 ( .CLK(n6268), .C(n6269) );
  CKBD0 U6151 ( .CLK(n6269), .C(n6270) );
  CKBD0 U6152 ( .CLK(n6270), .C(n6271) );
  CKBD0 U6153 ( .CLK(n6271), .C(n6272) );
  CKBD0 U6154 ( .CLK(n6272), .C(n6273) );
  CKBD0 U6155 ( .CLK(n6273), .C(n6274) );
  CKBD0 U6156 ( .CLK(n6274), .C(n6275) );
  CKBD0 U6157 ( .CLK(n6275), .C(n6276) );
  CKBD0 U6158 ( .CLK(n6276), .C(n6277) );
  CKBD0 U6159 ( .CLK(n6277), .C(n6278) );
  BUFFD0 U6160 ( .I(n6278), .Z(n6279) );
  CKBD0 U6161 ( .CLK(n6279), .C(n6280) );
  CKBD0 U6162 ( .CLK(n6280), .C(n6281) );
  CKBD0 U6163 ( .CLK(n6281), .C(n6282) );
  CKBD0 U6164 ( .CLK(n6282), .C(n6283) );
  CKBD0 U6165 ( .CLK(n6283), .C(n6284) );
  CKBD0 U6166 ( .CLK(n6284), .C(n6285) );
  CKBD0 U6167 ( .CLK(n6285), .C(n6286) );
  CKBD0 U6168 ( .CLK(n6286), .C(n6287) );
  CKBD0 U6169 ( .CLK(n6287), .C(n6288) );
  CKBD0 U6170 ( .CLK(n6288), .C(n6289) );
  BUFFD0 U6171 ( .I(n6289), .Z(n6290) );
  CKBD0 U6172 ( .CLK(n6290), .C(n6291) );
  CKBD0 U6173 ( .CLK(n6291), .C(n6292) );
  CKBD0 U6174 ( .CLK(n6292), .C(n6293) );
  CKBD0 U6175 ( .CLK(n6293), .C(n6294) );
  CKBD0 U6176 ( .CLK(n6294), .C(n6295) );
  CKBD0 U6177 ( .CLK(n6295), .C(n6296) );
  CKBD0 U6178 ( .CLK(n6296), .C(n6297) );
  CKBD0 U6179 ( .CLK(n6297), .C(n6298) );
  CKBD0 U6180 ( .CLK(n6298), .C(n6299) );
  CKBD0 U6181 ( .CLK(n6299), .C(n6300) );
  BUFFD0 U6182 ( .I(n6300), .Z(n6301) );
  CKBD0 U6183 ( .CLK(n6301), .C(n6302) );
  CKBD0 U6184 ( .CLK(n6302), .C(n6303) );
  CKBD0 U6185 ( .CLK(n6303), .C(n6304) );
  CKBD0 U6186 ( .CLK(n6304), .C(n6305) );
  CKBD0 U6187 ( .CLK(n6305), .C(n6306) );
  CKBD0 U6188 ( .CLK(n6306), .C(n6307) );
  CKBD0 U6189 ( .CLK(n6307), .C(n6308) );
  CKBD0 U6190 ( .CLK(n6308), .C(n6309) );
  CKBD0 U6191 ( .CLK(n6309), .C(n6310) );
  BUFFD0 U6192 ( .I(n6310), .Z(n6311) );
  CKBD0 U6193 ( .CLK(n6311), .C(n6312) );
  CKBD0 U6194 ( .CLK(n6312), .C(n6313) );
  CKBD0 U6195 ( .CLK(n6313), .C(n6314) );
  CKBD0 U6196 ( .CLK(n6314), .C(n6315) );
  CKBD0 U6197 ( .CLK(n6315), .C(n6316) );
  CKBD0 U6198 ( .CLK(n6316), .C(n6317) );
  CKBD0 U6199 ( .CLK(n6317), .C(n6318) );
  CKBD0 U6200 ( .CLK(n6318), .C(n6319) );
  CKBD0 U6201 ( .CLK(n6319), .C(n6320) );
  CKBD0 U6202 ( .CLK(n6320), .C(n6321) );
  BUFFD0 U6203 ( .I(n6321), .Z(n6322) );
  CKBD0 U6204 ( .CLK(n6322), .C(n6323) );
  CKBD0 U6205 ( .CLK(n6323), .C(n6324) );
  CKBD0 U6206 ( .CLK(n6324), .C(n6325) );
  CKBD0 U6207 ( .CLK(n6325), .C(n6326) );
  CKBD0 U6208 ( .CLK(n6326), .C(n6327) );
  CKBD0 U6209 ( .CLK(n6327), .C(n6328) );
  BUFFD0 U6210 ( .I(n6328), .Z(n6329) );
  CKBD0 U6211 ( .CLK(n6329), .C(n6330) );
  BUFFD0 U6212 ( .I(n6330), .Z(n6331) );
  CKBD0 U6213 ( .CLK(n6331), .C(n6332) );
  BUFFD0 U6214 ( .I(n6332), .Z(n6333) );
  CKBD0 U6215 ( .CLK(n6333), .C(n6334) );
  BUFFD0 U6216 ( .I(n6334), .Z(n6335) );
  CKBD0 U6217 ( .CLK(n6335), .C(n6336) );
  BUFFD0 U6218 ( .I(n6336), .Z(n6337) );
  CKBD0 U6219 ( .CLK(n6337), .C(n6338) );
  BUFFD0 U6220 ( .I(n6338), .Z(n6339) );
  CKBD0 U6221 ( .CLK(n6339), .C(n6340) );
  BUFFD0 U6222 ( .I(n6340), .Z(n6341) );
  CKBD0 U6223 ( .CLK(n6341), .C(n6342) );
  BUFFD0 U6224 ( .I(n6342), .Z(n6343) );
  BUFFD0 U6225 ( .I(n136), .Z(n6344) );
  BUFFD0 U6226 ( .I(n6346), .Z(n6345) );
  BUFFD0 U6227 ( .I(n6347), .Z(n6346) );
  BUFFD0 U6228 ( .I(Decoder[3]), .Z(n6347) );
  CKBD0 U6229 ( .CLK(n919), .C(n6348) );
  CKBD0 U6230 ( .CLK(n6348), .C(n6349) );
  CKBD0 U6231 ( .CLK(n6349), .C(n6350) );
  BUFFD0 U6232 ( .I(n6350), .Z(n6351) );
  CKBD0 U6233 ( .CLK(n6351), .C(n6352) );
  CKBD0 U6234 ( .CLK(n6352), .C(n6353) );
  CKBD0 U6235 ( .CLK(n6353), .C(n6354) );
  CKBD0 U6236 ( .CLK(n6354), .C(n6355) );
  CKBD0 U6237 ( .CLK(n6355), .C(n6356) );
  CKBD0 U6238 ( .CLK(n6356), .C(n6357) );
  CKBD0 U6239 ( .CLK(n6357), .C(n6358) );
  CKBD0 U6240 ( .CLK(n6358), .C(n6359) );
  CKBD0 U6241 ( .CLK(n6359), .C(n6360) );
  CKBD0 U6242 ( .CLK(n6360), .C(n6361) );
  BUFFD0 U6243 ( .I(n6361), .Z(n6362) );
  CKBD0 U6244 ( .CLK(n6362), .C(n6363) );
  CKBD0 U6245 ( .CLK(n6363), .C(n6364) );
  CKBD0 U6246 ( .CLK(n6364), .C(n6365) );
  CKBD0 U6247 ( .CLK(n6365), .C(n6366) );
  CKBD0 U6248 ( .CLK(n6366), .C(n6367) );
  CKBD0 U6249 ( .CLK(n6367), .C(n6368) );
  CKBD0 U6250 ( .CLK(n6368), .C(n6369) );
  CKBD0 U6251 ( .CLK(n6369), .C(n6370) );
  CKBD0 U6252 ( .CLK(n6370), .C(n6371) );
  BUFFD0 U6253 ( .I(n6371), .Z(n6372) );
  CKBD0 U6254 ( .CLK(n6372), .C(n6373) );
  CKBD0 U6255 ( .CLK(n6373), .C(n6374) );
  CKBD0 U6256 ( .CLK(n6374), .C(n6375) );
  CKBD0 U6257 ( .CLK(n6375), .C(n6376) );
  CKBD0 U6258 ( .CLK(n6376), .C(n6377) );
  CKBD0 U6259 ( .CLK(n6377), .C(n6378) );
  CKBD0 U6260 ( .CLK(n6378), .C(n6379) );
  CKBD0 U6261 ( .CLK(n6379), .C(n6380) );
  CKBD0 U6262 ( .CLK(n6380), .C(n6381) );
  CKBD0 U6263 ( .CLK(n6381), .C(n6382) );
  BUFFD0 U6264 ( .I(n6382), .Z(n6383) );
  CKBD0 U6265 ( .CLK(n6383), .C(n6384) );
  CKBD0 U6266 ( .CLK(n6384), .C(n6385) );
  CKBD0 U6267 ( .CLK(n6385), .C(n6386) );
  CKBD0 U6268 ( .CLK(n6386), .C(n6387) );
  CKBD0 U6269 ( .CLK(n6387), .C(n6388) );
  CKBD0 U6270 ( .CLK(n6388), .C(n6389) );
  CKBD0 U6271 ( .CLK(n6389), .C(n6390) );
  CKBD0 U6272 ( .CLK(n6390), .C(n6391) );
  CKBD0 U6273 ( .CLK(n6391), .C(n6392) );
  CKBD0 U6274 ( .CLK(n6392), .C(n6393) );
  BUFFD0 U6275 ( .I(n6393), .Z(n6394) );
  CKBD0 U6276 ( .CLK(n6394), .C(n6395) );
  CKBD0 U6277 ( .CLK(n6395), .C(n6396) );
  CKBD0 U6278 ( .CLK(n6396), .C(n6397) );
  CKBD0 U6279 ( .CLK(n6397), .C(n6398) );
  CKBD0 U6280 ( .CLK(n6398), .C(n6399) );
  CKBD0 U6281 ( .CLK(n6399), .C(n6400) );
  CKBD0 U6282 ( .CLK(n6400), .C(n6401) );
  CKBD0 U6283 ( .CLK(n6401), .C(n6402) );
  CKBD0 U6284 ( .CLK(n6402), .C(n6403) );
  CKBD0 U6285 ( .CLK(n6403), .C(n6404) );
  BUFFD0 U6286 ( .I(n6404), .Z(n6405) );
  CKBD0 U6287 ( .CLK(n6405), .C(n6406) );
  CKBD0 U6288 ( .CLK(n6406), .C(n6407) );
  CKBD0 U6289 ( .CLK(n6407), .C(n6408) );
  CKBD0 U6290 ( .CLK(n6408), .C(n6409) );
  CKBD0 U6291 ( .CLK(n6409), .C(n6410) );
  CKBD0 U6292 ( .CLK(n6410), .C(n6411) );
  CKBD0 U6293 ( .CLK(n6411), .C(n6412) );
  CKBD0 U6294 ( .CLK(n6412), .C(n6413) );
  CKBD0 U6295 ( .CLK(n6413), .C(n6414) );
  CKBD0 U6296 ( .CLK(n6414), .C(n6415) );
  BUFFD0 U6297 ( .I(n6415), .Z(n6416) );
  CKBD0 U6298 ( .CLK(n6416), .C(n6417) );
  CKBD0 U6299 ( .CLK(n6417), .C(n6418) );
  CKBD0 U6300 ( .CLK(n6418), .C(n6419) );
  CKBD0 U6301 ( .CLK(n6419), .C(n6420) );
  CKBD0 U6302 ( .CLK(n6420), .C(n6421) );
  CKBD0 U6303 ( .CLK(n6421), .C(n6422) );
  CKBD0 U6304 ( .CLK(n6422), .C(n6423) );
  CKBD0 U6305 ( .CLK(n6423), .C(n6424) );
  CKBD0 U6306 ( .CLK(n6424), .C(n6425) );
  CKBD0 U6307 ( .CLK(n6425), .C(n6426) );
  BUFFD0 U6308 ( .I(n6426), .Z(n6427) );
  CKBD0 U6309 ( .CLK(n6427), .C(n6428) );
  CKBD0 U6310 ( .CLK(n6428), .C(n6429) );
  CKBD0 U6311 ( .CLK(n6429), .C(n6430) );
  CKBD0 U6312 ( .CLK(n6430), .C(n6431) );
  CKBD0 U6313 ( .CLK(n6431), .C(n6432) );
  CKBD0 U6314 ( .CLK(n6432), .C(n6433) );
  CKBD0 U6315 ( .CLK(n6433), .C(n6434) );
  CKBD0 U6316 ( .CLK(n6434), .C(n6435) );
  CKBD0 U6317 ( .CLK(n6435), .C(n6436) );
  CKBD0 U6318 ( .CLK(n6436), .C(n6437) );
  BUFFD0 U6319 ( .I(n6437), .Z(n6438) );
  CKBD0 U6320 ( .CLK(n6438), .C(n6439) );
  CKBD0 U6321 ( .CLK(n6439), .C(n6440) );
  CKBD0 U6322 ( .CLK(n6440), .C(n6441) );
  CKBD0 U6323 ( .CLK(n6441), .C(n6442) );
  CKBD0 U6324 ( .CLK(n6442), .C(n6443) );
  CKBD0 U6325 ( .CLK(n6443), .C(n6444) );
  CKBD0 U6326 ( .CLK(n6444), .C(n6445) );
  CKBD0 U6327 ( .CLK(n6445), .C(n6446) );
  CKBD0 U6328 ( .CLK(n6446), .C(n6447) );
  BUFFD0 U6329 ( .I(n6447), .Z(n6448) );
  CKBD0 U6330 ( .CLK(n6448), .C(n6449) );
  CKBD0 U6331 ( .CLK(n6449), .C(n6450) );
  CKBD0 U6332 ( .CLK(n6450), .C(n6451) );
  CKBD0 U6333 ( .CLK(n6451), .C(n6452) );
  CKBD0 U6334 ( .CLK(n6452), .C(n6453) );
  CKBD0 U6335 ( .CLK(n6453), .C(n6454) );
  CKBD0 U6336 ( .CLK(n6454), .C(n6455) );
  CKBD0 U6337 ( .CLK(n6455), .C(n6456) );
  CKBD0 U6338 ( .CLK(n6456), .C(n6457) );
  CKBD0 U6339 ( .CLK(n6457), .C(n6458) );
  BUFFD0 U6340 ( .I(n6458), .Z(n6459) );
  CKBD0 U6341 ( .CLK(n6459), .C(n6460) );
  CKBD0 U6342 ( .CLK(n6460), .C(n6461) );
  CKBD0 U6343 ( .CLK(n6461), .C(n6462) );
  CKBD0 U6344 ( .CLK(n6462), .C(n6463) );
  CKBD0 U6345 ( .CLK(n6463), .C(n6464) );
  CKBD0 U6346 ( .CLK(n6464), .C(n6465) );
  BUFFD0 U6347 ( .I(n6465), .Z(n6466) );
  CKBD0 U6348 ( .CLK(n6466), .C(n6467) );
  BUFFD0 U6349 ( .I(n6467), .Z(n6468) );
  CKBD0 U6350 ( .CLK(n6468), .C(n6469) );
  BUFFD0 U6351 ( .I(n6469), .Z(n6470) );
  CKBD0 U6352 ( .CLK(n6470), .C(n6471) );
  BUFFD0 U6353 ( .I(n6471), .Z(n6472) );
  CKBD0 U6354 ( .CLK(n6472), .C(n6473) );
  BUFFD0 U6355 ( .I(n6473), .Z(n6474) );
  CKBD0 U6356 ( .CLK(n6474), .C(n6475) );
  BUFFD0 U6357 ( .I(n6475), .Z(n6476) );
  CKBD0 U6358 ( .CLK(n6476), .C(n6477) );
  BUFFD0 U6359 ( .I(n6477), .Z(n6478) );
  CKBD0 U6360 ( .CLK(n6478), .C(n6479) );
  BUFFD0 U6361 ( .I(n6479), .Z(n6480) );
  BUFFD0 U6362 ( .I(n135), .Z(n6481) );
  BUFFD0 U6363 ( .I(n6483), .Z(n6482) );
  BUFFD0 U6364 ( .I(n6484), .Z(n6483) );
  BUFFD0 U6365 ( .I(Decoder[2]), .Z(n6484) );
  CKBD0 U6366 ( .CLK(n917), .C(n6485) );
  CKBD0 U6367 ( .CLK(n6485), .C(n6486) );
  CKBD0 U6368 ( .CLK(n6486), .C(n6487) );
  BUFFD0 U6369 ( .I(n6487), .Z(n6488) );
  CKBD0 U6370 ( .CLK(n6488), .C(n6489) );
  CKBD0 U6371 ( .CLK(n6489), .C(n6490) );
  CKBD0 U6372 ( .CLK(n6490), .C(n6491) );
  CKBD0 U6373 ( .CLK(n6491), .C(n6492) );
  CKBD0 U6374 ( .CLK(n6492), .C(n6493) );
  CKBD0 U6375 ( .CLK(n6493), .C(n6494) );
  CKBD0 U6376 ( .CLK(n6494), .C(n6495) );
  CKBD0 U6377 ( .CLK(n6495), .C(n6496) );
  CKBD0 U6378 ( .CLK(n6496), .C(n6497) );
  CKBD0 U6379 ( .CLK(n6497), .C(n6498) );
  BUFFD0 U6380 ( .I(n6498), .Z(n6499) );
  CKBD0 U6381 ( .CLK(n6499), .C(n6500) );
  CKBD0 U6382 ( .CLK(n6500), .C(n6501) );
  CKBD0 U6383 ( .CLK(n6501), .C(n6502) );
  CKBD0 U6384 ( .CLK(n6502), .C(n6503) );
  CKBD0 U6385 ( .CLK(n6503), .C(n6504) );
  CKBD0 U6386 ( .CLK(n6504), .C(n6505) );
  CKBD0 U6387 ( .CLK(n6505), .C(n6506) );
  CKBD0 U6388 ( .CLK(n6506), .C(n6507) );
  CKBD0 U6389 ( .CLK(n6507), .C(n6508) );
  BUFFD0 U6390 ( .I(n6508), .Z(n6509) );
  CKBD0 U6391 ( .CLK(n6509), .C(n6510) );
  CKBD0 U6392 ( .CLK(n6510), .C(n6511) );
  CKBD0 U6393 ( .CLK(n6511), .C(n6512) );
  CKBD0 U6394 ( .CLK(n6512), .C(n6513) );
  CKBD0 U6395 ( .CLK(n6513), .C(n6514) );
  CKBD0 U6396 ( .CLK(n6514), .C(n6515) );
  CKBD0 U6397 ( .CLK(n6515), .C(n6516) );
  CKBD0 U6398 ( .CLK(n6516), .C(n6517) );
  CKBD0 U6399 ( .CLK(n6517), .C(n6518) );
  CKBD0 U6400 ( .CLK(n6518), .C(n6519) );
  BUFFD0 U6401 ( .I(n6519), .Z(n6520) );
  CKBD0 U6402 ( .CLK(n6520), .C(n6521) );
  CKBD0 U6403 ( .CLK(n6521), .C(n6522) );
  CKBD0 U6404 ( .CLK(n6522), .C(n6523) );
  CKBD0 U6405 ( .CLK(n6523), .C(n6524) );
  CKBD0 U6406 ( .CLK(n6524), .C(n6525) );
  CKBD0 U6407 ( .CLK(n6525), .C(n6526) );
  CKBD0 U6408 ( .CLK(n6526), .C(n6527) );
  CKBD0 U6409 ( .CLK(n6527), .C(n6528) );
  CKBD0 U6410 ( .CLK(n6528), .C(n6529) );
  CKBD0 U6411 ( .CLK(n6529), .C(n6530) );
  BUFFD0 U6412 ( .I(n6530), .Z(n6531) );
  CKBD0 U6413 ( .CLK(n6531), .C(n6532) );
  CKBD0 U6414 ( .CLK(n6532), .C(n6533) );
  CKBD0 U6415 ( .CLK(n6533), .C(n6534) );
  CKBD0 U6416 ( .CLK(n6534), .C(n6535) );
  CKBD0 U6417 ( .CLK(n6535), .C(n6536) );
  CKBD0 U6418 ( .CLK(n6536), .C(n6537) );
  CKBD0 U6419 ( .CLK(n6537), .C(n6538) );
  CKBD0 U6420 ( .CLK(n6538), .C(n6539) );
  CKBD0 U6421 ( .CLK(n6539), .C(n6540) );
  CKBD0 U6422 ( .CLK(n6540), .C(n6541) );
  BUFFD0 U6423 ( .I(n6541), .Z(n6542) );
  CKBD0 U6424 ( .CLK(n6542), .C(n6543) );
  CKBD0 U6425 ( .CLK(n6543), .C(n6544) );
  CKBD0 U6426 ( .CLK(n6544), .C(n6545) );
  CKBD0 U6427 ( .CLK(n6545), .C(n6546) );
  CKBD0 U6428 ( .CLK(n6546), .C(n6547) );
  CKBD0 U6429 ( .CLK(n6547), .C(n6548) );
  CKBD0 U6430 ( .CLK(n6548), .C(n6549) );
  CKBD0 U6431 ( .CLK(n6549), .C(n6550) );
  CKBD0 U6432 ( .CLK(n6550), .C(n6551) );
  CKBD0 U6433 ( .CLK(n6551), .C(n6552) );
  BUFFD0 U6434 ( .I(n6552), .Z(n6553) );
  CKBD0 U6435 ( .CLK(n6553), .C(n6554) );
  CKBD0 U6436 ( .CLK(n6554), .C(n6555) );
  CKBD0 U6437 ( .CLK(n6555), .C(n6556) );
  CKBD0 U6438 ( .CLK(n6556), .C(n6557) );
  CKBD0 U6439 ( .CLK(n6557), .C(n6558) );
  CKBD0 U6440 ( .CLK(n6558), .C(n6559) );
  CKBD0 U6441 ( .CLK(n6559), .C(n6560) );
  CKBD0 U6442 ( .CLK(n6560), .C(n6561) );
  CKBD0 U6443 ( .CLK(n6561), .C(n6562) );
  CKBD0 U6444 ( .CLK(n6562), .C(n6563) );
  BUFFD0 U6445 ( .I(n6563), .Z(n6564) );
  CKBD0 U6446 ( .CLK(n6564), .C(n6565) );
  CKBD0 U6447 ( .CLK(n6565), .C(n6566) );
  CKBD0 U6448 ( .CLK(n6566), .C(n6567) );
  CKBD0 U6449 ( .CLK(n6567), .C(n6568) );
  CKBD0 U6450 ( .CLK(n6568), .C(n6569) );
  CKBD0 U6451 ( .CLK(n6569), .C(n6570) );
  CKBD0 U6452 ( .CLK(n6570), .C(n6571) );
  CKBD0 U6453 ( .CLK(n6571), .C(n6572) );
  CKBD0 U6454 ( .CLK(n6572), .C(n6573) );
  BUFFD0 U6455 ( .I(n6573), .Z(n6574) );
  CKBD0 U6456 ( .CLK(n6574), .C(n6575) );
  CKBD0 U6457 ( .CLK(n6575), .C(n6576) );
  CKBD0 U6458 ( .CLK(n6576), .C(n6577) );
  CKBD0 U6459 ( .CLK(n6577), .C(n6578) );
  CKBD0 U6460 ( .CLK(n6578), .C(n6579) );
  CKBD0 U6461 ( .CLK(n6579), .C(n6580) );
  CKBD0 U6462 ( .CLK(n6580), .C(n6581) );
  CKBD0 U6463 ( .CLK(n6581), .C(n6582) );
  CKBD0 U6464 ( .CLK(n6582), .C(n6583) );
  CKBD0 U6465 ( .CLK(n6583), .C(n6584) );
  BUFFD0 U6466 ( .I(n6584), .Z(n6585) );
  CKBD0 U6467 ( .CLK(n6585), .C(n6586) );
  CKBD0 U6468 ( .CLK(n6586), .C(n6587) );
  CKBD0 U6469 ( .CLK(n6587), .C(n6588) );
  CKBD0 U6470 ( .CLK(n6588), .C(n6589) );
  CKBD0 U6471 ( .CLK(n6589), .C(n6590) );
  CKBD0 U6472 ( .CLK(n6590), .C(n6591) );
  CKBD0 U6473 ( .CLK(n6591), .C(n6592) );
  CKBD0 U6474 ( .CLK(n6592), .C(n6593) );
  CKBD0 U6475 ( .CLK(n6593), .C(n6594) );
  CKBD0 U6476 ( .CLK(n6594), .C(n6595) );
  BUFFD0 U6477 ( .I(n6595), .Z(n6596) );
  CKBD0 U6478 ( .CLK(n6596), .C(n6597) );
  CKBD0 U6479 ( .CLK(n6597), .C(n6598) );
  CKBD0 U6480 ( .CLK(n6598), .C(n6599) );
  CKBD0 U6481 ( .CLK(n6599), .C(n6600) );
  CKBD0 U6482 ( .CLK(n6600), .C(n6601) );
  CKBD0 U6483 ( .CLK(n6601), .C(n6602) );
  BUFFD0 U6484 ( .I(n6602), .Z(n6603) );
  CKBD0 U6485 ( .CLK(n6603), .C(n6604) );
  BUFFD0 U6486 ( .I(n6604), .Z(n6605) );
  CKBD0 U6487 ( .CLK(n6605), .C(n6606) );
  BUFFD0 U6488 ( .I(n6606), .Z(n6607) );
  CKBD0 U6489 ( .CLK(n6607), .C(n6608) );
  BUFFD0 U6490 ( .I(n6608), .Z(n6609) );
  CKBD0 U6491 ( .CLK(n6609), .C(n6610) );
  BUFFD0 U6492 ( .I(n6610), .Z(n6611) );
  CKBD0 U6493 ( .CLK(n6611), .C(n6612) );
  BUFFD0 U6494 ( .I(n6612), .Z(n6613) );
  CKBD0 U6495 ( .CLK(n6613), .C(n6614) );
  BUFFD0 U6496 ( .I(n6614), .Z(n6615) );
  CKBD0 U6497 ( .CLK(n6615), .C(n6616) );
  BUFFD0 U6498 ( .I(n6616), .Z(n6617) );
  BUFFD0 U6499 ( .I(n134), .Z(n6618) );
  BUFFD0 U6500 ( .I(n6620), .Z(n6619) );
  BUFFD0 U6501 ( .I(n6621), .Z(n6620) );
  BUFFD0 U6502 ( .I(Decoder[1]), .Z(n6621) );
  CKBD0 U6503 ( .CLK(n915), .C(n6622) );
  CKBD0 U6504 ( .CLK(n6622), .C(n6623) );
  CKBD0 U6505 ( .CLK(n6623), .C(n6624) );
  BUFFD0 U6506 ( .I(n6624), .Z(n6625) );
  CKBD0 U6507 ( .CLK(n6625), .C(n6626) );
  CKBD0 U6508 ( .CLK(n6626), .C(n6627) );
  CKBD0 U6509 ( .CLK(n6627), .C(n6628) );
  CKBD0 U6510 ( .CLK(n6628), .C(n6629) );
  CKBD0 U6511 ( .CLK(n6629), .C(n6630) );
  CKBD0 U6512 ( .CLK(n6630), .C(n6631) );
  CKBD0 U6513 ( .CLK(n6631), .C(n6632) );
  CKBD0 U6514 ( .CLK(n6632), .C(n6633) );
  CKBD0 U6515 ( .CLK(n6633), .C(n6634) );
  BUFFD0 U6516 ( .I(n6634), .Z(n6635) );
  CKBD0 U6517 ( .CLK(n6635), .C(n6636) );
  CKBD0 U6518 ( .CLK(n6636), .C(n6637) );
  CKBD0 U6519 ( .CLK(n6637), .C(n6638) );
  CKBD0 U6520 ( .CLK(n6638), .C(n6639) );
  CKBD0 U6521 ( .CLK(n6639), .C(n6640) );
  CKBD0 U6522 ( .CLK(n6640), .C(n6641) );
  CKBD0 U6523 ( .CLK(n6641), .C(n6642) );
  CKBD0 U6524 ( .CLK(n6642), .C(n6643) );
  CKBD0 U6525 ( .CLK(n6643), .C(n6644) );
  CKBD0 U6526 ( .CLK(n6644), .C(n6645) );
  BUFFD0 U6527 ( .I(n6645), .Z(n6646) );
  CKBD0 U6528 ( .CLK(n6646), .C(n6647) );
  CKBD0 U6529 ( .CLK(n6647), .C(n6648) );
  CKBD0 U6530 ( .CLK(n6648), .C(n6649) );
  CKBD0 U6531 ( .CLK(n6649), .C(n6650) );
  CKBD0 U6532 ( .CLK(n6650), .C(n6651) );
  CKBD0 U6533 ( .CLK(n6651), .C(n6652) );
  CKBD0 U6534 ( .CLK(n6652), .C(n6653) );
  CKBD0 U6535 ( .CLK(n6653), .C(n6654) );
  CKBD0 U6536 ( .CLK(n6654), .C(n6655) );
  CKBD0 U6537 ( .CLK(n6655), .C(n6656) );
  BUFFD0 U6538 ( .I(n6656), .Z(n6657) );
  CKBD0 U6539 ( .CLK(n6657), .C(n6658) );
  CKBD0 U6540 ( .CLK(n6658), .C(n6659) );
  CKBD0 U6541 ( .CLK(n6659), .C(n6660) );
  CKBD0 U6542 ( .CLK(n6660), .C(n6661) );
  CKBD0 U6543 ( .CLK(n6661), .C(n6662) );
  CKBD0 U6544 ( .CLK(n6662), .C(n6663) );
  CKBD0 U6545 ( .CLK(n6663), .C(n6664) );
  CKBD0 U6546 ( .CLK(n6664), .C(n6665) );
  CKBD0 U6547 ( .CLK(n6665), .C(n6666) );
  CKBD0 U6548 ( .CLK(n6666), .C(n6667) );
  BUFFD0 U6549 ( .I(n6667), .Z(n6668) );
  CKBD0 U6550 ( .CLK(n6668), .C(n6669) );
  CKBD0 U6551 ( .CLK(n6669), .C(n6670) );
  CKBD0 U6552 ( .CLK(n6670), .C(n6671) );
  CKBD0 U6553 ( .CLK(n6671), .C(n6672) );
  CKBD0 U6554 ( .CLK(n6672), .C(n6673) );
  CKBD0 U6555 ( .CLK(n6673), .C(n6674) );
  CKBD0 U6556 ( .CLK(n6674), .C(n6675) );
  CKBD0 U6557 ( .CLK(n6675), .C(n6676) );
  CKBD0 U6558 ( .CLK(n6676), .C(n6677) );
  CKBD0 U6559 ( .CLK(n6677), .C(n6678) );
  BUFFD0 U6560 ( .I(n6678), .Z(n6679) );
  CKBD0 U6561 ( .CLK(n6679), .C(n6680) );
  CKBD0 U6562 ( .CLK(n6680), .C(n6681) );
  CKBD0 U6563 ( .CLK(n6681), .C(n6682) );
  CKBD0 U6564 ( .CLK(n6682), .C(n6683) );
  CKBD0 U6565 ( .CLK(n6683), .C(n6684) );
  CKBD0 U6566 ( .CLK(n6684), .C(n6685) );
  CKBD0 U6567 ( .CLK(n6685), .C(n6686) );
  CKBD0 U6568 ( .CLK(n6686), .C(n6687) );
  CKBD0 U6569 ( .CLK(n6687), .C(n6688) );
  CKBD0 U6570 ( .CLK(n6688), .C(n6689) );
  BUFFD0 U6571 ( .I(n6689), .Z(n6690) );
  CKBD0 U6572 ( .CLK(n6690), .C(n6691) );
  CKBD0 U6573 ( .CLK(n6691), .C(n6692) );
  CKBD0 U6574 ( .CLK(n6692), .C(n6693) );
  CKBD0 U6575 ( .CLK(n6693), .C(n6694) );
  CKBD0 U6576 ( .CLK(n6694), .C(n6695) );
  CKBD0 U6577 ( .CLK(n6695), .C(n6696) );
  CKBD0 U6578 ( .CLK(n6696), .C(n6697) );
  CKBD0 U6579 ( .CLK(n6697), .C(n6698) );
  CKBD0 U6580 ( .CLK(n6698), .C(n6699) );
  CKBD0 U6581 ( .CLK(n6699), .C(n6700) );
  BUFFD0 U6582 ( .I(n6700), .Z(n6701) );
  CKBD0 U6583 ( .CLK(n6701), .C(n6702) );
  CKBD0 U6584 ( .CLK(n6702), .C(n6703) );
  CKBD0 U6585 ( .CLK(n6703), .C(n6704) );
  CKBD0 U6586 ( .CLK(n6704), .C(n6705) );
  CKBD0 U6587 ( .CLK(n6705), .C(n6706) );
  CKBD0 U6588 ( .CLK(n6706), .C(n6707) );
  CKBD0 U6589 ( .CLK(n6707), .C(n6708) );
  CKBD0 U6590 ( .CLK(n6708), .C(n6709) );
  CKBD0 U6591 ( .CLK(n6709), .C(n6710) );
  BUFFD0 U6592 ( .I(n6710), .Z(n6711) );
  CKBD0 U6593 ( .CLK(n6711), .C(n6712) );
  CKBD0 U6594 ( .CLK(n6712), .C(n6713) );
  CKBD0 U6595 ( .CLK(n6713), .C(n6714) );
  CKBD0 U6596 ( .CLK(n6714), .C(n6715) );
  CKBD0 U6597 ( .CLK(n6715), .C(n6716) );
  CKBD0 U6598 ( .CLK(n6716), .C(n6717) );
  CKBD0 U6599 ( .CLK(n6717), .C(n6718) );
  CKBD0 U6600 ( .CLK(n6718), .C(n6719) );
  CKBD0 U6601 ( .CLK(n6719), .C(n6720) );
  CKBD0 U6602 ( .CLK(n6720), .C(n6721) );
  BUFFD0 U6603 ( .I(n6721), .Z(n6722) );
  CKBD0 U6604 ( .CLK(n6722), .C(n6723) );
  CKBD0 U6605 ( .CLK(n6723), .C(n6724) );
  CKBD0 U6606 ( .CLK(n6724), .C(n6725) );
  CKBD0 U6607 ( .CLK(n6725), .C(n6726) );
  CKBD0 U6608 ( .CLK(n6726), .C(n6727) );
  CKBD0 U6609 ( .CLK(n6727), .C(n6728) );
  CKBD0 U6610 ( .CLK(n6728), .C(n6729) );
  CKBD0 U6611 ( .CLK(n6729), .C(n6730) );
  CKBD0 U6612 ( .CLK(n6730), .C(n6731) );
  CKBD0 U6613 ( .CLK(n6731), .C(n6732) );
  BUFFD0 U6614 ( .I(n6732), .Z(n6733) );
  CKBD0 U6615 ( .CLK(n6733), .C(n6734) );
  CKBD0 U6616 ( .CLK(n6734), .C(n6735) );
  CKBD0 U6617 ( .CLK(n6735), .C(n6736) );
  CKBD0 U6618 ( .CLK(n6736), .C(n6737) );
  CKBD0 U6619 ( .CLK(n6737), .C(n6738) );
  CKBD0 U6620 ( .CLK(n6738), .C(n6739) );
  BUFFD0 U6621 ( .I(n6739), .Z(n6740) );
  CKBD0 U6622 ( .CLK(n6740), .C(n6741) );
  BUFFD0 U6623 ( .I(n6741), .Z(n6742) );
  CKBD0 U6624 ( .CLK(n6742), .C(n6743) );
  BUFFD0 U6625 ( .I(n6743), .Z(n6744) );
  CKBD0 U6626 ( .CLK(n6744), .C(n6745) );
  BUFFD0 U6627 ( .I(n6745), .Z(n6746) );
  CKBD0 U6628 ( .CLK(n6746), .C(n6747) );
  BUFFD0 U6629 ( .I(n6747), .Z(n6748) );
  CKBD0 U6630 ( .CLK(n6748), .C(n6749) );
  BUFFD0 U6631 ( .I(n6749), .Z(n6750) );
  CKBD0 U6632 ( .CLK(n6750), .C(n6751) );
  BUFFD0 U6633 ( .I(n6751), .Z(n6752) );
  CKBD0 U6634 ( .CLK(n6752), .C(n6753) );
  BUFFD0 U6635 ( .I(n6753), .Z(n6754) );
  BUFFD0 U6636 ( .I(n133), .Z(n6755) );
  BUFFD0 U6637 ( .I(n6757), .Z(n6756) );
  BUFFD0 U6638 ( .I(n6758), .Z(n6757) );
  BUFFD0 U6639 ( .I(Decoder[0]), .Z(n6758) );
  CKBD0 U6640 ( .CLK(n913), .C(n6759) );
  CKBD0 U6641 ( .CLK(n6759), .C(n6760) );
  CKBD0 U6642 ( .CLK(n6760), .C(n6761) );
  BUFFD0 U6643 ( .I(n6761), .Z(n6762) );
  CKBD0 U6644 ( .CLK(n6762), .C(n6763) );
  CKBD0 U6645 ( .CLK(n6763), .C(n6764) );
  CKBD0 U6646 ( .CLK(n6764), .C(n6765) );
  CKBD0 U6647 ( .CLK(n6765), .C(n6766) );
  CKBD0 U6648 ( .CLK(n6766), .C(n6767) );
  CKBD0 U6649 ( .CLK(n6767), .C(n6768) );
  CKBD0 U6650 ( .CLK(n6768), .C(n6769) );
  CKBD0 U6651 ( .CLK(n6769), .C(n6770) );
  CKBD0 U6652 ( .CLK(n6770), .C(n6771) );
  CKBD0 U6653 ( .CLK(n6771), .C(n6772) );
  BUFFD0 U6654 ( .I(n6772), .Z(n6773) );
  CKBD0 U6655 ( .CLK(n6773), .C(n6774) );
  CKBD0 U6656 ( .CLK(n6774), .C(n6775) );
  CKBD0 U6657 ( .CLK(n6775), .C(n6776) );
  CKBD0 U6658 ( .CLK(n6776), .C(n6777) );
  CKBD0 U6659 ( .CLK(n6777), .C(n6778) );
  CKBD0 U6660 ( .CLK(n6778), .C(n6779) );
  CKBD0 U6661 ( .CLK(n6779), .C(n6780) );
  CKBD0 U6662 ( .CLK(n6780), .C(n6781) );
  CKBD0 U6663 ( .CLK(n6781), .C(n6782) );
  BUFFD0 U6664 ( .I(n6782), .Z(n6783) );
  CKBD0 U6665 ( .CLK(n6783), .C(n6784) );
  CKBD0 U6666 ( .CLK(n6784), .C(n6785) );
  CKBD0 U6667 ( .CLK(n6785), .C(n6786) );
  CKBD0 U6668 ( .CLK(n6786), .C(n6787) );
  CKBD0 U6669 ( .CLK(n6787), .C(n6788) );
  CKBD0 U6670 ( .CLK(n6788), .C(n6789) );
  CKBD0 U6671 ( .CLK(n6789), .C(n6790) );
  CKBD0 U6672 ( .CLK(n6790), .C(n6791) );
  CKBD0 U6673 ( .CLK(n6791), .C(n6792) );
  CKBD0 U6674 ( .CLK(n6792), .C(n6793) );
  BUFFD0 U6675 ( .I(n6793), .Z(n6794) );
  CKBD0 U6676 ( .CLK(n6794), .C(n6795) );
  CKBD0 U6677 ( .CLK(n6795), .C(n6796) );
  CKBD0 U6678 ( .CLK(n6796), .C(n6797) );
  CKBD0 U6679 ( .CLK(n6797), .C(n6798) );
  CKBD0 U6680 ( .CLK(n6798), .C(n6799) );
  CKBD0 U6681 ( .CLK(n6799), .C(n6800) );
  CKBD0 U6682 ( .CLK(n6800), .C(n6801) );
  CKBD0 U6683 ( .CLK(n6801), .C(n6802) );
  CKBD0 U6684 ( .CLK(n6802), .C(n6803) );
  CKBD0 U6685 ( .CLK(n6803), .C(n6804) );
  BUFFD0 U6686 ( .I(n6804), .Z(n6805) );
  CKBD0 U6687 ( .CLK(n6805), .C(n6806) );
  CKBD0 U6688 ( .CLK(n6806), .C(n6807) );
  CKBD0 U6689 ( .CLK(n6807), .C(n6808) );
  CKBD0 U6690 ( .CLK(n6808), .C(n6809) );
  CKBD0 U6691 ( .CLK(n6809), .C(n6810) );
  CKBD0 U6692 ( .CLK(n6810), .C(n6811) );
  CKBD0 U6693 ( .CLK(n6811), .C(n6812) );
  CKBD0 U6694 ( .CLK(n6812), .C(n6813) );
  CKBD0 U6695 ( .CLK(n6813), .C(n6814) );
  CKBD0 U6696 ( .CLK(n6814), .C(n6815) );
  BUFFD0 U6697 ( .I(n6815), .Z(n6816) );
  CKBD0 U6698 ( .CLK(n6816), .C(n6817) );
  CKBD0 U6699 ( .CLK(n6817), .C(n6818) );
  CKBD0 U6700 ( .CLK(n6818), .C(n6819) );
  CKBD0 U6701 ( .CLK(n6819), .C(n6820) );
  CKBD0 U6702 ( .CLK(n6820), .C(n6821) );
  CKBD0 U6703 ( .CLK(n6821), .C(n6822) );
  CKBD0 U6704 ( .CLK(n6822), .C(n6823) );
  CKBD0 U6705 ( .CLK(n6823), .C(n6824) );
  CKBD0 U6706 ( .CLK(n6824), .C(n6825) );
  CKBD0 U6707 ( .CLK(n6825), .C(n6826) );
  BUFFD0 U6708 ( .I(n6826), .Z(n6827) );
  CKBD0 U6709 ( .CLK(n6827), .C(n6828) );
  CKBD0 U6710 ( .CLK(n6828), .C(n6829) );
  CKBD0 U6711 ( .CLK(n6829), .C(n6830) );
  CKBD0 U6712 ( .CLK(n6830), .C(n6831) );
  CKBD0 U6713 ( .CLK(n6831), .C(n6832) );
  CKBD0 U6714 ( .CLK(n6832), .C(n6833) );
  CKBD0 U6715 ( .CLK(n6833), .C(n6834) );
  CKBD0 U6716 ( .CLK(n6834), .C(n6835) );
  CKBD0 U6717 ( .CLK(n6835), .C(n6836) );
  CKBD0 U6718 ( .CLK(n6836), .C(n6837) );
  BUFFD0 U6719 ( .I(n6837), .Z(n6838) );
  CKBD0 U6720 ( .CLK(n6838), .C(n6839) );
  CKBD0 U6721 ( .CLK(n6839), .C(n6840) );
  CKBD0 U6722 ( .CLK(n6840), .C(n6841) );
  CKBD0 U6723 ( .CLK(n6841), .C(n6842) );
  CKBD0 U6724 ( .CLK(n6842), .C(n6843) );
  CKBD0 U6725 ( .CLK(n6843), .C(n6844) );
  CKBD0 U6726 ( .CLK(n6844), .C(n6845) );
  CKBD0 U6727 ( .CLK(n6845), .C(n6846) );
  CKBD0 U6728 ( .CLK(n6846), .C(n6847) );
  BUFFD0 U6729 ( .I(n6847), .Z(n6848) );
  CKBD0 U6730 ( .CLK(n6848), .C(n6849) );
  CKBD0 U6731 ( .CLK(n6849), .C(n6850) );
  CKBD0 U6732 ( .CLK(n6850), .C(n6851) );
  CKBD0 U6733 ( .CLK(n6851), .C(n6852) );
  CKBD0 U6734 ( .CLK(n6852), .C(n6853) );
  CKBD0 U6735 ( .CLK(n6853), .C(n6854) );
  CKBD0 U6736 ( .CLK(n6854), .C(n6855) );
  CKBD0 U6737 ( .CLK(n6855), .C(n6856) );
  CKBD0 U6738 ( .CLK(n6856), .C(n6857) );
  CKBD0 U6739 ( .CLK(n6857), .C(n6858) );
  BUFFD0 U6740 ( .I(n6858), .Z(n6859) );
  CKBD0 U6741 ( .CLK(n6859), .C(n6860) );
  CKBD0 U6742 ( .CLK(n6860), .C(n6861) );
  CKBD0 U6743 ( .CLK(n6861), .C(n6862) );
  CKBD0 U6744 ( .CLK(n6862), .C(n6863) );
  CKBD0 U6745 ( .CLK(n6863), .C(n6864) );
  CKBD0 U6746 ( .CLK(n6864), .C(n6865) );
  CKBD0 U6747 ( .CLK(n6865), .C(n6866) );
  CKBD0 U6748 ( .CLK(n6866), .C(n6867) );
  CKBD0 U6749 ( .CLK(n6867), .C(n6868) );
  CKBD0 U6750 ( .CLK(n6868), .C(n6869) );
  BUFFD0 U6751 ( .I(n6869), .Z(n6870) );
  CKBD0 U6752 ( .CLK(n6870), .C(n6871) );
  CKBD0 U6753 ( .CLK(n6871), .C(n6872) );
  CKBD0 U6754 ( .CLK(n6872), .C(n6873) );
  CKBD0 U6755 ( .CLK(n6873), .C(n6874) );
  CKBD0 U6756 ( .CLK(n6874), .C(n6875) );
  CKBD0 U6757 ( .CLK(n6875), .C(n6876) );
  BUFFD0 U6758 ( .I(n6876), .Z(n6877) );
  CKBD0 U6759 ( .CLK(n6877), .C(n6878) );
  BUFFD0 U6760 ( .I(n6878), .Z(n6879) );
  CKBD0 U6761 ( .CLK(n6879), .C(n6880) );
  BUFFD0 U6762 ( .I(n6880), .Z(n6881) );
  CKBD0 U6763 ( .CLK(n6881), .C(n6882) );
  BUFFD0 U6764 ( .I(n6882), .Z(n6883) );
  CKBD0 U6765 ( .CLK(n6883), .C(n6884) );
  BUFFD0 U6766 ( .I(n6884), .Z(n6885) );
  CKBD0 U6767 ( .CLK(n6885), .C(n6886) );
  BUFFD0 U6768 ( .I(n6886), .Z(n6887) );
  CKBD0 U6769 ( .CLK(n6887), .C(n6888) );
  BUFFD0 U6770 ( .I(n6888), .Z(n6889) );
  CKBD0 U6771 ( .CLK(n6889), .C(n6890) );
  BUFFD0 U6772 ( .I(n6890), .Z(n6891) );
  BUFFD0 U6773 ( .I(n6893), .Z(n6892) );
  BUFFD0 U6774 ( .I(n99), .Z(n6893) );
  CKND2D0 U6775 ( .A1(n232), .A2(ParValidTimer[0]), .ZN(n10) );
  XOR2D0 U6776 ( .A1(n9021), .A2(n10), .Z(n11) );
  BUFFD0 U6777 ( .I(N39), .Z(n6894) );
  CKBD0 U6778 ( .CLK(Count32[0]), .C(n6903) );
  BUFFD0 U6779 ( .I(Count32[1]), .Z(n6895) );
  BUFFD0 U6780 ( .I(n100), .Z(n6896) );
  BUFFD0 U6781 ( .I(n12), .Z(n6897) );
  CKXOR2D0 U6782 ( .A1(n232), .A2(n6), .Z(n12) );
  BUFFD0 U6783 ( .I(n6899), .Z(n6898) );
  BUFFD0 U6784 ( .I(N41), .Z(n6899) );
  BUFFD0 U6785 ( .I(n6901), .Z(n6900) );
  BUFFD0 U6786 ( .I(N40), .Z(n6901) );
  BUFFD0 U6787 ( .I(N38), .Z(n6902) );
  BUFFD0 U6788 ( .I(n6905), .Z(n6904) );
  BUFFD0 U6789 ( .I(n6906), .Z(n6905) );
  BUFFD0 U6790 ( .I(n6907), .Z(n6906) );
  BUFFD0 U6791 ( .I(n132), .Z(n6907) );
  IOA22D0 U6792 ( .B1(n9128), .B2(n63), .A1(n1), .A2(Decoder[0]), .ZN(n132) );
  BUFFD0 U6793 ( .I(n6909), .Z(n6908) );
  BUFFD0 U6794 ( .I(n6910), .Z(n6909) );
  BUFFD0 U6795 ( .I(n6911), .Z(n6910) );
  BUFFD0 U6796 ( .I(n131), .Z(n6911) );
  IOA22D0 U6797 ( .B1(n9127), .B2(n62), .A1(n1), .A2(Decoder[1]), .ZN(n131) );
  BUFFD0 U6798 ( .I(n6913), .Z(n6912) );
  BUFFD0 U6799 ( .I(n6914), .Z(n6913) );
  BUFFD0 U6800 ( .I(n6915), .Z(n6914) );
  BUFFD0 U6801 ( .I(n130), .Z(n6915) );
  IOA22D0 U6802 ( .B1(n9127), .B2(n61), .A1(n1), .A2(Decoder[2]), .ZN(n130) );
  BUFFD0 U6803 ( .I(n6917), .Z(n6916) );
  BUFFD0 U6804 ( .I(n6918), .Z(n6917) );
  BUFFD0 U6805 ( .I(n6919), .Z(n6918) );
  BUFFD0 U6806 ( .I(n129), .Z(n6919) );
  IOA22D0 U6807 ( .B1(n9127), .B2(n60), .A1(n1), .A2(Decoder[3]), .ZN(n129) );
  BUFFD0 U6808 ( .I(n6921), .Z(n6920) );
  BUFFD0 U6809 ( .I(n6922), .Z(n6921) );
  BUFFD0 U6810 ( .I(n6923), .Z(n6922) );
  BUFFD0 U6811 ( .I(n128), .Z(n6923) );
  IOA22D0 U6812 ( .B1(n9127), .B2(n59), .A1(n1), .A2(Decoder[4]), .ZN(n128) );
  BUFFD0 U6813 ( .I(n6925), .Z(n6924) );
  BUFFD0 U6814 ( .I(n6926), .Z(n6925) );
  BUFFD0 U6815 ( .I(n6927), .Z(n6926) );
  BUFFD0 U6816 ( .I(n127), .Z(n6927) );
  IOA22D0 U6817 ( .B1(n9127), .B2(n58), .A1(n1), .A2(Decoder[5]), .ZN(n127) );
  CKBD0 U6818 ( .CLK(n126), .C(n6931) );
  MOAI22D1 U6819 ( .A1(n9127), .A2(n57), .B1(n9129), .B2(Decoder[6]), .ZN(n126) );
  BUFFD0 U6820 ( .I(n6929), .Z(n6928) );
  BUFFD0 U6821 ( .I(n6930), .Z(n6929) );
  BUFFD0 U6822 ( .I(n6931), .Z(n6930) );
  IOA22D4 U6823 ( .B1(n9127), .B2(n56), .A1(n1), .A2(Decoder[7]), .ZN(n125) );
  BUFFD0 U6824 ( .I(n6933), .Z(n6932) );
  BUFFD0 U6825 ( .I(n6934), .Z(n6933) );
  BUFFD0 U6826 ( .I(n6935), .Z(n6934) );
  BUFFD0 U6827 ( .I(n125), .Z(n6935) );
  CKBD0 U6828 ( .CLK(n124), .C(n6939) );
  BUFFD0 U6829 ( .I(n6937), .Z(n6936) );
  BUFFD0 U6830 ( .I(n6938), .Z(n6937) );
  BUFFD0 U6831 ( .I(n6939), .Z(n6938) );
  CKBD0 U6832 ( .CLK(n123), .C(n6943) );
  BUFFD0 U6833 ( .I(n6941), .Z(n6940) );
  BUFFD0 U6834 ( .I(n6942), .Z(n6941) );
  BUFFD0 U6835 ( .I(n6943), .Z(n6942) );
  IOA22D4 U6836 ( .B1(n9127), .B2(n53), .A1(n9129), .A2(Decoder[10]), .ZN(n122) );
  BUFFD0 U6837 ( .I(n6945), .Z(n6944) );
  BUFFD0 U6838 ( .I(n6946), .Z(n6945) );
  BUFFD0 U6839 ( .I(n6947), .Z(n6946) );
  BUFFD0 U6840 ( .I(n122), .Z(n6947) );
  IOA22D4 U6841 ( .B1(n9127), .B2(n52), .A1(n9129), .A2(Decoder[11]), .ZN(n121) );
  BUFFD0 U6842 ( .I(n6949), .Z(n6948) );
  BUFFD0 U6843 ( .I(n6950), .Z(n6949) );
  BUFFD0 U6844 ( .I(n6951), .Z(n6950) );
  BUFFD0 U6845 ( .I(n121), .Z(n6951) );
  IOA22D4 U6846 ( .B1(n9127), .B2(n51), .A1(n9129), .A2(Decoder[12]), .ZN(n120) );
  BUFFD0 U6847 ( .I(n6953), .Z(n6952) );
  BUFFD0 U6848 ( .I(n6954), .Z(n6953) );
  BUFFD0 U6849 ( .I(n6955), .Z(n6954) );
  BUFFD0 U6850 ( .I(n120), .Z(n6955) );
  IOA22D4 U6851 ( .B1(n9127), .B2(n50), .A1(n9129), .A2(Decoder[13]), .ZN(n119) );
  BUFFD0 U6852 ( .I(n6957), .Z(n6956) );
  BUFFD0 U6853 ( .I(n6958), .Z(n6957) );
  BUFFD0 U6854 ( .I(n6959), .Z(n6958) );
  BUFFD0 U6855 ( .I(n119), .Z(n6959) );
  IOA22D4 U6856 ( .B1(n9128), .B2(n49), .A1(n9129), .A2(Decoder[14]), .ZN(n118) );
  BUFFD0 U6857 ( .I(n6961), .Z(n6960) );
  BUFFD0 U6858 ( .I(n6962), .Z(n6961) );
  BUFFD0 U6859 ( .I(n6963), .Z(n6962) );
  BUFFD0 U6860 ( .I(n118), .Z(n6963) );
  IOA22D4 U6861 ( .B1(n9128), .B2(n48), .A1(n9129), .A2(Decoder[15]), .ZN(n117) );
  BUFFD0 U6862 ( .I(n6965), .Z(n6964) );
  BUFFD0 U6863 ( .I(n6966), .Z(n6965) );
  BUFFD0 U6864 ( .I(n6967), .Z(n6966) );
  BUFFD0 U6865 ( .I(n117), .Z(n6967) );
  IOA22D4 U6866 ( .B1(n9128), .B2(n47), .A1(n9129), .A2(Decoder[16]), .ZN(n116) );
  BUFFD0 U6867 ( .I(n6969), .Z(n6968) );
  BUFFD0 U6868 ( .I(n6970), .Z(n6969) );
  BUFFD0 U6869 ( .I(n6971), .Z(n6970) );
  BUFFD0 U6870 ( .I(n116), .Z(n6971) );
  IOA22D4 U6871 ( .B1(n9128), .B2(n46), .A1(n9129), .A2(Decoder[17]), .ZN(n115) );
  BUFFD0 U6872 ( .I(n6973), .Z(n6972) );
  BUFFD0 U6873 ( .I(n6974), .Z(n6973) );
  BUFFD0 U6874 ( .I(n6975), .Z(n6974) );
  BUFFD0 U6875 ( .I(n115), .Z(n6975) );
  IOA22D4 U6876 ( .B1(n9128), .B2(n45), .A1(n9129), .A2(Decoder[18]), .ZN(n114) );
  BUFFD0 U6877 ( .I(n6977), .Z(n6976) );
  BUFFD0 U6878 ( .I(n6978), .Z(n6977) );
  BUFFD0 U6879 ( .I(n6979), .Z(n6978) );
  BUFFD0 U6880 ( .I(n114), .Z(n6979) );
  IOA22D4 U6881 ( .B1(n9128), .B2(n44), .A1(n9129), .A2(Decoder[19]), .ZN(n113) );
  BUFFD0 U6882 ( .I(n6981), .Z(n6980) );
  BUFFD0 U6883 ( .I(n6982), .Z(n6981) );
  BUFFD0 U6884 ( .I(n6983), .Z(n6982) );
  BUFFD0 U6885 ( .I(n113), .Z(n6983) );
  IOA22D4 U6886 ( .B1(n9128), .B2(n43), .A1(n9128), .A2(Decoder[20]), .ZN(n112) );
  BUFFD0 U6887 ( .I(n6985), .Z(n6984) );
  BUFFD0 U6888 ( .I(n6986), .Z(n6985) );
  BUFFD0 U6889 ( .I(n6987), .Z(n6986) );
  BUFFD0 U6890 ( .I(n112), .Z(n6987) );
  IOA22D4 U6891 ( .B1(n9128), .B2(n42), .A1(n9129), .A2(Decoder[21]), .ZN(n111) );
  BUFFD0 U6892 ( .I(n6989), .Z(n6988) );
  BUFFD0 U6893 ( .I(n6990), .Z(n6989) );
  BUFFD0 U6894 ( .I(n6991), .Z(n6990) );
  BUFFD0 U6895 ( .I(n111), .Z(n6991) );
  IOA22D4 U6896 ( .B1(n9128), .B2(n41), .A1(n9129), .A2(Decoder[22]), .ZN(n110) );
  BUFFD0 U6897 ( .I(n6993), .Z(n6992) );
  BUFFD0 U6898 ( .I(n6994), .Z(n6993) );
  BUFFD0 U6899 ( .I(n6995), .Z(n6994) );
  BUFFD0 U6900 ( .I(n110), .Z(n6995) );
  IOA22D4 U6901 ( .B1(n9128), .B2(n40), .A1(n9129), .A2(Decoder[23]), .ZN(n109) );
  BUFFD0 U6902 ( .I(n6997), .Z(n6996) );
  BUFFD0 U6903 ( .I(n6998), .Z(n6997) );
  BUFFD0 U6904 ( .I(n6999), .Z(n6998) );
  BUFFD0 U6905 ( .I(n109), .Z(n6999) );
  IOA22D4 U6906 ( .B1(n9128), .B2(n39), .A1(n9129), .A2(Decoder[24]), .ZN(n108) );
  BUFFD0 U6907 ( .I(n7001), .Z(n7000) );
  BUFFD0 U6908 ( .I(n7002), .Z(n7001) );
  BUFFD0 U6909 ( .I(n7003), .Z(n7002) );
  BUFFD0 U6910 ( .I(n108), .Z(n7003) );
  IOA22D4 U6911 ( .B1(n9128), .B2(n38), .A1(n9129), .A2(Decoder[25]), .ZN(n107) );
  BUFFD0 U6912 ( .I(n7005), .Z(n7004) );
  BUFFD0 U6913 ( .I(n7006), .Z(n7005) );
  BUFFD0 U6914 ( .I(n7007), .Z(n7006) );
  BUFFD0 U6915 ( .I(n107), .Z(n7007) );
  IOA22D4 U6916 ( .B1(n9128), .B2(n37), .A1(n9129), .A2(Decoder[26]), .ZN(n106) );
  BUFFD0 U6917 ( .I(n7009), .Z(n7008) );
  BUFFD0 U6918 ( .I(n7010), .Z(n7009) );
  BUFFD0 U6919 ( .I(n7011), .Z(n7010) );
  BUFFD0 U6920 ( .I(n106), .Z(n7011) );
  IOA22D4 U6921 ( .B1(n9128), .B2(n36), .A1(n9129), .A2(Decoder[27]), .ZN(n105) );
  BUFFD0 U6922 ( .I(n7013), .Z(n7012) );
  BUFFD0 U6923 ( .I(n7014), .Z(n7013) );
  BUFFD0 U6924 ( .I(n7015), .Z(n7014) );
  BUFFD0 U6925 ( .I(n105), .Z(n7015) );
  IOA22D4 U6926 ( .B1(n9128), .B2(n35), .A1(n1), .A2(Decoder[28]), .ZN(n104)
         );
  BUFFD0 U6927 ( .I(n7017), .Z(n7016) );
  BUFFD0 U6928 ( .I(n7018), .Z(n7017) );
  BUFFD0 U6929 ( .I(n7019), .Z(n7018) );
  BUFFD0 U6930 ( .I(n104), .Z(n7019) );
  IOA22D4 U6931 ( .B1(n9128), .B2(n34), .A1(n1), .A2(Decoder[29]), .ZN(n103)
         );
  BUFFD0 U6932 ( .I(n7021), .Z(n7020) );
  BUFFD0 U6933 ( .I(n7022), .Z(n7021) );
  BUFFD0 U6934 ( .I(n7023), .Z(n7022) );
  BUFFD0 U6935 ( .I(n103), .Z(n7023) );
  IOA22D4 U6936 ( .B1(n9128), .B2(n33), .A1(n1), .A2(Decoder[30]), .ZN(n102)
         );
  BUFFD0 U6937 ( .I(n7025), .Z(n7024) );
  BUFFD0 U6938 ( .I(n7026), .Z(n7025) );
  BUFFD0 U6939 ( .I(n7027), .Z(n7026) );
  BUFFD0 U6940 ( .I(n102), .Z(n7027) );
  BUFFD0 U6941 ( .I(n7029), .Z(n7028) );
  BUFFD0 U6942 ( .I(n7030), .Z(n7029) );
  BUFFD0 U6943 ( .I(n7031), .Z(n7030) );
  BUFFD0 U6944 ( .I(n101), .Z(n7031) );
  BUFFD0 U6945 ( .I(n7033), .Z(n7032) );
  BUFFD0 U6946 ( .I(N37), .Z(n7033) );
  BUFFD0 U6947 ( .I(n7035), .Z(n7034) );
  BUFFD0 U6948 ( .I(N43), .Z(n7035) );
  OAI21D0 U6949 ( .A1(n3), .A2(n29), .B(n231), .ZN(n96) );
  BUFFD0 U6950 ( .I(n7037), .Z(n7036) );
  BUFFD0 U6951 ( .I(n7038), .Z(n7037) );
  BUFFD0 U6952 ( .I(n7039), .Z(n7038) );
  BUFFD0 U6953 ( .I(n96), .Z(n7039) );
  CKBD0 U6954 ( .CLK(n2145), .C(n7040) );
  CKND2D0 U6955 ( .A1(n16), .A2(n17), .ZN(n14) );
  CKBD0 U6956 ( .CLK(n2049), .C(n7041) );
  CKBD0 U6957 ( .CLK(n2241), .C(n7042) );
  CKBD0 U6958 ( .CLK(n1340), .C(n7043) );
  CKBD0 U6959 ( .CLK(n1953), .C(n7044) );
  CKBD0 U6960 ( .CLK(n2337), .C(n7045) );
  CKBD0 U6961 ( .CLK(n1642), .C(n7046) );
  CKBD0 U6962 ( .CLK(n1229), .C(n7047) );
  CKBD0 U6963 ( .CLK(n908), .C(n7048) );
  CKBD0 U6964 ( .CLK(n226), .C(n7049) );
  CKBD0 U6965 ( .CLK(n1546), .C(n7050) );
  CKBD0 U6966 ( .CLK(n1354), .C(n7051) );
  CKBD0 U6967 ( .CLK(n1842), .C(n7052) );
  CKBD0 U6968 ( .CLK(n811), .C(n7053) );
  CKBD0 U6969 ( .CLK(n1021), .C(n7054) );
  CKBD0 U6970 ( .CLK(n712), .C(n7055) );
  CKBD0 U6971 ( .CLK(n1745), .C(n7056) );
  CKBD0 U6972 ( .CLK(n1118), .C(n7057) );
  CKBD0 U6973 ( .CLK(n911), .C(n7058) );
  CKBD0 U6974 ( .CLK(n519), .C(n7059) );
  CKBD0 U6975 ( .CLK(n2529), .C(n7060) );
  BUFFD0 U6976 ( .I(n615), .Z(n7061) );
  BUFFD0 U6977 ( .I(n422), .Z(n7062) );
  CKBD0 U6978 ( .CLK(n326), .C(n7063) );
  BUFFD0 U6979 ( .I(n2433), .Z(n7064) );
  CKBD0 U6980 ( .CLK(n1450), .C(n7065) );
  CKBD0 U6981 ( .CLK(n1847), .C(n7066) );
  CKBD0 U6982 ( .CLK(n1645), .C(n7067) );
  CKBD0 U6983 ( .CLK(n1853), .C(n7068) );
  CKBD0 U6984 ( .CLK(n1649), .C(n7069) );
  CKBD0 U6985 ( .CLK(n1850), .C(n7070) );
  CKBD0 U6986 ( .CLK(n7040), .C(n7071) );
  CKBD0 U6987 ( .CLK(n1857), .C(n7072) );
  CKBD0 U6988 ( .CLK(n7041), .C(n7073) );
  CKBD0 U6989 ( .CLK(n7042), .C(n7074) );
  CKBD0 U6990 ( .CLK(n7043), .C(n7075) );
  CKBD0 U6991 ( .CLK(n7044), .C(n7076) );
  CKBD0 U6992 ( .CLK(n7045), .C(n7077) );
  CKBD0 U6993 ( .CLK(n7046), .C(n7078) );
  CKBD0 U6994 ( .CLK(n7047), .C(n7079) );
  CKBD0 U6995 ( .CLK(n7048), .C(n7080) );
  CKBD0 U6996 ( .CLK(n7049), .C(n7081) );
  CKBD0 U6997 ( .CLK(n7052), .C(n7082) );
  CKBD0 U6998 ( .CLK(n7050), .C(n7083) );
  CKBD0 U6999 ( .CLK(n7051), .C(n7084) );
  CKBD0 U7000 ( .CLK(n7053), .C(n7085) );
  CKBD0 U7001 ( .CLK(n7054), .C(n7086) );
  CKBD0 U7002 ( .CLK(n7055), .C(n7087) );
  CKBD0 U7003 ( .CLK(n7056), .C(n7088) );
  CKBD0 U7004 ( .CLK(n7057), .C(n7089) );
  CKBD0 U7005 ( .CLK(n7058), .C(n7090) );
  CKBD0 U7006 ( .CLK(n7059), .C(n7091) );
  CKBD0 U7007 ( .CLK(n7060), .C(n7092) );
  CKBD0 U7008 ( .CLK(n7061), .C(n7093) );
  CKBD0 U7009 ( .CLK(n7063), .C(n7094) );
  CKBD0 U7010 ( .CLK(n7062), .C(n7095) );
  CKBD0 U7011 ( .CLK(n7064), .C(n7096) );
  CKBD0 U7012 ( .CLK(n7065), .C(n7097) );
  CKBD0 U7013 ( .CLK(n7066), .C(n7098) );
  CKBD0 U7014 ( .CLK(n7067), .C(n7099) );
  CKBD0 U7015 ( .CLK(n7068), .C(n7100) );
  CKBD0 U7016 ( .CLK(n7069), .C(n7101) );
  CKBD0 U7017 ( .CLK(n7070), .C(n7102) );
  CKBD0 U7018 ( .CLK(n7071), .C(n7103) );
  CKBD0 U7019 ( .CLK(n7072), .C(n7104) );
  CKBD0 U7020 ( .CLK(n7073), .C(n7105) );
  CKBD0 U7021 ( .CLK(n7074), .C(n7106) );
  BUFFD0 U7022 ( .I(n7075), .Z(n7107) );
  CKBD0 U7023 ( .CLK(n7076), .C(n7108) );
  CKBD0 U7024 ( .CLK(n7077), .C(n7109) );
  CKBD0 U7025 ( .CLK(n7078), .C(n7110) );
  BUFFD0 U7026 ( .I(n7079), .Z(n7111) );
  CKBD0 U7027 ( .CLK(n7080), .C(n7112) );
  CKBD0 U7028 ( .CLK(n7081), .C(n7113) );
  CKBD0 U7029 ( .CLK(n7083), .C(n7114) );
  BUFFD0 U7030 ( .I(n7082), .Z(n7115) );
  CKBD0 U7031 ( .CLK(n7085), .C(n7116) );
  CKBD0 U7032 ( .CLK(n7084), .C(n7117) );
  CKBD0 U7033 ( .CLK(n7087), .C(n7118) );
  CKBD0 U7034 ( .CLK(n7086), .C(n7119) );
  CKBD0 U7035 ( .CLK(n7088), .C(n7120) );
  CKBD0 U7036 ( .CLK(n7089), .C(n7121) );
  CKBD0 U7037 ( .CLK(n7090), .C(n7122) );
  CKBD0 U7038 ( .CLK(n7091), .C(n7123) );
  CKBD0 U7039 ( .CLK(n7092), .C(n7124) );
  CKBD0 U7040 ( .CLK(n7094), .C(n7125) );
  CKBD0 U7041 ( .CLK(n7093), .C(n7126) );
  CKBD0 U7042 ( .CLK(n7095), .C(n7127) );
  CKBD0 U7043 ( .CLK(n7096), .C(n7128) );
  CKBD0 U7044 ( .CLK(n7097), .C(n7129) );
  CKBD0 U7045 ( .CLK(n7098), .C(n7130) );
  CKBD0 U7046 ( .CLK(n7099), .C(n7131) );
  CKBD0 U7047 ( .CLK(n7100), .C(n7132) );
  CKBD0 U7048 ( .CLK(n7101), .C(n7133) );
  CKBD0 U7049 ( .CLK(n7102), .C(n7134) );
  CKBD0 U7050 ( .CLK(n7103), .C(n7135) );
  CKBD0 U7051 ( .CLK(n7104), .C(n7136) );
  CKBD0 U7052 ( .CLK(n7105), .C(n7137) );
  CKBD0 U7053 ( .CLK(n7106), .C(n7138) );
  CKBD0 U7054 ( .CLK(n7107), .C(n7139) );
  CKBD0 U7055 ( .CLK(n7108), .C(n7140) );
  CKBD0 U7056 ( .CLK(n7109), .C(n7141) );
  CKBD0 U7057 ( .CLK(n7110), .C(n7142) );
  CKBD0 U7058 ( .CLK(n7111), .C(n7143) );
  BUFFD0 U7059 ( .I(n7112), .Z(n7144) );
  CKBD0 U7060 ( .CLK(n7113), .C(n7145) );
  CKBD0 U7061 ( .CLK(n7114), .C(n7146) );
  CKBD0 U7062 ( .CLK(n7115), .C(n7147) );
  BUFFD0 U7063 ( .I(n7116), .Z(n7148) );
  CKBD0 U7064 ( .CLK(n7117), .C(n7149) );
  CKBD0 U7065 ( .CLK(n7119), .C(n7150) );
  BUFFD0 U7066 ( .I(n7118), .Z(n7151) );
  CKBD0 U7067 ( .CLK(n7120), .C(n7152) );
  BUFFD0 U7068 ( .I(n7121), .Z(n7153) );
  BUFFD0 U7069 ( .I(n7123), .Z(n7154) );
  CKBD0 U7070 ( .CLK(n7122), .C(n7155) );
  CKBD0 U7071 ( .CLK(n7124), .C(n7156) );
  BUFFD0 U7072 ( .I(n7125), .Z(n7157) );
  CKBD0 U7073 ( .CLK(n7126), .C(n7158) );
  CKBD0 U7074 ( .CLK(n7127), .C(n7159) );
  CKBD0 U7075 ( .CLK(n7128), .C(n7160) );
  CKBD0 U7076 ( .CLK(n7129), .C(n7161) );
  CKBD0 U7077 ( .CLK(n7130), .C(n7162) );
  CKBD0 U7078 ( .CLK(n7131), .C(n7163) );
  CKBD0 U7079 ( .CLK(n7132), .C(n7164) );
  CKBD0 U7080 ( .CLK(n7133), .C(n7165) );
  CKBD0 U7081 ( .CLK(n7134), .C(n7166) );
  CKBD0 U7082 ( .CLK(n7135), .C(n7167) );
  CKBD0 U7083 ( .CLK(n7137), .C(n7168) );
  CKBD0 U7084 ( .CLK(n7136), .C(n7169) );
  CKBD0 U7085 ( .CLK(n7138), .C(n7170) );
  CKBD0 U7086 ( .CLK(n7139), .C(n7171) );
  CKBD0 U7087 ( .CLK(n7140), .C(n7172) );
  CKBD0 U7088 ( .CLK(n7141), .C(n7173) );
  CKBD0 U7089 ( .CLK(n7142), .C(n7174) );
  CKBD0 U7090 ( .CLK(n7143), .C(n7175) );
  CKBD0 U7091 ( .CLK(n7145), .C(n7176) );
  CKBD0 U7092 ( .CLK(n7144), .C(n7177) );
  CKBD0 U7093 ( .CLK(n7146), .C(n7178) );
  CKBD0 U7094 ( .CLK(n7147), .C(n7179) );
  CKBD0 U7095 ( .CLK(n7148), .C(n7180) );
  CKBD0 U7096 ( .CLK(n7150), .C(n7181) );
  CKBD0 U7097 ( .CLK(n7149), .C(n7182) );
  CKBD0 U7098 ( .CLK(n7151), .C(n7183) );
  BUFFD0 U7099 ( .I(n7152), .Z(n7184) );
  CKBD0 U7100 ( .CLK(n7153), .C(n7185) );
  CKBD0 U7101 ( .CLK(n7154), .C(n7186) );
  CKBD0 U7102 ( .CLK(n7155), .C(n7187) );
  BUFFD0 U7103 ( .I(n7156), .Z(n7188) );
  CKBD0 U7104 ( .CLK(n7157), .C(n7189) );
  CKBD0 U7105 ( .CLK(n7158), .C(n7190) );
  CKBD0 U7106 ( .CLK(n7159), .C(n7191) );
  CKBD0 U7107 ( .CLK(n7160), .C(n7192) );
  CKBD0 U7108 ( .CLK(n7161), .C(n7193) );
  CKBD0 U7109 ( .CLK(n7162), .C(n7194) );
  CKBD0 U7110 ( .CLK(n7163), .C(n7195) );
  CKBD0 U7111 ( .CLK(n7164), .C(n7196) );
  CKBD0 U7112 ( .CLK(n7165), .C(n7197) );
  CKBD0 U7113 ( .CLK(n7166), .C(n7198) );
  BUFFD0 U7114 ( .I(n7167), .Z(n7199) );
  BUFFD0 U7115 ( .I(n7168), .Z(n7200) );
  BUFFD0 U7116 ( .I(n7170), .Z(n7201) );
  CKBD0 U7117 ( .CLK(n7169), .C(n7202) );
  CKBD0 U7118 ( .CLK(n7171), .C(n7203) );
  BUFFD0 U7119 ( .I(n7172), .Z(n7204) );
  BUFFD0 U7120 ( .I(n7173), .Z(n7205) );
  BUFFD0 U7121 ( .I(n7174), .Z(n7206) );
  CKBD0 U7122 ( .CLK(n7175), .C(n7207) );
  CKBD0 U7123 ( .CLK(n7177), .C(n7208) );
  BUFFD0 U7124 ( .I(n7176), .Z(n7209) );
  BUFFD0 U7125 ( .I(n7178), .Z(n7210) );
  CKBD0 U7126 ( .CLK(n7179), .C(n7211) );
  CKBD0 U7127 ( .CLK(n7180), .C(n7212) );
  BUFFD0 U7128 ( .I(n7181), .Z(n7213) );
  CKBD0 U7129 ( .CLK(n7182), .C(n7214) );
  CKBD0 U7130 ( .CLK(n7183), .C(n7215) );
  CKBD0 U7131 ( .CLK(n7184), .C(n7216) );
  CKBD0 U7132 ( .CLK(n7185), .C(n7217) );
  CKBD0 U7133 ( .CLK(n7186), .C(n7218) );
  CKBD0 U7134 ( .CLK(n7187), .C(n7219) );
  CKBD0 U7135 ( .CLK(n7188), .C(n7220) );
  CKBD0 U7136 ( .CLK(n7189), .C(n7221) );
  CKBD0 U7137 ( .CLK(n7190), .C(n7222) );
  CKBD0 U7138 ( .CLK(n7191), .C(n7223) );
  CKBD0 U7139 ( .CLK(n7192), .C(n7224) );
  BUFFD0 U7140 ( .I(n7193), .Z(n7225) );
  CKBD0 U7141 ( .CLK(n7194), .C(n7226) );
  CKBD0 U7142 ( .CLK(n7195), .C(n7227) );
  CKBD0 U7143 ( .CLK(n7196), .C(n7228) );
  CKBD0 U7144 ( .CLK(n7197), .C(n7229) );
  CKBD0 U7145 ( .CLK(n7198), .C(n7230) );
  CKBD0 U7146 ( .CLK(n7199), .C(n7231) );
  CKBD0 U7147 ( .CLK(n7200), .C(n7232) );
  CKBD0 U7148 ( .CLK(n7201), .C(n7233) );
  CKBD0 U7149 ( .CLK(n7202), .C(n7234) );
  CKBD0 U7150 ( .CLK(n7203), .C(n7235) );
  CKBD0 U7151 ( .CLK(n7204), .C(n7236) );
  CKBD0 U7152 ( .CLK(n7205), .C(n7237) );
  CKBD0 U7153 ( .CLK(n7206), .C(n7238) );
  CKBD0 U7154 ( .CLK(n7207), .C(n7239) );
  CKBD0 U7155 ( .CLK(n7208), .C(n7240) );
  CKBD0 U7156 ( .CLK(n7209), .C(n7241) );
  CKBD0 U7157 ( .CLK(n7210), .C(n7242) );
  CKBD0 U7158 ( .CLK(n7211), .C(n7243) );
  CKBD0 U7159 ( .CLK(n7212), .C(n7244) );
  CKBD0 U7160 ( .CLK(n7213), .C(n7245) );
  CKBD0 U7161 ( .CLK(n7215), .C(n7246) );
  CKBD0 U7162 ( .CLK(n7214), .C(n7247) );
  CKBD0 U7163 ( .CLK(n7216), .C(n7248) );
  CKBD0 U7164 ( .CLK(n7217), .C(n7249) );
  CKBD0 U7165 ( .CLK(n7218), .C(n7250) );
  CKBD0 U7166 ( .CLK(n7220), .C(n7251) );
  CKBD0 U7167 ( .CLK(n7219), .C(n7252) );
  CKBD0 U7168 ( .CLK(n7221), .C(n7253) );
  CKBD0 U7169 ( .CLK(n7222), .C(n7254) );
  CKBD0 U7170 ( .CLK(n7223), .C(n7255) );
  CKBD0 U7171 ( .CLK(n7224), .C(n7256) );
  CKBD0 U7172 ( .CLK(n7225), .C(n7257) );
  CKBD0 U7173 ( .CLK(n7226), .C(n7258) );
  CKBD0 U7174 ( .CLK(n7227), .C(n7259) );
  CKBD0 U7175 ( .CLK(n7228), .C(n7260) );
  CKBD0 U7176 ( .CLK(n7229), .C(n7261) );
  CKBD0 U7177 ( .CLK(n7231), .C(n7262) );
  CKBD0 U7178 ( .CLK(n7230), .C(n7263) );
  CKBD0 U7179 ( .CLK(n7232), .C(n7264) );
  CKBD0 U7180 ( .CLK(n7233), .C(n7265) );
  CKBD0 U7181 ( .CLK(n7234), .C(n7266) );
  CKBD0 U7182 ( .CLK(n7235), .C(n7267) );
  CKBD0 U7183 ( .CLK(n7236), .C(n7268) );
  CKBD0 U7184 ( .CLK(n7237), .C(n7269) );
  CKBD0 U7185 ( .CLK(n7238), .C(n7270) );
  CKBD0 U7186 ( .CLK(n7239), .C(n7271) );
  CKBD0 U7187 ( .CLK(n7240), .C(n7272) );
  CKBD0 U7188 ( .CLK(n7241), .C(n7273) );
  CKBD0 U7189 ( .CLK(n7242), .C(n7274) );
  CKBD0 U7190 ( .CLK(n7243), .C(n7275) );
  CKBD0 U7191 ( .CLK(n7244), .C(n7276) );
  CKBD0 U7192 ( .CLK(n7245), .C(n7277) );
  CKBD0 U7193 ( .CLK(n7247), .C(n7278) );
  CKBD0 U7194 ( .CLK(n7246), .C(n7279) );
  CKBD0 U7195 ( .CLK(n7248), .C(n7280) );
  CKBD0 U7196 ( .CLK(n7249), .C(n7281) );
  CKBD0 U7197 ( .CLK(n7250), .C(n7282) );
  CKBD0 U7198 ( .CLK(n7251), .C(n7283) );
  CKBD0 U7199 ( .CLK(n7252), .C(n7284) );
  CKBD0 U7200 ( .CLK(n7253), .C(n7285) );
  CKBD0 U7201 ( .CLK(n7254), .C(n7286) );
  CKBD0 U7202 ( .CLK(n7255), .C(n7287) );
  CKBD0 U7203 ( .CLK(n7256), .C(n7288) );
  CKBD0 U7204 ( .CLK(n7257), .C(n7289) );
  BUFFD0 U7205 ( .I(n7258), .Z(n7290) );
  CKBD0 U7206 ( .CLK(n7259), .C(n7291) );
  CKBD0 U7207 ( .CLK(n7260), .C(n7292) );
  CKBD0 U7208 ( .CLK(n7261), .C(n7293) );
  CKBD0 U7209 ( .CLK(n7263), .C(n7294) );
  CKBD0 U7210 ( .CLK(n7262), .C(n7295) );
  CKBD0 U7211 ( .CLK(n7264), .C(n7296) );
  CKBD0 U7212 ( .CLK(n7265), .C(n7297) );
  CKBD0 U7213 ( .CLK(n7266), .C(n7298) );
  CKBD0 U7214 ( .CLK(n7267), .C(n7299) );
  CKBD0 U7215 ( .CLK(n7268), .C(n7300) );
  CKBD0 U7216 ( .CLK(n7269), .C(n7301) );
  CKBD0 U7217 ( .CLK(n7270), .C(n7302) );
  CKBD0 U7218 ( .CLK(n7271), .C(n7303) );
  CKBD0 U7219 ( .CLK(n7272), .C(n7304) );
  CKBD0 U7220 ( .CLK(n7273), .C(n7305) );
  BUFFD0 U7221 ( .I(n7278), .Z(n7306) );
  CKBD0 U7222 ( .CLK(n7274), .C(n7307) );
  CKBD0 U7223 ( .CLK(n7275), .C(n7308) );
  CKBD0 U7224 ( .CLK(n7276), .C(n7309) );
  CKBD0 U7225 ( .CLK(n7277), .C(n7310) );
  CKBD0 U7226 ( .CLK(n7279), .C(n7311) );
  CKBD0 U7227 ( .CLK(n7280), .C(n7312) );
  CKBD0 U7228 ( .CLK(n7281), .C(n7313) );
  CKBD0 U7229 ( .CLK(n7282), .C(n7314) );
  CKBD0 U7230 ( .CLK(n7283), .C(n7315) );
  CKBD0 U7231 ( .CLK(n7284), .C(n7316) );
  CKBD0 U7232 ( .CLK(n7285), .C(n7317) );
  CKBD0 U7233 ( .CLK(n7286), .C(n7318) );
  CKBD0 U7234 ( .CLK(n7287), .C(n7319) );
  CKBD0 U7235 ( .CLK(n7288), .C(n7320) );
  CKBD0 U7236 ( .CLK(n7289), .C(n7321) );
  CKBD0 U7237 ( .CLK(n7290), .C(n7322) );
  BUFFD0 U7238 ( .I(n7291), .Z(n7323) );
  BUFFD0 U7239 ( .I(n7292), .Z(n7324) );
  CKBD0 U7240 ( .CLK(n7293), .C(n7325) );
  BUFFD0 U7241 ( .I(n7294), .Z(n7326) );
  CKBD0 U7242 ( .CLK(n7295), .C(n7327) );
  CKBD0 U7243 ( .CLK(n7296), .C(n7328) );
  CKBD0 U7244 ( .CLK(n7297), .C(n7329) );
  CKBD0 U7245 ( .CLK(n7298), .C(n7330) );
  CKBD0 U7246 ( .CLK(n7299), .C(n7331) );
  CKBD0 U7247 ( .CLK(n7300), .C(n7332) );
  CKBD0 U7248 ( .CLK(n7301), .C(n7333) );
  CKBD0 U7249 ( .CLK(n7302), .C(n7334) );
  CKBD0 U7250 ( .CLK(n7303), .C(n7335) );
  CKBD0 U7251 ( .CLK(n7304), .C(n7336) );
  CKBD0 U7252 ( .CLK(n7305), .C(n7337) );
  CKBD0 U7253 ( .CLK(n7306), .C(n7338) );
  CKBD0 U7254 ( .CLK(n7307), .C(n7339) );
  CKBD0 U7255 ( .CLK(n7308), .C(n7340) );
  CKBD0 U7256 ( .CLK(n7309), .C(n7341) );
  CKBD0 U7257 ( .CLK(n7310), .C(n7342) );
  CKBD0 U7258 ( .CLK(n7311), .C(n7343) );
  CKBD0 U7259 ( .CLK(n7312), .C(n7344) );
  CKBD0 U7260 ( .CLK(n7313), .C(n7345) );
  CKBD0 U7261 ( .CLK(n7314), .C(n7346) );
  CKBD0 U7262 ( .CLK(n7315), .C(n7347) );
  CKBD0 U7263 ( .CLK(n7316), .C(n7348) );
  CKBD0 U7264 ( .CLK(n7317), .C(n7349) );
  CKBD0 U7265 ( .CLK(n7318), .C(n7350) );
  CKBD0 U7266 ( .CLK(n7319), .C(n7351) );
  CKBD0 U7267 ( .CLK(n7320), .C(n7352) );
  CKBD0 U7268 ( .CLK(n7321), .C(n7353) );
  CKBD0 U7269 ( .CLK(n7322), .C(n7354) );
  CKBD0 U7270 ( .CLK(n7323), .C(n7355) );
  CKBD0 U7271 ( .CLK(n7324), .C(n7356) );
  CKBD0 U7272 ( .CLK(n7325), .C(n7357) );
  CKBD0 U7273 ( .CLK(n7326), .C(n7358) );
  CKBD0 U7274 ( .CLK(n7327), .C(n7359) );
  CKBD0 U7275 ( .CLK(n7328), .C(n7360) );
  CKBD0 U7276 ( .CLK(n7329), .C(n7361) );
  CKBD0 U7277 ( .CLK(n7330), .C(n7362) );
  CKBD0 U7278 ( .CLK(n7331), .C(n7363) );
  CKBD0 U7279 ( .CLK(n7332), .C(n7364) );
  CKBD0 U7280 ( .CLK(n7333), .C(n7365) );
  CKBD0 U7281 ( .CLK(n7334), .C(n7366) );
  CKBD0 U7282 ( .CLK(n7335), .C(n7367) );
  CKBD0 U7283 ( .CLK(n7336), .C(n7368) );
  CKBD0 U7284 ( .CLK(n7337), .C(n7369) );
  CKBD0 U7285 ( .CLK(n7339), .C(n7370) );
  CKBD0 U7286 ( .CLK(n7338), .C(n7371) );
  CKBD0 U7287 ( .CLK(n7340), .C(n7372) );
  CKBD0 U7288 ( .CLK(n7341), .C(n7373) );
  CKBD0 U7289 ( .CLK(n7342), .C(n7374) );
  CKBD0 U7290 ( .CLK(n7343), .C(n7375) );
  CKBD0 U7291 ( .CLK(n7344), .C(n7376) );
  BUFFD0 U7292 ( .I(n7348), .Z(n7377) );
  CKBD0 U7293 ( .CLK(n7345), .C(n7378) );
  CKBD0 U7294 ( .CLK(n7346), .C(n7379) );
  CKBD0 U7295 ( .CLK(n7347), .C(n7380) );
  CKBD0 U7296 ( .CLK(n7349), .C(n7381) );
  CKBD0 U7297 ( .CLK(n7350), .C(n7382) );
  CKBD0 U7298 ( .CLK(n7351), .C(n7383) );
  CKBD0 U7299 ( .CLK(n7352), .C(n7384) );
  CKBD0 U7300 ( .CLK(n7353), .C(n7385) );
  CKBD0 U7301 ( .CLK(n7354), .C(n7386) );
  CKBD0 U7302 ( .CLK(n7355), .C(n7387) );
  CKBD0 U7303 ( .CLK(n7356), .C(n7388) );
  BUFFD0 U7304 ( .I(n7357), .Z(n7389) );
  CKBD0 U7305 ( .CLK(n7358), .C(n7390) );
  CKBD0 U7306 ( .CLK(n7359), .C(n7391) );
  BUFFD0 U7307 ( .I(n7362), .Z(n7392) );
  CKBD0 U7308 ( .CLK(n7360), .C(n7393) );
  CKBD0 U7309 ( .CLK(n7361), .C(n7394) );
  CKBD0 U7310 ( .CLK(n7363), .C(n7395) );
  CKBD0 U7311 ( .CLK(n7364), .C(n7396) );
  CKBD0 U7312 ( .CLK(n7365), .C(n7397) );
  CKBD0 U7313 ( .CLK(n7366), .C(n7398) );
  CKBD0 U7314 ( .CLK(n7367), .C(n7399) );
  CKBD0 U7315 ( .CLK(n7368), .C(n7400) );
  CKBD0 U7316 ( .CLK(n7369), .C(n7401) );
  CKBD0 U7317 ( .CLK(n7370), .C(n7402) );
  CKBD0 U7318 ( .CLK(n7371), .C(n7403) );
  CKBD0 U7319 ( .CLK(n7372), .C(n7404) );
  CKBD0 U7320 ( .CLK(n7373), .C(n7405) );
  CKBD0 U7321 ( .CLK(n7374), .C(n7406) );
  CKBD0 U7322 ( .CLK(n7375), .C(n7407) );
  CKBD0 U7323 ( .CLK(n7376), .C(n7408) );
  CKBD0 U7324 ( .CLK(n7378), .C(n7409) );
  CKBD0 U7325 ( .CLK(n7377), .C(n7410) );
  CKBD0 U7326 ( .CLK(n7379), .C(n7411) );
  CKBD0 U7327 ( .CLK(n7380), .C(n7412) );
  CKBD0 U7328 ( .CLK(n7381), .C(n7413) );
  CKBD0 U7329 ( .CLK(n7382), .C(n7414) );
  CKBD0 U7330 ( .CLK(n7383), .C(n7415) );
  CKBD0 U7331 ( .CLK(n7384), .C(n7416) );
  CKBD0 U7332 ( .CLK(n7385), .C(n7417) );
  CKBD0 U7333 ( .CLK(n7391), .C(n7418) );
  CKBD0 U7334 ( .CLK(n7393), .C(n7419) );
  CKBD0 U7335 ( .CLK(n7394), .C(n7420) );
  CKBD0 U7336 ( .CLK(n7395), .C(n7421) );
  CKBD0 U7337 ( .CLK(n7396), .C(n7422) );
  CKBD0 U7338 ( .CLK(n7397), .C(n7423) );
  CKBD0 U7339 ( .CLK(n7398), .C(n7424) );
  CKBD0 U7340 ( .CLK(n7399), .C(n7425) );
  CKBD0 U7341 ( .CLK(n7400), .C(n7426) );
  CKBD0 U7342 ( .CLK(n7401), .C(n7427) );
  CKBD0 U7343 ( .CLK(n7404), .C(n7428) );
  CKBD0 U7344 ( .CLK(n7402), .C(n7429) );
  CKBD0 U7345 ( .CLK(n7405), .C(n7430) );
  CKBD0 U7346 ( .CLK(n7406), .C(n7431) );
  CKBD0 U7347 ( .CLK(n7407), .C(n7432) );
  CKBD0 U7348 ( .CLK(n7408), .C(n7433) );
  CKBD0 U7349 ( .CLK(n7409), .C(n7434) );
  CKBD0 U7350 ( .CLK(n7411), .C(n7435) );
  CKBD0 U7351 ( .CLK(n7412), .C(n7436) );
  CKBD0 U7352 ( .CLK(n7413), .C(n7437) );
  BUFFD0 U7353 ( .I(n7416), .Z(n7438) );
  CKBD0 U7354 ( .CLK(n7414), .C(n7439) );
  CKBD0 U7355 ( .CLK(n7386), .C(n7440) );
  CKBD0 U7356 ( .CLK(n7387), .C(n7441) );
  CKBD0 U7357 ( .CLK(n7388), .C(n7442) );
  CKBD0 U7358 ( .CLK(n7389), .C(n7443) );
  CKBD0 U7359 ( .CLK(n7390), .C(n7444) );
  CKBD0 U7360 ( .CLK(n7392), .C(n7445) );
  CKBD0 U7361 ( .CLK(n7403), .C(n7446) );
  CKBD0 U7362 ( .CLK(n7410), .C(n7447) );
  CKBD0 U7363 ( .CLK(n7440), .C(n7448) );
  CKBD0 U7364 ( .CLK(n7441), .C(n7449) );
  CKBD0 U7365 ( .CLK(n7442), .C(n7450) );
  CKBD0 U7366 ( .CLK(n7443), .C(n7451) );
  CKBD0 U7367 ( .CLK(n7444), .C(n7452) );
  CKBD0 U7368 ( .CLK(n7445), .C(n7453) );
  CKBD0 U7369 ( .CLK(n7446), .C(n7454) );
  CKBD0 U7370 ( .CLK(n7447), .C(n7455) );
  CKBD0 U7371 ( .CLK(n7448), .C(n7456) );
  CKBD0 U7372 ( .CLK(n7415), .C(n7457) );
  CKBD0 U7373 ( .CLK(n7449), .C(n7458) );
  CKBD0 U7374 ( .CLK(n7450), .C(n7459) );
  CKBD0 U7375 ( .CLK(n7417), .C(n7460) );
  CKBD0 U7376 ( .CLK(n7451), .C(n7461) );
  CKBD0 U7377 ( .CLK(n7452), .C(n7462) );
  CKBD0 U7378 ( .CLK(n7453), .C(n7463) );
  CKBD0 U7379 ( .CLK(n7418), .C(n7464) );
  CKBD0 U7380 ( .CLK(n7454), .C(n7465) );
  CKBD0 U7381 ( .CLK(n7419), .C(n7466) );
  CKBD0 U7382 ( .CLK(n7420), .C(n7467) );
  BUFFD0 U7383 ( .I(n7421), .Z(n7468) );
  CKBD0 U7384 ( .CLK(n7455), .C(n7469) );
  CKBD0 U7385 ( .CLK(n7422), .C(n7470) );
  CKBD0 U7386 ( .CLK(n7456), .C(n7471) );
  CKBD0 U7387 ( .CLK(n7458), .C(n7472) );
  CKBD0 U7388 ( .CLK(n7459), .C(n7473) );
  CKBD0 U7389 ( .CLK(n7461), .C(n7474) );
  CKBD0 U7390 ( .CLK(n7462), .C(n7475) );
  CKBD0 U7391 ( .CLK(n7463), .C(n7476) );
  CKBD0 U7392 ( .CLK(n7465), .C(n7477) );
  CKBD0 U7393 ( .CLK(n7423), .C(n7478) );
  CKBD0 U7394 ( .CLK(n7424), .C(n7479) );
  BUFFD0 U7395 ( .I(n7425), .Z(n7480) );
  CKBD0 U7396 ( .CLK(n7426), .C(n7481) );
  CKBD0 U7397 ( .CLK(n7427), .C(n7482) );
  CKBD0 U7398 ( .CLK(n7429), .C(n7483) );
  BUFFD0 U7399 ( .I(n7428), .Z(n7484) );
  CKBD0 U7400 ( .CLK(n7469), .C(n7485) );
  CKBD0 U7401 ( .CLK(n7471), .C(n7486) );
  CKBD0 U7402 ( .CLK(n7472), .C(n7487) );
  CKBD0 U7403 ( .CLK(n7473), .C(n7488) );
  CKBD0 U7404 ( .CLK(n7474), .C(n7489) );
  CKBD0 U7405 ( .CLK(n7475), .C(n7490) );
  CKBD0 U7406 ( .CLK(n7476), .C(n7491) );
  CKBD0 U7407 ( .CLK(n7477), .C(n7492) );
  CKBD0 U7408 ( .CLK(n7430), .C(n7493) );
  CKBD0 U7409 ( .CLK(n7432), .C(n7494) );
  CKBD0 U7410 ( .CLK(n7431), .C(n7495) );
  CKBD0 U7411 ( .CLK(n7433), .C(n7496) );
  CKBD0 U7412 ( .CLK(n7434), .C(n7497) );
  CKBD0 U7413 ( .CLK(n7485), .C(n7498) );
  CKBD0 U7414 ( .CLK(n7486), .C(n7499) );
  CKBD0 U7415 ( .CLK(n7487), .C(n7500) );
  CKBD0 U7416 ( .CLK(n7488), .C(n7501) );
  CKBD0 U7417 ( .CLK(n7489), .C(n7502) );
  CKBD0 U7418 ( .CLK(n7490), .C(n7503) );
  CKBD0 U7419 ( .CLK(n7491), .C(n7504) );
  CKBD0 U7420 ( .CLK(n7492), .C(n7505) );
  CKBD0 U7421 ( .CLK(n7435), .C(n7506) );
  CKBD0 U7422 ( .CLK(n7436), .C(n7507) );
  CKBD0 U7423 ( .CLK(n7437), .C(n7508) );
  BUFFD0 U7424 ( .I(n7439), .Z(n7509) );
  BUFFD0 U7425 ( .I(n7457), .Z(n7510) );
  CKBD0 U7426 ( .CLK(n7498), .C(n7511) );
  CKBD0 U7427 ( .CLK(n7438), .C(n7512) );
  CKBD0 U7428 ( .CLK(n7460), .C(n7513) );
  CKBD0 U7429 ( .CLK(n7499), .C(n7514) );
  CKBD0 U7430 ( .CLK(n7500), .C(n7515) );
  CKBD0 U7431 ( .CLK(n7501), .C(n7516) );
  CKBD0 U7432 ( .CLK(n7502), .C(n7517) );
  CKBD0 U7433 ( .CLK(n7464), .C(n7518) );
  CKBD0 U7434 ( .CLK(n7503), .C(n7519) );
  CKBD0 U7435 ( .CLK(n7466), .C(n7520) );
  CKBD0 U7436 ( .CLK(n7467), .C(n7521) );
  CKBD0 U7437 ( .CLK(n7468), .C(n7522) );
  CKBD0 U7438 ( .CLK(n7470), .C(n7523) );
  CKBD0 U7439 ( .CLK(n7504), .C(n7524) );
  CKBD0 U7440 ( .CLK(n7478), .C(n7525) );
  CKBD0 U7441 ( .CLK(n7479), .C(n7526) );
  CKBD0 U7442 ( .CLK(n7480), .C(n7527) );
  BUFFD0 U7443 ( .I(n7481), .Z(n7528) );
  CKBD0 U7444 ( .CLK(n7482), .C(n7529) );
  CKBD0 U7445 ( .CLK(n7483), .C(n7530) );
  CKBD0 U7446 ( .CLK(n7484), .C(n7531) );
  CKBD0 U7447 ( .CLK(n7505), .C(n7532) );
  CKBD0 U7448 ( .CLK(n7511), .C(n7533) );
  CKBD0 U7449 ( .CLK(n7514), .C(n7534) );
  BUFFD0 U7450 ( .I(n7515), .Z(n7535) );
  BUFFD0 U7451 ( .I(n7516), .Z(n7536) );
  CKBD0 U7452 ( .CLK(n7517), .C(n7537) );
  BUFFD0 U7453 ( .I(n7519), .Z(n7538) );
  CKBD0 U7454 ( .CLK(n7524), .C(n7539) );
  BUFFD0 U7455 ( .I(n7493), .Z(n7540) );
  CKBD0 U7456 ( .CLK(n7495), .C(n7541) );
  BUFFD0 U7457 ( .I(n7494), .Z(n7542) );
  CKBD0 U7458 ( .CLK(n7496), .C(n7543) );
  BUFFD0 U7459 ( .I(n7497), .Z(n7544) );
  BUFFD0 U7460 ( .I(n7506), .Z(n7545) );
  BUFFD0 U7461 ( .I(n7532), .Z(n7546) );
  CKBD0 U7462 ( .CLK(n7533), .C(n7547) );
  BUFFD0 U7463 ( .I(n7534), .Z(n7548) );
  CKBD0 U7464 ( .CLK(n7535), .C(n7549) );
  CKBD0 U7465 ( .CLK(n7536), .C(n7550) );
  CKBD0 U7466 ( .CLK(n7537), .C(n7551) );
  CKBD0 U7467 ( .CLK(n7538), .C(n7552) );
  CKBD0 U7468 ( .CLK(n7539), .C(n7553) );
  CKBD0 U7469 ( .CLK(n7507), .C(n7554) );
  BUFFD0 U7470 ( .I(n7508), .Z(n7555) );
  CKBD0 U7471 ( .CLK(n7509), .C(n7556) );
  CKBD0 U7472 ( .CLK(n7546), .C(n7557) );
  CKBD0 U7473 ( .CLK(n7547), .C(n7558) );
  CKBD0 U7474 ( .CLK(n7548), .C(n7559) );
  CKBD0 U7475 ( .CLK(n7549), .C(n7560) );
  CKBD0 U7476 ( .CLK(n7550), .C(n7561) );
  CKBD0 U7477 ( .CLK(n7551), .C(n7562) );
  CKBD0 U7478 ( .CLK(n7552), .C(n7563) );
  CKBD0 U7479 ( .CLK(n7553), .C(n7564) );
  CKBD0 U7480 ( .CLK(n7510), .C(n7565) );
  CKBD0 U7481 ( .CLK(n7512), .C(n7566) );
  CKBD0 U7482 ( .CLK(n7557), .C(n7567) );
  CKBD0 U7483 ( .CLK(n7513), .C(n7568) );
  BUFFD0 U7484 ( .I(n7558), .Z(n7569) );
  CKBD0 U7485 ( .CLK(n7559), .C(n7570) );
  BUFFD0 U7486 ( .I(n7518), .Z(n7571) );
  CKBD0 U7487 ( .CLK(n7560), .C(n7572) );
  CKBD0 U7488 ( .CLK(n7561), .C(n7573) );
  BUFFD0 U7489 ( .I(n7520), .Z(n7574) );
  BUFFD0 U7490 ( .I(n7562), .Z(n7575) );
  CKBD0 U7491 ( .CLK(n7563), .C(n7576) );
  BUFFD0 U7492 ( .I(n7564), .Z(n7577) );
  CKBD0 U7493 ( .CLK(n7567), .C(n7578) );
  CKBD0 U7494 ( .CLK(n7569), .C(n7579) );
  CKBD0 U7495 ( .CLK(n7570), .C(n7580) );
  BUFFD0 U7496 ( .I(n7521), .Z(n7581) );
  CKBD0 U7497 ( .CLK(n7522), .C(n7582) );
  CKBD0 U7498 ( .CLK(n7523), .C(n7583) );
  CKBD0 U7499 ( .CLK(n7525), .C(n7584) );
  CKBD0 U7500 ( .CLK(n7526), .C(n7585) );
  CKBD0 U7501 ( .CLK(n7572), .C(n7586) );
  CKBD0 U7502 ( .CLK(n7573), .C(n7587) );
  CKBD0 U7503 ( .CLK(n7575), .C(n7588) );
  CKBD0 U7504 ( .CLK(n7576), .C(n7589) );
  CKBD0 U7505 ( .CLK(n7577), .C(n7590) );
  CKBD0 U7506 ( .CLK(n7578), .C(n7591) );
  CKBD0 U7507 ( .CLK(n7579), .C(n7592) );
  CKBD0 U7508 ( .CLK(n7580), .C(n7593) );
  CKBD0 U7509 ( .CLK(n7527), .C(n7594) );
  CKBD0 U7510 ( .CLK(n7529), .C(n7595) );
  CKBD0 U7511 ( .CLK(n7528), .C(n7596) );
  CKBD0 U7512 ( .CLK(n7530), .C(n7597) );
  CKBD0 U7513 ( .CLK(n7531), .C(n7598) );
  CKBD0 U7514 ( .CLK(n7540), .C(n7599) );
  CKBD0 U7515 ( .CLK(n7586), .C(n7600) );
  CKBD0 U7516 ( .CLK(n7587), .C(n7601) );
  BUFFD0 U7517 ( .I(n7541), .Z(n7602) );
  CKBD0 U7518 ( .CLK(n7588), .C(n7603) );
  CKBD0 U7519 ( .CLK(n7589), .C(n7604) );
  CKBD0 U7520 ( .CLK(n7590), .C(n7605) );
  CKBD0 U7521 ( .CLK(n7591), .C(n7606) );
  CKBD0 U7522 ( .CLK(n7592), .C(n7607) );
  CKBD0 U7523 ( .CLK(n7593), .C(n7608) );
  CKBD0 U7524 ( .CLK(n7542), .C(n7609) );
  BUFFD0 U7525 ( .I(n7543), .Z(n7610) );
  CKBD0 U7526 ( .CLK(n7544), .C(n7611) );
  CKBD0 U7527 ( .CLK(n7545), .C(n7612) );
  CKBD0 U7528 ( .CLK(n7600), .C(n7613) );
  CKBD0 U7529 ( .CLK(n7601), .C(n7614) );
  CKBD0 U7530 ( .CLK(n7603), .C(n7615) );
  CKBD0 U7531 ( .CLK(n7604), .C(n7616) );
  CKBD0 U7532 ( .CLK(n7605), .C(n7617) );
  CKBD0 U7533 ( .CLK(n7606), .C(n7618) );
  CKBD0 U7534 ( .CLK(n7607), .C(n7619) );
  CKBD0 U7535 ( .CLK(n7608), .C(n7620) );
  BUFFD0 U7536 ( .I(n7554), .Z(n7621) );
  CKBD0 U7537 ( .CLK(n7555), .C(n7622) );
  CKBD0 U7538 ( .CLK(n7556), .C(n7623) );
  CKBD0 U7539 ( .CLK(n7565), .C(n7624) );
  CKBD0 U7540 ( .CLK(n7613), .C(n7625) );
  CKBD0 U7541 ( .CLK(n7614), .C(n7626) );
  CKBD0 U7542 ( .CLK(n7615), .C(n7627) );
  CKBD0 U7543 ( .CLK(n7616), .C(n7628) );
  CKBD0 U7544 ( .CLK(n7617), .C(n7629) );
  CKBD0 U7545 ( .CLK(n7618), .C(n7630) );
  CKBD0 U7546 ( .CLK(n7619), .C(n7631) );
  CKBD0 U7547 ( .CLK(n7620), .C(n7632) );
  CKBD0 U7548 ( .CLK(n7566), .C(n7633) );
  CKBD0 U7549 ( .CLK(n7625), .C(n7634) );
  CKBD0 U7550 ( .CLK(n7626), .C(n7635) );
  CKBD0 U7551 ( .CLK(n7627), .C(n7636) );
  CKBD0 U7552 ( .CLK(n7628), .C(n7637) );
  CKBD0 U7553 ( .CLK(n7629), .C(n7638) );
  CKBD0 U7554 ( .CLK(n7630), .C(n7639) );
  CKBD0 U7555 ( .CLK(n7631), .C(n7640) );
  CKBD0 U7556 ( .CLK(n7632), .C(n7641) );
  CKBD0 U7557 ( .CLK(n7568), .C(n7642) );
  CKBD0 U7558 ( .CLK(n7634), .C(n7643) );
  CKBD0 U7559 ( .CLK(n7635), .C(n7644) );
  CKBD0 U7560 ( .CLK(n7636), .C(n7645) );
  CKBD0 U7561 ( .CLK(n7637), .C(n7646) );
  CKBD0 U7562 ( .CLK(n7638), .C(n7647) );
  CKBD0 U7563 ( .CLK(n7639), .C(n7648) );
  CKBD0 U7564 ( .CLK(n7640), .C(n7649) );
  CKBD0 U7565 ( .CLK(n7641), .C(n7650) );
  CKBD0 U7566 ( .CLK(n7643), .C(n7651) );
  CKBD0 U7567 ( .CLK(n7644), .C(n7652) );
  CKBD0 U7568 ( .CLK(n7645), .C(n7653) );
  CKBD0 U7569 ( .CLK(n7646), .C(n7654) );
  CKBD0 U7570 ( .CLK(n7571), .C(n7655) );
  CKBD0 U7571 ( .CLK(n7647), .C(n7656) );
  CKBD0 U7572 ( .CLK(n7574), .C(n7657) );
  CKBD0 U7573 ( .CLK(n7581), .C(n7658) );
  CKBD0 U7574 ( .CLK(n7582), .C(n7659) );
  CKBD0 U7575 ( .CLK(n7648), .C(n7660) );
  CKBD0 U7576 ( .CLK(n7649), .C(n7661) );
  BUFFD0 U7577 ( .I(n7650), .Z(n7662) );
  BUFFD0 U7578 ( .I(n7651), .Z(n7663) );
  BUFFD0 U7579 ( .I(n7652), .Z(n7664) );
  CKBD0 U7580 ( .CLK(n7653), .C(n7665) );
  BUFFD0 U7581 ( .I(n7654), .Z(n7666) );
  CKBD0 U7582 ( .CLK(n7656), .C(n7667) );
  BUFFD0 U7583 ( .I(n7583), .Z(n7668) );
  BUFFD0 U7584 ( .I(n7584), .Z(n7669) );
  BUFFD0 U7585 ( .I(n7585), .Z(n7670) );
  CKBD0 U7586 ( .CLK(n7594), .C(n7671) );
  CKBD0 U7587 ( .CLK(n7596), .C(n7672) );
  BUFFD0 U7588 ( .I(n7595), .Z(n7673) );
  BUFFD0 U7589 ( .I(n7660), .Z(n7674) );
  CKBD0 U7590 ( .CLK(n7661), .C(n7675) );
  CKBD0 U7591 ( .CLK(n7662), .C(n7676) );
  CKBD0 U7592 ( .CLK(n7663), .C(n7677) );
  CKBD0 U7593 ( .CLK(n7664), .C(n7678) );
  CKBD0 U7594 ( .CLK(n7665), .C(n7679) );
  CKBD0 U7595 ( .CLK(n7666), .C(n7680) );
  CKBD0 U7596 ( .CLK(n7667), .C(n7681) );
  BUFFD0 U7597 ( .I(n7597), .Z(n7682) );
  CKBD0 U7598 ( .CLK(n7598), .C(n7683) );
  CKBD0 U7599 ( .CLK(n7599), .C(n7684) );
  CKBD0 U7600 ( .CLK(n7602), .C(n7685) );
  CKBD0 U7601 ( .CLK(n7609), .C(n7686) );
  CKBD0 U7602 ( .CLK(n7610), .C(n7687) );
  CKBD0 U7603 ( .CLK(n7611), .C(n7688) );
  CKBD0 U7604 ( .CLK(n7674), .C(n7689) );
  CKBD0 U7605 ( .CLK(n7612), .C(n7690) );
  CKBD0 U7606 ( .CLK(n7621), .C(n7691) );
  CKBD0 U7607 ( .CLK(n7622), .C(n7692) );
  CKBD0 U7608 ( .CLK(n7675), .C(n7693) );
  CKBD0 U7609 ( .CLK(n7676), .C(n7694) );
  CKBD0 U7610 ( .CLK(n7677), .C(n7695) );
  CKBD0 U7611 ( .CLK(n7678), .C(n7696) );
  CKBD0 U7612 ( .CLK(n7679), .C(n7697) );
  CKBD0 U7613 ( .CLK(n7680), .C(n7698) );
  BUFFD0 U7614 ( .I(n7681), .Z(n7699) );
  CKBD0 U7615 ( .CLK(n7689), .C(n7700) );
  CKBD0 U7616 ( .CLK(n7623), .C(n7701) );
  CKBD0 U7617 ( .CLK(n7624), .C(n7702) );
  BUFFD0 U7618 ( .I(n7693), .Z(n7703) );
  CKBD0 U7619 ( .CLK(n7694), .C(n7704) );
  CKBD0 U7620 ( .CLK(n7695), .C(n7705) );
  CKBD0 U7621 ( .CLK(n7696), .C(n7706) );
  BUFFD0 U7622 ( .I(n7697), .Z(n7707) );
  CKBD0 U7623 ( .CLK(n7698), .C(n7708) );
  CKBD0 U7624 ( .CLK(n7699), .C(n7709) );
  CKBD0 U7625 ( .CLK(n7633), .C(n7710) );
  CKBD0 U7626 ( .CLK(n7700), .C(n7711) );
  BUFFD0 U7627 ( .I(n7642), .Z(n7712) );
  CKBD0 U7628 ( .CLK(n7703), .C(n7713) );
  CKBD0 U7629 ( .CLK(n7704), .C(n7714) );
  CKBD0 U7630 ( .CLK(n7705), .C(n7715) );
  CKBD0 U7631 ( .CLK(n7706), .C(n7716) );
  CKBD0 U7632 ( .CLK(n7707), .C(n7717) );
  CKBD0 U7633 ( .CLK(n7708), .C(n7718) );
  CKBD0 U7634 ( .CLK(n7709), .C(n7719) );
  CKBD0 U7635 ( .CLK(n7711), .C(n7720) );
  CKBD0 U7636 ( .CLK(n7713), .C(n7721) );
  CKBD0 U7637 ( .CLK(n7655), .C(n7722) );
  CKBD0 U7638 ( .CLK(n7714), .C(n7723) );
  CKBD0 U7639 ( .CLK(n7657), .C(n7724) );
  CKBD0 U7640 ( .CLK(n7658), .C(n7725) );
  CKBD0 U7641 ( .CLK(n7659), .C(n7726) );
  CKBD0 U7642 ( .CLK(n7668), .C(n7727) );
  CKBD0 U7643 ( .CLK(n7715), .C(n7728) );
  CKBD0 U7644 ( .CLK(n7716), .C(n7729) );
  CKBD0 U7645 ( .CLK(n7669), .C(n7730) );
  CKBD0 U7646 ( .CLK(n7717), .C(n7731) );
  CKBD0 U7647 ( .CLK(n7718), .C(n7732) );
  CKBD0 U7648 ( .CLK(n7719), .C(n7733) );
  CKBD0 U7649 ( .CLK(n7720), .C(n7734) );
  CKBD0 U7650 ( .CLK(n7721), .C(n7735) );
  CKBD0 U7651 ( .CLK(n7723), .C(n7736) );
  CKBD0 U7652 ( .CLK(n7670), .C(n7737) );
  CKBD0 U7653 ( .CLK(n7671), .C(n7738) );
  CKBD0 U7654 ( .CLK(n7672), .C(n7739) );
  CKBD0 U7655 ( .CLK(n7673), .C(n7740) );
  CKBD0 U7656 ( .CLK(n7682), .C(n7741) );
  CKBD0 U7657 ( .CLK(n7728), .C(n7742) );
  CKBD0 U7658 ( .CLK(n7729), .C(n7743) );
  CKBD0 U7659 ( .CLK(n7683), .C(n7744) );
  CKBD0 U7660 ( .CLK(n7731), .C(n7745) );
  CKBD0 U7661 ( .CLK(n7732), .C(n7746) );
  CKBD0 U7662 ( .CLK(n7733), .C(n7747) );
  CKBD0 U7663 ( .CLK(n7734), .C(n7748) );
  CKBD0 U7664 ( .CLK(n7735), .C(n7749) );
  CKBD0 U7665 ( .CLK(n7736), .C(n7750) );
  CKBD0 U7666 ( .CLK(n7684), .C(n7751) );
  CKBD0 U7667 ( .CLK(n7685), .C(n7752) );
  CKBD0 U7668 ( .CLK(n7686), .C(n7753) );
  CKBD0 U7669 ( .CLK(n7687), .C(n7754) );
  CKBD0 U7670 ( .CLK(n7688), .C(n7755) );
  CKBD0 U7671 ( .CLK(n7742), .C(n7756) );
  CKBD0 U7672 ( .CLK(n7743), .C(n7757) );
  CKBD0 U7673 ( .CLK(n7745), .C(n7758) );
  CKBD0 U7674 ( .CLK(n7746), .C(n7759) );
  CKBD0 U7675 ( .CLK(n7747), .C(n7760) );
  CKBD0 U7676 ( .CLK(n7748), .C(n7761) );
  CKBD0 U7677 ( .CLK(n7749), .C(n7762) );
  CKBD0 U7678 ( .CLK(n7750), .C(n7763) );
  CKBD0 U7679 ( .CLK(n7690), .C(n7764) );
  CKBD0 U7680 ( .CLK(n7691), .C(n7765) );
  CKBD0 U7681 ( .CLK(n7692), .C(n7766) );
  CKBD0 U7682 ( .CLK(n7756), .C(n7767) );
  CKBD0 U7683 ( .CLK(n7757), .C(n7768) );
  CKBD0 U7684 ( .CLK(n7701), .C(n7769) );
  CKBD0 U7685 ( .CLK(n7758), .C(n7770) );
  CKBD0 U7686 ( .CLK(n7759), .C(n7771) );
  CKBD0 U7687 ( .CLK(n7760), .C(n7772) );
  CKBD0 U7688 ( .CLK(n7761), .C(n7773) );
  CKBD0 U7689 ( .CLK(n7762), .C(n7774) );
  CKBD0 U7690 ( .CLK(n7763), .C(n7775) );
  CKBD0 U7691 ( .CLK(n7702), .C(n7776) );
  CKBD0 U7692 ( .CLK(n7767), .C(n7777) );
  CKBD0 U7693 ( .CLK(n7768), .C(n7778) );
  CKBD0 U7694 ( .CLK(n7770), .C(n7779) );
  CKBD0 U7695 ( .CLK(n7771), .C(n7780) );
  CKBD0 U7696 ( .CLK(n7772), .C(n7781) );
  CKBD0 U7697 ( .CLK(n7773), .C(n7782) );
  CKBD0 U7698 ( .CLK(n7774), .C(n7783) );
  CKBD0 U7699 ( .CLK(n7775), .C(n7784) );
  CKBD0 U7700 ( .CLK(n7710), .C(n7785) );
  CKBD0 U7701 ( .CLK(n7712), .C(n7786) );
  CKBD0 U7702 ( .CLK(n7777), .C(n7787) );
  CKBD0 U7703 ( .CLK(n7778), .C(n7788) );
  CKBD0 U7704 ( .CLK(n7779), .C(n7789) );
  CKBD0 U7705 ( .CLK(n7780), .C(n7790) );
  CKBD0 U7706 ( .CLK(n7781), .C(n7791) );
  BUFFD0 U7707 ( .I(n7782), .Z(n7792) );
  CKBD0 U7708 ( .CLK(n7783), .C(n7793) );
  BUFFD0 U7709 ( .I(n7784), .Z(n7794) );
  BUFFD0 U7710 ( .I(n7787), .Z(n7795) );
  BUFFD0 U7711 ( .I(n7788), .Z(n7796) );
  CKBD0 U7712 ( .CLK(n7789), .C(n7797) );
  BUFFD0 U7713 ( .I(n7790), .Z(n7798) );
  CKBD0 U7714 ( .CLK(n7791), .C(n7799) );
  CKBD0 U7715 ( .CLK(n7792), .C(n7800) );
  CKBD0 U7716 ( .CLK(n7793), .C(n7801) );
  CKBD0 U7717 ( .CLK(n7794), .C(n7802) );
  CKBD0 U7718 ( .CLK(n7795), .C(n7803) );
  CKBD0 U7719 ( .CLK(n7796), .C(n7804) );
  CKBD0 U7720 ( .CLK(n7797), .C(n7805) );
  CKBD0 U7721 ( .CLK(n7798), .C(n7806) );
  CKBD0 U7722 ( .CLK(n7722), .C(n7807) );
  CKBD0 U7723 ( .CLK(n7799), .C(n7808) );
  CKBD0 U7724 ( .CLK(n7724), .C(n7809) );
  CKBD0 U7725 ( .CLK(n7725), .C(n7810) );
  CKBD0 U7726 ( .CLK(n7726), .C(n7811) );
  CKBD0 U7727 ( .CLK(n7727), .C(n7812) );
  CKBD0 U7728 ( .CLK(n7730), .C(n7813) );
  CKBD0 U7729 ( .CLK(n7737), .C(n7814) );
  CKBD0 U7730 ( .CLK(n7738), .C(n7815) );
  CKBD0 U7731 ( .CLK(n7800), .C(n7816) );
  CKBD0 U7732 ( .CLK(n7739), .C(n7817) );
  CKBD0 U7733 ( .CLK(n7740), .C(n7818) );
  CKBD0 U7734 ( .CLK(n7741), .C(n7819) );
  CKBD0 U7735 ( .CLK(n7744), .C(n7820) );
  CKBD0 U7736 ( .CLK(n7751), .C(n7821) );
  CKBD0 U7737 ( .CLK(n7752), .C(n7822) );
  CKBD0 U7738 ( .CLK(n7801), .C(n7823) );
  CKBD0 U7739 ( .CLK(n7802), .C(n7824) );
  CKBD0 U7740 ( .CLK(n7803), .C(n7825) );
  CKBD0 U7741 ( .CLK(n7804), .C(n7826) );
  BUFFD0 U7742 ( .I(n7805), .Z(n7827) );
  CKBD0 U7743 ( .CLK(n7806), .C(n7828) );
  BUFFD0 U7744 ( .I(n7808), .Z(n7829) );
  CKBD0 U7745 ( .CLK(n7816), .C(n7830) );
  CKBD0 U7746 ( .CLK(n7753), .C(n7831) );
  CKBD0 U7747 ( .CLK(n7754), .C(n7832) );
  CKBD0 U7748 ( .CLK(n7755), .C(n7833) );
  CKBD0 U7749 ( .CLK(n7764), .C(n7834) );
  BUFFD0 U7750 ( .I(n7823), .Z(n7835) );
  CKBD0 U7751 ( .CLK(n7765), .C(n7836) );
  CKBD0 U7752 ( .CLK(n7824), .C(n7837) );
  CKBD0 U7753 ( .CLK(n7825), .C(n7838) );
  CKBD0 U7754 ( .CLK(n7826), .C(n7839) );
  CKBD0 U7755 ( .CLK(n7827), .C(n7840) );
  CKBD0 U7756 ( .CLK(n7828), .C(n7841) );
  CKBD0 U7757 ( .CLK(n7829), .C(n7842) );
  CKBD0 U7758 ( .CLK(n7830), .C(n7843) );
  CKBD0 U7759 ( .CLK(n7766), .C(n7844) );
  CKBD0 U7760 ( .CLK(n7769), .C(n7845) );
  CKBD0 U7761 ( .CLK(n7776), .C(n7846) );
  CKBD0 U7762 ( .CLK(n7835), .C(n7847) );
  CKBD0 U7763 ( .CLK(n7837), .C(n7848) );
  CKBD0 U7764 ( .CLK(n7838), .C(n7849) );
  CKBD0 U7765 ( .CLK(n7839), .C(n7850) );
  CKBD0 U7766 ( .CLK(n7840), .C(n7851) );
  CKBD0 U7767 ( .CLK(n7841), .C(n7852) );
  CKBD0 U7768 ( .CLK(n7842), .C(n7853) );
  CKBD0 U7769 ( .CLK(n7843), .C(n7854) );
  CKBD0 U7770 ( .CLK(n7785), .C(n7855) );
  CKBD0 U7771 ( .CLK(n7786), .C(n7856) );
  CKBD0 U7772 ( .CLK(n7847), .C(n7857) );
  CKBD0 U7773 ( .CLK(n7848), .C(n7858) );
  CKBD0 U7774 ( .CLK(n7849), .C(n7859) );
  CKBD0 U7775 ( .CLK(n7850), .C(n7860) );
  CKBD0 U7776 ( .CLK(n7851), .C(n7861) );
  CKBD0 U7777 ( .CLK(n7852), .C(n7862) );
  CKBD0 U7778 ( .CLK(n7853), .C(n7863) );
  CKBD0 U7779 ( .CLK(n7854), .C(n7864) );
  CKBD0 U7780 ( .CLK(n7857), .C(n7865) );
  CKBD0 U7781 ( .CLK(n7807), .C(n7866) );
  CKBD0 U7782 ( .CLK(n7858), .C(n7867) );
  CKBD0 U7783 ( .CLK(n7809), .C(n7868) );
  CKBD0 U7784 ( .CLK(n7810), .C(n7869) );
  CKBD0 U7785 ( .CLK(n7859), .C(n7870) );
  CKBD0 U7786 ( .CLK(n7860), .C(n7871) );
  CKBD0 U7787 ( .CLK(n7861), .C(n7872) );
  CKBD0 U7788 ( .CLK(n7862), .C(n7873) );
  CKBD0 U7789 ( .CLK(n7863), .C(n7874) );
  CKBD0 U7790 ( .CLK(n7864), .C(n7875) );
  CKBD0 U7791 ( .CLK(n7865), .C(n7876) );
  CKBD0 U7792 ( .CLK(n7867), .C(n7877) );
  CKBD0 U7793 ( .CLK(n7811), .C(n7878) );
  CKBD0 U7794 ( .CLK(n7812), .C(n7879) );
  CKBD0 U7795 ( .CLK(n7813), .C(n7880) );
  CKBD0 U7796 ( .CLK(n7814), .C(n7881) );
  CKBD0 U7797 ( .CLK(n7815), .C(n7882) );
  CKBD0 U7798 ( .CLK(n7817), .C(n7883) );
  CKBD0 U7799 ( .CLK(n7870), .C(n7884) );
  CKBD0 U7800 ( .CLK(n7818), .C(n7885) );
  CKBD0 U7801 ( .CLK(n7871), .C(n7886) );
  CKBD0 U7802 ( .CLK(n7872), .C(n7887) );
  CKBD0 U7803 ( .CLK(n7873), .C(n7888) );
  CKBD0 U7804 ( .CLK(n7874), .C(n7889) );
  CKBD0 U7805 ( .CLK(n7875), .C(n7890) );
  CKBD0 U7806 ( .CLK(n7876), .C(n7891) );
  CKBD0 U7807 ( .CLK(n7877), .C(n7892) );
  CKBD0 U7808 ( .CLK(n7819), .C(n7893) );
  CKBD0 U7809 ( .CLK(n7820), .C(n7894) );
  CKBD0 U7810 ( .CLK(n7821), .C(n7895) );
  CKBD0 U7811 ( .CLK(n7822), .C(n7896) );
  CKBD0 U7812 ( .CLK(n7831), .C(n7897) );
  CKBD0 U7813 ( .CLK(n7832), .C(n7898) );
  CKBD0 U7814 ( .CLK(n7884), .C(n7899) );
  CKBD0 U7815 ( .CLK(n7886), .C(n7900) );
  CKBD0 U7816 ( .CLK(n7887), .C(n7901) );
  CKBD0 U7817 ( .CLK(n7888), .C(n7902) );
  CKBD0 U7818 ( .CLK(n7889), .C(n7903) );
  CKBD0 U7819 ( .CLK(n7890), .C(n7904) );
  CKBD0 U7820 ( .CLK(n7891), .C(n7905) );
  CKBD0 U7821 ( .CLK(n7892), .C(n7906) );
  CKBD0 U7822 ( .CLK(n7833), .C(n7907) );
  CKBD0 U7823 ( .CLK(n7834), .C(n7908) );
  CKBD0 U7824 ( .CLK(n7836), .C(n7909) );
  CKBD0 U7825 ( .CLK(n7899), .C(n7910) );
  CKBD0 U7826 ( .CLK(n7900), .C(n7911) );
  CKBD0 U7827 ( .CLK(n7901), .C(n7912) );
  CKBD0 U7828 ( .CLK(n7902), .C(n7913) );
  CKBD0 U7829 ( .CLK(n7903), .C(n7914) );
  CKBD0 U7830 ( .CLK(n7904), .C(n7915) );
  CKBD0 U7831 ( .CLK(n7905), .C(n7916) );
  CKBD0 U7832 ( .CLK(n7906), .C(n7917) );
  CKBD0 U7833 ( .CLK(n7910), .C(n7918) );
  CKBD0 U7834 ( .CLK(n7911), .C(n7919) );
  CKBD0 U7835 ( .CLK(n7912), .C(n7920) );
  CKBD0 U7836 ( .CLK(n7913), .C(n7921) );
  CKBD0 U7837 ( .CLK(n7914), .C(n7922) );
  BUFFD0 U7838 ( .I(n7915), .Z(n7923) );
  CKBD0 U7839 ( .CLK(n7916), .C(n7924) );
  BUFFD0 U7840 ( .I(n7917), .Z(n7925) );
  CKBD0 U7841 ( .CLK(n7844), .C(n7926) );
  CKBD0 U7842 ( .CLK(n7845), .C(n7927) );
  CKBD0 U7843 ( .CLK(n7846), .C(n7928) );
  BUFFD0 U7844 ( .I(n7918), .Z(n7929) );
  BUFFD0 U7845 ( .I(n7919), .Z(n7930) );
  CKBD0 U7846 ( .CLK(n7920), .C(n7931) );
  BUFFD0 U7847 ( .I(n7921), .Z(n7932) );
  CKBD0 U7848 ( .CLK(n7922), .C(n7933) );
  CKBD0 U7849 ( .CLK(n7923), .C(n7934) );
  CKBD0 U7850 ( .CLK(n7924), .C(n7935) );
  CKBD0 U7851 ( .CLK(n7925), .C(n7936) );
  CKBD0 U7852 ( .CLK(n7855), .C(n7937) );
  CKBD0 U7853 ( .CLK(n7856), .C(n7938) );
  CKBD0 U7854 ( .CLK(n7929), .C(n7939) );
  CKBD0 U7855 ( .CLK(n7930), .C(n7940) );
  CKBD0 U7856 ( .CLK(n7931), .C(n7941) );
  CKBD0 U7857 ( .CLK(n7932), .C(n7942) );
  CKBD0 U7858 ( .CLK(n7933), .C(n7943) );
  CKBD0 U7859 ( .CLK(n7866), .C(n7944) );
  CKBD0 U7860 ( .CLK(n7934), .C(n7945) );
  CKBD0 U7861 ( .CLK(n7868), .C(n7946) );
  CKBD0 U7862 ( .CLK(n7869), .C(n7947) );
  CKBD0 U7863 ( .CLK(n7878), .C(n7948) );
  CKBD0 U7864 ( .CLK(n7879), .C(n7949) );
  BUFFD0 U7865 ( .I(n7935), .Z(n7950) );
  CKBD0 U7866 ( .CLK(n7880), .C(n7951) );
  CKBD0 U7867 ( .CLK(n7936), .C(n7952) );
  CKBD0 U7868 ( .CLK(n7939), .C(n7953) );
  CKBD0 U7869 ( .CLK(n7940), .C(n7954) );
  BUFFD0 U7870 ( .I(n7941), .Z(n7955) );
  CKBD0 U7871 ( .CLK(n7942), .C(n7956) );
  BUFFD0 U7872 ( .I(n7943), .Z(n7957) );
  CKBD0 U7873 ( .CLK(n7945), .C(n7958) );
  CKBD0 U7874 ( .CLK(n7881), .C(n7959) );
  CKBD0 U7875 ( .CLK(n7882), .C(n7960) );
  CKBD0 U7876 ( .CLK(n7883), .C(n7961) );
  CKBD0 U7877 ( .CLK(n7885), .C(n7962) );
  CKBD0 U7878 ( .CLK(n7893), .C(n7963) );
  CKBD0 U7879 ( .CLK(n7894), .C(n7964) );
  CKBD0 U7880 ( .CLK(n7950), .C(n7965) );
  CKBD0 U7881 ( .CLK(n7952), .C(n7966) );
  CKBD0 U7882 ( .CLK(n7953), .C(n7967) );
  CKBD0 U7883 ( .CLK(n7954), .C(n7968) );
  CKBD0 U7884 ( .CLK(n7955), .C(n7969) );
  CKBD0 U7885 ( .CLK(n7956), .C(n7970) );
  CKBD0 U7886 ( .CLK(n7957), .C(n7971) );
  CKBD0 U7887 ( .CLK(n7958), .C(n7972) );
  CKBD0 U7888 ( .CLK(n7895), .C(n7973) );
  CKBD0 U7889 ( .CLK(n7896), .C(n7974) );
  CKBD0 U7890 ( .CLK(n7897), .C(n7975) );
  CKBD0 U7891 ( .CLK(n7898), .C(n7976) );
  CKBD0 U7892 ( .CLK(n7907), .C(n7977) );
  CKBD0 U7893 ( .CLK(n7965), .C(n7978) );
  CKBD0 U7894 ( .CLK(n7908), .C(n7979) );
  CKBD0 U7895 ( .CLK(n7966), .C(n7980) );
  CKBD0 U7896 ( .CLK(n7967), .C(n7981) );
  CKBD0 U7897 ( .CLK(n7968), .C(n7982) );
  CKBD0 U7898 ( .CLK(n7969), .C(n7983) );
  CKBD0 U7899 ( .CLK(n7970), .C(n7984) );
  CKBD0 U7900 ( .CLK(n7971), .C(n7985) );
  CKBD0 U7901 ( .CLK(n7972), .C(n7986) );
  CKBD0 U7902 ( .CLK(n7909), .C(n7987) );
  CKBD0 U7903 ( .CLK(n7926), .C(n7988) );
  CKBD0 U7904 ( .CLK(n7978), .C(n7989) );
  CKBD0 U7905 ( .CLK(n7980), .C(n7990) );
  CKBD0 U7906 ( .CLK(n7981), .C(n7991) );
  CKBD0 U7907 ( .CLK(n7982), .C(n7992) );
  CKBD0 U7908 ( .CLK(n7983), .C(n7993) );
  CKBD0 U7909 ( .CLK(n7984), .C(n7994) );
  CKBD0 U7910 ( .CLK(n7985), .C(n7995) );
  CKBD0 U7911 ( .CLK(n7986), .C(n7996) );
  CKBD0 U7912 ( .CLK(n7927), .C(n7997) );
  CKBD0 U7913 ( .CLK(n7928), .C(n7998) );
  CKBD0 U7914 ( .CLK(n7989), .C(n7999) );
  CKBD0 U7915 ( .CLK(n7990), .C(n8000) );
  CKBD0 U7916 ( .CLK(n7991), .C(n8001) );
  CKBD0 U7917 ( .CLK(n7992), .C(n8002) );
  CKBD0 U7918 ( .CLK(n7993), .C(n8003) );
  CKBD0 U7919 ( .CLK(n7994), .C(n8004) );
  CKBD0 U7920 ( .CLK(n7995), .C(n8005) );
  CKBD0 U7921 ( .CLK(n7937), .C(n8006) );
  CKBD0 U7922 ( .CLK(n7996), .C(n8007) );
  CKBD0 U7923 ( .CLK(n7938), .C(n8008) );
  CKBD0 U7924 ( .CLK(n7999), .C(n8009) );
  CKBD0 U7925 ( .CLK(n8000), .C(n8010) );
  CKBD0 U7926 ( .CLK(n7944), .C(n8011) );
  CKBD0 U7927 ( .CLK(n8001), .C(n8012) );
  CKBD0 U7928 ( .CLK(n8002), .C(n8013) );
  CKBD0 U7929 ( .CLK(n7946), .C(n8014) );
  CKBD0 U7930 ( .CLK(n8003), .C(n8015) );
  CKBD0 U7931 ( .CLK(n8004), .C(n8016) );
  CKBD0 U7932 ( .CLK(n8005), .C(n8017) );
  CKBD0 U7933 ( .CLK(n8007), .C(n8018) );
  CKBD0 U7934 ( .CLK(n8009), .C(n8019) );
  CKBD0 U7935 ( .CLK(n8010), .C(n8020) );
  CKBD0 U7936 ( .CLK(n7947), .C(n8021) );
  CKBD0 U7937 ( .CLK(n7948), .C(n8022) );
  CKBD0 U7938 ( .CLK(n7949), .C(n8023) );
  CKBD0 U7939 ( .CLK(n7951), .C(n8024) );
  CKBD0 U7940 ( .CLK(n7959), .C(n8025) );
  CKBD0 U7941 ( .CLK(n8012), .C(n8026) );
  CKBD0 U7942 ( .CLK(n8013), .C(n8027) );
  CKBD0 U7943 ( .CLK(n8015), .C(n8028) );
  CKBD0 U7944 ( .CLK(n8016), .C(n8029) );
  CKBD0 U7945 ( .CLK(n8017), .C(n8030) );
  CKBD0 U7946 ( .CLK(n8018), .C(n8031) );
  CKBD0 U7947 ( .CLK(n8019), .C(n8032) );
  CKBD0 U7948 ( .CLK(n8020), .C(n8033) );
  CKBD0 U7949 ( .CLK(n7960), .C(n8034) );
  CKBD0 U7950 ( .CLK(n7961), .C(n8035) );
  CKBD0 U7951 ( .CLK(n7962), .C(n8036) );
  CKBD0 U7952 ( .CLK(n7963), .C(n8037) );
  CKBD0 U7953 ( .CLK(n7964), .C(n8038) );
  CKBD0 U7954 ( .CLK(n8026), .C(n8039) );
  CKBD0 U7955 ( .CLK(n8027), .C(n8040) );
  CKBD0 U7956 ( .CLK(n8028), .C(n8041) );
  CKBD0 U7957 ( .CLK(n8029), .C(n8042) );
  CKBD0 U7958 ( .CLK(n8030), .C(n8043) );
  CKBD0 U7959 ( .CLK(n8031), .C(n8044) );
  CKBD0 U7960 ( .CLK(n8032), .C(n8045) );
  CKBD0 U7961 ( .CLK(n8033), .C(n8046) );
  CKBD0 U7962 ( .CLK(n7973), .C(n8047) );
  CKBD0 U7963 ( .CLK(n8039), .C(n8048) );
  CKBD0 U7964 ( .CLK(n8040), .C(n8049) );
  CKBD0 U7965 ( .CLK(n8041), .C(n8050) );
  CKBD0 U7966 ( .CLK(n8042), .C(n8051) );
  CKBD0 U7967 ( .CLK(n8043), .C(n8052) );
  BUFFD0 U7968 ( .I(n8044), .Z(n8053) );
  CKBD0 U7969 ( .CLK(n8045), .C(n8054) );
  BUFFD0 U7970 ( .I(n8046), .Z(n8055) );
  CKBD0 U7971 ( .CLK(n7974), .C(n8056) );
  CKBD0 U7972 ( .CLK(n7975), .C(n8057) );
  CKBD0 U7973 ( .CLK(n7976), .C(n8058) );
  CKBD0 U7974 ( .CLK(n7977), .C(n8059) );
  CKBD0 U7975 ( .CLK(n7979), .C(n8060) );
  BUFFD0 U7976 ( .I(n8048), .Z(n8061) );
  BUFFD0 U7977 ( .I(n8049), .Z(n8062) );
  CKBD0 U7978 ( .CLK(n8050), .C(n8063) );
  BUFFD0 U7979 ( .I(n8051), .Z(n8064) );
  CKBD0 U7980 ( .CLK(n8052), .C(n8065) );
  CKBD0 U7981 ( .CLK(n8053), .C(n8066) );
  CKBD0 U7982 ( .CLK(n8054), .C(n8067) );
  CKBD0 U7983 ( .CLK(n8055), .C(n8068) );
  CKBD0 U7984 ( .CLK(n7987), .C(n8069) );
  CKBD0 U7985 ( .CLK(n7988), .C(n8070) );
  CKBD0 U7986 ( .CLK(n8061), .C(n8071) );
  CKBD0 U7987 ( .CLK(n8062), .C(n8072) );
  CKBD0 U7988 ( .CLK(n8063), .C(n8073) );
  CKBD0 U7989 ( .CLK(n8064), .C(n8074) );
  CKBD0 U7990 ( .CLK(n8065), .C(n8075) );
  CKBD0 U7991 ( .CLK(n8066), .C(n8076) );
  BUFFD0 U7992 ( .I(n8067), .Z(n8077) );
  CKBD0 U7993 ( .CLK(n8068), .C(n8078) );
  CKBD0 U7994 ( .CLK(n7997), .C(n8079) );
  CKBD0 U7995 ( .CLK(n7998), .C(n8080) );
  CKBD0 U7996 ( .CLK(n8006), .C(n8081) );
  CKBD0 U7997 ( .CLK(n8071), .C(n8082) );
  CKBD0 U7998 ( .CLK(n8072), .C(n8083) );
  CKBD0 U7999 ( .CLK(n8008), .C(n8084) );
  BUFFD0 U8000 ( .I(n8073), .Z(n8085) );
  CKBD0 U8001 ( .CLK(n8074), .C(n8086) );
  BUFFD0 U8002 ( .I(n8075), .Z(n8087) );
  CKBD0 U8003 ( .CLK(n8011), .C(n8088) );
  CKBD0 U8004 ( .CLK(n8076), .C(n8089) );
  CKBD0 U8005 ( .CLK(n8014), .C(n8090) );
  CKBD0 U8006 ( .CLK(n8021), .C(n8091) );
  CKBD0 U8007 ( .CLK(n8022), .C(n8092) );
  CKBD0 U8008 ( .CLK(n8077), .C(n8093) );
  CKBD0 U8009 ( .CLK(n8078), .C(n8094) );
  CKBD0 U8010 ( .CLK(n8082), .C(n8095) );
  CKBD0 U8011 ( .CLK(n8083), .C(n8096) );
  CKBD0 U8012 ( .CLK(n8085), .C(n8097) );
  CKBD0 U8013 ( .CLK(n8086), .C(n8098) );
  CKBD0 U8014 ( .CLK(n8087), .C(n8099) );
  CKBD0 U8015 ( .CLK(n8089), .C(n8100) );
  CKBD0 U8016 ( .CLK(n8023), .C(n8101) );
  CKBD0 U8017 ( .CLK(n8024), .C(n8102) );
  CKBD0 U8018 ( .CLK(n8025), .C(n8103) );
  CKBD0 U8019 ( .CLK(n8034), .C(n8104) );
  CKBD0 U8020 ( .CLK(n8035), .C(n8105) );
  CKBD0 U8021 ( .CLK(n8036), .C(n8106) );
  CKBD0 U8022 ( .CLK(n8093), .C(n8107) );
  CKBD0 U8023 ( .CLK(n8038), .C(n8108) );
  CKBD0 U8024 ( .CLK(n8094), .C(n8109) );
  CKBD0 U8025 ( .CLK(n8095), .C(n8110) );
  CKBD0 U8026 ( .CLK(n8096), .C(n8111) );
  CKBD0 U8027 ( .CLK(n8097), .C(n8112) );
  CKBD0 U8028 ( .CLK(n8098), .C(n8113) );
  CKBD0 U8029 ( .CLK(n8099), .C(n8114) );
  CKBD0 U8030 ( .CLK(n8100), .C(n8115) );
  CKBD0 U8031 ( .CLK(n8037), .C(n8116) );
  CKBD0 U8032 ( .CLK(n8047), .C(n8117) );
  CKBD0 U8033 ( .CLK(n8057), .C(n8118) );
  CKBD0 U8034 ( .CLK(n8056), .C(n8119) );
  CKBD0 U8035 ( .CLK(n8058), .C(n8120) );
  CKBD0 U8036 ( .CLK(n8059), .C(n8121) );
  CKBD0 U8037 ( .CLK(n8107), .C(n8122) );
  CKBD0 U8038 ( .CLK(n8109), .C(n8123) );
  CKBD0 U8039 ( .CLK(n8110), .C(n8124) );
  CKBD0 U8040 ( .CLK(n8111), .C(n8125) );
  CKBD0 U8041 ( .CLK(n8112), .C(n8126) );
  CKBD0 U8042 ( .CLK(n8113), .C(n8127) );
  CKBD0 U8043 ( .CLK(n8114), .C(n8128) );
  CKBD0 U8044 ( .CLK(n8115), .C(n8129) );
  CKBD0 U8045 ( .CLK(n8060), .C(n8130) );
  CKBD0 U8046 ( .CLK(n8069), .C(n8131) );
  CKBD0 U8047 ( .CLK(n8070), .C(n8132) );
  CKBD0 U8048 ( .CLK(n8122), .C(n8133) );
  CKBD0 U8049 ( .CLK(n8123), .C(n8134) );
  CKBD0 U8050 ( .CLK(n8124), .C(n8135) );
  CKBD0 U8051 ( .CLK(n8125), .C(n8136) );
  CKBD0 U8052 ( .CLK(n8126), .C(n8137) );
  CKBD0 U8053 ( .CLK(n8127), .C(n8138) );
  CKBD0 U8054 ( .CLK(n8128), .C(n8139) );
  CKBD0 U8055 ( .CLK(n8129), .C(n8140) );
  CKBD0 U8056 ( .CLK(n8079), .C(n8141) );
  CKBD0 U8057 ( .CLK(n8080), .C(n8142) );
  CKBD0 U8058 ( .CLK(n8133), .C(n8143) );
  CKBD0 U8059 ( .CLK(n8134), .C(n8144) );
  CKBD0 U8060 ( .CLK(n8135), .C(n8145) );
  CKBD0 U8061 ( .CLK(n8136), .C(n8146) );
  CKBD0 U8062 ( .CLK(n8137), .C(n8147) );
  CKBD0 U8063 ( .CLK(n8138), .C(n8148) );
  CKBD0 U8064 ( .CLK(n8139), .C(n8149) );
  CKBD0 U8065 ( .CLK(n8140), .C(n8150) );
  CKBD0 U8066 ( .CLK(n8081), .C(n8151) );
  CKBD0 U8067 ( .CLK(n8084), .C(n8152) );
  CKBD0 U8068 ( .CLK(n8143), .C(n8153) );
  CKBD0 U8069 ( .CLK(n8144), .C(n8154) );
  CKBD0 U8070 ( .CLK(n8145), .C(n8155) );
  CKBD0 U8071 ( .CLK(n8146), .C(n8156) );
  CKBD0 U8072 ( .CLK(n8147), .C(n8157) );
  CKBD0 U8073 ( .CLK(n8148), .C(n8158) );
  CKBD0 U8074 ( .CLK(n8149), .C(n8159) );
  CKBD0 U8075 ( .CLK(n8150), .C(n8160) );
  CKBD0 U8076 ( .CLK(n8153), .C(n8161) );
  CKBD0 U8077 ( .CLK(n8088), .C(n8162) );
  CKBD0 U8078 ( .CLK(n8154), .C(n8163) );
  CKBD0 U8079 ( .CLK(n8090), .C(n8164) );
  CKBD0 U8080 ( .CLK(n8091), .C(n8165) );
  BUFFD0 U8081 ( .I(n8092), .Z(n8166) );
  CKBD0 U8082 ( .CLK(n8101), .C(n8167) );
  CKBD0 U8083 ( .CLK(n8102), .C(n8168) );
  CKBD0 U8084 ( .CLK(n8155), .C(n8169) );
  CKBD0 U8085 ( .CLK(n8156), .C(n8170) );
  CKBD0 U8086 ( .CLK(n8103), .C(n8171) );
  BUFFD0 U8087 ( .I(n8104), .Z(n8172) );
  CKBD0 U8088 ( .CLK(n8106), .C(n8173) );
  BUFFD0 U8089 ( .I(n8105), .Z(n8174) );
  CKBD0 U8090 ( .CLK(n8116), .C(n8175) );
  CKBD0 U8091 ( .CLK(n8157), .C(n8176) );
  BUFFD0 U8092 ( .I(n8108), .Z(n8177) );
  BUFFD0 U8093 ( .I(n8117), .Z(n8178) );
  CKBD0 U8094 ( .CLK(n8119), .C(n8179) );
  BUFFD0 U8095 ( .I(n8118), .Z(n8180) );
  CKBD0 U8096 ( .CLK(n8120), .C(n8181) );
  BUFFD0 U8097 ( .I(n8121), .Z(n8182) );
  CKBD0 U8098 ( .CLK(n8158), .C(n8183) );
  BUFFD0 U8099 ( .I(n8130), .Z(n8184) );
  CKBD0 U8100 ( .CLK(n8131), .C(n8185) );
  BUFFD0 U8101 ( .I(n8132), .Z(n8186) );
  CKBD0 U8102 ( .CLK(n8159), .C(n8187) );
  BUFFD0 U8103 ( .I(n8151), .Z(n8188) );
  CKBD0 U8104 ( .CLK(n8141), .C(n8189) );
  CKBD0 U8105 ( .CLK(n8142), .C(n8190) );
  CKBD0 U8106 ( .CLK(n8152), .C(n8191) );
  CKBD0 U8107 ( .CLK(n8160), .C(n8192) );
  CKBD0 U8108 ( .CLK(n8161), .C(n8193) );
  BUFFD0 U8109 ( .I(n8162), .Z(n8194) );
  CKBD0 U8110 ( .CLK(n8163), .C(n8195) );
  BUFFD0 U8111 ( .I(n8164), .Z(n8196) );
  BUFFD0 U8112 ( .I(n8165), .Z(n8197) );
  CKBD0 U8113 ( .CLK(n8166), .C(n8198) );
  BUFFD0 U8114 ( .I(n8167), .Z(n8199) );
  CKBD0 U8115 ( .CLK(n8169), .C(n8200) );
  CKBD0 U8116 ( .CLK(n8170), .C(n8201) );
  BUFFD0 U8117 ( .I(n8168), .Z(n8202) );
  BUFFD0 U8118 ( .I(n8171), .Z(n8203) );
  CKBD0 U8119 ( .CLK(n8172), .C(n8204) );
  CKBD0 U8120 ( .CLK(n8174), .C(n8205) );
  BUFFD0 U8121 ( .I(n8173), .Z(n8206) );
  CKBD0 U8122 ( .CLK(n8177), .C(n8207) );
  BUFFD0 U8123 ( .I(n8175), .Z(n8208) );
  CKBD0 U8124 ( .CLK(n8176), .C(n8209) );
  CKBD0 U8125 ( .CLK(n8178), .C(n8210) );
  CKBD0 U8126 ( .CLK(n8180), .C(n8211) );
  BUFFD0 U8127 ( .I(n8179), .Z(n8212) );
  BUFFD0 U8128 ( .I(n8181), .Z(n8213) );
  CKBD0 U8129 ( .CLK(n8182), .C(n8214) );
  CKBD0 U8130 ( .CLK(n8184), .C(n8215) );
  CKBD0 U8131 ( .CLK(n8183), .C(n8216) );
  BUFFD0 U8132 ( .I(n8185), .Z(n8217) );
  CKBD0 U8133 ( .CLK(n8186), .C(n8218) );
  BUFFD0 U8134 ( .I(n8189), .Z(n8219) );
  BUFFD0 U8135 ( .I(n8190), .Z(n8220) );
  CKBD0 U8136 ( .CLK(n8187), .C(n8221) );
  CKBD0 U8137 ( .CLK(n8188), .C(n8222) );
  BUFFD0 U8138 ( .I(n8191), .Z(n8223) );
  BUFFD0 U8139 ( .I(n8192), .Z(n8224) );
  CKBD0 U8140 ( .CLK(n8193), .C(n8225) );
  BUFFD0 U8141 ( .I(n8195), .Z(n8226) );
  CKBD0 U8142 ( .CLK(n8194), .C(n8227) );
  CKBD0 U8143 ( .CLK(n8196), .C(n8228) );
  BUFFD0 U8144 ( .I(n8200), .Z(n8229) );
  BUFFD0 U8145 ( .I(n8201), .Z(n8230) );
  CKBD0 U8146 ( .CLK(n8197), .C(n8231) );
  CKBD0 U8147 ( .CLK(n8209), .C(n8232) );
  BUFFD0 U8148 ( .I(n8216), .Z(n8233) );
  CKBD0 U8149 ( .CLK(n8221), .C(n8234) );
  CKBD0 U8150 ( .CLK(n8224), .C(n8235) );
  CKBD0 U8151 ( .CLK(n8225), .C(n8236) );
  CKBD0 U8152 ( .CLK(n8226), .C(n8237) );
  BUFFD0 U8153 ( .I(n8198), .Z(n8238) );
  CKBD0 U8154 ( .CLK(n8199), .C(n8239) );
  CKBD0 U8155 ( .CLK(n8202), .C(n8240) );
  CKBD0 U8156 ( .CLK(n8203), .C(n8241) );
  CKBD0 U8157 ( .CLK(n8229), .C(n8242) );
  CKBD0 U8158 ( .CLK(n8230), .C(n8243) );
  BUFFD0 U8159 ( .I(n8204), .Z(n8244) );
  CKBD0 U8160 ( .CLK(n8232), .C(n8245) );
  CKBD0 U8161 ( .CLK(n8233), .C(n8246) );
  CKBD0 U8162 ( .CLK(n8234), .C(n8247) );
  CKBD0 U8163 ( .CLK(n8235), .C(n8248) );
  BUFFD0 U8164 ( .I(n8236), .Z(n8249) );
  CKBD0 U8165 ( .CLK(n8237), .C(n8250) );
  CKBD0 U8166 ( .CLK(n8206), .C(n8251) );
  BUFFD0 U8167 ( .I(n8205), .Z(n8252) );
  CKBD0 U8168 ( .CLK(n8208), .C(n8253) );
  BUFFD0 U8169 ( .I(n8207), .Z(n8254) );
  BUFFD0 U8170 ( .I(n8210), .Z(n8255) );
  CKBD0 U8171 ( .CLK(n8242), .C(n8256) );
  CKBD0 U8172 ( .CLK(n8212), .C(n8257) );
  CKBD0 U8173 ( .CLK(n8243), .C(n8258) );
  BUFFD0 U8174 ( .I(n8245), .Z(n8259) );
  CKBD0 U8175 ( .CLK(n8246), .C(n8260) );
  BUFFD0 U8176 ( .I(n8247), .Z(n8261) );
  CKBD0 U8177 ( .CLK(n8248), .C(n8262) );
  CKBD0 U8178 ( .CLK(n8249), .C(n8263) );
  CKBD0 U8179 ( .CLK(n8250), .C(n8264) );
  BUFFD0 U8180 ( .I(n8211), .Z(n8265) );
  CKBD0 U8181 ( .CLK(n8213), .C(n8266) );
  BUFFD0 U8182 ( .I(n8214), .Z(n8267) );
  BUFFD0 U8183 ( .I(n8215), .Z(n8268) );
  CKBD0 U8184 ( .CLK(n8256), .C(n8269) );
  CKBD0 U8185 ( .CLK(n8217), .C(n8270) );
  CKBD0 U8186 ( .CLK(n8258), .C(n8271) );
  CKBD0 U8187 ( .CLK(n8259), .C(n8272) );
  CKBD0 U8188 ( .CLK(n8260), .C(n8273) );
  CKBD0 U8189 ( .CLK(n8261), .C(n8274) );
  CKBD0 U8190 ( .CLK(n8262), .C(n8275) );
  CKBD0 U8191 ( .CLK(n8263), .C(n8276) );
  CKBD0 U8192 ( .CLK(n8264), .C(n8277) );
  BUFFD0 U8193 ( .I(n8218), .Z(n8278) );
  CKBD0 U8194 ( .CLK(n8219), .C(n8279) );
  CKBD0 U8195 ( .CLK(n8220), .C(n8280) );
  CKBD0 U8196 ( .CLK(n8269), .C(n8281) );
  CKBD0 U8197 ( .CLK(n8271), .C(n8282) );
  CKBD0 U8198 ( .CLK(n8272), .C(n8283) );
  CKBD0 U8199 ( .CLK(n8273), .C(n8284) );
  CKBD0 U8200 ( .CLK(n8274), .C(n8285) );
  CKBD0 U8201 ( .CLK(n8275), .C(n8286) );
  CKBD0 U8202 ( .CLK(n8276), .C(n8287) );
  CKBD0 U8203 ( .CLK(n8277), .C(n8288) );
  CKBD0 U8204 ( .CLK(n8222), .C(n8289) );
  CKBD0 U8205 ( .CLK(n8223), .C(n8290) );
  CKBD0 U8206 ( .CLK(n8281), .C(n8291) );
  CKBD0 U8207 ( .CLK(n8282), .C(n8292) );
  CKBD0 U8208 ( .CLK(n8283), .C(n8293) );
  CKBD0 U8209 ( .CLK(n8284), .C(n8294) );
  CKBD0 U8210 ( .CLK(n8285), .C(n8295) );
  BUFFD0 U8211 ( .I(n8227), .Z(n8296) );
  CKBD0 U8212 ( .CLK(n8286), .C(n8297) );
  BUFFD0 U8213 ( .I(n8228), .Z(n8298) );
  BUFFD0 U8214 ( .I(n8231), .Z(n8299) );
  CKBD0 U8215 ( .CLK(n8238), .C(n8300) );
  CKBD0 U8216 ( .CLK(n8287), .C(n8301) );
  BUFFD0 U8217 ( .I(n8239), .Z(n8302) );
  CKBD0 U8218 ( .CLK(n8288), .C(n8303) );
  CKBD0 U8219 ( .CLK(n8291), .C(n8304) );
  CKBD0 U8220 ( .CLK(n8292), .C(n8305) );
  CKBD0 U8221 ( .CLK(n8293), .C(n8306) );
  CKBD0 U8222 ( .CLK(n8294), .C(n8307) );
  CKBD0 U8223 ( .CLK(n8295), .C(n8308) );
  CKBD0 U8224 ( .CLK(n8297), .C(n8309) );
  BUFFD0 U8225 ( .I(n8240), .Z(n8310) );
  BUFFD0 U8226 ( .I(n8241), .Z(n8311) );
  CKBD0 U8227 ( .CLK(n8244), .C(n8312) );
  CKBD0 U8228 ( .CLK(n8252), .C(n8313) );
  BUFFD0 U8229 ( .I(n8251), .Z(n8314) );
  CKBD0 U8230 ( .CLK(n8254), .C(n8315) );
  CKBD0 U8231 ( .CLK(n8301), .C(n8316) );
  BUFFD0 U8232 ( .I(n8253), .Z(n8317) );
  CKBD0 U8233 ( .CLK(n8303), .C(n8318) );
  CKBD0 U8234 ( .CLK(n8304), .C(n8319) );
  CKBD0 U8235 ( .CLK(n8305), .C(n8320) );
  CKBD0 U8236 ( .CLK(n8306), .C(n8321) );
  CKBD0 U8237 ( .CLK(n8307), .C(n8322) );
  CKBD0 U8238 ( .CLK(n8308), .C(n8323) );
  CKBD0 U8239 ( .CLK(n8309), .C(n8324) );
  CKBD0 U8240 ( .CLK(n8255), .C(n8325) );
  CKBD0 U8241 ( .CLK(n8265), .C(n8326) );
  BUFFD0 U8242 ( .I(n8257), .Z(n8327) );
  BUFFD0 U8243 ( .I(n8266), .Z(n8328) );
  CKBD0 U8244 ( .CLK(n8267), .C(n8329) );
  CKBD0 U8245 ( .CLK(n8316), .C(n8330) );
  CKBD0 U8246 ( .CLK(n8318), .C(n8331) );
  CKBD0 U8247 ( .CLK(n8319), .C(n8332) );
  CKBD0 U8248 ( .CLK(n8320), .C(n8333) );
  CKBD0 U8249 ( .CLK(n8321), .C(n8334) );
  CKBD0 U8250 ( .CLK(n8322), .C(n8335) );
  CKBD0 U8251 ( .CLK(n8323), .C(n8336) );
  CKBD0 U8252 ( .CLK(n8324), .C(n8337) );
  CKBD0 U8253 ( .CLK(n8268), .C(n8338) );
  BUFFD0 U8254 ( .I(n8279), .Z(n8339) );
  BUFFD0 U8255 ( .I(n8280), .Z(n8340) );
  BUFFD0 U8256 ( .I(n8270), .Z(n8341) );
  CKBD0 U8257 ( .CLK(n8278), .C(n8342) );
  CKBD0 U8258 ( .CLK(n8330), .C(n8343) );
  CKBD0 U8259 ( .CLK(n8331), .C(n8344) );
  CKBD0 U8260 ( .CLK(n8333), .C(n8345) );
  CKBD0 U8261 ( .CLK(n8332), .C(n8346) );
  CKBD0 U8262 ( .CLK(n8334), .C(n8347) );
  CKBD0 U8263 ( .CLK(n8335), .C(n8348) );
  CKBD0 U8264 ( .CLK(n8336), .C(n8349) );
  CKBD0 U8265 ( .CLK(n8337), .C(n8350) );
  BUFFD0 U8266 ( .I(n8289), .Z(n8351) );
  BUFFD0 U8267 ( .I(n8290), .Z(n8352) );
  CKBD0 U8268 ( .CLK(n8343), .C(n8353) );
  CKBD0 U8269 ( .CLK(n8344), .C(n8354) );
  BUFFD0 U8270 ( .I(n8345), .Z(n8355) );
  CKBD0 U8271 ( .CLK(n8346), .C(n8356) );
  CKBD0 U8272 ( .CLK(n8296), .C(n8357) );
  CKBD0 U8273 ( .CLK(n8347), .C(n8358) );
  CKBD0 U8274 ( .CLK(n8298), .C(n8359) );
  CKBD0 U8275 ( .CLK(n8299), .C(n8360) );
  BUFFD0 U8276 ( .I(n8300), .Z(n8361) );
  CKBD0 U8277 ( .CLK(n8302), .C(n8362) );
  CKBD0 U8278 ( .CLK(n8310), .C(n8363) );
  CKBD0 U8279 ( .CLK(n8348), .C(n8364) );
  CKBD0 U8280 ( .CLK(n8311), .C(n8365) );
  BUFFD0 U8281 ( .I(n8312), .Z(n8366) );
  CKBD0 U8282 ( .CLK(n8314), .C(n8367) );
  BUFFD0 U8283 ( .I(n8313), .Z(n8368) );
  CKBD0 U8284 ( .CLK(n8317), .C(n8369) );
  BUFFD0 U8285 ( .I(n8315), .Z(n8370) );
  CKBD0 U8286 ( .CLK(n8349), .C(n8371) );
  BUFFD0 U8287 ( .I(n8325), .Z(n8372) );
  CKBD0 U8288 ( .CLK(n8327), .C(n8373) );
  BUFFD0 U8289 ( .I(n8326), .Z(n8374) );
  CKBD0 U8290 ( .CLK(n8328), .C(n8375) );
  BUFFD0 U8291 ( .I(n8329), .Z(n8376) );
  CKBD0 U8292 ( .CLK(n8339), .C(n8377) );
  BUFFD0 U8293 ( .I(n8350), .Z(n8378) );
  CKBD0 U8294 ( .CLK(n8353), .C(n8379) );
  BUFFD0 U8295 ( .I(n8354), .Z(n8380) );
  BUFFD0 U8296 ( .I(n8356), .Z(n8381) );
  CKBD0 U8297 ( .CLK(n8355), .C(n8382) );
  CKBD0 U8298 ( .CLK(n8358), .C(n8383) );
  BUFFD0 U8299 ( .I(n8364), .Z(n8384) );
  CKBD0 U8300 ( .CLK(n8371), .C(n8385) );
  BUFFD0 U8301 ( .I(n8338), .Z(n8386) );
  CKBD0 U8302 ( .CLK(n8340), .C(n8387) );
  CKBD0 U8303 ( .CLK(n8341), .C(n8388) );
  BUFFD0 U8304 ( .I(n8342), .Z(n8389) );
  CKBD0 U8305 ( .CLK(n8351), .C(n8390) );
  CKBD0 U8306 ( .CLK(n8352), .C(n8391) );
  CKBD0 U8307 ( .CLK(n8378), .C(n8392) );
  CKBD0 U8308 ( .CLK(n8379), .C(n8393) );
  CKBD0 U8309 ( .CLK(n8380), .C(n8394) );
  CKBD0 U8310 ( .CLK(n8381), .C(n8395) );
  CKBD0 U8311 ( .CLK(n8382), .C(n8396) );
  CKBD0 U8312 ( .CLK(n8383), .C(n8397) );
  CKBD0 U8313 ( .CLK(n8384), .C(n8398) );
  CKBD0 U8314 ( .CLK(n8385), .C(n8399) );
  CKBD0 U8315 ( .CLK(n8392), .C(n8400) );
  BUFFD0 U8316 ( .I(n8393), .Z(n8401) );
  CKBD0 U8317 ( .CLK(n8394), .C(n8402) );
  BUFFD0 U8318 ( .I(n8357), .Z(n8403) );
  CKBD0 U8319 ( .CLK(n8395), .C(n8404) );
  CKBD0 U8320 ( .CLK(n8396), .C(n8405) );
  BUFFD0 U8321 ( .I(n8359), .Z(n8406) );
  BUFFD0 U8322 ( .I(n8397), .Z(n8407) );
  CKBD0 U8323 ( .CLK(n8398), .C(n8408) );
  BUFFD0 U8324 ( .I(n8399), .Z(n8409) );
  CKBD0 U8325 ( .CLK(n8400), .C(n8410) );
  CKBD0 U8326 ( .CLK(n8401), .C(n8411) );
  CKBD0 U8327 ( .CLK(n8402), .C(n8412) );
  BUFFD0 U8328 ( .I(n8360), .Z(n8413) );
  CKBD0 U8329 ( .CLK(n8361), .C(n8414) );
  BUFFD0 U8330 ( .I(n8362), .Z(n8415) );
  BUFFD0 U8331 ( .I(n8363), .Z(n8416) );
  BUFFD0 U8332 ( .I(n8365), .Z(n8417) );
  CKBD0 U8333 ( .CLK(n8404), .C(n8418) );
  CKBD0 U8334 ( .CLK(n8366), .C(n8419) );
  CKBD0 U8335 ( .CLK(n8405), .C(n8420) );
  CKBD0 U8336 ( .CLK(n8407), .C(n8421) );
  CKBD0 U8337 ( .CLK(n8408), .C(n8422) );
  CKBD0 U8338 ( .CLK(n8409), .C(n8423) );
  CKBD0 U8339 ( .CLK(n8410), .C(n8424) );
  CKBD0 U8340 ( .CLK(n8411), .C(n8425) );
  CKBD0 U8341 ( .CLK(n8412), .C(n8426) );
  CKBD0 U8342 ( .CLK(n8368), .C(n8427) );
  BUFFD0 U8343 ( .I(n8367), .Z(n8428) );
  CKBD0 U8344 ( .CLK(n8370), .C(n8429) );
  BUFFD0 U8345 ( .I(n8369), .Z(n8430) );
  CKBD0 U8346 ( .CLK(n8372), .C(n8431) );
  CKBD0 U8347 ( .CLK(n8418), .C(n8432) );
  CKBD0 U8348 ( .CLK(n8420), .C(n8433) );
  BUFFD0 U8349 ( .I(n8377), .Z(n8434) );
  CKBD0 U8350 ( .CLK(n8374), .C(n8435) );
  CKBD0 U8351 ( .CLK(n8421), .C(n8436) );
  CKBD0 U8352 ( .CLK(n8422), .C(n8437) );
  CKBD0 U8353 ( .CLK(n8423), .C(n8438) );
  CKBD0 U8354 ( .CLK(n8424), .C(n8439) );
  CKBD0 U8355 ( .CLK(n8425), .C(n8440) );
  CKBD0 U8356 ( .CLK(n8426), .C(n8441) );
  BUFFD0 U8357 ( .I(n8373), .Z(n8442) );
  BUFFD0 U8358 ( .I(n8387), .Z(n8443) );
  BUFFD0 U8359 ( .I(n8375), .Z(n8444) );
  CKBD0 U8360 ( .CLK(n8376), .C(n8445) );
  CKBD0 U8361 ( .CLK(n8386), .C(n8446) );
  BUFFD0 U8362 ( .I(n8390), .Z(n8447) );
  BUFFD0 U8363 ( .I(n8391), .Z(n8448) );
  CKBD0 U8364 ( .CLK(n8432), .C(n8449) );
  CKBD0 U8365 ( .CLK(n8433), .C(n8450) );
  CKBD0 U8366 ( .CLK(n8436), .C(n8451) );
  CKBD0 U8367 ( .CLK(n8437), .C(n8452) );
  CKBD0 U8368 ( .CLK(n8438), .C(n8453) );
  CKBD0 U8369 ( .CLK(n8439), .C(n8454) );
  CKBD0 U8370 ( .CLK(n8440), .C(n8455) );
  CKBD0 U8371 ( .CLK(n8441), .C(n8456) );
  BUFFD0 U8372 ( .I(n8388), .Z(n8457) );
  CKBD0 U8373 ( .CLK(n8389), .C(n8458) );
  CKBD0 U8374 ( .CLK(n8449), .C(n8459) );
  CKBD0 U8375 ( .CLK(n8450), .C(n8460) );
  CKBD0 U8376 ( .CLK(n8451), .C(n8461) );
  CKBD0 U8377 ( .CLK(n8452), .C(n8462) );
  CKBD0 U8378 ( .CLK(n8453), .C(n8463) );
  CKBD0 U8379 ( .CLK(n8454), .C(n8464) );
  CKBD0 U8380 ( .CLK(n8455), .C(n8465) );
  CKBD0 U8381 ( .CLK(n8456), .C(n8466) );
  CKBD0 U8382 ( .CLK(n8459), .C(n8467) );
  CKBD0 U8383 ( .CLK(n8460), .C(n8468) );
  CKBD0 U8384 ( .CLK(n8461), .C(n8469) );
  CKBD0 U8385 ( .CLK(n8462), .C(n8470) );
  CKBD0 U8386 ( .CLK(n8463), .C(n8471) );
  CKBD0 U8387 ( .CLK(n8403), .C(n8472) );
  CKBD0 U8388 ( .CLK(n8464), .C(n8473) );
  CKBD0 U8389 ( .CLK(n8406), .C(n8474) );
  CKBD0 U8390 ( .CLK(n8413), .C(n8475) );
  BUFFD0 U8391 ( .I(n8414), .Z(n8476) );
  CKBD0 U8392 ( .CLK(n8465), .C(n8477) );
  CKBD0 U8393 ( .CLK(n8415), .C(n8478) );
  CKBD0 U8394 ( .CLK(n8466), .C(n8479) );
  CKBD0 U8395 ( .CLK(n8467), .C(n8480) );
  CKBD0 U8396 ( .CLK(n8468), .C(n8481) );
  CKBD0 U8397 ( .CLK(n8469), .C(n8482) );
  CKBD0 U8398 ( .CLK(n8470), .C(n8483) );
  CKBD0 U8399 ( .CLK(n8471), .C(n8484) );
  CKBD0 U8400 ( .CLK(n8473), .C(n8485) );
  CKBD0 U8401 ( .CLK(n8477), .C(n8486) );
  BUFFD0 U8402 ( .I(n8480), .Z(n8487) );
  CKBD0 U8403 ( .CLK(n8479), .C(n8488) );
  CKBD0 U8404 ( .CLK(n8481), .C(n8489) );
  CKBD0 U8405 ( .CLK(n8482), .C(n8490) );
  CKBD0 U8406 ( .CLK(n8483), .C(n8491) );
  CKBD0 U8407 ( .CLK(n8484), .C(n8492) );
  CKBD0 U8408 ( .CLK(n8485), .C(n8493) );
  CKBD0 U8409 ( .CLK(n8486), .C(n8494) );
  CKBD0 U8410 ( .CLK(n8488), .C(n8495) );
  CKBD0 U8411 ( .CLK(n8487), .C(n8496) );
  BUFFD0 U8412 ( .I(n8489), .Z(n8497) );
  CKBD0 U8413 ( .CLK(n8490), .C(n8498) );
  BUFFD0 U8414 ( .I(n8491), .Z(n8499) );
  CKBD0 U8415 ( .CLK(n8492), .C(n8500) );
  CKBD0 U8416 ( .CLK(n8416), .C(n8501) );
  CKBD0 U8417 ( .CLK(n8417), .C(n8502) );
  BUFFD0 U8418 ( .I(n8419), .Z(n8503) );
  CKBD0 U8419 ( .CLK(n8428), .C(n8504) );
  BUFFD0 U8420 ( .I(n8427), .Z(n8505) );
  CKBD0 U8421 ( .CLK(n8430), .C(n8506) );
  BUFFD0 U8422 ( .I(n8493), .Z(n8507) );
  CKBD0 U8423 ( .CLK(n8494), .C(n8508) );
  BUFFD0 U8424 ( .I(n8495), .Z(n8509) );
  CKBD0 U8425 ( .CLK(n8496), .C(n8510) );
  CKBD0 U8426 ( .CLK(n8497), .C(n8511) );
  CKBD0 U8427 ( .CLK(n8498), .C(n8512) );
  CKBD0 U8428 ( .CLK(n8499), .C(n8513) );
  CKBD0 U8429 ( .CLK(n8500), .C(n8514) );
  BUFFD0 U8430 ( .I(n8429), .Z(n8515) );
  BUFFD0 U8431 ( .I(n8431), .Z(n8516) );
  CKBD0 U8432 ( .CLK(n8434), .C(n8517) );
  CKBD0 U8433 ( .CLK(n8442), .C(n8518) );
  BUFFD0 U8434 ( .I(n8435), .Z(n8519) );
  CKBD0 U8435 ( .CLK(n8443), .C(n8520) );
  CKBD0 U8436 ( .CLK(n8444), .C(n8521) );
  CKBD0 U8437 ( .CLK(n8507), .C(n8522) );
  CKBD0 U8438 ( .CLK(n8508), .C(n8523) );
  CKBD0 U8439 ( .CLK(n8509), .C(n8524) );
  CKBD0 U8440 ( .CLK(n8510), .C(n8525) );
  CKBD0 U8441 ( .CLK(n8511), .C(n8526) );
  CKBD0 U8442 ( .CLK(n8512), .C(n8527) );
  CKBD0 U8443 ( .CLK(n8513), .C(n8528) );
  CKBD0 U8444 ( .CLK(n8514), .C(n8529) );
  BUFFD0 U8445 ( .I(n8445), .Z(n8530) );
  CKBD0 U8446 ( .CLK(n8447), .C(n8531) );
  BUFFD0 U8447 ( .I(n8446), .Z(n8532) );
  CKBD0 U8448 ( .CLK(n8448), .C(n8533) );
  CKBD0 U8449 ( .CLK(n8457), .C(n8534) );
  BUFFD0 U8450 ( .I(n8458), .Z(n8535) );
  CKBD0 U8451 ( .CLK(n8522), .C(n8536) );
  BUFFD0 U8452 ( .I(n8523), .Z(n8537) );
  CKBD0 U8453 ( .CLK(n8524), .C(n8538) );
  CKBD0 U8454 ( .CLK(n8525), .C(n8539) );
  CKBD0 U8455 ( .CLK(n8526), .C(n8540) );
  BUFFD0 U8456 ( .I(n8472), .Z(n8541) );
  BUFFD0 U8457 ( .I(n8527), .Z(n8542) );
  BUFFD0 U8458 ( .I(n8474), .Z(n8543) );
  BUFFD0 U8459 ( .I(n8475), .Z(n8544) );
  CKBD0 U8460 ( .CLK(n8476), .C(n8545) );
  BUFFD0 U8461 ( .I(n8478), .Z(n8546) );
  BUFFD0 U8462 ( .I(n8501), .Z(n8547) );
  CKBD0 U8463 ( .CLK(n8528), .C(n8548) );
  BUFFD0 U8464 ( .I(n8502), .Z(n8549) );
  CKBD0 U8465 ( .CLK(n8503), .C(n8550) );
  CKBD0 U8466 ( .CLK(n8505), .C(n8551) );
  BUFFD0 U8467 ( .I(n8517), .Z(n8552) );
  BUFFD0 U8468 ( .I(n8504), .Z(n8553) );
  BUFFD0 U8469 ( .I(n8520), .Z(n8554) );
  CKBD0 U8470 ( .CLK(n8515), .C(n8555) );
  BUFFD0 U8471 ( .I(n8529), .Z(n8556) );
  CKBD0 U8472 ( .CLK(n8536), .C(n8557) );
  CKBD0 U8473 ( .CLK(n8537), .C(n8558) );
  CKBD0 U8474 ( .CLK(n8538), .C(n8559) );
  CKBD0 U8475 ( .CLK(n8539), .C(n8560) );
  CKBD0 U8476 ( .CLK(n8540), .C(n8561) );
  CKBD0 U8477 ( .CLK(n8542), .C(n8562) );
  BUFFD0 U8478 ( .I(n8506), .Z(n8563) );
  CKBD0 U8479 ( .CLK(n8516), .C(n8564) );
  CKBD0 U8480 ( .CLK(n8548), .C(n8565) );
  CKBD0 U8481 ( .CLK(n8519), .C(n8566) );
  BUFFD0 U8482 ( .I(n8531), .Z(n8567) );
  BUFFD0 U8483 ( .I(n8518), .Z(n8568) );
  BUFFD0 U8484 ( .I(n8533), .Z(n8569) );
  BUFFD0 U8485 ( .I(n8521), .Z(n8570) );
  CKBD0 U8486 ( .CLK(n8530), .C(n8571) );
  CKBD0 U8487 ( .CLK(n8532), .C(n8572) );
  CKBD0 U8488 ( .CLK(n8556), .C(n8573) );
  BUFFD0 U8489 ( .I(n8534), .Z(n8574) );
  CKBD0 U8490 ( .CLK(n8535), .C(n8575) );
  CKBD0 U8491 ( .CLK(n8557), .C(n8576) );
  CKBD0 U8492 ( .CLK(n8558), .C(n8577) );
  CKBD0 U8493 ( .CLK(n8559), .C(n8578) );
  CKBD0 U8494 ( .CLK(n8541), .C(n8579) );
  CKBD0 U8495 ( .CLK(n8560), .C(n8580) );
  CKBD0 U8496 ( .CLK(n8561), .C(n8581) );
  CKBD0 U8497 ( .CLK(n8543), .C(n8582) );
  CKBD0 U8498 ( .CLK(n8544), .C(n8583) );
  CKBD0 U8499 ( .CLK(n8562), .C(n8584) );
  CKBD0 U8500 ( .CLK(n8565), .C(n8585) );
  CKBD0 U8501 ( .CLK(n8573), .C(n8586) );
  CKBD0 U8502 ( .CLK(n8576), .C(n8587) );
  CKBD0 U8503 ( .CLK(n8577), .C(n8588) );
  CKBD0 U8504 ( .CLK(n8578), .C(n8589) );
  BUFFD0 U8505 ( .I(n8545), .Z(n8590) );
  CKBD0 U8506 ( .CLK(n8546), .C(n8591) );
  CKBD0 U8507 ( .CLK(n8547), .C(n8592) );
  CKBD0 U8508 ( .CLK(n8549), .C(n8593) );
  CKBD0 U8509 ( .CLK(n8580), .C(n8594) );
  CKBD0 U8510 ( .CLK(n8581), .C(n8595) );
  CKBD0 U8511 ( .CLK(n8584), .C(n8596) );
  CKBD0 U8512 ( .CLK(n8585), .C(n8597) );
  CKBD0 U8513 ( .CLK(n8586), .C(n8598) );
  CKBD0 U8514 ( .CLK(n8587), .C(n8599) );
  CKBD0 U8515 ( .CLK(n8588), .C(n8600) );
  CKBD0 U8516 ( .CLK(n8589), .C(n8601) );
  BUFFD0 U8517 ( .I(n8550), .Z(n8602) );
  CKBD0 U8518 ( .CLK(n8552), .C(n8603) );
  CKBD0 U8519 ( .CLK(n8553), .C(n8604) );
  BUFFD0 U8520 ( .I(n8551), .Z(n8605) );
  CKBD0 U8521 ( .CLK(n8563), .C(n8606) );
  CKBD0 U8522 ( .CLK(n8554), .C(n8607) );
  BUFFD0 U8523 ( .I(n8555), .Z(n8608) );
  BUFFD0 U8524 ( .I(n8564), .Z(n8609) );
  CKBD0 U8525 ( .CLK(n8594), .C(n8610) );
  CKBD0 U8526 ( .CLK(n8595), .C(n8611) );
  CKBD0 U8527 ( .CLK(n8568), .C(n8612) );
  CKBD0 U8528 ( .CLK(n8596), .C(n8613) );
  CKBD0 U8529 ( .CLK(n8597), .C(n8614) );
  CKBD0 U8530 ( .CLK(n8598), .C(n8615) );
  CKBD0 U8531 ( .CLK(n8599), .C(n8616) );
  CKBD0 U8532 ( .CLK(n8600), .C(n8617) );
  CKBD0 U8533 ( .CLK(n8601), .C(n8618) );
  CKBD0 U8534 ( .CLK(n8567), .C(n8619) );
  CKBD0 U8535 ( .CLK(n8569), .C(n8620) );
  BUFFD0 U8536 ( .I(n8566), .Z(n8621) );
  CKBD0 U8537 ( .CLK(n8570), .C(n8622) );
  BUFFD0 U8538 ( .I(n8571), .Z(n8623) );
  BUFFD0 U8539 ( .I(n8572), .Z(n8624) );
  CKBD0 U8540 ( .CLK(n8610), .C(n8625) );
  CKBD0 U8541 ( .CLK(n8611), .C(n8626) );
  CKBD0 U8542 ( .CLK(n8574), .C(n8627) );
  CKBD0 U8543 ( .CLK(n8613), .C(n8628) );
  CKBD0 U8544 ( .CLK(n8614), .C(n8629) );
  CKBD0 U8545 ( .CLK(n8615), .C(n8630) );
  CKBD0 U8546 ( .CLK(n8616), .C(n8631) );
  CKBD0 U8547 ( .CLK(n8617), .C(n8632) );
  CKBD0 U8548 ( .CLK(n8618), .C(n8633) );
  BUFFD0 U8549 ( .I(n8575), .Z(n8634) );
  CKBD0 U8550 ( .CLK(n8625), .C(n8635) );
  CKBD0 U8551 ( .CLK(n8626), .C(n8636) );
  CKBD0 U8552 ( .CLK(n8628), .C(n8637) );
  CKBD0 U8553 ( .CLK(n8629), .C(n8638) );
  CKBD0 U8554 ( .CLK(n8630), .C(n8639) );
  CKBD0 U8555 ( .CLK(n8631), .C(n8640) );
  BUFFD0 U8556 ( .I(n8579), .Z(n8641) );
  CKBD0 U8557 ( .CLK(n8632), .C(n8642) );
  BUFFD0 U8558 ( .I(n8582), .Z(n8643) );
  BUFFD0 U8559 ( .I(n8583), .Z(n8644) );
  CKBD0 U8560 ( .CLK(n8590), .C(n8645) );
  CKBD0 U8561 ( .CLK(n8633), .C(n8646) );
  CKBD0 U8562 ( .CLK(n8635), .C(n8647) );
  CKBD0 U8563 ( .CLK(n8636), .C(n8648) );
  CKBD0 U8564 ( .CLK(n8637), .C(n8649) );
  CKBD0 U8565 ( .CLK(n8638), .C(n8650) );
  CKBD0 U8566 ( .CLK(n8639), .C(n8651) );
  BUFFD0 U8567 ( .I(n8640), .Z(n8652) );
  CKBD0 U8568 ( .CLK(n8642), .C(n8653) );
  BUFFD0 U8569 ( .I(n8603), .Z(n8654) );
  BUFFD0 U8570 ( .I(n8591), .Z(n8655) );
  BUFFD0 U8571 ( .I(n8607), .Z(n8656) );
  BUFFD0 U8572 ( .I(n8592), .Z(n8657) );
  BUFFD0 U8573 ( .I(n8593), .Z(n8658) );
  CKBD0 U8574 ( .CLK(n8602), .C(n8659) );
  CKBD0 U8575 ( .CLK(n8605), .C(n8660) );
  BUFFD0 U8576 ( .I(n8604), .Z(n8661) );
  BUFFD0 U8577 ( .I(n8619), .Z(n8662) );
  BUFFD0 U8578 ( .I(n8620), .Z(n8663) );
  BUFFD0 U8579 ( .I(n8646), .Z(n8664) );
  BUFFD0 U8580 ( .I(n8647), .Z(n8665) );
  BUFFD0 U8581 ( .I(n8648), .Z(n8666) );
  CKBD0 U8582 ( .CLK(n8649), .C(n8667) );
  BUFFD0 U8583 ( .I(n8650), .Z(n8668) );
  CKBD0 U8584 ( .CLK(n8651), .C(n8669) );
  CKBD0 U8585 ( .CLK(n8652), .C(n8670) );
  CKBD0 U8586 ( .CLK(n8653), .C(n8671) );
  CKBD0 U8587 ( .CLK(n8608), .C(n8672) );
  CKBD0 U8588 ( .CLK(n8664), .C(n8673) );
  CKBD0 U8589 ( .CLK(n8665), .C(n8674) );
  CKBD0 U8590 ( .CLK(n8666), .C(n8675) );
  CKBD0 U8591 ( .CLK(n8667), .C(n8676) );
  CKBD0 U8592 ( .CLK(n8668), .C(n8677) );
  CKBD0 U8593 ( .CLK(n8669), .C(n8678) );
  CKBD0 U8594 ( .CLK(n8670), .C(n8679) );
  CKBD0 U8595 ( .CLK(n8671), .C(n8680) );
  CKBD0 U8596 ( .CLK(n8673), .C(n8681) );
  CKBD0 U8597 ( .CLK(n8674), .C(n8682) );
  CKBD0 U8598 ( .CLK(n8675), .C(n8683) );
  BUFFD0 U8599 ( .I(n8676), .Z(n8684) );
  CKBD0 U8600 ( .CLK(n8677), .C(n8685) );
  BUFFD0 U8601 ( .I(n8678), .Z(n8686) );
  CKBD0 U8602 ( .CLK(n8679), .C(n8687) );
  BUFFD0 U8603 ( .I(n8606), .Z(n8688) );
  CKBD0 U8604 ( .CLK(n8609), .C(n8689) );
  CKBD0 U8605 ( .CLK(n8621), .C(n8690) );
  BUFFD0 U8606 ( .I(n8612), .Z(n8691) );
  BUFFD0 U8607 ( .I(n8622), .Z(n8692) );
  CKBD0 U8608 ( .CLK(n8623), .C(n8693) );
  BUFFD0 U8609 ( .I(n8680), .Z(n8694) );
  CKBD0 U8610 ( .CLK(n8681), .C(n8695) );
  CKBD0 U8611 ( .CLK(n8682), .C(n8696) );
  CKBD0 U8612 ( .CLK(n8683), .C(n8697) );
  CKBD0 U8613 ( .CLK(n8684), .C(n8698) );
  CKBD0 U8614 ( .CLK(n8685), .C(n8699) );
  CKBD0 U8615 ( .CLK(n8686), .C(n8700) );
  CKBD0 U8616 ( .CLK(n8687), .C(n8701) );
  CKBD0 U8617 ( .CLK(n8624), .C(n8702) );
  CKBD0 U8618 ( .CLK(n8634), .C(n8703) );
  CKBD0 U8619 ( .CLK(n8694), .C(n8704) );
  BUFFD0 U8620 ( .I(n8627), .Z(n8705) );
  CKBD0 U8621 ( .CLK(n8695), .C(n8706) );
  CKBD0 U8622 ( .CLK(n8696), .C(n8707) );
  CKBD0 U8623 ( .CLK(n8697), .C(n8708) );
  CKBD0 U8624 ( .CLK(n8698), .C(n8709) );
  CKBD0 U8625 ( .CLK(n8641), .C(n8710) );
  CKBD0 U8626 ( .CLK(n8699), .C(n8711) );
  CKBD0 U8627 ( .CLK(n8643), .C(n8712) );
  CKBD0 U8628 ( .CLK(n8644), .C(n8713) );
  BUFFD0 U8629 ( .I(n8645), .Z(n8714) );
  CKBD0 U8630 ( .CLK(n8654), .C(n8715) );
  CKBD0 U8631 ( .CLK(n8655), .C(n8716) );
  CKBD0 U8632 ( .CLK(n8700), .C(n8717) );
  CKBD0 U8633 ( .CLK(n8657), .C(n8718) );
  CKBD0 U8634 ( .CLK(n8656), .C(n8719) );
  CKBD0 U8635 ( .CLK(n8701), .C(n8720) );
  CKBD0 U8636 ( .CLK(n8704), .C(n8721) );
  CKBD0 U8637 ( .CLK(n8706), .C(n8722) );
  CKBD0 U8638 ( .CLK(n8707), .C(n8723) );
  CKBD0 U8639 ( .CLK(n8708), .C(n8724) );
  CKBD0 U8640 ( .CLK(n8709), .C(n8725) );
  CKBD0 U8641 ( .CLK(n8711), .C(n8726) );
  BUFFD0 U8642 ( .I(n8659), .Z(n8727) );
  CKBD0 U8643 ( .CLK(n8661), .C(n8728) );
  BUFFD0 U8644 ( .I(n8660), .Z(n8729) );
  CKBD0 U8645 ( .CLK(n8662), .C(n8730) );
  CKBD0 U8646 ( .CLK(n8663), .C(n8731) );
  BUFFD0 U8647 ( .I(n8672), .Z(n8732) );
  CKBD0 U8648 ( .CLK(n8717), .C(n8733) );
  CKBD0 U8649 ( .CLK(n8658), .C(n8734) );
  BUFFD0 U8650 ( .I(n8689), .Z(n8735) );
  CKBD0 U8651 ( .CLK(n8691), .C(n8736) );
  BUFFD0 U8652 ( .I(n8690), .Z(n8737) );
  CKBD0 U8653 ( .CLK(n8692), .C(n8738) );
  CKBD0 U8654 ( .CLK(n8688), .C(n8739) );
  BUFFD0 U8655 ( .I(n8693), .Z(n8740) );
  BUFFD0 U8656 ( .I(n8702), .Z(n8741) );
  BUFFD0 U8657 ( .I(n8703), .Z(n8742) );
  CKBD0 U8658 ( .CLK(n8720), .C(n8743) );
  CKBD0 U8659 ( .CLK(n8721), .C(n8744) );
  CKBD0 U8660 ( .CLK(n8705), .C(n8745) );
  CKBD0 U8661 ( .CLK(n8722), .C(n8746) );
  CKBD0 U8662 ( .CLK(n8723), .C(n8747) );
  CKBD0 U8663 ( .CLK(n8724), .C(n8748) );
  BUFFD0 U8664 ( .I(n8710), .Z(n8749) );
  CKBD0 U8665 ( .CLK(n8725), .C(n8750) );
  BUFFD0 U8666 ( .I(n8715), .Z(n8751) );
  BUFFD0 U8667 ( .I(n8719), .Z(n8752) );
  BUFFD0 U8668 ( .I(n8712), .Z(n8753) );
  BUFFD0 U8669 ( .I(n8713), .Z(n8754) );
  CKBD0 U8670 ( .CLK(n8714), .C(n8755) );
  BUFFD0 U8671 ( .I(n8730), .Z(n8756) );
  BUFFD0 U8672 ( .I(n8716), .Z(n8757) );
  BUFFD0 U8673 ( .I(n8731), .Z(n8758) );
  BUFFD0 U8674 ( .I(n8718), .Z(n8759) );
  CKBD0 U8675 ( .CLK(n8726), .C(n8760) );
  CKBD0 U8676 ( .CLK(n8727), .C(n8761) );
  BUFFD0 U8677 ( .I(n8734), .Z(n8762) );
  CKBD0 U8678 ( .CLK(n8729), .C(n8763) );
  BUFFD0 U8679 ( .I(n8728), .Z(n8764) );
  CKBD0 U8680 ( .CLK(n8732), .C(n8765) );
  BUFFD0 U8681 ( .I(n8739), .Z(n8766) );
  CKBD0 U8682 ( .CLK(n8735), .C(n8767) );
  CKBD0 U8683 ( .CLK(n8733), .C(n8768) );
  CKBD0 U8684 ( .CLK(n8737), .C(n8769) );
  BUFFD0 U8685 ( .I(n8736), .Z(n8770) );
  BUFFD0 U8686 ( .I(n8738), .Z(n8771) );
  CKBD0 U8687 ( .CLK(n8740), .C(n8772) );
  CKBD0 U8688 ( .CLK(n8741), .C(n8773) );
  CKBD0 U8689 ( .CLK(n8742), .C(n8774) );
  CKBD0 U8690 ( .CLK(n8743), .C(n8775) );
  BUFFD0 U8691 ( .I(n8745), .Z(n8776) );
  CKBD0 U8692 ( .CLK(n8744), .C(n8777) );
  CKBD0 U8693 ( .CLK(n8746), .C(n8778) );
  CKBD0 U8694 ( .CLK(n8747), .C(n8779) );
  CKBD0 U8695 ( .CLK(n8748), .C(n8780) );
  CKBD0 U8696 ( .CLK(n8749), .C(n8781) );
  CKBD0 U8697 ( .CLK(n8751), .C(n8782) );
  CKBD0 U8698 ( .CLK(n8750), .C(n8783) );
  CKBD0 U8699 ( .CLK(n8753), .C(n8784) );
  CKBD0 U8700 ( .CLK(n8752), .C(n8785) );
  CKBD0 U8701 ( .CLK(n8754), .C(n8786) );
  BUFFD0 U8702 ( .I(n8755), .Z(n8787) );
  CKBD0 U8703 ( .CLK(n8757), .C(n8788) );
  CKBD0 U8704 ( .CLK(n8756), .C(n8789) );
  CKBD0 U8705 ( .CLK(n8758), .C(n8790) );
  CKBD0 U8706 ( .CLK(n8759), .C(n8791) );
  CKBD0 U8707 ( .CLK(n8762), .C(n8792) );
  BUFFD0 U8708 ( .I(n8761), .Z(n8793) );
  CKBD0 U8709 ( .CLK(n8760), .C(n8794) );
  CKBD0 U8710 ( .CLK(n8764), .C(n8795) );
  BUFFD0 U8711 ( .I(n8763), .Z(n8796) );
  CKBD0 U8712 ( .CLK(n8766), .C(n8797) );
  BUFFD0 U8713 ( .I(n8765), .Z(n8798) );
  BUFFD0 U8714 ( .I(n8767), .Z(n8799) );
  CKBD0 U8715 ( .CLK(n8768), .C(n8800) );
  CKBD0 U8716 ( .CLK(n8770), .C(n8801) );
  BUFFD0 U8717 ( .I(n8769), .Z(n8802) );
  CKBD0 U8718 ( .CLK(n8771), .C(n8803) );
  BUFFD0 U8719 ( .I(n8772), .Z(n8804) );
  BUFFD0 U8720 ( .I(n8773), .Z(n8805) );
  BUFFD0 U8721 ( .I(n8774), .Z(n8806) );
  CKBD0 U8722 ( .CLK(n8775), .C(n8807) );
  CKBD0 U8723 ( .CLK(n8776), .C(n8808) );
  CKBD0 U8724 ( .CLK(n8777), .C(n8809) );
  CKBD0 U8725 ( .CLK(n8778), .C(n8810) );
  BUFFD0 U8726 ( .I(n8782), .Z(n8811) );
  CKBD0 U8727 ( .CLK(n8779), .C(n8812) );
  CKBD0 U8728 ( .CLK(n8780), .C(n8813) );
  BUFFD0 U8729 ( .I(n8785), .Z(n8814) );
  CKBD0 U8730 ( .CLK(n8783), .C(n8815) );
  CKBD0 U8731 ( .CLK(n8794), .C(n8816) );
  CKBD0 U8732 ( .CLK(n8800), .C(n8817) );
  CKBD0 U8733 ( .CLK(n8807), .C(n8818) );
  CKBD0 U8734 ( .CLK(n8809), .C(n8819) );
  CKBD0 U8735 ( .CLK(n8810), .C(n8820) );
  BUFFD0 U8736 ( .I(n8781), .Z(n8821) );
  BUFFD0 U8737 ( .I(n8789), .Z(n8822) );
  BUFFD0 U8738 ( .I(n8790), .Z(n8823) );
  CKBD0 U8739 ( .CLK(n8812), .C(n8824) );
  CKBD0 U8740 ( .CLK(n8813), .C(n8825) );
  CKBD0 U8741 ( .CLK(n8815), .C(n8826) );
  CKBD0 U8742 ( .CLK(n8816), .C(n8827) );
  CKBD0 U8743 ( .CLK(n8817), .C(n8828) );
  CKBD0 U8744 ( .CLK(n8818), .C(n8829) );
  CKBD0 U8745 ( .CLK(n8819), .C(n8830) );
  CKBD0 U8746 ( .CLK(n8820), .C(n8831) );
  CKBD0 U8747 ( .CLK(n8824), .C(n8832) );
  CKBD0 U8748 ( .CLK(n8825), .C(n8833) );
  CKBD0 U8749 ( .CLK(n8826), .C(n8834) );
  CKBD0 U8750 ( .CLK(n8827), .C(n8835) );
  CKBD0 U8751 ( .CLK(n8828), .C(n8836) );
  BUFFD0 U8752 ( .I(n8829), .Z(n8837) );
  CKBD0 U8753 ( .CLK(n8830), .C(n8838) );
  BUFFD0 U8754 ( .I(n8831), .Z(n8839) );
  CKBD0 U8755 ( .CLK(n8787), .C(n8840) );
  CKBD0 U8756 ( .CLK(n8793), .C(n8841) );
  BUFFD0 U8757 ( .I(n8832), .Z(n8842) );
  BUFFD0 U8758 ( .I(n8833), .Z(n8843) );
  BUFFD0 U8759 ( .I(n8834), .Z(n8844) );
  BUFFD0 U8760 ( .I(n8835), .Z(n8845) );
  BUFFD0 U8761 ( .I(n8836), .Z(n8846) );
  CKBD0 U8762 ( .CLK(n8837), .C(n8847) );
  BUFFD0 U8763 ( .I(n8838), .Z(n8848) );
  CKBD0 U8764 ( .CLK(n8839), .C(n8849) );
  CKBD0 U8765 ( .CLK(n8796), .C(n8850) );
  CKBD0 U8766 ( .CLK(n8842), .C(n8851) );
  CKBD0 U8767 ( .CLK(n8843), .C(n8852) );
  CKBD0 U8768 ( .CLK(n8844), .C(n8853) );
  CKBD0 U8769 ( .CLK(n8845), .C(n8854) );
  CKBD0 U8770 ( .CLK(n8846), .C(n8855) );
  CKBD0 U8771 ( .CLK(n8847), .C(n8856) );
  CKBD0 U8772 ( .CLK(n8848), .C(n8857) );
  BUFFD0 U8773 ( .I(n8849), .Z(n8858) );
  CKBD0 U8774 ( .CLK(n8798), .C(n8859) );
  BUFFD0 U8775 ( .I(n8851), .Z(n8860) );
  BUFFD0 U8776 ( .I(n8852), .Z(n8861) );
  BUFFD0 U8777 ( .I(n8853), .Z(n8862) );
  BUFFD0 U8778 ( .I(n8854), .Z(n8863) );
  BUFFD0 U8779 ( .I(n8855), .Z(n8864) );
  BUFFD0 U8780 ( .I(n8856), .Z(n8865) );
  BUFFD0 U8781 ( .I(n8857), .Z(n8866) );
  CKBD0 U8782 ( .CLK(n8858), .C(n8867) );
  CKBD0 U8783 ( .CLK(n8860), .C(n8868) );
  CKBD0 U8784 ( .CLK(n8861), .C(n8869) );
  CKBD0 U8785 ( .CLK(n8862), .C(n8870) );
  CKBD0 U8786 ( .CLK(n8863), .C(n8871) );
  CKBD0 U8787 ( .CLK(n8864), .C(n8872) );
  CKBD0 U8788 ( .CLK(n8865), .C(n8873) );
  CKBD0 U8789 ( .CLK(n8866), .C(n8874) );
  BUFFD0 U8790 ( .I(n8867), .Z(n8875) );
  CKBD0 U8791 ( .CLK(n8804), .C(n8876) );
  BUFFD0 U8792 ( .I(n8868), .Z(n8877) );
  BUFFD0 U8793 ( .I(n8869), .Z(n8878) );
  BUFFD0 U8794 ( .I(n8870), .Z(n8879) );
  BUFFD0 U8795 ( .I(n8871), .Z(n8880) );
  BUFFD0 U8796 ( .I(n8872), .Z(n8881) );
  BUFFD0 U8797 ( .I(n8873), .Z(n8882) );
  BUFFD0 U8798 ( .I(n8874), .Z(n8883) );
  CKBD0 U8799 ( .CLK(n8875), .C(n8884) );
  CKBD0 U8800 ( .CLK(n8877), .C(n8885) );
  CKBD0 U8801 ( .CLK(n8878), .C(n8886) );
  CKBD0 U8802 ( .CLK(n8879), .C(n8887) );
  CKBD0 U8803 ( .CLK(n8880), .C(n8888) );
  CKBD0 U8804 ( .CLK(n8881), .C(n8889) );
  CKBD0 U8805 ( .CLK(n8882), .C(n8890) );
  CKBD0 U8806 ( .CLK(n8883), .C(n8891) );
  BUFFD0 U8807 ( .I(n8884), .Z(n8892) );
  CKBD0 U8808 ( .CLK(n8799), .C(n8893) );
  BUFFD0 U8809 ( .I(n8788), .Z(n8894) );
  BUFFD0 U8810 ( .I(n8784), .Z(n8895) );
  BUFFD0 U8811 ( .I(n8786), .Z(n8896) );
  BUFFD0 U8812 ( .I(n8885), .Z(n8897) );
  BUFFD0 U8813 ( .I(n8886), .Z(n8898) );
  BUFFD0 U8814 ( .I(n8795), .Z(n8899) );
  BUFFD0 U8815 ( .I(n8791), .Z(n8900) );
  CKBD0 U8816 ( .CLK(n8802), .C(n8901) );
  BUFFD0 U8817 ( .I(n8887), .Z(n8902) );
  CKBD0 U8818 ( .CLK(n8806), .C(n8903) );
  CKBD0 U8819 ( .CLK(n8805), .C(n8904) );
  BUFFD0 U8820 ( .I(n8792), .Z(n8905) );
  BUFFD0 U8821 ( .I(n8888), .Z(n8906) );
  BUFFD0 U8822 ( .I(n8803), .Z(n8907) );
  BUFFD0 U8823 ( .I(n8801), .Z(n8908) );
  BUFFD0 U8824 ( .I(n8797), .Z(n8909) );
  BUFFD0 U8825 ( .I(n8889), .Z(n8910) );
  BUFFD0 U8826 ( .I(n8890), .Z(n8911) );
  CKBD0 U8827 ( .CLK(n8811), .C(n8912) );
  CKBD0 U8828 ( .CLK(n8814), .C(n8913) );
  BUFFD0 U8829 ( .I(n8891), .Z(n8914) );
  CKBD0 U8830 ( .CLK(n8892), .C(n8915) );
  CKBD0 U8831 ( .CLK(n8897), .C(n8916) );
  CKBD0 U8832 ( .CLK(n8898), .C(n8917) );
  CKBD0 U8833 ( .CLK(n8902), .C(n8918) );
  CKBD0 U8834 ( .CLK(n8906), .C(n8919) );
  CKBD0 U8835 ( .CLK(n8910), .C(n8920) );
  CKBD0 U8836 ( .CLK(n8911), .C(n8921) );
  CKBD0 U8837 ( .CLK(n8914), .C(n8922) );
  BUFFD0 U8838 ( .I(n8915), .Z(n8923) );
  BUFFD0 U8839 ( .I(n8916), .Z(n8924) );
  BUFFD0 U8840 ( .I(n8917), .Z(n8925) );
  BUFFD0 U8841 ( .I(n8918), .Z(n8926) );
  BUFFD0 U8842 ( .I(n8919), .Z(n8927) );
  BUFFD0 U8843 ( .I(n8920), .Z(n8928) );
  BUFFD0 U8844 ( .I(n8921), .Z(n8929) );
  CKBD0 U8845 ( .CLK(n8822), .C(n8930) );
  CKBD0 U8846 ( .CLK(n8823), .C(n8931) );
  BUFFD0 U8847 ( .I(n8922), .Z(n8932) );
  CKBD0 U8848 ( .CLK(n8923), .C(n8933) );
  CKBD0 U8849 ( .CLK(n8924), .C(n8934) );
  CKBD0 U8850 ( .CLK(n8925), .C(n8935) );
  CKBD0 U8851 ( .CLK(n8926), .C(n8936) );
  CKBD0 U8852 ( .CLK(n8927), .C(n8937) );
  CKBD0 U8853 ( .CLK(n8928), .C(n8938) );
  CKBD0 U8854 ( .CLK(n8929), .C(n8939) );
  CKBD0 U8855 ( .CLK(n8932), .C(n8940) );
  BUFFD0 U8856 ( .I(n8933), .Z(n8941) );
  BUFFD0 U8857 ( .I(n8934), .Z(n8942) );
  BUFFD0 U8858 ( .I(n8935), .Z(n8943) );
  BUFFD0 U8859 ( .I(n8936), .Z(n8944) );
  BUFFD0 U8860 ( .I(n8937), .Z(n8945) );
  BUFFD0 U8861 ( .I(n8938), .Z(n8946) );
  BUFFD0 U8862 ( .I(n8939), .Z(n8947) );
  BUFFD0 U8863 ( .I(n8940), .Z(n8948) );
  BUFFD0 U8864 ( .I(n8808), .Z(n8949) );
  CKBD0 U8865 ( .CLK(n8941), .C(n8950) );
  CKBD0 U8866 ( .CLK(n8821), .C(n8951) );
  CKBD0 U8867 ( .CLK(n8942), .C(n8952) );
  CKBD0 U8868 ( .CLK(n8943), .C(n8953) );
  CKBD0 U8869 ( .CLK(n8894), .C(n8954) );
  CKBD0 U8870 ( .CLK(n8895), .C(n8955) );
  CKBD0 U8871 ( .CLK(n8896), .C(n8956) );
  CKBD0 U8872 ( .CLK(n8944), .C(n8957) );
  CKBD0 U8873 ( .CLK(n8899), .C(n8958) );
  CKBD0 U8874 ( .CLK(n8900), .C(n8959) );
  BUFFD0 U8875 ( .I(n8840), .Z(n8960) );
  CKBD0 U8876 ( .CLK(n8945), .C(n8961) );
  BUFFD0 U8877 ( .I(n8841), .Z(n8962) );
  BUFFD0 U8878 ( .I(n8850), .Z(n8963) );
  BUFFD0 U8879 ( .I(n8859), .Z(n8964) );
  CKBD0 U8880 ( .CLK(n8905), .C(n8965) );
  BUFFD0 U8881 ( .I(n8893), .Z(n8966) );
  CKBD0 U8882 ( .CLK(n8907), .C(n8967) );
  CKBD0 U8883 ( .CLK(n8946), .C(n8968) );
  CKBD0 U8884 ( .CLK(n8908), .C(n8969) );
  BUFFD0 U8885 ( .I(n8876), .Z(n8970) );
  CKBD0 U8886 ( .CLK(n8909), .C(n8971) );
  BUFFD0 U8887 ( .I(n8901), .Z(n8972) );
  BUFFD0 U8888 ( .I(n8903), .Z(n8973) );
  BUFFD0 U8889 ( .I(n8904), .Z(n8974) );
  CKBD0 U8890 ( .CLK(n8947), .C(n8975) );
  CKBD0 U8891 ( .CLK(n8948), .C(n8976) );
  CKBD0 U8892 ( .CLK(n8949), .C(n8977) );
  BUFFD0 U8893 ( .I(n8912), .Z(n8978) );
  BUFFD0 U8894 ( .I(n8913), .Z(n8979) );
  BUFFD0 U8895 ( .I(n8930), .Z(n8980) );
  BUFFD0 U8896 ( .I(n8950), .Z(n8981) );
  BUFFD0 U8897 ( .I(n8931), .Z(n8982) );
  BUFFD0 U8898 ( .I(n8952), .Z(n8983) );
  BUFFD0 U8899 ( .I(n8953), .Z(n8984) );
  BUFFD0 U8900 ( .I(n8957), .Z(n8985) );
  BUFFD0 U8901 ( .I(n8961), .Z(n8986) );
  BUFFD0 U8902 ( .I(n8968), .Z(n8987) );
  BUFFD0 U8903 ( .I(n8951), .Z(n8988) );
  BUFFD0 U8904 ( .I(n8954), .Z(n8989) );
  BUFFD0 U8905 ( .I(n8955), .Z(n8990) );
  BUFFD0 U8906 ( .I(n8956), .Z(n8991) );
  BUFFD0 U8907 ( .I(n8958), .Z(n8992) );
  BUFFD0 U8908 ( .I(n8959), .Z(n8993) );
  BUFFD0 U8909 ( .I(n8975), .Z(n8994) );
  BUFFD0 U8910 ( .I(n8976), .Z(n8995) );
  BUFFD0 U8911 ( .I(n8965), .Z(n8996) );
  BUFFD0 U8912 ( .I(n8971), .Z(n8997) );
  CKBD0 U8913 ( .CLK(n8981), .C(n8998) );
  CKBD0 U8914 ( .CLK(n8983), .C(n8999) );
  CKBD0 U8915 ( .CLK(n8984), .C(n9000) );
  CKBD0 U8916 ( .CLK(n8985), .C(n9001) );
  CKBD0 U8917 ( .CLK(n8986), .C(n9002) );
  CKBD0 U8918 ( .CLK(n8987), .C(n9003) );
  CKBD0 U8919 ( .CLK(n8994), .C(n9004) );
  CKBD0 U8920 ( .CLK(n8995), .C(n9005) );
  BUFFD0 U8921 ( .I(n8998), .Z(n9006) );
  BUFFD0 U8922 ( .I(n8969), .Z(n9007) );
  BUFFD0 U8923 ( .I(n8967), .Z(n9008) );
  BUFFD0 U8924 ( .I(n8999), .Z(n9009) );
  BUFFD0 U8925 ( .I(n9000), .Z(n9010) );
  BUFFD0 U8926 ( .I(n9001), .Z(n9011) );
  BUFFD0 U8927 ( .I(n8977), .Z(n9012) );
  BUFFD0 U8928 ( .I(n9002), .Z(n9013) );
  BUFFD0 U8929 ( .I(n9003), .Z(n9014) );
  BUFFD0 U8930 ( .I(n9004), .Z(n9015) );
  BUFFD0 U8931 ( .I(n9005), .Z(n9016) );
  BUFFD0 U8932 ( .I(n9126), .Z(n9017) );
  BUFFD0 U8933 ( .I(n13), .Z(n9018) );
  INR2XD0 U8934 ( .A1(n9027), .B1(n9127), .ZN(n97) );
  BUFFD0 U8935 ( .I(n9020), .Z(n9019) );
  BUFFD0 U8936 ( .I(n97), .Z(n9020) );
  CKBD0 U8937 ( .CLK(ParValidTimer[1]), .C(n9021) );
  BUFFD0 U8938 ( .I(n98), .Z(n9022) );
  BUFFD0 U8939 ( .I(n9024), .Z(n9023) );
  BUFFD0 U8940 ( .I(n8), .Z(n9024) );
  BUFFD1 U8941 ( .I(n9147), .Z(n9150) );
  BUFFD1 U8942 ( .I(n9151), .Z(n9149) );
  BUFFD1 U8943 ( .I(n9151), .Z(n9148) );
  BUFFD1 U8944 ( .I(n9152), .Z(n9147) );
  BUFFD1 U8945 ( .I(n9153), .Z(n9151) );
  BUFFD1 U8946 ( .I(n9153), .Z(n9152) );
  BUFFD1 U8947 ( .I(n9154), .Z(n9153) );
  INVD1 U8948 ( .I(Reset), .ZN(n9154) );
  INVD1 U8949 ( .I(n9018), .ZN(n9126) );
  BUFFD1 U8950 ( .I(n9130), .Z(n9137) );
  BUFFD1 U8951 ( .I(n9130), .Z(n9138) );
  BUFFD1 U8952 ( .I(n9131), .Z(n9139) );
  BUFFD1 U8953 ( .I(n9131), .Z(n9140) );
  BUFFD1 U8954 ( .I(n9132), .Z(n9141) );
  BUFFD1 U8955 ( .I(n9132), .Z(n9142) );
  BUFFD1 U8956 ( .I(n9133), .Z(n9143) );
  BUFFD1 U8957 ( .I(n9133), .Z(n9144) );
  BUFFD1 U8958 ( .I(n9134), .Z(n9145) );
  BUFFD1 U8959 ( .I(n9134), .Z(n9146) );
  INVD1 U8960 ( .I(n231), .ZN(n9127) );
  INVD1 U8961 ( .I(n231), .ZN(n9128) );
  INVD1 U8962 ( .I(n231), .ZN(n9129) );
  BUFFD1 U8963 ( .I(n9135), .Z(n9132) );
  BUFFD1 U8964 ( .I(n9135), .Z(n9133) );
  BUFFD1 U8965 ( .I(n9131), .Z(n9134) );
  BUFFD1 U8966 ( .I(n9136), .Z(n9130) );
  BUFFD1 U8967 ( .I(n9136), .Z(n9131) );
  IND2D1 U8968 ( .A1(n14), .B1(n15), .ZN(n13) );
  NR2D1 U8969 ( .A1(n15), .A2(n14), .ZN(N47) );
  BUFFD1 U8970 ( .I(SerClock), .Z(n9135) );
  BUFFD1 U8971 ( .I(SerClock), .Z(n9136) );
  NR2D1 U8972 ( .A1(ParClk), .A2(n232), .ZN(n3) );
  NR2D1 U8973 ( .A1(ParClk), .A2(n27), .ZN(N37) );
  NR4D0 U8974 ( .A1(n28), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n26) );
  AN2D1 U8975 ( .A1(N34), .A2(n2), .Z(N42) );
  AN2D1 U8976 ( .A1(N33), .A2(n2), .Z(N41) );
  AN2D1 U8977 ( .A1(N32), .A2(n2), .Z(N40) );
  AN2D1 U8978 ( .A1(N31), .A2(n2), .Z(N39) );
  INVD1 U8979 ( .I(n9021), .ZN(n7) );
  AO22D0 U8980 ( .A1(n6891), .A2(n9126), .B1(n6756), .B2(n9018), .Z(n133) );
  AO22D0 U8981 ( .A1(n6754), .A2(n9126), .B1(n6619), .B2(n9018), .Z(n134) );
  AO22D0 U8982 ( .A1(n6617), .A2(n9017), .B1(n6482), .B2(n9018), .Z(n135) );
  AO22D0 U8983 ( .A1(n6480), .A2(n9017), .B1(n6345), .B2(n9018), .Z(n136) );
  AO22D0 U8984 ( .A1(n6343), .A2(n9017), .B1(n6208), .B2(n9018), .Z(n137) );
  AO22D0 U8985 ( .A1(n6206), .A2(n9017), .B1(n6071), .B2(n9018), .Z(n138) );
  AO22D0 U8986 ( .A1(n6069), .A2(n9017), .B1(n5933), .B2(n9018), .Z(n139) );
  AO22D0 U8987 ( .A1(n5932), .A2(n9017), .B1(Decoder[7]), .B2(n9018), .Z(n140)
         );
  AO22D0 U8988 ( .A1(n5796), .A2(n9126), .B1(n5660), .B2(n9018), .Z(n141) );
  AO22D0 U8989 ( .A1(n5659), .A2(n9017), .B1(n5523), .B2(n13), .Z(n142) );
  AO22D0 U8990 ( .A1(n5522), .A2(n9017), .B1(Decoder[10]), .B2(n13), .Z(n143)
         );
  AO22D0 U8991 ( .A1(n5386), .A2(n9126), .B1(Decoder[11]), .B2(n9018), .Z(n144) );
  AO22D0 U8992 ( .A1(n5250), .A2(n9017), .B1(Decoder[12]), .B2(n13), .Z(n145)
         );
  AO22D0 U8993 ( .A1(n5114), .A2(n9017), .B1(Decoder[13]), .B2(n13), .Z(n146)
         );
  AO22D0 U8994 ( .A1(n4978), .A2(n9017), .B1(Decoder[14]), .B2(n13), .Z(n147)
         );
  AO22D0 U8995 ( .A1(n4842), .A2(n9126), .B1(Decoder[15]), .B2(n13), .Z(n148)
         );
  AO22D0 U8996 ( .A1(n4706), .A2(n9126), .B1(Decoder[16]), .B2(n13), .Z(n149)
         );
  AO22D0 U8997 ( .A1(n4570), .A2(n9126), .B1(Decoder[17]), .B2(n9018), .Z(n150) );
  AO22D0 U8998 ( .A1(n4434), .A2(n9126), .B1(Decoder[18]), .B2(n9018), .Z(n151) );
  AO22D0 U8999 ( .A1(n4298), .A2(n9126), .B1(Decoder[19]), .B2(n13), .Z(n152)
         );
  AO22D0 U9000 ( .A1(n4162), .A2(n9126), .B1(Decoder[20]), .B2(n9018), .Z(n153) );
  AO22D0 U9001 ( .A1(n4026), .A2(n9126), .B1(Decoder[21]), .B2(n13), .Z(n154)
         );
  AO22D0 U9002 ( .A1(n3890), .A2(n9017), .B1(Decoder[22]), .B2(n13), .Z(n155)
         );
  AO22D0 U9003 ( .A1(n3754), .A2(n9126), .B1(Decoder[23]), .B2(n13), .Z(n156)
         );
  AO22D0 U9004 ( .A1(n3618), .A2(n9126), .B1(Decoder[24]), .B2(n13), .Z(n157)
         );
  AO22D0 U9005 ( .A1(n3482), .A2(n9126), .B1(Decoder[25]), .B2(n13), .Z(n158)
         );
  AO22D0 U9006 ( .A1(n3346), .A2(n9126), .B1(Decoder[26]), .B2(n13), .Z(n159)
         );
  AO22D0 U9007 ( .A1(n3210), .A2(n9126), .B1(Decoder[27]), .B2(n13), .Z(n160)
         );
  AO22D0 U9008 ( .A1(n3074), .A2(n9017), .B1(Decoder[28]), .B2(n13), .Z(n161)
         );
  AO22D0 U9009 ( .A1(n2938), .A2(n9126), .B1(Decoder[29]), .B2(n13), .Z(n162)
         );
  AO22D0 U9010 ( .A1(n2802), .A2(n9126), .B1(Decoder[30]), .B2(n13), .Z(n163)
         );
  AO22D0 U9011 ( .A1(n2663), .A2(n9126), .B1(Decoder[31]), .B2(n13), .Z(n164)
         );
  OAI31D0 U9012 ( .A1(n6), .A2(n230), .A3(n7), .B(n232), .ZN(n9027) );
  NR2D1 U9013 ( .A1(n11), .A2(n9127), .ZN(n99) );
  NR2D1 U9014 ( .A1(n6897), .A2(n9127), .ZN(n100) );
  NR2D1 U9015 ( .A1(n9127), .A2(n9023), .ZN(n98) );
  XOR2D1 U9016 ( .A1(n230), .A2(n9), .Z(n8) );
  NR2D1 U9017 ( .A1(n7), .A2(n10), .ZN(n9) );
  NR4D0 U9018 ( .A1(n22), .A2(n8996), .A3(n8991), .A4(n8988), .ZN(n21) );
  NR4D0 U9019 ( .A1(n9015), .A2(n9013), .A3(n9009), .A4(n9006), .ZN(n16) );
  NR4D0 U9020 ( .A1(n9016), .A2(n9014), .A3(n9011), .A4(n9010), .ZN(n17) );
  AN4D1 U9021 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .Z(n15) );
  INR4D0 U9022 ( .A1(n8982), .B1(n25), .B2(n9008), .B3(n9012), .ZN(n18) );
  NR4D0 U9023 ( .A1(n24), .A2(n9007), .A3(n8992), .A4(n8989), .ZN(n19) );
  NR4D0 U9024 ( .A1(n23), .A2(n8997), .A3(n8993), .A4(n8990), .ZN(n20) );
  ND3D1 U9025 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n25) );
  AN2D1 U9026 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_0 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_3 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N46, N47, N48, N49, N63, N64, N65, N66,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n115, n121, n122, n124,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n140, n141, n142, n143, n144, n8;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n128), .CPN(StateClock), .Q(FullFIFO), .QN(n115) );
  DFND1 EmptyFIFOr_reg ( .D(n127), .CPN(StateClock), .Q(EmptyFIFO) );
  IAO21D1 U6 ( .A1(n39), .A2(n40), .B(Reset), .ZN(n38) );
  MOAI22D1 U7 ( .A1(n142), .A2(n41), .B1(n41), .B2(OldReadAr[1]), .ZN(n129) );
  MOAI22D1 U8 ( .A1(n141), .A2(n41), .B1(n41), .B2(OldReadAr[2]), .ZN(n130) );
  MOAI22D1 U9 ( .A1(n42), .A2(n43), .B1(n42), .B2(OldWriteAr[1]), .ZN(n131) );
  MOAI22D1 U10 ( .A1(n42), .A2(n44), .B1(n42), .B2(OldWriteAr[2]), .ZN(n132)
         );
  MOAI22D1 U11 ( .A1(n144), .A2(n42), .B1(n42), .B2(OldWriteAr[0]), .ZN(n133)
         );
  MOAI22D1 U70 ( .A1(n143), .A2(n41), .B1(n41), .B2(OldReadAr[0]), .ZN(n140)
         );
  DFNCND1 \NextState_reg[0]  ( .D(n137), .CPN(StateClock), .CDN(n8), .Q(
        NextState[0]), .QN(n124) );
  DFNCND1 \NextState_reg[1]  ( .D(n135), .CPN(StateClock), .CDN(n8), .Q(
        NextState[1]), .QN(n122) );
  DFNCND1 \NextState_reg[2]  ( .D(n134), .CPN(StateClock), .CDN(n8), .Q(
        NextState[2]), .QN(n121) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n8), .Q(
        CurState[2]) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n8), .Q(
        CurState[1]) );
  EDFCNQD1 \WriteAr_reg[2]  ( .D(N65), .E(N66), .CP(StateClock), .CDN(n8), .Q(
        WriteAddr[2]) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n8), .Q(
        CurState[0]) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(N64), .E(N66), .CP(StateClock), .CDN(n8), .Q(
        WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N48), .CP(StateClock), .CDN(n8), .Q(
        ReadAddr[2]), .QN(n141) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N47), .E(N48), .CP(StateClock), .CDN(n8), .Q(
        ReadAddr[1]), .QN(n142) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N46), .E(N48), .CP(StateClock), .CDN(n8), .Q(
        ReadAddr[0]), .QN(n143) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N63), .E(N66), .CP(StateClock), .CDN(n8), .Q(
        WriteAddr[0]), .QN(n144) );
  DFNCND1 WriteCmdr_reg ( .D(n136), .CPN(StateClock), .CDN(n8), .Q(WriteCmd), 
        .QN(n85) );
  DFNCND1 ReadCmdr_reg ( .D(n138), .CPN(StateClock), .CDN(n8), .Q(ReadCmd) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n131), .CPN(StateClock), .CDN(n8), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n132), .CPN(StateClock), .CDN(n8), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n133), .CPN(StateClock), .CDN(n8), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n130), .CPN(StateClock), .CDN(n8), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n129), .CPN(StateClock), .CDN(n8), .Q(
        OldReadAr[1]) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n140), .CPN(StateClock), .CDN(n8), .Q(
        OldReadAr[0]) );
  INVD1 U3 ( .I(Reset), .ZN(n8) );
  INVD1 U4 ( .I(n77), .ZN(n84) );
  MAOI22D0 U5 ( .A1(ReadAddr[0]), .A2(n75), .B1(n43), .B2(n98), .ZN(n101) );
  INVD1 U12 ( .I(n40), .ZN(n35) );
  ND2D1 U13 ( .A1(n83), .A2(n37), .ZN(n86) );
  ND2D1 U14 ( .A1(WriteReq), .A2(n45), .ZN(n42) );
  ND2D1 U15 ( .A1(ReadReq), .A2(n86), .ZN(n41) );
  INVD1 U16 ( .I(n46), .ZN(n52) );
  NR2D1 U17 ( .A1(n68), .A2(n79), .ZN(n39) );
  ND2D1 U18 ( .A1(n83), .A2(n35), .ZN(n45) );
  XNR2D1 U19 ( .A1(n44), .A2(n75), .ZN(n77) );
  INVD1 U20 ( .I(n75), .ZN(n81) );
  XNR2D1 U21 ( .A1(n84), .A2(ReadAddr[2]), .ZN(n56) );
  ND3D1 U22 ( .A1(n37), .A2(n35), .A3(n112), .ZN(N66) );
  NR2D1 U23 ( .A1(ReadAddr[0]), .A2(n109), .ZN(N46) );
  NR2D1 U24 ( .A1(n99), .A2(n109), .ZN(N49) );
  NR2D1 U25 ( .A1(n113), .A2(n109), .ZN(N47) );
  XNR2D1 U26 ( .A1(ReadAddr[0]), .A2(ReadAddr[1]), .ZN(n113) );
  INVD1 U27 ( .I(ReadReq), .ZN(n106) );
  MAOI22D0 U28 ( .A1(WriteAddr[0]), .A2(n103), .B1(n142), .B2(n98), .ZN(n102)
         );
  OAI222D0 U29 ( .A1(n44), .A2(ReadAddr[2]), .B1(n43), .B2(ReadAddr[1]), .C1(
        n144), .C2(ReadAddr[0]), .ZN(n73) );
  OAI33D1 U30 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n101), .B1(n44), .B2(
        WriteAddr[1]), .B3(n102), .ZN(n54) );
  OAI33D1 U31 ( .A1(ReadAddr[1]), .A2(n101), .A3(n44), .B1(n102), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n55) );
  AOI22D0 U32 ( .A1(n68), .A2(CurState[1]), .B1(n51), .B2(n39), .ZN(n83) );
  NR3D0 U33 ( .A1(CurState[1]), .A2(CurState[2]), .A3(CurState[0]), .ZN(n40)
         );
  OAI211D1 U34 ( .A1(CurState[1]), .A2(n79), .B(n83), .C(n104), .ZN(n46) );
  AOI21D1 U35 ( .A1(WriteReq), .A2(n40), .B(n105), .ZN(n104) );
  AOI21D1 U36 ( .A1(CurState[0]), .A2(n106), .B(n68), .ZN(n105) );
  ND2D1 U37 ( .A1(CurState[1]), .A2(n39), .ZN(n37) );
  INVD1 U38 ( .I(WriteAddr[2]), .ZN(n44) );
  OAI33D1 U39 ( .A1(n85), .A2(n40), .A3(n86), .B1(n87), .B2(n88), .B3(n89), 
        .ZN(n136) );
  XNR2D1 U40 ( .A1(n44), .A2(OldWriteAr[2]), .ZN(n89) );
  XNR2D1 U41 ( .A1(n43), .A2(OldWriteAr[1]), .ZN(n88) );
  INVD1 U42 ( .I(WriteAddr[1]), .ZN(n43) );
  NR2D1 U43 ( .A1(n43), .A2(n144), .ZN(n75) );
  OAI211D1 U44 ( .A1(n144), .A2(ReadAddr[1]), .B(n80), .C(n81), .ZN(n78) );
  OAI21D1 U45 ( .A1(WriteAddr[1]), .A2(n142), .B(n143), .ZN(n80) );
  OAI21D1 U46 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n81), .ZN(n100) );
  INVD1 U47 ( .I(CurState[0]), .ZN(n79) );
  OAI32D1 U48 ( .A1(n107), .A2(n108), .A3(n106), .B1(n86), .B2(n109), .ZN(n138) );
  XNR2D1 U49 ( .A1(n142), .A2(OldReadAr[1]), .ZN(n108) );
  ND3D1 U50 ( .A1(n110), .A2(n86), .A3(n111), .ZN(n107) );
  XNR2D1 U51 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .ZN(n110) );
  XOR2D1 U52 ( .A1(n100), .A2(n142), .Z(n57) );
  INVD1 U53 ( .I(CurState[2]), .ZN(n68) );
  ND2D1 U54 ( .A1(n144), .A2(n143), .ZN(n98) );
  AOI31D0 U55 ( .A1(n65), .A2(n66), .A3(n67), .B(n68), .ZN(n64) );
  AOI22D0 U56 ( .A1(n69), .A2(ReadAddr[1]), .B1(n144), .B2(ReadAddr[0]), .ZN(
        n67) );
  OAI21D1 U57 ( .A1(n69), .A2(n73), .B(n43), .ZN(n65) );
  OAI21D1 U58 ( .A1(ReadAddr[1]), .A2(n72), .B(n73), .ZN(n66) );
  OAI22D0 U59 ( .A1(n46), .A2(n122), .B1(n52), .B2(n59), .ZN(n135) );
  AOI31D0 U60 ( .A1(n60), .A2(n61), .A3(n62), .B(n40), .ZN(n59) );
  IIND4D1 U61 ( .A1(n69), .A2(n73), .B1(n78), .B2(n79), .ZN(n61) );
  AOI31D0 U62 ( .A1(n143), .A2(CurState[0]), .A3(n63), .B(n64), .ZN(n62) );
  OAI22D0 U63 ( .A1(n46), .A2(n124), .B1(n52), .B2(n92), .ZN(n137) );
  AOI21D1 U64 ( .A1(CurState[1]), .A2(n93), .B(n39), .ZN(n92) );
  OAI21D1 U65 ( .A1(CurState[2]), .A2(n94), .B(n95), .ZN(n93) );
  AOI22D0 U66 ( .A1(n55), .A2(ReadAddr[2]), .B1(n141), .B2(n54), .ZN(n94) );
  OAI31D0 U67 ( .A1(n96), .A2(n97), .A3(n58), .B(CurState[0]), .ZN(n95) );
  XNR2D1 U68 ( .A1(WriteAddr[2]), .A2(n99), .ZN(n97) );
  INVD1 U69 ( .I(n57), .ZN(n96) );
  OAI21D1 U71 ( .A1(n46), .A2(n121), .B(n47), .ZN(n134) );
  OAI211D1 U72 ( .A1(CurState[2]), .A2(n48), .B(CurState[0]), .C(n49), .ZN(n47) );
  AOI21D1 U73 ( .A1(n50), .A2(n51), .B(n52), .ZN(n49) );
  NR4D0 U74 ( .A1(n56), .A2(n57), .A3(n51), .A4(n58), .ZN(n48) );
  INVD1 U75 ( .I(CurState[1]), .ZN(n51) );
  NR3D0 U76 ( .A1(n57), .A2(n144), .A3(n74), .ZN(n63) );
  AOI21D1 U77 ( .A1(n69), .A2(n75), .B(n76), .ZN(n74) );
  OAI32D1 U78 ( .A1(n44), .A2(n141), .A3(n75), .B1(ReadAddr[2]), .B2(n77), 
        .ZN(n76) );
  AOI31D0 U79 ( .A1(n144), .A2(CurState[0]), .A3(n82), .B(n83), .ZN(n60) );
  NR3D0 U80 ( .A1(n57), .A2(n143), .A3(n56), .ZN(n82) );
  NR2D1 U81 ( .A1(n143), .A2(n142), .ZN(n103) );
  XOR2D1 U82 ( .A1(n103), .A2(n141), .Z(n99) );
  AO22D0 U83 ( .A1(ReadAddr[2]), .A2(n54), .B1(n55), .B2(n141), .Z(n50) );
  XNR2D1 U84 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n72) );
  ND2D1 U85 ( .A1(ReadCmd), .A2(n35), .ZN(n109) );
  OAI21D1 U86 ( .A1(n144), .A2(n143), .B(n98), .ZN(n58) );
  OAI32D1 U87 ( .A1(n37), .A2(Reset), .A3(ReadReq), .B1(n38), .B2(n115), .ZN(
        n128) );
  ND2D1 U88 ( .A1(WriteCmd), .A2(n37), .ZN(n112) );
  NR2D1 U89 ( .A1(WriteAddr[2]), .A2(n141), .ZN(n69) );
  OAI22D0 U90 ( .A1(n143), .A2(n37), .B1(WriteAddr[0]), .B2(n112), .ZN(N63) );
  OAI22D0 U91 ( .A1(n141), .A2(n37), .B1(n84), .B2(n112), .ZN(N65) );
  OAI22D0 U92 ( .A1(n142), .A2(n37), .B1(n100), .B2(n112), .ZN(N64) );
  OAI31D0 U93 ( .A1(n35), .A2(WriteReq), .A3(Reset), .B(n36), .ZN(n127) );
  OAI31D0 U94 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(EmptyFIFO), 
        .ZN(n36) );
  ND3D1 U95 ( .A1(n90), .A2(n45), .A3(WriteReq), .ZN(n87) );
  XNR2D1 U96 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n90) );
  IND2D1 U97 ( .A1(ReadCmd), .B1(n35), .ZN(N48) );
  XNR2D1 U98 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n111) );
  ND2D1 U99 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid3_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockW, Dreadyr, \Storage[7][32] , \Storage[7][31] ,
         \Storage[7][30] , \Storage[7][29] , \Storage[7][28] ,
         \Storage[7][27] , \Storage[7][26] , \Storage[7][25] ,
         \Storage[7][24] , \Storage[7][23] , \Storage[7][22] ,
         \Storage[7][21] , \Storage[7][20] , \Storage[7][19] ,
         \Storage[7][18] , \Storage[7][17] , \Storage[7][16] ,
         \Storage[7][15] , \Storage[7][14] , \Storage[7][13] ,
         \Storage[7][12] , \Storage[7][11] , \Storage[7][10] , \Storage[7][9] ,
         \Storage[7][8] , \Storage[7][7] , \Storage[7][6] , \Storage[7][5] ,
         \Storage[7][4] , \Storage[7][3] , \Storage[7][2] , \Storage[7][1] ,
         \Storage[7][0] , \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N87, N99, N161, N194, N227, N260, N293,
         N326, N359, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n78) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n77) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n74) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n71) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n68) );
  XOR4D1 U21 ( .A1(n83), .A2(N74), .A3(n84), .A4(N77), .Z(n82) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n84) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n90) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n89) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n86) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n80) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(N194), .CP(n179), .CDN(
        n197), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n164), .CP(n175), .CDN(
        n203), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n164), .CP(n175), .CDN(
        n200), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n164), .CP(n175), .CDN(
        n206), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n164), .CP(n179), .CDN(
        n203), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n164), .CP(n182), .CDN(
        n206), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n164), .CP(n186), .CDN(
        n203), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n164), .CP(n174), .CDN(
        n200), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n164), .CP(n179), .CDN(
        n206), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n164), .CP(n178), .CDN(
        n203), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n164), .CP(n184), .CDN(n196), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n164), .CP(n185), .CDN(n192), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n164), .CP(ClockW), .CDN(
        n203), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n164), .CP(n184), .CDN(n192), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n164), .CP(ClockW), .CDN(
        n197), .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n164), .CP(n184), .CDN(n195), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n164), .CP(n177), .CDN(n194), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n162), .CP(n182), .CDN(n206), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(N194), .CP(n174), .CDN(n192), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(N194), .CP(n175), .CDN(n195), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n170), .CP(n181), .CDN(
        n205), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(N99), .CP(n181), .CDN(n207), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n170), .CP(n182), .CDN(
        n193), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n170), .CP(n182), .CDN(
        n202), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n170), .CP(n182), .CDN(
        n205), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n170), .CP(n182), .CDN(
        n193), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n170), .CP(n182), .CDN(
        n206), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n172), .CP(n182), .CDN(
        n201), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n172), .CP(n177), .CDN(
        n199), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n172), .CP(n184), .CDN(
        n206), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n172), .CP(n179), .CDN(n192), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n172), .CP(n180), .CDN(n192), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n172), .CP(n181), .CDN(n192), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n172), .CP(n177), .CDN(n192), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n172), .CP(n174), .CDN(n192), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n172), .CP(n186), .CDN(n192), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n172), .CP(n185), .CDN(n192), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n170), .CP(n183), .CDN(n192), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n170), .CP(n183), .CDN(n192), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n170), .CP(n183), .CDN(n192), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n146), .CP(n175), .CDN(
        n200), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n148), .CP(ClockW), .CDN(
        n200), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n148), .CP(n177), .CDN(
        n202), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n148), .CP(n178), .CDN(
        n200), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n148), .CP(n174), .CDN(
        n200), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n148), .CP(ClockW), .CDN(
        n194), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n148), .CP(n185), .CDN(
        n201), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n148), .CP(n183), .CDN(
        n202), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n148), .CP(n183), .CDN(
        n204), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n148), .CP(n184), .CDN(
        n201), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n148), .CP(n186), .CDN(n192), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n148), .CP(n185), .CDN(n206), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n148), .CP(n174), .CDN(n206), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n148), .CP(n177), .CDN(n206), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n148), .CP(n182), .CDN(n201), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n148), .CP(n179), .CDN(n207), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n148), .CP(n180), .CDN(n204), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(N326), .CP(n178), .CDN(n205), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(N326), .CP(n178), .CDN(n202), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(N326), .CP(n178), .CDN(n207), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(N293), .CP(n185), .CDN(
        n197), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n152), .CP(n184), .CDN(
        n196), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n152), .CP(n179), .CDN(
        n199), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n152), .CP(n176), .CDN(
        n199), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n152), .CP(n186), .CDN(
        n199), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n152), .CP(n184), .CDN(
        n199), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n152), .CP(ClockW), .CDN(
        n199), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n152), .CP(n176), .CDN(
        n199), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n152), .CP(n179), .CDN(
        n199), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n152), .CP(n176), .CDN(
        n199), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n152), .CP(n182), .CDN(n205), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n152), .CP(n174), .CDN(n198), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n152), .CP(n174), .CDN(n201), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n152), .CP(n180), .CDN(n205), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n152), .CP(n183), .CDN(n205), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n152), .CP(n176), .CDN(n197), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n152), .CP(n186), .CDN(n192), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n150), .CP(n178), .CDN(n206), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(N293), .CP(n185), .CDN(n205), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(N293), .CP(n179), .CDN(n207), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(N260), .CP(n176), .CDN(
        n198), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n156), .CP(n181), .CDN(
        n198), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n156), .CP(n178), .CDN(
        n206), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n156), .CP(n178), .CDN(
        n198), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n156), .CP(n176), .CDN(
        n198), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n156), .CP(n183), .CDN(
        n198), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n156), .CP(n182), .CDN(
        n205), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n156), .CP(n175), .CDN(
        n202), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n156), .CP(n181), .CDN(
        n207), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n156), .CP(n178), .CDN(
        n199), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n156), .CP(n183), .CDN(n197), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n156), .CP(n186), .CDN(n197), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n156), .CP(ClockW), .CDN(
        n197), .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n156), .CP(n175), .CDN(n197), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n156), .CP(n174), .CDN(n197), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n156), .CP(n185), .CDN(n197), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n156), .CP(n175), .CDN(n197), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n154), .CP(n181), .CDN(n197), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(N260), .CP(n185), .CDN(n197), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(N260), .CP(ClockW), .CDN(
        n197), .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(N227), .CP(n178), .CDN(
        n196), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n160), .CP(n184), .CDN(
        n196), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n160), .CP(n185), .CDN(
        n195), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n160), .CP(n181), .CDN(
        n195), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n160), .CP(ClockW), .CDN(
        n195), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n160), .CP(n178), .CDN(
        n195), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n160), .CP(n183), .CDN(
        n195), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n160), .CP(n179), .CDN(
        n195), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n160), .CP(n174), .CDN(
        n195), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n160), .CP(n175), .CDN(
        n195), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n160), .CP(n184), .CDN(n194), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n160), .CP(n186), .CDN(n194), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n160), .CP(n175), .CDN(n194), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n160), .CP(n183), .CDN(n194), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n160), .CP(n185), .CDN(n194), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n160), .CP(n174), .CDN(n194), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n160), .CP(n186), .CDN(n194), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n158), .CP(n185), .CDN(n194), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(N227), .CP(n184), .CDN(n194), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(N227), .CP(n183), .CDN(n194), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n166), .CP(n174), .CDN(
        n196), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n168), .CP(n181), .CDN(
        n193), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n168), .CP(n174), .CDN(
        n193), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n168), .CP(n181), .CDN(
        n193), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n168), .CP(n182), .CDN(
        n193), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n168), .CP(n179), .CDN(
        n193), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n168), .CP(n179), .CDN(
        n193), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n168), .CP(n179), .CDN(
        n193), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n166), .CP(n179), .CDN(
        n193), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n166), .CP(n179), .CDN(
        n193), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n166), .CP(n179), .CDN(n207), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n166), .CP(n179), .CDN(n198), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n166), .CP(n179), .CDN(n207), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n168), .CP(n179), .CDN(n198), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n168), .CP(n180), .CDN(n193), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n168), .CP(n180), .CDN(n196), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n168), .CP(n180), .CDN(n195), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(N161), .CP(n180), .CDN(n207), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n166), .CP(n180), .CDN(n204), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n166), .CP(n180), .CDN(n196), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(N359), .CP(n177), .CDN(
        n202), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n144), .CP(n177), .CDN(
        n202), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n144), .CP(n177), .CDN(
        n201), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(N359), .CP(n177), .CDN(
        n201), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(N359), .CP(n177), .CDN(
        n201), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(N359), .CP(n183), .CDN(
        n201), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(N359), .CP(n177), .CDN(
        n201), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n144), .CP(n182), .CDN(
        n201), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n144), .CP(n176), .CDN(
        n201), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n144), .CP(n175), .CDN(
        n201), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n144), .CP(n181), .CDN(n199), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n144), .CP(n182), .CDN(n200), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n144), .CP(n179), .CDN(n193), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n144), .CP(n180), .CDN(n199), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n144), .CP(n176), .CDN(n206), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n144), .CP(n184), .CDN(n204), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n144), .CP(n174), .CDN(n205), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n144), .CP(n182), .CDN(n195), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n142), .CP(n183), .CDN(n198), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n142), .CP(n184), .CDN(n199), 
        .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n2), .CP(n187), .CDN(n192), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N87), .E(N194), .CP(n177), .CDN(n194), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(N194), .CP(n174), .CDN(
        n192), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(N194), .CP(n180), .CDN(
        n204), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(N194), .CP(n180), .CDN(
        n200), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n162), .CP(ClockW), .CDN(
        n207), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n162), .CP(n186), .CDN(
        n192), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n162), .CP(n180), .CDN(
        n207), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n162), .CP(n184), .CDN(
        n205), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n162), .CP(n186), .CDN(
        n196), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n164), .CP(n185), .CDN(
        n193), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n164), .CP(n184), .CDN(
        n197), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n164), .CP(ClockW), .CDN(
        n206), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n164), .CP(n174), .CDN(
        n203), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N87), .E(n170), .CP(n180), .CDN(n195), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n170), .CP(n180), .CDN(
        n207), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n170), .CP(n180), .CDN(
        n207), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(N99), .CP(n181), .CDN(n207), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(N99), .CP(n181), .CDN(n207), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n170), .CP(n181), .CDN(
        n205), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N99), .CP(n181), .CDN(n199), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n170), .CP(n181), .CDN(
        n207), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n170), .CP(n181), .CDN(
        n194), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n170), .CP(n181), .CDN(
        n203), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(N99), .CP(n182), .CDN(n197), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(N99), .CP(n182), .CDN(n193), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(N99), .CP(n182), .CDN(n206), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N87), .E(N326), .CP(n175), .CDN(n206), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(N326), .CP(ClockW), .CDN(
        n200), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(N326), .CP(n185), .CDN(
        n200), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n146), .CP(n186), .CDN(
        n200), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n146), .CP(n185), .CDN(
        n200), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n146), .CP(n176), .CDN(
        n200), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(N326), .CP(n178), .CDN(
        n200), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n146), .CP(n182), .CDN(
        n200), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n146), .CP(n176), .CDN(
        n200), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n148), .CP(n175), .CDN(
        n200), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n148), .CP(n184), .CDN(
        n204), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n148), .CP(n175), .CDN(
        n192), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n148), .CP(n186), .CDN(
        n203), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N87), .E(N293), .CP(n178), .CDN(n200), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(N293), .CP(n178), .CDN(
        n206), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(N293), .CP(n178), .CDN(
        n192), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(N293), .CP(n178), .CDN(
        n202), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n150), .CP(n178), .CDN(
        n200), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n150), .CP(n178), .CDN(
        n194), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n150), .CP(n183), .CDN(
        n196), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n150), .CP(n181), .CDN(
        n206), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n150), .CP(n174), .CDN(
        n193), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n152), .CP(n174), .CDN(
        n196), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n152), .CP(n181), .CDN(
        n199), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n152), .CP(ClockW), .CDN(
        n199), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n152), .CP(n175), .CDN(
        n199), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N87), .E(N260), .CP(n177), .CDN(n205), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(N260), .CP(ClockW), .CDN(
        n198), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(N260), .CP(n184), .CDN(
        n198), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(N260), .CP(n183), .CDN(
        n198), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n154), .CP(n178), .CDN(
        n198), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n154), .CP(n186), .CDN(
        n198), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n154), .CP(n175), .CDN(
        n198), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n154), .CP(n185), .CDN(
        n198), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n154), .CP(n186), .CDN(
        n198), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n156), .CP(n175), .CDN(
        n198), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n156), .CP(n186), .CDN(
        n195), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n156), .CP(n183), .CDN(
        n202), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n156), .CP(n181), .CDN(
        n201), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N87), .E(N227), .CP(n185), .CDN(n197), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(N227), .CP(n182), .CDN(
        n196), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(N227), .CP(n184), .CDN(
        n196), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(N227), .CP(n179), .CDN(
        n196), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n158), .CP(ClockW), .CDN(
        n196), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n158), .CP(n184), .CDN(
        n196), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n158), .CP(n185), .CDN(
        n196), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n158), .CP(n180), .CDN(
        n196), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n158), .CP(n175), .CDN(
        n196), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n160), .CP(n183), .CDN(
        n196), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n160), .CP(n186), .CDN(
        n195), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n160), .CP(n177), .CDN(
        n195), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n160), .CP(n183), .CDN(
        n195), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N87), .E(n166), .CP(n177), .CDN(n204), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(N161), .CP(n176), .CDN(
        n195), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(N161), .CP(n185), .CDN(
        n195), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(N161), .CP(n186), .CDN(
        n196), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(N161), .CP(n180), .CDN(
        n194), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(N161), .CP(n180), .CDN(
        n204), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(N161), .CP(n177), .CDN(
        n207), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n166), .CP(n184), .CDN(
        n205), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n166), .CP(n180), .CDN(
        n204), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n168), .CP(n175), .CDN(
        n195), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n168), .CP(n186), .CDN(
        n193), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n168), .CP(n183), .CDN(
        n193), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n168), .CP(ClockW), .CDN(
        n193), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N87), .E(n142), .CP(n176), .CDN(n201), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n142), .CP(n176), .CDN(
        n202), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(N359), .CP(n177), .CDN(
        n202), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(N359), .CP(n177), .CDN(
        n201), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n144), .CP(n177), .CDN(
        n201), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n144), .CP(n177), .CDN(
        n201), .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N53), .E(n189), .CP(n187), .CDN(n197), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N54), .E(n189), .CP(n187), .CDN(n206), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N55), .E(n189), .CP(n188), .CDN(n193), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N56), .E(n189), .CP(n187), .CDN(n198), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N57), .E(n189), .CP(n188), .CDN(n206), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N58), .E(n189), .CP(n188), .CDN(n194), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N59), .E(n189), .CP(n188), .CDN(n197), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N60), .E(n189), .CP(n187), .CDN(n205), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N61), .E(n189), .CP(n188), .CDN(n199), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N62), .E(n189), .CP(n187), .CDN(n194), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N63), .E(n189), .CP(n187), .CDN(n205), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N64), .E(n189), .CP(n187), .CDN(n198), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N65), .E(n189), .CP(n187), .CDN(n203), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N66), .E(n189), .CP(n187), .CDN(n203), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N67), .E(n189), .CP(n187), .CDN(n203), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N68), .E(n189), .CP(n187), .CDN(n203), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N69), .E(n189), .CP(n187), .CDN(n203), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N70), .E(Read), .CP(n187), .CDN(n203), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N71), .E(Read), .CP(n188), .CDN(n203), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N72), .E(Read), .CP(n188), .CDN(n203), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N73), .E(Read), .CP(n188), .CDN(n203), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N74), .E(Read), .CP(n188), .CDN(n203), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N75), .E(Read), .CP(n188), .CDN(n203), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N76), .E(Read), .CP(n188), .CDN(n204), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N77), .E(Read), .CP(n188), .CDN(n205), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N78), .E(Read), .CP(n188), .CDN(n204), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N79), .E(Read), .CP(n188), .CDN(n200), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N80), .E(Read), .CP(n188), .CDN(n201), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N81), .E(Read), .CP(n187), .CDN(n202), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N82), .E(Read), .CP(n188), .CDN(n202), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N83), .E(Read), .CP(n188), .CDN(n201), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N84), .E(Read), .CP(n187), .CDN(n205), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N85), .E(Read), .CP(n187), .CDN(n199), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  INVD0 U3 ( .I(n142), .ZN(n145) );
  CKND0 U4 ( .CLK(n143), .CN(n142) );
  CKBD0 U5 ( .CLK(N49), .C(n136) );
  CKBXD0 U6 ( .I(n191), .Z(n137) );
  CKBD0 U7 ( .CLK(N48), .C(n191) );
  INVD0 U8 ( .I(N99), .ZN(n171) );
  CKND2D0 U9 ( .A1(ClkR), .A2(ChipEna), .ZN(n1) );
  INVD0 U10 ( .I(N161), .ZN(n167) );
  CKNXD0 U11 ( .I(n167), .ZN(n166) );
  CKNXD0 U12 ( .I(n155), .ZN(n154) );
  CKNXD0 U18 ( .I(n151), .ZN(n150) );
  CKNXD0 U19 ( .I(n159), .ZN(n158) );
  INVD0 U20 ( .I(N326), .ZN(n147) );
  CKNXD0 U23 ( .I(n147), .ZN(n146) );
  CKNXD0 U24 ( .I(n163), .ZN(n162) );
  CKAN2D0 U25 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U26 ( .I(N50), .ZN(n130) );
  BUFFD1 U31 ( .I(n206), .Z(n194) );
  BUFFD1 U32 ( .I(n204), .Z(n195) );
  BUFFD1 U33 ( .I(n204), .Z(n196) );
  BUFFD1 U34 ( .I(n205), .Z(n197) );
  BUFFD1 U35 ( .I(n204), .Z(n198) );
  BUFFD1 U36 ( .I(n205), .Z(n199) );
  BUFFD1 U37 ( .I(n204), .Z(n200) );
  BUFFD1 U38 ( .I(n204), .Z(n201) );
  BUFFD1 U39 ( .I(n204), .Z(n202) );
  BUFFD1 U40 ( .I(n205), .Z(n203) );
  BUFFD1 U41 ( .I(n207), .Z(n192) );
  BUFFD1 U42 ( .I(n204), .Z(n193) );
  BUFFD1 U43 ( .I(n207), .Z(n206) );
  BUFFD1 U44 ( .I(n207), .Z(n205) );
  BUFFD1 U45 ( .I(n207), .Z(n204) );
  INVD1 U46 ( .I(Reset), .ZN(n207) );
  BUFFD1 U47 ( .I(ClockW), .Z(n178) );
  BUFFD1 U48 ( .I(n183), .Z(n177) );
  BUFFD1 U49 ( .I(n178), .Z(n176) );
  INVD1 U50 ( .I(n165), .ZN(n164) );
  INVD1 U51 ( .I(n161), .ZN(n160) );
  INVD1 U52 ( .I(n149), .ZN(n148) );
  INVD1 U53 ( .I(n145), .ZN(n144) );
  BUFFD1 U54 ( .I(n185), .Z(n182) );
  BUFFD1 U55 ( .I(n185), .Z(n181) );
  BUFFD1 U56 ( .I(n186), .Z(n180) );
  BUFFD1 U57 ( .I(n186), .Z(n179) );
  BUFFD1 U58 ( .I(n184), .Z(n183) );
  BUFFD1 U59 ( .I(n138), .Z(n140) );
  BUFFD1 U60 ( .I(n133), .Z(n135) );
  BUFFD1 U61 ( .I(N49), .Z(n134) );
  BUFFD1 U62 ( .I(n136), .Z(n133) );
  INVD1 U63 ( .I(n158), .ZN(n161) );
  INVD1 U64 ( .I(n146), .ZN(n149) );
  INVD1 U65 ( .I(n162), .ZN(n165) );
  INVD1 U66 ( .I(n173), .ZN(n172) );
  INVD1 U67 ( .I(n169), .ZN(n168) );
  INVD1 U68 ( .I(n157), .ZN(n156) );
  INVD1 U69 ( .I(n153), .ZN(n152) );
  BUFFD1 U70 ( .I(n174), .Z(n184) );
  BUFFD1 U71 ( .I(n174), .Z(n185) );
  BUFFD1 U72 ( .I(n174), .Z(n186) );
  INVD1 U73 ( .I(n1), .ZN(n188) );
  INVD1 U74 ( .I(n1), .ZN(n187) );
  XOR3D1 U75 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n76), .Z(n75) );
  XOR3D1 U76 ( .A1(n77), .A2(DataI[17]), .A3(n78), .Z(n76) );
  XOR3D1 U77 ( .A1(n71), .A2(DataI[3]), .A3(n72), .Z(n70) );
  XOR3D1 U78 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n73), .Z(n72) );
  XOR3D1 U79 ( .A1(n74), .A2(DataI[10]), .A3(n75), .Z(n73) );
  XOR3D1 U80 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n67), .Z(N87) );
  XOR3D1 U81 ( .A1(DataI[0]), .A2(n68), .A3(n69), .Z(n67) );
  XOR3D1 U82 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n70), .Z(n69) );
  XOR3D1 U83 ( .A1(N69), .A2(N68), .A3(n85), .Z(n83) );
  XOR3D1 U84 ( .A1(N67), .A2(n86), .A3(n87), .Z(n85) );
  BUFFD1 U85 ( .I(n137), .Z(n141) );
  XOR3D1 U86 ( .A1(N62), .A2(N61), .A3(n88), .Z(n87) );
  XOR3D1 U87 ( .A1(n89), .A2(N60), .A3(n90), .Z(n88) );
  XOR3D1 U88 ( .A1(N81), .A2(N76), .A3(n79), .Z(N85) );
  XOR3D1 U89 ( .A1(N75), .A2(n80), .A3(n81), .Z(n79) );
  XOR3D1 U90 ( .A1(N79), .A2(N78), .A3(n82), .Z(n81) );
  BUFFD1 U91 ( .I(n191), .Z(n138) );
  BUFFD1 U92 ( .I(n191), .Z(n139) );
  INVD1 U93 ( .I(n130), .ZN(n131) );
  INVD1 U94 ( .I(n130), .ZN(n132) );
  INVD1 U95 ( .I(AddrW[0]), .ZN(n93) );
  INVD1 U96 ( .I(n170), .ZN(n173) );
  INVD1 U97 ( .I(n166), .ZN(n169) );
  INVD1 U98 ( .I(n154), .ZN(n157) );
  INVD1 U99 ( .I(n150), .ZN(n153) );
  INVD1 U100 ( .I(N194), .ZN(n163) );
  NR3D0 U101 ( .A1(n91), .A2(AddrW[0]), .A3(n66), .ZN(N194) );
  INVD1 U102 ( .I(N227), .ZN(n159) );
  NR3D0 U103 ( .A1(n91), .A2(n66), .A3(n93), .ZN(N227) );
  NR3D0 U104 ( .A1(n91), .A2(AddrW[0]), .A3(n92), .ZN(N326) );
  INVD1 U105 ( .I(N359), .ZN(n143) );
  NR3D0 U106 ( .A1(n91), .A2(n92), .A3(n93), .ZN(N359) );
  INVD1 U107 ( .I(n190), .ZN(n189) );
  BUFFD1 U108 ( .I(n175), .Z(n174) );
  BUFFD1 U109 ( .I(ClockW), .Z(n175) );
  MUX4ND0 U110 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n141), .S1(n135), .ZN(n8)
         );
  MUX4ND0 U111 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n141), .S1(n135), .ZN(n11)
         );
  MUX4ND0 U112 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n141), .S1(n133), .ZN(n26)
         );
  MUX4ND0 U113 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n191), .S1(n133), .ZN(
        n41) );
  MUX4ND0 U114 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n141), .S1(n133), .ZN(
        n44) );
  MUX4ND0 U115 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n139), .S1(N49), .ZN(n62) );
  MUX4ND0 U116 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n141), .S1(N49), .ZN(n65) );
  MUX4ND0 U117 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n139), .S1(n136), .ZN(
        n111) );
  MUX4ND0 U118 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n141), .S1(N49), .ZN(
        n114) );
  MUX4ND0 U119 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n141), .S1(n134), .ZN(
        n123) );
  MUX4ND0 U120 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n141), .S1(N49), .ZN(
        n126) );
  MUX4ND0 U121 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n138), .S1(n133), .ZN(n23)
         );
  MUX4ND0 U122 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(N48), .S1(n133), .ZN(n29)
         );
  MUX4ND0 U123 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n191), .S1(n133), .ZN(
        n53) );
  MUX4ND0 U124 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n139), .S1(N49), .ZN(
        n102) );
  MUX4ND0 U125 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n141), .S1(N49), .ZN(
        n105) );
  MUX4ND0 U126 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n141), .S1(n135), .ZN(n5)
         );
  MUX4ND0 U127 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n137), .S1(n135), .ZN(n17)
         );
  MUX4ND0 U128 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n137), .S1(n133), .ZN(
        n35) );
  MUX4ND0 U129 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n137), .S1(n133), .ZN(
        n38) );
  MUX4ND0 U130 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n191), .S1(n133), .ZN(
        n47) );
  MUX4ND0 U131 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n139), .S1(n133), .ZN(
        n59) );
  MUX4ND0 U132 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n139), .S1(N49), .ZN(n96) );
  MUX4ND0 U133 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n139), .S1(n136), .ZN(
        n108) );
  MUX4ND0 U134 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n141), .S1(N49), .ZN(
        n117) );
  MUX4ND0 U135 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n141), .S1(N49), .ZN(
        n120) );
  MUX4ND0 U136 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n141), .S1(n135), .ZN(n14)
         );
  MUX4ND0 U137 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n137), .S1(n135), .ZN(n20)
         );
  MUX4ND0 U138 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n137), .S1(n133), .ZN(n32)
         );
  MUX4ND0 U139 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n191), .S1(n133), .ZN(
        n50) );
  MUX4ND0 U140 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n139), .S1(n133), .ZN(
        n56) );
  MUX4ND0 U141 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(N48), .S1(N49), .ZN(n99)
         );
  MUX4ND0 U142 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n141), .S1(n133), .ZN(
        n129) );
  INVD1 U143 ( .I(n171), .ZN(n170) );
  NR3D0 U144 ( .A1(n66), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N99) );
  INVD1 U145 ( .I(AddrW[1]), .ZN(n91) );
  ND2D1 U146 ( .A1(AddrW[2]), .A2(Write), .ZN(n92) );
  IND2D1 U147 ( .A1(AddrW[2]), .B1(Write), .ZN(n66) );
  INVD1 U148 ( .I(N260), .ZN(n155) );
  NR3D0 U149 ( .A1(n92), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N260) );
  NR3D0 U150 ( .A1(n93), .A2(AddrW[1]), .A3(n66), .ZN(N161) );
  INVD1 U151 ( .I(N293), .ZN(n151) );
  NR3D0 U152 ( .A1(n93), .A2(AddrW[1]), .A3(n92), .ZN(N293) );
  INVD1 U153 ( .I(Read), .ZN(n190) );
  OR2D1 U154 ( .A1(Read), .A2(Dreadyr), .Z(n2) );
  CKAN2D0 U155 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX3ND0 U156 ( .I0(n3), .I1(n4), .I2(n5), .S0(n135), .S1(n131), .ZN(N84) );
  MUX3ND0 U157 ( .I0(n6), .I1(n7), .I2(n8), .S0(n135), .S1(n131), .ZN(N83) );
  MUX3ND0 U158 ( .I0(n9), .I1(n10), .I2(n11), .S0(n135), .S1(n131), .ZN(N82)
         );
  MUX3ND0 U159 ( .I0(n12), .I1(n13), .I2(n14), .S0(n135), .S1(n131), .ZN(N81)
         );
  MUX3ND0 U160 ( .I0(n15), .I1(n16), .I2(n17), .S0(n135), .S1(n131), .ZN(N80)
         );
  MUX3ND0 U161 ( .I0(n18), .I1(n19), .I2(n20), .S0(n135), .S1(n131), .ZN(N79)
         );
  MUX3ND0 U162 ( .I0(n21), .I1(n22), .I2(n23), .S0(n135), .S1(n131), .ZN(N78)
         );
  MUX3ND0 U163 ( .I0(n24), .I1(n25), .I2(n26), .S0(n135), .S1(n131), .ZN(N77)
         );
  MUX3ND0 U164 ( .I0(n27), .I1(n28), .I2(n29), .S0(n135), .S1(n131), .ZN(N76)
         );
  MUX3ND0 U165 ( .I0(n30), .I1(n31), .I2(n32), .S0(n135), .S1(n131), .ZN(N75)
         );
  MUX3ND0 U166 ( .I0(n33), .I1(n34), .I2(n35), .S0(n135), .S1(n131), .ZN(N74)
         );
  MUX3ND0 U167 ( .I0(n36), .I1(n37), .I2(n38), .S0(n135), .S1(n131), .ZN(N73)
         );
  MUX3ND0 U168 ( .I0(n39), .I1(n40), .I2(n41), .S0(n135), .S1(n131), .ZN(N72)
         );
  MUX3ND0 U169 ( .I0(n42), .I1(n43), .I2(n44), .S0(n134), .S1(n131), .ZN(N71)
         );
  MUX3ND0 U170 ( .I0(n45), .I1(n46), .I2(n47), .S0(n134), .S1(n131), .ZN(N70)
         );
  MUX3ND0 U171 ( .I0(n48), .I1(n49), .I2(n50), .S0(n134), .S1(n131), .ZN(N69)
         );
  MUX3ND0 U172 ( .I0(n51), .I1(n52), .I2(n53), .S0(n134), .S1(n131), .ZN(N68)
         );
  MUX3ND0 U173 ( .I0(n54), .I1(n55), .I2(n56), .S0(n134), .S1(n131), .ZN(N67)
         );
  MUX3ND0 U174 ( .I0(n57), .I1(n58), .I2(n59), .S0(n134), .S1(n131), .ZN(N66)
         );
  MUX3ND0 U175 ( .I0(n60), .I1(n61), .I2(n62), .S0(n134), .S1(n131), .ZN(N65)
         );
  MUX3ND0 U176 ( .I0(n63), .I1(n64), .I2(n65), .S0(n134), .S1(n132), .ZN(N64)
         );
  MUX3ND0 U177 ( .I0(n94), .I1(n95), .I2(n96), .S0(n134), .S1(n132), .ZN(N63)
         );
  MUX3ND0 U178 ( .I0(n97), .I1(n98), .I2(n99), .S0(n134), .S1(n132), .ZN(N62)
         );
  MUX3ND0 U179 ( .I0(n100), .I1(n101), .I2(n102), .S0(n134), .S1(n132), .ZN(
        N61) );
  MUX3ND0 U180 ( .I0(n103), .I1(n104), .I2(n105), .S0(n134), .S1(n132), .ZN(
        N60) );
  MUX3ND0 U181 ( .I0(n106), .I1(n107), .I2(n108), .S0(n134), .S1(n132), .ZN(
        N59) );
  MUX3ND0 U182 ( .I0(n109), .I1(n110), .I2(n111), .S0(n134), .S1(n132), .ZN(
        N58) );
  MUX3ND0 U183 ( .I0(n112), .I1(n113), .I2(n114), .S0(n134), .S1(n132), .ZN(
        N57) );
  MUX3ND0 U184 ( .I0(n115), .I1(n116), .I2(n117), .S0(n134), .S1(n132), .ZN(
        N56) );
  MUX3ND0 U185 ( .I0(n118), .I1(n119), .I2(n120), .S0(n136), .S1(n132), .ZN(
        N55) );
  MUX3ND0 U186 ( .I0(n121), .I1(n122), .I2(n123), .S0(n133), .S1(n132), .ZN(
        N54) );
  MUX3ND0 U187 ( .I0(n124), .I1(n125), .I2(n126), .S0(N49), .S1(n132), .ZN(N53) );
  MUX3ND0 U188 ( .I0(n127), .I1(n128), .I2(n129), .S0(n134), .S1(n132), .ZN(
        N52) );
  MUX2ND0 U189 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n140), .ZN(n4)
         );
  MUX2ND0 U190 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n140), .ZN(n3)
         );
  MUX2ND0 U191 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(N48), .ZN(n7)
         );
  MUX2ND0 U192 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n140), .ZN(n6)
         );
  MUX2ND0 U193 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n137), .ZN(n10) );
  MUX2ND0 U194 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n140), .ZN(n9)
         );
  MUX2ND0 U195 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n141), .ZN(n13) );
  MUX2ND0 U196 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n141), .ZN(n12) );
  MUX2ND0 U197 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n140), .ZN(n16) );
  MUX2ND0 U198 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n138), .ZN(n15) );
  MUX2ND0 U199 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n140), .ZN(n19) );
  MUX2ND0 U200 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n140), .ZN(n18) );
  MUX2ND0 U201 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n137), .ZN(n22) );
  MUX2ND0 U202 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n140), .ZN(n21) );
  MUX2ND0 U203 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n140), .ZN(n25) );
  MUX2ND0 U204 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n140), .ZN(n24) );
  MUX2ND0 U205 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n140), .ZN(n28) );
  MUX2ND0 U206 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n140), .ZN(n27) );
  MUX2ND0 U207 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n140), .ZN(n31) );
  MUX2ND0 U208 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n140), .ZN(n30) );
  MUX2ND0 U209 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n140), .ZN(
        n34) );
  MUX2ND0 U210 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n140), .ZN(
        n33) );
  MUX2ND0 U211 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n140), .ZN(
        n37) );
  MUX2ND0 U212 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n140), .ZN(
        n36) );
  MUX2ND0 U213 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n140), .ZN(
        n40) );
  MUX2ND0 U214 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n138), .ZN(
        n39) );
  MUX2ND0 U215 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(N48), .ZN(
        n43) );
  MUX2ND0 U216 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n138), .ZN(
        n42) );
  MUX2ND0 U217 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(N48), .ZN(
        n46) );
  MUX2ND0 U218 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n138), .ZN(
        n45) );
  MUX2ND0 U219 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(N48), .ZN(
        n49) );
  MUX2ND0 U220 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(N48), .ZN(
        n48) );
  MUX2ND0 U221 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(N48), .ZN(
        n52) );
  MUX2ND0 U222 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(N48), .ZN(
        n51) );
  MUX2ND0 U223 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n138), .ZN(
        n55) );
  MUX2ND0 U224 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n139), .ZN(
        n54) );
  MUX2ND0 U225 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n138), .ZN(
        n58) );
  MUX2ND0 U226 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n139), .ZN(
        n57) );
  MUX2ND0 U227 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(n139), .ZN(
        n61) );
  MUX2ND0 U228 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n139), .ZN(
        n60) );
  MUX2ND0 U229 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n139), .ZN(
        n64) );
  MUX2ND0 U230 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(n139), .ZN(
        n63) );
  MUX2ND0 U231 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(n139), .ZN(
        n95) );
  MUX2ND0 U232 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(n191), .ZN(
        n94) );
  MUX2ND0 U233 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(N48), .ZN(
        n98) );
  MUX2ND0 U234 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(N48), .ZN(
        n97) );
  MUX2ND0 U235 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(N48), .ZN(
        n101) );
  MUX2ND0 U236 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(N48), .ZN(
        n100) );
  MUX2ND0 U237 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n191), .ZN(
        n104) );
  MUX2ND0 U238 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n191), .ZN(
        n103) );
  MUX2ND0 U239 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n139), .ZN(
        n107) );
  MUX2ND0 U240 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n139), .ZN(
        n106) );
  MUX2ND0 U241 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n139), .ZN(
        n110) );
  MUX2ND0 U242 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n139), .ZN(
        n109) );
  MUX2ND0 U243 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n137), .ZN(
        n113) );
  MUX2ND0 U244 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n137), .ZN(
        n112) );
  MUX2ND0 U245 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n139), .ZN(
        n116) );
  MUX2ND0 U246 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n137), .ZN(
        n115) );
  MUX2ND0 U247 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n191), .ZN(
        n119) );
  MUX2ND0 U248 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n138), .ZN(
        n118) );
  MUX2ND0 U249 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(n138), .ZN(
        n122) );
  MUX2ND0 U250 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n138), .ZN(
        n121) );
  MUX2ND0 U251 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(n191), .ZN(
        n125) );
  MUX2ND0 U252 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n138), .ZN(
        n124) );
  MUX2ND0 U253 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n140), .ZN(
        n128) );
  MUX2ND0 U254 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n139), .ZN(
        n127) );
endmodule


module PLLTop_0 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_0 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_0 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_0 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N47, N48, N49, N50, N51, N67, N68, N69,
         N70, N71, n35, n36, n37, n38, n40, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n83, n84, n85, n86, n87, n90, n92, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n141, n143, n144, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n1, n2, n13, n14;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n151), .CPN(StateClock), .Q(FullFIFO) );
  DFND1 EmptyFIFOr_reg ( .D(n147), .CPN(StateClock), .Q(EmptyFIFO), .QN(n132)
         );
  MOAI22D1 U6 ( .A1(n165), .A2(n40), .B1(n40), .B2(OldReadAr[1]), .ZN(n149) );
  OA21D1 U11 ( .A1(n172), .A2(n170), .B(n35), .Z(n44) );
  MOAI22D1 U12 ( .A1(n168), .A2(n45), .B1(n45), .B2(OldWriteAr[2]), .ZN(n152)
         );
  MOAI22D1 U13 ( .A1(n169), .A2(n45), .B1(n45), .B2(OldWriteAr[0]), .ZN(n153)
         );
  MOAI22D1 U14 ( .A1(n45), .A2(n46), .B1(n45), .B2(OldWriteAr[1]), .ZN(n154)
         );
  MOAI22D1 U15 ( .A1(n167), .A2(n45), .B1(n45), .B2(OldWriteAr[3]), .ZN(n155)
         );
  IAO21D1 U31 ( .A1(n73), .A2(n74), .B(n55), .ZN(n72) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n76), .B(n75), .Z(n81) );
  MOAI22D1 U88 ( .A1(n166), .A2(n40), .B1(n40), .B2(OldReadAr[0]), .ZN(n162)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n150), .CPN(StateClock), .CDN(n13), .QN(n2)
         );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n148), .CPN(StateClock), .CDN(n14), .QN(n1)
         );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n162), .CPN(StateClock), .CDN(n13), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n155), .CPN(StateClock), .CDN(n13), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n154), .CPN(StateClock), .CDN(n14), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n153), .CPN(StateClock), .CDN(n14), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n152), .CPN(StateClock), .CDN(n13), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n149), .CPN(StateClock), .CDN(n14), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n159), .CPN(StateClock), .CDN(n13), .Q(
        NextState[0]), .QN(n144) );
  DFNCND1 \NextState_reg[1]  ( .D(n158), .CPN(StateClock), .CDN(n13), .Q(
        NextState[1]), .QN(n143) );
  DFNCND1 \NextState_reg[2]  ( .D(n156), .CPN(StateClock), .CDN(n13), .Q(
        NextState[2]), .QN(n141) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n13), 
        .QN(n170) );
  DFNCND1 WriteCmdr_reg ( .D(n157), .CPN(StateClock), .CDN(n13), .Q(WriteCmd)
         );
  DFNCND1 ReadCmdr_reg ( .D(n160), .CPN(StateClock), .CDN(n13), .Q(ReadCmd) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n13), 
        .QN(n171) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n13), .Q(
        n52), .QN(n172) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N68), .E(N71), .CP(StateClock), .CDN(n14), .Q(
        WriteAddr[1]), .QN(n46) );
  EDFCND1 \ReadAr_reg[3]  ( .D(N51), .E(N50), .CP(StateClock), .CDN(n14), .Q(
        ReadAddr[3]), .QN(n163) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N50), .CP(StateClock), .CDN(n14), .Q(
        ReadAddr[2]), .QN(n164) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N48), .E(N50), .CP(StateClock), .CDN(n14), .Q(
        ReadAddr[1]), .QN(n165) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N47), .E(N50), .CP(StateClock), .CDN(n14), .Q(
        ReadAddr[0]), .QN(n166) );
  EDFCND1 \WriteAr_reg[3]  ( .D(N70), .E(N71), .CP(StateClock), .CDN(n14), .Q(
        WriteAddr[3]), .QN(n167) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N69), .E(N71), .CP(StateClock), .CDN(n14), .Q(
        WriteAddr[2]), .QN(n168) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N67), .E(N71), .CP(StateClock), .CDN(n14), .Q(
        WriteAddr[0]), .QN(n169) );
  CKNXD0 U3 ( .I(Reset), .ZN(n14) );
  CKNXD0 U4 ( .I(Reset), .ZN(n13) );
  INVD1 U5 ( .I(n48), .ZN(n49) );
  ND2D1 U7 ( .A1(n66), .A2(n42), .ZN(n119) );
  OAI211D1 U8 ( .A1(n35), .A2(n63), .B(n66), .C(n115), .ZN(n48) );
  INR2D1 U9 ( .A1(n71), .B1(n116), .ZN(n115) );
  AOI21D1 U10 ( .A1(n52), .A2(n117), .B(n170), .ZN(n116) );
  MAOI22D0 U16 ( .A1(n69), .A2(n170), .B1(n170), .B2(n71), .ZN(n66) );
  ND2D1 U17 ( .A1(n66), .A2(n35), .ZN(n47) );
  INVD1 U18 ( .I(n106), .ZN(n76) );
  OA211D0 U19 ( .A1(n75), .A2(n76), .B(n77), .C(n78), .Z(n55) );
  INVD1 U20 ( .I(n85), .ZN(n77) );
  NR3D0 U21 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n78) );
  NR3D0 U22 ( .A1(WriteAddr[2]), .A2(n46), .A3(ReadAddr[2]), .ZN(n80) );
  ND2D1 U23 ( .A1(n130), .A2(ReadAddr[2]), .ZN(n129) );
  INVD1 U24 ( .I(n40), .ZN(n38) );
  ND2D1 U25 ( .A1(n107), .A2(n108), .ZN(n85) );
  XNR2D1 U26 ( .A1(ReadAddr[1]), .A2(n46), .ZN(n107) );
  INVD1 U27 ( .I(n90), .ZN(n84) );
  INVD1 U28 ( .I(n97), .ZN(n108) );
  INVD1 U29 ( .I(n53), .ZN(n42) );
  OAI21D1 U30 ( .A1(n130), .A2(ReadAddr[2]), .B(n129), .ZN(n114) );
  ND3D1 U32 ( .A1(n42), .A2(n35), .A3(n56), .ZN(N71) );
  AOI21D1 U33 ( .A1(n76), .A2(n83), .B(ReadAddr[1]), .ZN(n105) );
  ND2D1 U35 ( .A1(n35), .A2(n118), .ZN(N50) );
  NR3D0 U36 ( .A1(n117), .A2(n124), .A3(n125), .ZN(n123) );
  XNR2D1 U37 ( .A1(ReadAddr[3]), .A2(n2), .ZN(n125) );
  XNR2D1 U38 ( .A1(ReadAddr[2]), .A2(n1), .ZN(n124) );
  XNR2D1 U39 ( .A1(n126), .A2(WriteAddr[3]), .ZN(n99) );
  XNR2D1 U40 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n104) );
  NR2D1 U41 ( .A1(n114), .A2(n118), .ZN(N49) );
  NR2D1 U42 ( .A1(n131), .A2(n118), .ZN(N48) );
  XNR2D1 U43 ( .A1(ReadAddr[1]), .A2(ReadAddr[0]), .ZN(n131) );
  NR2D1 U44 ( .A1(n112), .A2(n118), .ZN(N51) );
  NR2D1 U45 ( .A1(ReadAddr[0]), .A2(n118), .ZN(N47) );
  ND2D1 U46 ( .A1(WriteReq), .A2(n47), .ZN(n45) );
  OAI32D1 U47 ( .A1(n35), .A2(WriteReq), .A3(Reset), .B1(n36), .B2(n132), .ZN(
        n147) );
  AOI21D1 U48 ( .A1(n37), .A2(n35), .B(Reset), .ZN(n36) );
  OAI22D0 U49 ( .A1(n48), .A2(n141), .B1(n49), .B2(n50), .ZN(n156) );
  AOI21D1 U50 ( .A1(n51), .A2(n52), .B(n53), .ZN(n50) );
  OAI22D0 U51 ( .A1(n171), .A2(n54), .B1(n170), .B2(n55), .ZN(n51) );
  OAI22D0 U52 ( .A1(n48), .A2(n143), .B1(n49), .B2(n67), .ZN(n158) );
  AOI31D0 U53 ( .A1(n68), .A2(n69), .A3(n170), .B(n70), .ZN(n67) );
  IOA21D1 U54 ( .A1(n52), .A2(n54), .B(n86), .ZN(n68) );
  OAI31D0 U55 ( .A1(n71), .A2(n170), .A3(n72), .B(n35), .ZN(n70) );
  OAI22D0 U56 ( .A1(n48), .A2(n144), .B1(n49), .B2(n100), .ZN(n159) );
  AOI22D0 U57 ( .A1(n101), .A2(n52), .B1(n102), .B2(n103), .ZN(n100) );
  AOI211D1 U58 ( .A1(n164), .A2(n106), .B(n37), .C(n85), .ZN(n102) );
  AOI221D0 U59 ( .A1(n90), .A2(n76), .B1(n104), .B2(ReadAddr[1]), .C(n105), 
        .ZN(n103) );
  NR3D0 U60 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n60) );
  XNR2D1 U61 ( .A1(n167), .A2(OldWriteAr[3]), .ZN(n62) );
  XNR2D1 U62 ( .A1(n46), .A2(OldWriteAr[1]), .ZN(n61) );
  OAI21D1 U63 ( .A1(n56), .A2(n47), .B(n57), .ZN(n157) );
  ND4D1 U64 ( .A1(n58), .A2(n47), .A3(n59), .A4(n60), .ZN(n57) );
  XNR2D1 U65 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n58) );
  XNR2D1 U66 ( .A1(WriteAddr[2]), .A2(OldWriteAr[2]), .ZN(n59) );
  INVD1 U67 ( .I(WriteReq), .ZN(n63) );
  CKND2D0 U68 ( .A1(ReadReq), .A2(n119), .ZN(n40) );
  ND2D1 U69 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n128) );
  AOI21D1 U70 ( .A1(n128), .A2(n168), .B(n126), .ZN(n98) );
  ND2D1 U71 ( .A1(n171), .A2(n52), .ZN(n71) );
  OAI22D0 U72 ( .A1(n38), .A2(n1), .B1(n164), .B2(n40), .ZN(n148) );
  OAI22D0 U73 ( .A1(n38), .A2(n2), .B1(n163), .B2(n40), .ZN(n150) );
  AOI21D1 U74 ( .A1(n83), .A2(n84), .B(WriteAddr[1]), .ZN(n79) );
  NR2D1 U75 ( .A1(WriteAddr[2]), .A2(n164), .ZN(n90) );
  OAI21D1 U76 ( .A1(n171), .A2(n109), .B(n170), .ZN(n101) );
  NR4D0 U77 ( .A1(n108), .A2(n110), .A3(n95), .A4(n111), .ZN(n109) );
  XNR2D1 U78 ( .A1(WriteAddr[2]), .A2(n114), .ZN(n110) );
  XNR2D1 U79 ( .A1(WriteAddr[3]), .A2(n112), .ZN(n111) );
  ND4D1 U80 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n54) );
  XNR2D1 U81 ( .A1(n99), .A2(n163), .ZN(n94) );
  XNR2D1 U82 ( .A1(ReadAddr[2]), .A2(n98), .ZN(n96) );
  NR2D1 U83 ( .A1(n128), .A2(n168), .ZN(n126) );
  NR2D1 U84 ( .A1(n46), .A2(n168), .ZN(n75) );
  XNR2D1 U85 ( .A1(ReadAddr[3]), .A2(n167), .ZN(n106) );
  XNR2D1 U86 ( .A1(WriteAddr[0]), .A2(n166), .ZN(n97) );
  XNR2D1 U87 ( .A1(n163), .A2(n129), .ZN(n112) );
  ND2D1 U89 ( .A1(ReadCmd), .A2(n35), .ZN(n118) );
  ND2D1 U90 ( .A1(WriteCmd), .A2(n42), .ZN(n56) );
  OAI211D1 U91 ( .A1(n46), .A2(ReadAddr[1]), .B(n83), .C(n92), .ZN(n74) );
  AOI22D0 U92 ( .A1(n163), .A2(WriteAddr[3]), .B1(n166), .B2(WriteAddr[0]), 
        .ZN(n92) );
  OAI21D1 U93 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n128), .ZN(n113) );
  ND3D1 U94 ( .A1(n171), .A2(n170), .A3(n172), .ZN(n35) );
  OAI211D1 U95 ( .A1(n165), .A2(WriteAddr[1]), .B(n84), .C(n87), .ZN(n73) );
  AOI22D0 U96 ( .A1(n167), .A2(ReadAddr[3]), .B1(n169), .B2(ReadAddr[0]), .ZN(
        n87) );
  OAI22D0 U97 ( .A1(n165), .A2(n42), .B1(n113), .B2(n56), .ZN(N68) );
  OAI22D0 U98 ( .A1(n163), .A2(n42), .B1(n99), .B2(n56), .ZN(N70) );
  OAI22D0 U99 ( .A1(n164), .A2(n42), .B1(n127), .B2(n56), .ZN(N69) );
  INVD1 U100 ( .I(n98), .ZN(n127) );
  OAI22D0 U101 ( .A1(n166), .A2(n42), .B1(WriteAddr[0]), .B2(n56), .ZN(N67) );
  NR3D0 U102 ( .A1(n171), .A2(n172), .A3(n170), .ZN(n53) );
  ND2D1 U103 ( .A1(n164), .A2(WriteAddr[2]), .ZN(n83) );
  INVD1 U104 ( .I(n171), .ZN(n69) );
  ND3D1 U105 ( .A1(n170), .A2(n69), .A3(n172), .ZN(n37) );
  OAI21D1 U106 ( .A1(n118), .A2(n119), .B(n120), .ZN(n160) );
  ND4D1 U107 ( .A1(n121), .A2(n119), .A3(n122), .A4(n123), .ZN(n120) );
  XNR2D1 U108 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n121) );
  XNR2D1 U109 ( .A1(ReadAddr[1]), .A2(OldReadAr[1]), .ZN(n122) );
  OAI21D1 U110 ( .A1(n74), .A2(n73), .B(n172), .ZN(n86) );
  NR2D1 U111 ( .A1(n166), .A2(n165), .ZN(n130) );
  XNR2D1 U112 ( .A1(n113), .A2(n165), .ZN(n95) );
  OAI31D0 U113 ( .A1(n42), .A2(Reset), .A3(ReadReq), .B(n43), .ZN(n151) );
  OAI21D1 U114 ( .A1(n44), .A2(Reset), .B(FullFIFO), .ZN(n43) );
  ND2D1 U115 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U116 ( .I(ReadReq), .ZN(n117) );
endmodule


module DPMem1kx32_AWid4_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, N133, N166, N199, N232, N265, N298, N331, N364, N397,
         N430, N463, N496, N529, N562, N595, N628, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n103, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n102,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  OR2D1 U3 ( .A1(Read), .A2(Dreadyr), .Z(n103) );
  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n76) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n75) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n72) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n69) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n66) );
  XOR4D1 U21 ( .A1(n81), .A2(N71), .A3(n82), .A4(N74), .Z(n80) );
  XNR4D1 U22 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n82) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n88) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n87) );
  XNR4D1 U29 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .ZN(n84) );
  XNR4D1 U30 ( .A1(N79), .A2(N77), .A3(N81), .A4(N80), .ZN(n78) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N84), .E(N595), .CP(n257), .CDN(n298), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(N595), .CP(n257), .CDN(
        n297), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(N595), .CP(n257), .CDN(
        n297), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(N595), .CP(n258), .CDN(
        n297), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(n194), .CP(n258), .CDN(
        n297), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(n194), .CP(n259), .CDN(
        n296), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(n192), .CP(n259), .CDN(
        n296), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(N595), .CP(n259), .CDN(
        n296), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(n194), .CP(n259), .CDN(
        n296), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(n194), .CP(n260), .CDN(
        n296), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(n194), .CP(n260), .CDN(
        n296), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(n194), .CP(n260), .CDN(n295), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(n192), .CP(n261), .CDN(n295), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(n192), .CP(n261), .CDN(n295), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(n192), .CP(n261), .CDN(n295), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N84), .E(N562), .CP(n261), .CDN(n295), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(n198), .CP(n261), .CDN(
        n294), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(n198), .CP(n261), .CDN(
        n294), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(n198), .CP(n261), .CDN(
        n294), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(n198), .CP(n262), .CDN(
        n294), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(n198), .CP(n262), .CDN(
        n294), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(N562), .CP(n262), .CDN(
        n294), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(N562), .CP(n262), .CDN(
        n294), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(n196), .CP(n262), .CDN(
        n293), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(n196), .CP(n262), .CDN(
        n293), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(n196), .CP(n262), .CDN(
        n293), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(n198), .CP(n263), .CDN(
        n293), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(n196), .CP(n263), .CDN(
        n293), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(N562), .CP(n263), .CDN(n292), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(DataI[6]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(N562), .CP(n264), .CDN(n292), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(n198), .CP(n264), .CDN(n292), .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(n198), .CP(n264), .CDN(n292), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(n198), .CP(n264), .CDN(n292), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N84), .E(N463), .CP(n254), .CDN(n288), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(n210), .CP(n254), .CDN(
        n287), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(n210), .CP(n257), .CDN(
        n287), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(n210), .CP(n258), .CDN(
        n287), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(n210), .CP(n268), .CDN(
        n287), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(n210), .CP(n267), .CDN(
        n287), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(N463), .CP(n265), .CDN(
        n287), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(N463), .CP(n266), .CDN(
        n287), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(n208), .CP(n273), .CDN(
        n314), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(n208), .CP(n270), .CDN(
        n288), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(n208), .CP(n269), .CDN(
        n290), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(n208), .CP(n261), .CDN(
        n315), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(n208), .CP(n262), .CDN(
        n291), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(DataI[15]), .E(n208), .CP(n260), .CDN(
        n289), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(DataI[14]), .E(n208), .CP(n259), .CDN(
        n311), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(DataI[13]), .E(n208), .CP(n264), .CDN(
        n293), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(n210), .CP(n263), .CDN(
        n288), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(n208), .CP(n265), .CDN(
        n288), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(n208), .CP(n266), .CDN(
        n288), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(N463), .CP(n270), .CDN(n315), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(N463), .CP(n262), .CDN(n314), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(DataI[7]), .E(N463), .CP(n265), .CDN(n291), .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(DataI[6]), .E(N463), .CP(n268), .CDN(n287), .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(DataI[5]), .E(N463), .CP(n277), .CDN(n287), .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(N463), .CP(n278), .CDN(n287), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(N463), .CP(n255), .CDN(n287), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(n210), .CP(n259), .CDN(n287), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(n210), .CP(n253), .CDN(n287), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(n210), .CP(n252), .CDN(n287), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N84), .E(n212), .CP(n268), .CDN(n288), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(n214), .CP(n273), .CDN(
        n310), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(N430), .CP(n270), .CDN(
        n314), .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(N430), .CP(n269), .CDN(
        n305), .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(N430), .CP(n264), .CDN(
        n292), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(N430), .CP(n275), .CDN(
        n308), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(n214), .CP(n259), .CDN(
        n309), .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(n214), .CP(n252), .CDN(
        n290), .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(n214), .CP(n275), .CDN(
        n315), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(n214), .CP(n274), .CDN(
        n289), .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(n214), .CP(n273), .CDN(
        n294), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(n214), .CP(n272), .CDN(
        n289), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(n214), .CP(n271), .CDN(
        n290), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(DataI[15]), .E(n214), .CP(n256), .CDN(
        n292), .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(n214), .CP(n260), .CDN(
        n291), .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(n214), .CP(n252), .CDN(
        n293), .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(n212), .CP(n276), .CDN(
        n294), .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(n212), .CP(n254), .CDN(
        n289), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(N430), .CP(n256), .CDN(
        n290), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(N430), .CP(n255), .CDN(n307), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(N430), .CP(n258), .CDN(n310), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(DataI[7]), .E(n212), .CP(n257), .CDN(n316), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(n212), .CP(n263), .CDN(n305), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(n212), .CP(n257), .CDN(n307), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(n212), .CP(n260), .CDN(n306), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(n212), .CP(n262), .CDN(n305), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(n212), .CP(n261), .CDN(n308), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(n212), .CP(n264), .CDN(n308), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(n214), .CP(n263), .CDN(n291), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N84), .E(N331), .CP(n270), .CDN(n309), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n226), .CP(n271), .CDN(
        n305), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n226), .CP(n275), .CDN(
        n292), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n226), .CP(n253), .CDN(
        n312), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n226), .CP(ClockW), .CDN(
        n306), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n226), .CP(n274), .CDN(
        n306), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(N331), .CP(n277), .CDN(
        n310), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(N331), .CP(n266), .CDN(
        n307), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n224), .CP(n257), .CDN(
        n307), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n224), .CP(n252), .CDN(
        n301), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n224), .CP(n271), .CDN(
        n295), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n224), .CP(n272), .CDN(
        n312), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n224), .CP(n273), .CDN(
        n289), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n224), .CP(n275), .CDN(
        n309), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n224), .CP(ClockW), .CDN(
        n307), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n224), .CP(n262), .CDN(
        n310), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n226), .CP(n258), .CDN(
        n316), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n224), .CP(n255), .CDN(
        n311), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n224), .CP(n264), .CDN(
        n306), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(N331), .CP(n274), .CDN(n308), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(N331), .CP(n264), .CDN(n316), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(N331), .CP(n263), .CDN(n298), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(N331), .CP(n263), .CDN(n301), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(N331), .CP(n253), .CDN(n312), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(N331), .CP(n256), .CDN(n294), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(N331), .CP(n255), .CDN(n309), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n226), .CP(n258), .CDN(n311), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n226), .CP(n257), .CDN(n305), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n226), .CP(n261), .CDN(n295), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N84), .E(N298), .CP(n277), .CDN(n311), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n230), .CP(n252), .CDN(
        n314), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n230), .CP(n278), .CDN(
        n310), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n230), .CP(n274), .CDN(
        n308), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n230), .CP(n256), .CDN(
        n287), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n230), .CP(n270), .CDN(
        n307), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(N298), .CP(n269), .CDN(
        n306), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(N298), .CP(n267), .CDN(
        n313), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n228), .CP(n273), .CDN(
        n296), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n228), .CP(n278), .CDN(
        n313), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n228), .CP(n261), .CDN(
        n294), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n228), .CP(n271), .CDN(
        n308), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n228), .CP(n266), .CDN(
        n301), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n228), .CP(n257), .CDN(
        n288), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n228), .CP(n267), .CDN(
        n306), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n228), .CP(n259), .CDN(
        n305), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n230), .CP(n269), .CDN(
        n298), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n228), .CP(n265), .CDN(
        n315), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n228), .CP(n274), .CDN(
        n306), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(N298), .CP(n277), .CDN(n300), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(N298), .CP(n263), .CDN(n296), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(N298), .CP(n278), .CDN(n307), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(N298), .CP(n270), .CDN(n291), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(N298), .CP(n253), .CDN(n307), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(N298), .CP(n266), .CDN(n298), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(N298), .CP(n253), .CDN(n299), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n230), .CP(n270), .CDN(n310), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n230), .CP(n278), .CDN(n290), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n230), .CP(n252), .CDN(n295), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N84), .E(N199), .CP(n276), .CDN(n308), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n242), .CP(n253), .CDN(
        n303), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n242), .CP(n273), .CDN(
        n302), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(n242), .CP(n258), .CDN(
        n313), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n242), .CP(ClockW), .CDN(
        n304), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n242), .CP(n271), .CDN(
        n315), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(N199), .CP(n267), .CDN(
        n312), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(N199), .CP(n260), .CDN(
        n304), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n240), .CP(n275), .CDN(
        n303), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n240), .CP(n277), .CDN(
        n302), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n240), .CP(n271), .CDN(
        n304), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n240), .CP(n271), .CDN(
        n314), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n240), .CP(n277), .CDN(
        n303), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n240), .CP(n268), .CDN(
        n314), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n240), .CP(n266), .CDN(
        n302), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n240), .CP(n271), .CDN(
        n304), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n242), .CP(n271), .CDN(
        n306), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n240), .CP(n274), .CDN(
        n303), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n240), .CP(n272), .CDN(
        n302), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(N199), .CP(n274), .CDN(n304), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(N199), .CP(n276), .CDN(n303), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(N199), .CP(n259), .CDN(n302), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(N199), .CP(n266), .CDN(n299), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(N199), .CP(ClockW), .CDN(
        n304), .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(N199), .CP(n261), .CDN(n303), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(N199), .CP(n271), .CDN(n302), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n242), .CP(n253), .CDN(n301), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n242), .CP(n278), .CDN(n304), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n242), .CP(n271), .CDN(n303), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N84), .E(N166), .CP(n267), .CDN(n302), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n246), .CP(n269), .CDN(
        n299), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n246), .CP(n270), .CDN(
        n288), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n246), .CP(n276), .CDN(
        n293), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n246), .CP(n277), .CDN(
        n297), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n246), .CP(n254), .CDN(
        n300), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(N166), .CP(n270), .CDN(
        n300), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(N166), .CP(n275), .CDN(
        n287), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n244), .CP(n277), .CDN(
        n293), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n244), .CP(ClockW), .CDN(
        n312), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n244), .CP(n265), .CDN(
        n316), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n244), .CP(n253), .CDN(
        n314), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n244), .CP(n272), .CDN(
        n300), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n244), .CP(n274), .CDN(
        n310), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n244), .CP(n273), .CDN(
        n293), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n244), .CP(n257), .CDN(
        n316), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n246), .CP(n272), .CDN(
        n312), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n244), .CP(n269), .CDN(
        n305), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n244), .CP(n278), .CDN(
        n311), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(N166), .CP(n252), .CDN(n315), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(N166), .CP(n269), .CDN(n316), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(N166), .CP(n276), .CDN(n307), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(N166), .CP(n252), .CDN(n310), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(N166), .CP(n272), .CDN(n311), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(N166), .CP(n278), .CDN(n309), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(N166), .CP(n260), .CDN(n315), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n246), .CP(n278), .CDN(n314), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n246), .CP(n271), .CDN(n316), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n246), .CP(n268), .CDN(n315), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N84), .E(n188), .CP(n254), .CDN(n301), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(n190), .CP(n254), .CDN(
        n300), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(n188), .CP(n254), .CDN(
        n300), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(N628), .CP(n255), .CDN(
        n300), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(n190), .CP(n255), .CDN(
        n300), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(n190), .CP(n255), .CDN(
        n300), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(n190), .CP(n255), .CDN(
        n299), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(n190), .CP(n256), .CDN(
        n299), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(n190), .CP(n256), .CDN(
        n299), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(n188), .CP(n256), .CDN(
        n299), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(n188), .CP(n256), .CDN(
        n299), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(N628), .CP(n256), .CDN(
        n299), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(N628), .CP(n256), .CDN(n298), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(N628), .CP(n256), .CDN(n298), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(N628), .CP(n256), .CDN(n298), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(n188), .CP(n256), .CDN(n298), .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(n188), .CP(n257), .CDN(n298), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(n188), .CP(n257), .CDN(n298), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(n188), .CP(n257), .CDN(n298), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(n188), .CP(n257), .CDN(n298), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(n188), .CP(n257), .CDN(n298), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(n190), .CP(n257), .CDN(n298), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N84), .E(N529), .CP(n265), .CDN(n292), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(n202), .CP(n266), .CDN(
        n291), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(N529), .CP(n266), .CDN(
        n291), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(n202), .CP(n266), .CDN(
        n291), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(n202), .CP(n266), .CDN(
        n290), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(n200), .CP(n266), .CDN(
        n290), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(N529), .CP(n266), .CDN(
        n290), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(N529), .CP(n266), .CDN(
        n290), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(N529), .CP(n266), .CDN(
        n290), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(DataI[15]), .E(N529), .CP(n266), .CDN(
        n290), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(DataI[14]), .E(N529), .CP(n267), .CDN(
        n290), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(N529), .CP(n267), .CDN(
        n290), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(N529), .CP(n267), .CDN(
        n290), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(n200), .CP(n267), .CDN(
        n290), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(n200), .CP(n267), .CDN(
        n290), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(n200), .CP(n267), .CDN(n289), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(n200), .CP(n267), .CDN(n289), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(DataI[7]), .E(n200), .CP(n267), .CDN(n289), .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(DataI[6]), .E(n200), .CP(n267), .CDN(n289), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(DataI[5]), .E(n200), .CP(n268), .CDN(n289), .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(n200), .CP(n268), .CDN(n289), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(n200), .CP(n268), .CDN(n289), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(n202), .CP(n268), .CDN(n289), .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(n202), .CP(n268), .CDN(n289), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(n202), .CP(n268), .CDN(n289), .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N84), .E(N496), .CP(n268), .CDN(n289), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(n206), .CP(n268), .CDN(
        n315), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(n206), .CP(n268), .CDN(
        n295), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(n206), .CP(n272), .CDN(
        n293), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(n206), .CP(n264), .CDN(
        n298), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(n206), .CP(n265), .CDN(
        n292), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(N496), .CP(n267), .CDN(
        n297), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(N496), .CP(n268), .CDN(
        n294), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(n204), .CP(n254), .CDN(
        n315), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(n204), .CP(n258), .CDN(
        n315), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(n204), .CP(n257), .CDN(
        n315), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(n204), .CP(n256), .CDN(
        n315), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(n204), .CP(n255), .CDN(
        n315), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(DataI[15]), .E(n204), .CP(n259), .CDN(
        n314), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(DataI[14]), .E(n204), .CP(n276), .CDN(
        n314), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(n204), .CP(ClockW), .CDN(
        n306), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(n206), .CP(n253), .CDN(
        n300), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(n204), .CP(n277), .CDN(
        n299), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(n204), .CP(n270), .CDN(
        n293), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(N496), .CP(n277), .CDN(n288), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(N496), .CP(n252), .CDN(n288), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(DataI[7]), .E(N496), .CP(n275), .CDN(n288), .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(DataI[6]), .E(N496), .CP(n274), .CDN(n288), .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(DataI[5]), .E(N496), .CP(n272), .CDN(n288), .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(N496), .CP(n271), .CDN(n288), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(N496), .CP(n252), .CDN(n288), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(n206), .CP(n256), .CDN(n288), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(n206), .CP(n264), .CDN(n288), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(n206), .CP(n263), .CDN(n288), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N84), .E(N397), .CP(n269), .CDN(n298), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(n218), .CP(n259), .CDN(
        n307), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(n218), .CP(n262), .CDN(
        n296), .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(n218), .CP(n264), .CDN(
        n313), .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(n218), .CP(n270), .CDN(
        n311), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(n218), .CP(n269), .CDN(
        n313), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(N397), .CP(n265), .CDN(
        n291), .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(N397), .CP(n273), .CDN(
        n309), .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(n216), .CP(n252), .CDN(
        n313), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(n216), .CP(n253), .CDN(
        n288), .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(n216), .CP(n274), .CDN(
        n306), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(n216), .CP(n268), .CDN(
        n294), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(n216), .CP(n269), .CDN(
        n308), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(DataI[15]), .E(n216), .CP(n274), .CDN(
        n305), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(n216), .CP(n258), .CDN(
        n313), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(n216), .CP(n278), .CDN(
        n308), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(n218), .CP(n255), .CDN(
        n316), .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(n216), .CP(n263), .CDN(
        n310), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(n216), .CP(n257), .CDN(
        n316), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(N397), .CP(n258), .CDN(n295), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(N397), .CP(n255), .CDN(n292), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(DataI[7]), .E(N397), .CP(n256), .CDN(n314), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(N397), .CP(n254), .CDN(n294), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(N397), .CP(n259), .CDN(n308), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(N397), .CP(n260), .CDN(n316), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(N397), .CP(n261), .CDN(n307), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(n218), .CP(n274), .CDN(n305), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(n218), .CP(n275), .CDN(n308), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(n218), .CP(n256), .CDN(n315), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N84), .E(N364), .CP(ClockW), .CDN(n306), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n222), .CP(n276), .CDN(
        n316), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n222), .CP(n255), .CDN(
        n292), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n222), .CP(n256), .CDN(
        n294), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n222), .CP(n261), .CDN(
        n299), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(n222), .CP(n262), .CDN(
        n311), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(N364), .CP(n259), .CDN(
        n298), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(N364), .CP(n260), .CDN(
        n316), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n220), .CP(n263), .CDN(
        n310), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n220), .CP(n269), .CDN(
        n316), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n220), .CP(n254), .CDN(
        n306), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n220), .CP(n264), .CDN(
        n292), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n220), .CP(n278), .CDN(
        n313), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n220), .CP(n278), .CDN(
        n305), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n220), .CP(n258), .CDN(
        n310), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n220), .CP(n256), .CDN(
        n290), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n222), .CP(n277), .CDN(
        n310), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n220), .CP(n253), .CDN(
        n313), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n220), .CP(n253), .CDN(
        n305), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(N364), .CP(n270), .CDN(n314), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(N364), .CP(n276), .CDN(n314), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(N364), .CP(n268), .CDN(n313), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(N364), .CP(n275), .CDN(n307), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(N364), .CP(n274), .CDN(n314), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(N364), .CP(n254), .CDN(n308), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(N364), .CP(n268), .CDN(n308), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n222), .CP(n277), .CDN(n307), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n222), .CP(n276), .CDN(n312), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n222), .CP(n275), .CDN(n306), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N84), .E(N265), .CP(n254), .CDN(n308), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n234), .CP(n269), .CDN(
        n296), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n234), .CP(n267), .CDN(
        n298), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n234), .CP(n260), .CDN(
        n311), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n234), .CP(n260), .CDN(
        n316), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n234), .CP(n265), .CDN(
        n316), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(N265), .CP(n276), .CDN(
        n301), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(N265), .CP(n269), .CDN(
        n294), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n232), .CP(n277), .CDN(
        n312), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n232), .CP(n275), .CDN(
        n293), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n232), .CP(n278), .CDN(
        n305), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n232), .CP(n265), .CDN(
        n313), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n232), .CP(n272), .CDN(
        n312), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n232), .CP(n262), .CDN(
        n312), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n232), .CP(n252), .CDN(
        n301), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n232), .CP(n253), .CDN(
        n301), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n234), .CP(ClockW), .CDN(
        n310), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n232), .CP(n266), .CDN(
        n311), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n232), .CP(n258), .CDN(
        n313), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(N265), .CP(ClockW), .CDN(
        n313), .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(N265), .CP(n276), .CDN(n301), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(N265), .CP(n275), .CDN(n311), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(N265), .CP(n274), .CDN(n296), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(N265), .CP(n253), .CDN(n305), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(N265), .CP(n267), .CDN(n306), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(N265), .CP(n270), .CDN(n309), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n234), .CP(n278), .CDN(n310), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n234), .CP(n257), .CDN(n307), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n234), .CP(n272), .CDN(n307), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N84), .E(N232), .CP(n276), .CDN(n309), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n238), .CP(ClockW), .CDN(
        n306), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n238), .CP(n273), .CDN(
        n297), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n238), .CP(n272), .CDN(
        n288), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n238), .CP(n271), .CDN(
        n297), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(n238), .CP(n253), .CDN(
        n313), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(N232), .CP(n273), .CDN(
        n308), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(N232), .CP(n274), .CDN(
        n307), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n236), .CP(n271), .CDN(
        n304), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n236), .CP(n272), .CDN(
        n311), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n236), .CP(n278), .CDN(
        n302), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n236), .CP(n278), .CDN(
        n304), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n236), .CP(n254), .CDN(
        n289), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n236), .CP(ClockW), .CDN(
        n302), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n236), .CP(n252), .CDN(
        n304), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n236), .CP(n252), .CDN(
        n295), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n238), .CP(n255), .CDN(
        n306), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n236), .CP(n270), .CDN(
        n304), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n236), .CP(n269), .CDN(
        n314), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(N232), .CP(n252), .CDN(n304), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(N232), .CP(n261), .CDN(n303), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(N232), .CP(n262), .CDN(n297), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(N232), .CP(n269), .CDN(n304), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(N232), .CP(n276), .CDN(n304), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(N232), .CP(n268), .CDN(n315), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(N232), .CP(n262), .CDN(n304), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n238), .CP(ClockW), .CDN(
        n304), .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n238), .CP(n273), .CDN(n313), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n238), .CP(n277), .CDN(n304), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N84), .E(N133), .CP(n272), .CDN(n305), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(N133), .CP(n267), .CDN(
        n292), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n248), .CP(ClockW), .CDN(
        n289), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n248), .CP(n253), .CDN(
        n314), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n248), .CP(n252), .CDN(
        n297), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n248), .CP(n271), .CDN(
        n312), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n250), .CP(n252), .CDN(
        n313), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n250), .CP(n273), .CDN(
        n306), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n250), .CP(n270), .CDN(
        n309), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n250), .CP(n269), .CDN(
        n310), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n250), .CP(n273), .CDN(
        n311), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n250), .CP(n259), .CDN(
        n309), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n250), .CP(n263), .CDN(
        n312), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n250), .CP(n254), .CDN(
        n312), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n250), .CP(n267), .CDN(
        n312), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n250), .CP(n258), .CDN(
        n312), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(N133), .CP(n271), .CDN(
        n312), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(N133), .CP(n277), .CDN(
        n310), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(N133), .CP(n272), .CDN(
        n309), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(N133), .CP(n276), .CDN(n293), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(N133), .CP(n272), .CDN(n289), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(N133), .CP(n275), .CDN(n311), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(N133), .CP(n277), .CDN(n309), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n248), .CP(n268), .CDN(n292), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n248), .CP(n273), .CDN(n311), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(N133), .CP(n260), .CDN(n309), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n248), .CP(n265), .CDN(n310), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n248), .CP(n273), .CDN(n311), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n248), .CP(ClockW), .CDN(
        n309), .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n103), .CP(ClockR), .CDN(n290), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(n192), .CP(n258), .CDN(
        n297), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(N595), .CP(n258), .CDN(
        n297), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(n198), .CP(n261), .CDN(
        n294), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(n198), .CP(n261), .CDN(
        n294), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(n196), .CP(n262), .CDN(
        n294), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(N562), .CP(n262), .CDN(
        n294), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(n210), .CP(n261), .CDN(
        n287), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(n210), .CP(n262), .CDN(
        n287), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(n208), .CP(n253), .CDN(
        n287), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(N463), .CP(n276), .CDN(
        n287), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(N430), .CP(n255), .CDN(
        n316), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(N430), .CP(n274), .CDN(
        n311), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(N430), .CP(ClockW), .CDN(
        n296), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(N430), .CP(n276), .CDN(
        n316), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n226), .CP(n277), .CDN(
        n313), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n226), .CP(n276), .CDN(
        n299), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n224), .CP(n255), .CDN(
        n309), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(N331), .CP(n269), .CDN(
        n308), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n230), .CP(n272), .CDN(
        n291), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n230), .CP(n261), .CDN(
        n289), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n228), .CP(n262), .CDN(
        n315), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(N298), .CP(n275), .CDN(
        n305), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n242), .CP(n253), .CDN(
        n303), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n242), .CP(n252), .CDN(
        n297), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n240), .CP(n270), .CDN(
        n304), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(N199), .CP(n276), .CDN(
        n316), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n246), .CP(n264), .CDN(
        n297), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n246), .CP(n263), .CDN(
        n296), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n244), .CP(n275), .CDN(
        n290), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(N166), .CP(n273), .CDN(
        n295), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(N628), .CP(n254), .CDN(
        n300), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(n202), .CP(n265), .CDN(
        n291), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(n200), .CP(n265), .CDN(
        n291), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(N529), .CP(n265), .CDN(
        n291), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(n206), .CP(n261), .CDN(
        n300), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(n206), .CP(n275), .CDN(
        n290), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(n204), .CP(n273), .CDN(
        n299), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(N496), .CP(n278), .CDN(
        n295), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(n218), .CP(n267), .CDN(
        n305), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(n218), .CP(n275), .CDN(
        n315), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(n216), .CP(n274), .CDN(
        n291), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(N397), .CP(n272), .CDN(
        n307), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n222), .CP(n270), .CDN(
        n309), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n222), .CP(n257), .CDN(
        n310), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n220), .CP(n256), .CDN(
        n311), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(N364), .CP(n265), .CDN(
        n309), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n234), .CP(n266), .CDN(
        n305), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n234), .CP(n269), .CDN(
        n300), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n232), .CP(n259), .CDN(
        n309), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(N265), .CP(n266), .CDN(
        n300), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n238), .CP(n270), .CDN(
        n306), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n238), .CP(n253), .CDN(
        n301), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n236), .CP(n260), .CDN(
        n291), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(N232), .CP(n264), .CDN(
        n308), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(n248), .CP(n274), .CDN(
        n307), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n250), .CP(n275), .CDN(
        n308), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N133), .CP(n276), .CDN(
        n298), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n250), .CP(n273), .CDN(
        n299), .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N50), .E(n283), .CP(n279), .CDN(n304), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N51), .E(n281), .CP(ClockR), .CDN(n303), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N52), .E(Read), .CP(n279), .CDN(n303), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N53), .E(n283), .CP(ClockR), .CDN(n303), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N54), .E(Read), .CP(n279), .CDN(n303), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N55), .E(Read), .CP(ClockR), .CDN(n303), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N56), .E(Read), .CP(n279), .CDN(n303), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N57), .E(Read), .CP(n279), .CDN(n303), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N58), .E(Read), .CP(ClockR), .CDN(n303), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N59), .E(Read), .CP(n279), .CDN(n303), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N60), .E(n281), .CP(ClockR), .CDN(n303), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N61), .E(n281), .CP(n279), .CDN(n303), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N62), .E(n281), .CP(ClockR), .CDN(n302), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N63), .E(n281), .CP(n279), .CDN(n302), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N64), .E(n281), .CP(ClockR), .CDN(n302), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N65), .E(n281), .CP(n279), .CDN(n302), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N66), .E(n281), .CP(ClockR), .CDN(n302), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N67), .E(n281), .CP(n279), .CDN(n302), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N68), .E(n281), .CP(n279), .CDN(n302), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N69), .E(n281), .CP(n279), .CDN(n302), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N70), .E(Read), .CP(n279), .CDN(n302), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N71), .E(Read), .CP(n279), .CDN(n302), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N72), .E(Read), .CP(n279), .CDN(n302), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N73), .E(Read), .CP(n279), .CDN(n301), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N74), .E(Read), .CP(n279), .CDN(n301), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N75), .E(Read), .CP(n279), .CDN(n301), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N76), .E(Read), .CP(n279), .CDN(n301), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N77), .E(n283), .CP(ClockR), .CDN(n301), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N78), .E(Read), .CP(ClockR), .CDN(n301), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N79), .E(Read), .CP(ClockR), .CDN(n301), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N80), .E(n283), .CP(ClockR), .CDN(n301), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N81), .E(Read), .CP(ClockR), .CDN(n301), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N82), .E(Read), .CP(ClockR), .CDN(n301), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKBD0 U4 ( .CLK(N45), .C(n176) );
  CKBD0 U5 ( .CLK(N45), .C(n175) );
  CKBD0 U6 ( .CLK(N44), .C(n285) );
  CKNXD0 U7 ( .I(n192), .ZN(n195) );
  CKNXD0 U8 ( .I(n248), .ZN(n251) );
  NR2XD0 U9 ( .A1(n94), .A2(n98), .ZN(N133) );
  INVD0 U10 ( .I(n236), .ZN(n239) );
  INVD0 U11 ( .I(n237), .ZN(n236) );
  CKNXD0 U12 ( .I(n239), .ZN(n238) );
  INVD0 U18 ( .I(n232), .ZN(n235) );
  INVD0 U19 ( .I(n233), .ZN(n232) );
  CKNXD0 U20 ( .I(n235), .ZN(n234) );
  INVD0 U23 ( .I(n220), .ZN(n223) );
  INVD0 U24 ( .I(n221), .ZN(n220) );
  CKNXD0 U25 ( .I(n223), .ZN(n222) );
  INVD0 U26 ( .I(n216), .ZN(n219) );
  INVD0 U31 ( .I(n217), .ZN(n216) );
  CKNXD0 U32 ( .I(n219), .ZN(n218) );
  INVD0 U33 ( .I(n204), .ZN(n207) );
  INVD0 U34 ( .I(n205), .ZN(n204) );
  CKNXD0 U35 ( .I(n207), .ZN(n206) );
  INVD0 U36 ( .I(n244), .ZN(n247) );
  INVD0 U37 ( .I(n245), .ZN(n244) );
  CKNXD0 U38 ( .I(n247), .ZN(n246) );
  INVD0 U39 ( .I(n240), .ZN(n243) );
  INVD0 U40 ( .I(n241), .ZN(n240) );
  CKNXD0 U41 ( .I(n243), .ZN(n242) );
  INVD0 U42 ( .I(n228), .ZN(n231) );
  INVD0 U43 ( .I(n229), .ZN(n228) );
  CKNXD0 U44 ( .I(n231), .ZN(n230) );
  INVD0 U45 ( .I(n224), .ZN(n227) );
  INVD0 U46 ( .I(n225), .ZN(n224) );
  CKNXD0 U47 ( .I(n227), .ZN(n226) );
  INVD0 U48 ( .I(n208), .ZN(n211) );
  INVD0 U49 ( .I(n209), .ZN(n208) );
  CKNXD0 U50 ( .I(n211), .ZN(n210) );
  INVD0 U51 ( .I(n196), .ZN(n199) );
  INVD0 U52 ( .I(n197), .ZN(n196) );
  CKNXD0 U53 ( .I(n199), .ZN(n198) );
  INVD0 U54 ( .I(n200), .ZN(n203) );
  CKNXD0 U55 ( .I(n201), .ZN(n200) );
  INVD0 U56 ( .I(n195), .ZN(n194) );
  CKNXD0 U57 ( .I(n193), .ZN(n192) );
  INVD0 U58 ( .I(n249), .ZN(n248) );
  INVD0 U59 ( .I(n282), .ZN(n281) );
  CKNXD0 U60 ( .I(n284), .ZN(n283) );
  NR2XD0 U61 ( .A1(n92), .A2(n98), .ZN(N265) );
  NR2XD0 U62 ( .A1(n90), .A2(n97), .ZN(N364) );
  NR2XD0 U63 ( .A1(n89), .A2(n93), .ZN(N496) );
  NR2XD0 U64 ( .A1(n92), .A2(n97), .ZN(N298) );
  NR2XD0 U65 ( .A1(n90), .A2(n98), .ZN(N331) );
  NR2XD0 U66 ( .A1(n89), .A2(n92), .ZN(N562) );
  INVD0 U67 ( .I(N595), .ZN(n193) );
  NR2XD0 U68 ( .A1(n90), .A2(n91), .ZN(N595) );
  NR2XD0 U69 ( .A1(n93), .A2(n97), .ZN(N232) );
  INVD0 U70 ( .I(N529), .ZN(n201) );
  CKNXD0 U71 ( .I(n203), .ZN(n202) );
  NR2XD0 U72 ( .A1(n91), .A2(n92), .ZN(N529) );
  NR2XD0 U73 ( .A1(n93), .A2(n98), .ZN(N199) );
  INVD0 U74 ( .I(N133), .ZN(n249) );
  CKNXD0 U75 ( .I(n251), .ZN(n250) );
  NR2XD0 U76 ( .A1(n91), .A2(n94), .ZN(N397) );
  NR2XD0 U77 ( .A1(n94), .A2(n97), .ZN(N166) );
  NR2XD0 U78 ( .A1(n91), .A2(n93), .ZN(N463) );
  INVD0 U79 ( .I(n188), .ZN(n191) );
  INVD0 U80 ( .I(n191), .ZN(n190) );
  INVD0 U81 ( .I(n189), .ZN(n188) );
  NR2XD0 U82 ( .A1(n89), .A2(n90), .ZN(N628) );
  INVD0 U83 ( .I(n212), .ZN(n215) );
  INVD0 U84 ( .I(n215), .ZN(n214) );
  INVD0 U85 ( .I(n213), .ZN(n212) );
  NR2XD0 U86 ( .A1(n89), .A2(n94), .ZN(N430) );
  INVD0 U87 ( .I(n286), .ZN(n173) );
  CKBD0 U88 ( .CLK(N46), .C(n286) );
  CKAN2D0 U89 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  INVD1 U90 ( .I(N47), .ZN(n171) );
  BUFFD1 U91 ( .I(n305), .Z(n287) );
  BUFFD1 U92 ( .I(n312), .Z(n288) );
  BUFFD1 U93 ( .I(n311), .Z(n289) );
  BUFFD1 U94 ( .I(n311), .Z(n290) );
  BUFFD1 U95 ( .I(n310), .Z(n291) );
  BUFFD1 U96 ( .I(n310), .Z(n292) );
  BUFFD1 U97 ( .I(n309), .Z(n293) );
  BUFFD1 U98 ( .I(n309), .Z(n294) );
  BUFFD1 U99 ( .I(n308), .Z(n295) );
  BUFFD1 U100 ( .I(n308), .Z(n296) );
  BUFFD1 U101 ( .I(n307), .Z(n297) );
  BUFFD1 U102 ( .I(n307), .Z(n298) );
  BUFFD1 U103 ( .I(n306), .Z(n299) );
  BUFFD1 U104 ( .I(n306), .Z(n300) );
  BUFFD1 U105 ( .I(n305), .Z(n301) );
  BUFFD1 U106 ( .I(n305), .Z(n302) );
  BUFFD1 U107 ( .I(n304), .Z(n303) );
  BUFFD1 U108 ( .I(n312), .Z(n311) );
  BUFFD1 U109 ( .I(n312), .Z(n310) );
  BUFFD1 U110 ( .I(n312), .Z(n309) );
  BUFFD1 U111 ( .I(n313), .Z(n308) );
  BUFFD1 U112 ( .I(n313), .Z(n307) );
  BUFFD1 U113 ( .I(n313), .Z(n306) );
  BUFFD1 U114 ( .I(n314), .Z(n305) );
  BUFFD1 U115 ( .I(n314), .Z(n304) );
  BUFFD1 U116 ( .I(n316), .Z(n312) );
  BUFFD1 U117 ( .I(n315), .Z(n313) );
  BUFFD1 U118 ( .I(n315), .Z(n314) );
  BUFFD1 U119 ( .I(n316), .Z(n315) );
  INVD1 U120 ( .I(Reset), .ZN(n316) );
  BUFFD1 U121 ( .I(n269), .Z(n268) );
  BUFFD1 U122 ( .I(n269), .Z(n267) );
  BUFFD1 U123 ( .I(n270), .Z(n266) );
  BUFFD1 U124 ( .I(n270), .Z(n265) );
  BUFFD1 U125 ( .I(n271), .Z(n264) );
  BUFFD1 U126 ( .I(n271), .Z(n263) );
  BUFFD1 U127 ( .I(n272), .Z(n262) );
  BUFFD1 U128 ( .I(n272), .Z(n261) );
  BUFFD1 U129 ( .I(n273), .Z(n260) );
  BUFFD1 U130 ( .I(n273), .Z(n259) );
  BUFFD1 U131 ( .I(n274), .Z(n258) );
  BUFFD1 U132 ( .I(n274), .Z(n257) );
  BUFFD1 U133 ( .I(n275), .Z(n256) );
  BUFFD1 U134 ( .I(n275), .Z(n255) );
  BUFFD1 U135 ( .I(n276), .Z(n254) );
  BUFFD1 U136 ( .I(n277), .Z(n276) );
  BUFFD1 U137 ( .I(n272), .Z(n269) );
  BUFFD1 U138 ( .I(n271), .Z(n270) );
  BUFFD1 U139 ( .I(n278), .Z(n271) );
  BUFFD1 U140 ( .I(n278), .Z(n272) );
  BUFFD1 U141 ( .I(n278), .Z(n273) );
  BUFFD1 U142 ( .I(n277), .Z(n274) );
  BUFFD1 U143 ( .I(n277), .Z(n275) );
  BUFFD1 U144 ( .I(n252), .Z(n278) );
  BUFFD1 U145 ( .I(n252), .Z(n277) );
  BUFFD1 U146 ( .I(n182), .Z(n183) );
  BUFFD1 U147 ( .I(n182), .Z(n184) );
  BUFFD1 U148 ( .I(n182), .Z(n185) );
  BUFFD1 U149 ( .I(n182), .Z(n186) );
  BUFFD1 U150 ( .I(n285), .Z(n187) );
  BUFFD1 U151 ( .I(n176), .Z(n177) );
  BUFFD1 U152 ( .I(n175), .Z(n178) );
  BUFFD1 U153 ( .I(n175), .Z(n179) );
  BUFFD1 U154 ( .I(n175), .Z(n180) );
  BUFFD1 U155 ( .I(N45), .Z(n181) );
  INVD1 U156 ( .I(N397), .ZN(n217) );
  BUFFD1 U157 ( .I(n253), .Z(n252) );
  INVD1 U158 ( .I(n280), .ZN(n279) );
  XOR3D1 U159 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n65), .Z(N84) );
  XOR3D1 U160 ( .A1(DataI[0]), .A2(n66), .A3(n67), .Z(n65) );
  XOR3D1 U161 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n68), .Z(n67) );
  XOR3D1 U162 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n74), .Z(n73) );
  XOR3D1 U163 ( .A1(n75), .A2(DataI[17]), .A3(n76), .Z(n74) );
  XOR3D1 U164 ( .A1(n69), .A2(DataI[3]), .A3(n70), .Z(n68) );
  XOR3D1 U165 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n71), .Z(n70) );
  XOR3D1 U166 ( .A1(n72), .A2(DataI[10]), .A3(n73), .Z(n71) );
  XOR3D1 U167 ( .A1(N59), .A2(N58), .A3(n86), .Z(n85) );
  XOR3D1 U168 ( .A1(n87), .A2(N57), .A3(n88), .Z(n86) );
  XOR3D1 U169 ( .A1(N66), .A2(N65), .A3(n83), .Z(n81) );
  XOR3D1 U170 ( .A1(N64), .A2(n84), .A3(n85), .Z(n83) );
  XOR3D1 U171 ( .A1(N78), .A2(N73), .A3(n77), .Z(N82) );
  XOR3D1 U172 ( .A1(N72), .A2(n78), .A3(n79), .Z(n77) );
  XOR3D1 U173 ( .A1(N76), .A2(N75), .A3(n80), .Z(n79) );
  BUFFD1 U174 ( .I(n285), .Z(n182) );
  INVD1 U175 ( .I(n171), .ZN(n172) );
  INVD1 U176 ( .I(n173), .ZN(n174) );
  INVD1 U177 ( .I(N199), .ZN(n241) );
  INVD1 U178 ( .I(N232), .ZN(n237) );
  ND2D1 U179 ( .A1(n101), .A2(n96), .ZN(n98) );
  ND2D1 U180 ( .A1(n99), .A2(n100), .ZN(n94) );
  ND2D1 U181 ( .A1(n95), .A2(n96), .ZN(n91) );
  INVD1 U182 ( .I(N265), .ZN(n233) );
  INVD1 U183 ( .I(N298), .ZN(n229) );
  INVD1 U184 ( .I(N331), .ZN(n225) );
  INVD1 U185 ( .I(N364), .ZN(n221) );
  INVD1 U186 ( .I(N166), .ZN(n245) );
  INVD1 U187 ( .I(N430), .ZN(n213) );
  INVD1 U188 ( .I(N463), .ZN(n209) );
  INVD1 U189 ( .I(N496), .ZN(n205) );
  INVD1 U190 ( .I(N562), .ZN(n197) );
  INVD1 U191 ( .I(N628), .ZN(n189) );
  INVD1 U192 ( .I(n283), .ZN(n282) );
  INVD1 U193 ( .I(ClockR), .ZN(n280) );
  BUFFD1 U194 ( .I(ClockW), .Z(n253) );
  MUX4D0 U195 ( .I0(n8), .I1(n6), .I2(n7), .I3(n5), .S0(n172), .S1(n174), .Z(
        N80) );
  MUX4D0 U196 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n186), .S1(n176), .Z(n7)
         );
  MUX4D0 U197 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(N44), .S1(n177), .Z(n6)
         );
  MUX4D0 U198 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(N44), .S1(n180), .Z(n8) );
  MUX4D0 U199 ( .I0(n12), .I1(n10), .I2(n11), .I3(n9), .S0(n172), .S1(n174), 
        .Z(N79) );
  MUX4D0 U200 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(N44), .S1(n176), .Z(n11)
         );
  MUX4D0 U201 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n184), .S1(n176), .Z(n10) );
  MUX4D0 U202 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n186), .S1(n175), .Z(n12)
         );
  MUX4D0 U203 ( .I0(n32), .I1(n30), .I2(n31), .I3(n29), .S0(n172), .S1(n174), 
        .Z(N74) );
  MUX4D0 U204 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n285), .S1(n176), .Z(n31)
         );
  MUX4D0 U205 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n285), .S1(n181), .Z(n30) );
  MUX4D0 U206 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(N44), .S1(n175), .Z(n32)
         );
  MUX4D0 U207 ( .I0(n52), .I1(n50), .I2(n51), .I3(n49), .S0(n172), .S1(n174), 
        .Z(N69) );
  MUX4D0 U208 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n187), .S1(n176), .Z(n51) );
  MUX4D0 U209 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n183), .S1(n179), .Z(
        n50) );
  MUX4D0 U210 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n182), .S1(n178), .Z(n52) );
  MUX4D0 U211 ( .I0(n56), .I1(n54), .I2(n55), .I3(n53), .S0(n172), .S1(n174), 
        .Z(N68) );
  MUX4D0 U212 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n285), .S1(n179), .Z(n55) );
  MUX4D0 U213 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n182), .S1(n176), .Z(
        n54) );
  MUX4D0 U214 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(N44), .S1(n179), .Z(n56)
         );
  MUX4D0 U215 ( .I0(n118), .I1(n116), .I2(n117), .I3(n115), .S0(n172), .S1(
        n174), .Z(N62) );
  MUX4D0 U216 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n184), .S1(n178), .Z(
        n117) );
  MUX4D0 U217 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n184), .S1(n178), .Z(
        n116) );
  MUX4D0 U218 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n184), .S1(n178), .Z(
        n118) );
  MUX4D0 U219 ( .I0(n122), .I1(n120), .I2(n121), .I3(n119), .S0(n172), .S1(
        n174), .Z(N61) );
  MUX4D0 U220 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n184), .S1(n178), .Z(
        n121) );
  MUX4D0 U221 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n184), .S1(n178), .Z(
        n120) );
  MUX4D0 U222 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n184), .S1(n178), .Z(
        n122) );
  MUX4D0 U223 ( .I0(n146), .I1(n144), .I2(n145), .I3(n143), .S0(N47), .S1(n286), .Z(N55) );
  MUX4D0 U224 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n186), .S1(n180), .Z(
        n145) );
  MUX4D0 U225 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n186), .S1(n180), .Z(
        n144) );
  MUX4D0 U226 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n186), .S1(n180), .Z(
        n146) );
  MUX4D0 U227 ( .I0(n150), .I1(n148), .I2(n149), .I3(n147), .S0(N47), .S1(n286), .Z(N54) );
  MUX4D0 U228 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n187), .S1(N45), .Z(n149) );
  MUX4D0 U229 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n187), .S1(n180), .Z(
        n148) );
  MUX4D0 U230 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n187), .S1(N45), .Z(n150) );
  MUX4D0 U231 ( .I0(n162), .I1(n160), .I2(n161), .I3(n159), .S0(N47), .S1(N46), 
        .Z(N51) );
  MUX4D0 U232 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n182), .S1(n181), .Z(
        n161) );
  MUX4D0 U233 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n182), .S1(n181), .Z(
        n160) );
  MUX4D0 U234 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n187), .S1(n181), .Z(
        n162) );
  MUX4D0 U235 ( .I0(n166), .I1(n164), .I2(n165), .I3(n163), .S0(N47), .S1(N46), 
        .Z(N50) );
  MUX4D0 U236 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n182), .S1(n181), .Z(
        n165) );
  MUX4D0 U237 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n186), .S1(n181), .Z(
        n164) );
  MUX4D0 U238 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n182), .S1(n181), .Z(
        n166) );
  MUX4D0 U239 ( .I0(n28), .I1(n26), .I2(n27), .I3(n25), .S0(n172), .S1(n174), 
        .Z(N75) );
  MUX4D0 U240 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(N44), .S1(n175), .Z(n27)
         );
  MUX4D0 U241 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(N44), .S1(n175), .Z(n26)
         );
  MUX4D0 U242 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(N44), .S1(n176), .Z(n28)
         );
  MUX4D0 U243 ( .I0(n106), .I1(n104), .I2(n105), .I3(n102), .S0(n172), .S1(
        n174), .Z(N65) );
  MUX4D0 U244 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n183), .S1(n179), .Z(
        n105) );
  MUX4D0 U245 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n183), .S1(n178), .Z(
        n104) );
  MUX4D0 U246 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n183), .S1(n178), .Z(
        n106) );
  MUX4D0 U247 ( .I0(n134), .I1(n132), .I2(n133), .I3(n131), .S0(N47), .S1(N46), 
        .Z(N58) );
  MUX4D0 U248 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n185), .S1(n179), .Z(
        n133) );
  MUX4D0 U249 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n185), .S1(n179), .Z(
        n132) );
  MUX4D0 U250 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n185), .S1(n179), .Z(
        n134) );
  MUX4D0 U251 ( .I0(n138), .I1(n136), .I2(n137), .I3(n135), .S0(N47), .S1(N46), 
        .Z(N57) );
  MUX4D0 U252 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n186), .S1(n180), .Z(
        n137) );
  MUX4D0 U253 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n186), .S1(n180), .Z(
        n136) );
  MUX4D0 U254 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n186), .S1(n180), .Z(
        n138) );
  MUX4D0 U255 ( .I0(n4), .I1(n2), .I2(n3), .I3(n1), .S0(n172), .S1(n174), .Z(
        N81) );
  MUX4D0 U256 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n185), .S1(n181), .Z(n3)
         );
  MUX4D0 U257 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n184), .S1(n177), .Z(n2)
         );
  MUX4D0 U258 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n185), .S1(n177), .Z(n4)
         );
  MUX4D0 U259 ( .I0(n20), .I1(n18), .I2(n19), .I3(n17), .S0(n172), .S1(n174), 
        .Z(N77) );
  MUX4D0 U260 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n285), .S1(n177), .Z(n19)
         );
  MUX4D0 U261 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n185), .S1(n177), .Z(n18) );
  MUX4D0 U262 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n184), .S1(n177), .Z(n20)
         );
  MUX4D0 U263 ( .I0(n44), .I1(n42), .I2(n43), .I3(n41), .S0(n172), .S1(n174), 
        .Z(N71) );
  MUX4D0 U264 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n185), .S1(n175), .Z(n43) );
  MUX4D0 U265 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(N44), .S1(n175), .Z(
        n42) );
  MUX4D0 U266 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n285), .S1(n175), .Z(n44) );
  MUX4D0 U267 ( .I0(n48), .I1(n46), .I2(n47), .I3(n45), .S0(n172), .S1(n174), 
        .Z(N70) );
  MUX4D0 U268 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n182), .S1(n180), .Z(n47) );
  MUX4D0 U269 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n285), .S1(n181), .Z(
        n46) );
  MUX4D0 U270 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n183), .S1(n181), .Z(n48) );
  MUX4D0 U271 ( .I0(n60), .I1(n58), .I2(n59), .I3(n57), .S0(n172), .S1(n174), 
        .Z(N67) );
  MUX4D0 U272 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n182), .S1(n178), .Z(n59) );
  MUX4D0 U273 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n183), .S1(n179), .Z(
        n58) );
  MUX4D0 U274 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n183), .S1(n178), .Z(n60) );
  MUX4D0 U275 ( .I0(n114), .I1(n112), .I2(n113), .I3(n111), .S0(n172), .S1(
        n174), .Z(N63) );
  MUX4D0 U276 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n184), .S1(n178), .Z(
        n113) );
  MUX4D0 U277 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n184), .S1(n178), .Z(
        n112) );
  MUX4D0 U278 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n184), .S1(n178), .Z(
        n114) );
  MUX4D0 U279 ( .I0(n126), .I1(n124), .I2(n125), .I3(n123), .S0(N47), .S1(N46), 
        .Z(N60) );
  MUX4D0 U280 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n185), .S1(n179), .Z(
        n125) );
  MUX4D0 U281 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n185), .S1(n179), .Z(
        n124) );
  MUX4D0 U282 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n185), .S1(n179), .Z(
        n126) );
  MUX4D0 U283 ( .I0(n142), .I1(n140), .I2(n141), .I3(n139), .S0(N47), .S1(n286), .Z(N56) );
  MUX4D0 U284 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n186), .S1(n180), .Z(
        n141) );
  MUX4D0 U285 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n186), .S1(n180), .Z(
        n140) );
  MUX4D0 U286 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n186), .S1(n180), .Z(
        n142) );
  MUX4D0 U287 ( .I0(n154), .I1(n152), .I2(n153), .I3(n151), .S0(N47), .S1(n286), .Z(N53) );
  MUX4D0 U288 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n187), .S1(N45), .Z(n153) );
  MUX4D0 U289 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n187), .S1(n176), .Z(
        n152) );
  MUX4D0 U290 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n187), .S1(n176), .Z(
        n154) );
  MUX4D0 U291 ( .I0(n158), .I1(n156), .I2(n157), .I3(n155), .S0(N47), .S1(n286), .Z(N52) );
  MUX4D0 U292 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n187), .S1(n181), .Z(
        n157) );
  MUX4D0 U293 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n187), .S1(N45), .Z(
        n156) );
  MUX4D0 U294 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n187), .S1(N45), .Z(n158) );
  MUX4D0 U295 ( .I0(n24), .I1(n22), .I2(n23), .I3(n21), .S0(n172), .S1(n174), 
        .Z(N76) );
  MUX4D0 U296 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n186), .S1(n177), .Z(n23)
         );
  MUX4D0 U297 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n185), .S1(n177), .Z(n22) );
  MUX4D0 U298 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n184), .S1(n177), .Z(n24)
         );
  MUX4D0 U299 ( .I0(n40), .I1(n38), .I2(n39), .I3(n37), .S0(n172), .S1(n174), 
        .Z(N72) );
  MUX4D0 U300 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n186), .S1(n180), .Z(n39)
         );
  MUX4D0 U301 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(N44), .S1(n175), .Z(n38)
         );
  MUX4D0 U302 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n184), .S1(n175), .Z(n40)
         );
  MUX4D0 U303 ( .I0(n64), .I1(n62), .I2(n63), .I3(n61), .S0(n172), .S1(n174), 
        .Z(N66) );
  MUX4D0 U304 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n183), .S1(n178), .Z(n63) );
  MUX4D0 U305 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n183), .S1(n177), .Z(
        n62) );
  MUX4D0 U306 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n183), .S1(n178), .Z(n64) );
  MUX4D0 U307 ( .I0(n110), .I1(n108), .I2(n109), .I3(n107), .S0(n172), .S1(
        n174), .Z(N64) );
  MUX4D0 U308 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n183), .S1(n176), .Z(
        n109) );
  MUX4D0 U309 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n183), .S1(n177), .Z(
        n108) );
  MUX4D0 U310 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n183), .S1(n177), .Z(
        n110) );
  MUX4D0 U311 ( .I0(n130), .I1(n128), .I2(n129), .I3(n127), .S0(N47), .S1(N46), 
        .Z(N59) );
  MUX4D0 U312 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n185), .S1(n179), .Z(
        n129) );
  MUX4D0 U313 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n185), .S1(n179), .Z(
        n128) );
  MUX4D0 U314 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n185), .S1(n179), .Z(
        n130) );
  MUX4D0 U315 ( .I0(n170), .I1(n168), .I2(n169), .I3(n167), .S0(N47), .S1(N46), 
        .Z(N49) );
  MUX4D0 U316 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n182), .S1(n181), .Z(
        n169) );
  MUX4D0 U317 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n182), .S1(n181), .Z(
        n168) );
  MUX4D0 U318 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n186), .S1(n181), .Z(
        n170) );
  MUX4D0 U319 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n182), .S1(n181), .Z(
        n167) );
  MUX4D0 U320 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n184), .S1(n177), .Z(n1)
         );
  MUX4D0 U321 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(N44), .S1(n181), .Z(n5)
         );
  MUX4D0 U322 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(N44), .S1(n181), .Z(n9)
         );
  MUX4D0 U323 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n183), .S1(n177), .Z(n17) );
  MUX4D0 U324 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n185), .S1(n177), .Z(n21) );
  MUX4D0 U325 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n182), .S1(n175), .Z(n25) );
  MUX4D0 U326 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n285), .S1(n181), .Z(n29) );
  MUX4D0 U327 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n185), .S1(n180), .Z(n37) );
  MUX4D0 U328 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(N44), .S1(n175), .Z(
        n41) );
  MUX4D0 U329 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(N44), .S1(n176), .Z(
        n45) );
  MUX4D0 U330 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n182), .S1(n179), .Z(
        n49) );
  MUX4D0 U331 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n183), .S1(n178), .Z(
        n53) );
  MUX4D0 U332 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n183), .S1(n176), .Z(
        n57) );
  MUX4D0 U333 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n183), .S1(n177), .Z(
        n61) );
  MUX4D0 U334 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n183), .S1(n179), .Z(
        n102) );
  MUX4D0 U335 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n183), .S1(n179), .Z(
        n107) );
  MUX4D0 U336 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n184), .S1(n178), .Z(
        n111) );
  MUX4D0 U337 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n184), .S1(n178), .Z(
        n115) );
  MUX4D0 U338 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n184), .S1(n178), .Z(
        n119) );
  MUX4D0 U339 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n185), .S1(n179), .Z(
        n123) );
  MUX4D0 U340 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n185), .S1(n179), .Z(
        n127) );
  MUX4D0 U341 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n185), .S1(n179), .Z(
        n131) );
  MUX4D0 U342 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n186), .S1(n180), .Z(
        n135) );
  MUX4D0 U343 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n186), .S1(n180), .Z(
        n139) );
  MUX4D0 U344 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n186), .S1(n180), .Z(
        n143) );
  MUX4D0 U345 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n187), .S1(N45), .Z(
        n147) );
  MUX4D0 U346 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n187), .S1(n176), .Z(
        n151) );
  MUX4D0 U347 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n187), .S1(N45), .Z(
        n155) );
  MUX4D0 U348 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n182), .S1(n181), .Z(
        n159) );
  MUX4D0 U349 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n182), .S1(n181), .Z(
        n163) );
  MUX4D0 U350 ( .I0(n36), .I1(n34), .I2(n35), .I3(n33), .S0(n172), .S1(n174), 
        .Z(N73) );
  MUX4D0 U351 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n285), .S1(N45), .Z(n35)
         );
  MUX4D0 U352 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(N44), .S1(N45), .Z(n34)
         );
  MUX4D0 U353 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n185), .S1(N45), .Z(n36)
         );
  MUX4D0 U354 ( .I0(n16), .I1(n14), .I2(n15), .I3(n13), .S0(N47), .S1(n286), 
        .Z(N78) );
  MUX4D0 U355 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n184), .S1(n177), .Z(n15)
         );
  MUX4D0 U356 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n182), .S1(n177), .Z(n14) );
  MUX4D0 U357 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n183), .S1(n177), .Z(n16)
         );
  MUX4D0 U358 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n285), .S1(n177), .Z(n13) );
  MUX4D0 U359 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n184), .S1(N45), .Z(n33)
         );
  ND2D1 U360 ( .A1(AddrW[1]), .A2(n100), .ZN(n93) );
  ND2D1 U361 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n90) );
  ND2D1 U362 ( .A1(n101), .A2(AddrW[0]), .ZN(n97) );
  ND2D1 U363 ( .A1(AddrW[2]), .A2(n99), .ZN(n92) );
  ND2D1 U364 ( .A1(AddrW[0]), .A2(n95), .ZN(n89) );
  INR2D1 U365 ( .A1(Write), .B1(AddrW[3]), .ZN(n101) );
  INVD1 U366 ( .I(AddrW[1]), .ZN(n99) );
  INVD1 U367 ( .I(AddrW[0]), .ZN(n96) );
  INVD1 U368 ( .I(AddrW[2]), .ZN(n100) );
  AN2D1 U369 ( .A1(Write), .A2(AddrW[3]), .Z(n95) );
  INVD1 U370 ( .I(Read), .ZN(n284) );
  INR2D1 U371 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INR2D1 U372 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U373 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_0 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n5,
         n7, n8, n9, n4;

  AO211D1 U8 ( .A1(n7), .A2(n8), .B(N8), .C(N5), .Z(n9) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n5), .QN(N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n5), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n4), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n4), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n5), .Q(\ClockInN[0] ), 
        .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n5), .QN(n7) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n4), .QN(n5) );
  INVD1 U3 ( .I(Reset), .ZN(n4) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n7), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n8), .A2(n7), .B(n9), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n8) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_0 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n17, n18, n19, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n20, n22, n23, n24, n25, n26, n27, n28,
         n29;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_0_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_0_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_0_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n17), .CP(FastClock), .CDN(n1), .Q(ClockOut) );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n1), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n1), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n19), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[4]), .QN(n13) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n18), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[1]), .QN(n29) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n21), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[0]), .QN(n27) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n1), .Q(
        DivideFactor[3]), .QN(n22) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
  AO222D0 U4 ( .A1(N27), .A2(n2), .B1(N35), .B2(n3), .C1(DivideFactor[0]), 
        .C2(n4), .Z(n21) );
  AO222D0 U5 ( .A1(N31), .A2(n2), .B1(N39), .B2(n3), .C1(DivideFactor[4]), 
        .C2(n4), .Z(n19) );
  AO222D0 U6 ( .A1(N28), .A2(n2), .B1(N36), .B2(n3), .C1(DivideFactor[1]), 
        .C2(n4), .Z(n18) );
  CKND0 U7 ( .CLK(N54), .CN(n4) );
  AN2D0 U8 ( .A1(n5), .A2(n6), .Z(n3) );
  AN3D0 U9 ( .A1(n7), .A2(n8), .A3(n9), .Z(n2) );
  CKXOR2D0 U10 ( .A1(ClockOut), .A2(n10), .Z(n17) );
  AO22D0 U11 ( .A1(N32), .A2(n9), .B1(N40), .B2(n5), .Z(N55) );
  MUX2ND0 U12 ( .I0(n11), .I1(n12), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U13 ( .A1(AdjustFreq[1]), .A2(n6), .ZN(n12) );
  ND3D0 U14 ( .A1(n13), .A2(n8), .A3(n14), .ZN(n6) );
  ND4D0 U15 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n14) );
  IND3D0 U16 ( .A1(AdjustFreq[1]), .B1(n8), .B2(n7), .ZN(n11) );
  CKND2D0 U17 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n7) );
  AO22D0 U18 ( .A1(N30), .A2(n9), .B1(N38), .B2(n5), .Z(N51) );
  AO22D0 U19 ( .A1(N29), .A2(n9), .B1(N37), .B2(n5), .Z(N49) );
  AN2D0 U20 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n5) );
  NR2D0 U21 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n9) );
  INR2D0 U22 ( .A1(N14), .B1(n10), .ZN(N21) );
  INR2D0 U23 ( .A1(N13), .B1(n10), .ZN(N20) );
  INR2D0 U24 ( .A1(N12), .B1(n10), .ZN(N19) );
  INR2D0 U25 ( .A1(N11), .B1(n10), .ZN(N18) );
  INR2D0 U26 ( .A1(N10), .B1(n10), .ZN(N17) );
  INR2D0 U27 ( .A1(N9), .B1(n10), .ZN(N16) );
  OA21D0 U28 ( .A1(FastDivvy[5]), .A2(n8), .B(n15), .Z(n10) );
  IOA22D0 U29 ( .B1(n16), .B2(n20), .A1(n8), .A2(FastDivvy[5]), .ZN(n15) );
  AOI221D0 U30 ( .A1(FastDivvy[4]), .A2(n13), .B1(FastDivvy[3]), .B2(n22), .C(
        n23), .ZN(n20) );
  AOI221D0 U31 ( .A1(DivideFactor[3]), .A2(n24), .B1(DivideFactor[2]), .B2(n25), .C(n26), .ZN(n23) );
  IAO21D0 U32 ( .A1(n25), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n26) );
  OAI32D0 U33 ( .A1(n27), .A2(FastDivvy[0]), .A3(n28), .B1(FastDivvy[1]), .B2(
        n29), .ZN(n25) );
  AN2D0 U34 ( .A1(FastDivvy[1]), .A2(n29), .Z(n28) );
  CKND0 U35 ( .CLK(FastDivvy[3]), .CN(n24) );
  NR2D0 U36 ( .A1(FastDivvy[4]), .A2(n13), .ZN(n16) );
  CKND0 U37 ( .CLK(DivideFactor[5]), .CN(n8) );
  CKND0 U38 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U39 ( .A1(WireD[5]), .A2(n1), .ZN(WireD[0]) );
endmodule


module MultiCounter_0 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_0_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module FIFOTop_AWid3_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(n1), .ClkW(ClkW), .Reset(n3) );
  DPMem1kx32_AWid3_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(n1), .ClkW(ClkW), .ChipEna(
        \*Logic1* ), .Read(n2), .Write(SM_MemWriteCmd), .Reset(n3) );
  INVD0 U2 ( .I(n4), .ZN(n3) );
  BUFFD0 U3 ( .I(ClkR), .Z(n1) );
  INVD1 U4 ( .I(Reseter), .ZN(n4) );
  BUFFD1 U5 ( .I(SM_MemReadCmd), .Z(n2) );
  TIEH U6 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_1 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_1_DW01_dec_0 \ShifterBlock/sub_132  ( .A({\Sh_N[5] , N6, 
        N5, N4, N3, N2}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n18), .CP(n23), .CDN(n29), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n24), .CP(ParClk), .CDN(n27), .Q(HalfParClkr)
         );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(n23), .CDN(n27), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n23), .CDN(n27), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n23), .CDN(n28), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n22), .CDN(n29), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n22), .CDN(n27), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(n22), .CDN(n29), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(n22), .CDN(n28), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(n22), .CDN(n28), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(n21), .CDN(n28), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n21), .CDN(n28), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n21), .CDN(n28), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(n21), .CDN(n28), .Q(InBuf[9]) );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n23), .CDN(n29), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(n23), .CDN(n29), .Q(InBuf[5]) );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n23), .CDN(n29), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(n22), .CDN(n29), .Q(InBuf[1]) );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(n23), .CDN(n27), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n23), .CDN(n28), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(n23), .CDN(n27), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(n22), .CDN(n29), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(n22), .CDN(n28), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n22), .CDN(n27), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n22), .CDN(n29), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(n21), .CDN(n28), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(n21), .CDN(n28), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(n21), .CDN(n28), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(n21), .CDN(n28), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(n21), .CDN(n29), .Q(InBuf[8]) );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n21), .CDN(n29), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(n23), .CDN(n29), .Q(InBuf[4]) );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n22), .CDN(n29), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(n21), .CDN(n29), .Q(InBuf[0]) );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n27), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n27), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n27), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n27), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n27), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n27), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(N31), .CP(SerClk), .CDN(n28), .Q(SerOut) );
  INR2D1 U3 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
  CKBD0 U4 ( .CLK(Reset), .C(n25) );
  CKBXD0 U5 ( .I(Reset), .Z(n26) );
  MUX2ND0 U6 ( .I0(n11), .I1(n12), .S(N4), .ZN(n1) );
  MUX2ND0 U7 ( .I0(n7), .I1(n8), .S(N4), .ZN(n2) );
  INVD0 U8 ( .I(n19), .ZN(n24) );
  MUX2ND0 U9 ( .I0(n9), .I1(n10), .S(N4), .ZN(n3) );
  MUX2ND0 U10 ( .I0(n5), .I1(n6), .S(N4), .ZN(n4) );
  INVD0 U11 ( .I(n20), .ZN(n19) );
  INVD0 U12 ( .I(HalfParClkr), .ZN(n20) );
  INVD1 U13 ( .I(n25), .ZN(n29) );
  INVD1 U14 ( .I(n26), .ZN(n28) );
  INVD1 U15 ( .I(n26), .ZN(n27) );
  INVD1 U16 ( .I(n24), .ZN(n21) );
  INVD1 U17 ( .I(n20), .ZN(n22) );
  INVD1 U18 ( .I(n20), .ZN(n23) );
  INVD1 U19 ( .I(n31), .ZN(n30) );
  ND2D1 U20 ( .A1(N3), .A2(N2), .ZN(n32) );
  AN2D1 U21 ( .A1(N4), .A2(n30), .Z(N26) );
  MUX4ND0 U22 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n5) );
  MUX4ND0 U23 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n6) );
  MUX4ND0 U24 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n7) );
  MUX4ND0 U25 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n8) );
  MUX4ND0 U26 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n9) );
  MUX4ND0 U27 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n10) );
  MUX4ND0 U28 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n11) );
  MUX4ND0 U29 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n12) );
  NR2D1 U30 ( .A1(n32), .A2(N4), .ZN(N24) );
  INVD1 U31 ( .I(n17), .ZN(n18) );
  INVD1 U32 ( .I(N85), .ZN(n17) );
  MUX2ND0 U33 ( .I0(n13), .I1(n14), .S(N6), .ZN(N29) );
  MUX2ND0 U34 ( .I0(n15), .I1(n16), .S(N6), .ZN(N27) );
  MUX2ND0 U35 ( .I0(n14), .I1(n13), .S(N6), .ZN(N25) );
  MUX2ND0 U36 ( .I0(n16), .I1(n15), .S(N6), .ZN(N23) );
  MUX2ND0 U37 ( .I0(n2), .I1(n3), .S(N5), .ZN(n14) );
  MUX2ND0 U38 ( .I0(n1), .I1(n4), .S(N5), .ZN(n13) );
  MUX2ND0 U39 ( .I0(n3), .I1(n1), .S(N5), .ZN(n16) );
  MUX2ND0 U40 ( .I0(n4), .I1(n2), .S(N5), .ZN(n15) );
  OR2D1 U41 ( .A1(N2), .A2(N3), .Z(n31) );
  MUX2ND0 U42 ( .I0(n32), .I1(n31), .S(N4), .ZN(N28) );
  AN2D0 U43 ( .A1(ParIn[31]), .A2(n18), .Z(N84) );
  AN2D0 U44 ( .A1(ParIn[30]), .A2(n18), .Z(N83) );
  AN2D0 U45 ( .A1(ParIn[29]), .A2(N85), .Z(N82) );
  AN2D0 U46 ( .A1(ParIn[28]), .A2(N85), .Z(N81) );
  AN2D0 U47 ( .A1(ParIn[27]), .A2(n18), .Z(N80) );
  AN2D0 U48 ( .A1(ParIn[26]), .A2(N85), .Z(N79) );
  AN2D0 U49 ( .A1(ParIn[25]), .A2(N85), .Z(N78) );
  AN2D0 U50 ( .A1(ParIn[24]), .A2(N85), .Z(N77) );
  AN2D0 U51 ( .A1(ParIn[23]), .A2(N85), .Z(N76) );
  AN2D0 U52 ( .A1(ParIn[22]), .A2(N85), .Z(N75) );
  AN2D0 U53 ( .A1(ParIn[21]), .A2(N85), .Z(N74) );
  AN2D0 U54 ( .A1(ParIn[20]), .A2(N85), .Z(N73) );
  AN2D0 U55 ( .A1(ParIn[19]), .A2(n18), .Z(N72) );
  AN2D0 U56 ( .A1(ParIn[18]), .A2(n18), .Z(N71) );
  AN2D0 U57 ( .A1(ParIn[17]), .A2(N85), .Z(N70) );
  AN2D0 U58 ( .A1(ParIn[16]), .A2(n18), .Z(N69) );
  AN2D0 U59 ( .A1(ParIn[15]), .A2(N85), .Z(N68) );
  AN2D0 U60 ( .A1(ParIn[14]), .A2(n18), .Z(N67) );
  AN2D0 U61 ( .A1(ParIn[13]), .A2(N85), .Z(N66) );
  AN2D0 U62 ( .A1(ParIn[12]), .A2(n18), .Z(N65) );
  AN2D0 U63 ( .A1(ParIn[11]), .A2(N85), .Z(N64) );
  AN2D0 U64 ( .A1(ParIn[10]), .A2(n18), .Z(N63) );
  AN2D0 U65 ( .A1(ParIn[9]), .A2(n18), .Z(N62) );
  AN2D0 U66 ( .A1(ParIn[8]), .A2(n18), .Z(N61) );
  AN2D0 U67 ( .A1(ParIn[7]), .A2(n18), .Z(N60) );
  AN2D0 U68 ( .A1(ParIn[6]), .A2(N85), .Z(N59) );
  AN2D0 U69 ( .A1(ParIn[5]), .A2(n18), .Z(N58) );
  AN2D0 U70 ( .A1(ParIn[4]), .A2(n18), .Z(N57) );
  AN2D0 U71 ( .A1(ParIn[3]), .A2(n18), .Z(N56) );
  AN2D0 U72 ( .A1(ParIn[2]), .A2(n18), .Z(N55) );
  AN2D0 U73 ( .A1(ParIn[1]), .A2(n18), .Z(N54) );
  AN2D0 U74 ( .A1(ParIn[0]), .A2(n18), .Z(N53) );
  IND2D0 U75 ( .A1(n33), .B1(n34), .ZN(N31) );
  OAI21D0 U76 ( .A1(N23), .A2(n35), .B(n36), .ZN(n34) );
  MUX2ND0 U77 ( .I0(n37), .I1(n38), .S(n35), .ZN(n36) );
  MUX3ND0 U78 ( .I0(N25), .I1(n39), .I2(N24), .S0(\Sh_N[5] ), .S1(n40), .ZN(
        n38) );
  NR2D0 U79 ( .A1(\Sh_N[5] ), .A2(N5), .ZN(n40) );
  MUX2D0 U80 ( .I0(n41), .I1(N26), .S(n42), .Z(n39) );
  NR2D0 U81 ( .A1(N6), .A2(N5), .ZN(n42) );
  INR2D0 U82 ( .A1(N27), .B1(N6), .ZN(n41) );
  CKND0 U83 ( .CLK(N5), .CN(n37) );
  CKND2D0 U84 ( .A1(n43), .A2(n44), .ZN(n35) );
  MUX2ND0 U85 ( .I0(n45), .I1(n46), .S(N5), .ZN(n33) );
  CKND2D0 U86 ( .A1(N29), .A2(n47), .ZN(n46) );
  CKND2D0 U87 ( .A1(N28), .A2(n47), .ZN(n45) );
  NR2D0 U88 ( .A1(n44), .A2(n43), .ZN(n47) );
  CKND0 U89 ( .CLK(N6), .CN(n43) );
  CKND0 U90 ( .CLK(\Sh_N[5] ), .CN(n44) );
  INR3D0 U91 ( .A1(n18), .B1(Reset), .B2(n24), .ZN(FIFO_ReadReq) );
endmodule


module SerialTx_1 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_2 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid4_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD0 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_1 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n1, n4, n5, n30, n31, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9027,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U29 ( .A1(n9128), .A2(n9246), .B1(n9129), .B2(Decoder[19]), .ZN(
        n9209) );
  MOAI22D1 U36 ( .A1(n9127), .A2(n9239), .B1(n9129), .B2(Decoder[12]), .ZN(
        n9202) );
  OR3D1 U92 ( .A1(n8960), .A2(n8963), .A3(n8972), .Z(n9266) );
  OR3D1 U94 ( .A1(n8962), .A2(n8966), .A3(n8974), .Z(n9265) );
  OR3D1 U96 ( .A1(n8964), .A2(n8970), .A3(n8973), .Z(n9264) );
  OA21D1 U99 ( .A1(n9262), .A2(n9261), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n9260) );
  DesDecoder_DWid32_1_DW01_inc_0 \ClkGen/add_206  ( .A({Count32[4:2], n6919, 
        n6927}), .SUM({N34, N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(n4), .CPN(n9135), .CDN(n9152), .Q(FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(n30), .CPN(n9132), .CDN(n9148), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(n228), .CPN(n9130), .CDN(n9147), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(n329), .CPN(n9130), .CDN(n9149), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(n426), .CPN(SerClock), .CDN(n9149), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(n524), .CPN(n9136), .CDN(n9150), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(n621), .CPN(n9134), .CDN(n9150), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(n719), .CPN(n9136), .CDN(n9149), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(n721), .CPN(n9134), .CDN(n9149), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(n819), .CPN(n9135), .CDN(n9150), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(n917), .CPN(n9145), .CDN(n9147), .Q(FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(n920), .CPN(n9145), .CDN(n9147), .Q(FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(n922), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(n924), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(n926), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(n928), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(n930), .CPN(n9145), .CDN(n9148), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(n932), .CPN(n9136), .CDN(n9148), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(n934), .CPN(n9131), .CDN(n9148), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(n1031), .CPN(n9131), .CDN(n9150), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(n1129), .CPN(n9135), .CDN(n9153), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(n1131), .CPN(n9133), .CDN(n9152), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(n1133), .CPN(SerClock), .CDN(n9149), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(n1135), .CPN(n9135), .CDN(n9151), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(n1137), .CPN(n9133), .CDN(n9154), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(n1139), .CPN(n9132), .CDN(n9149), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(n1141), .CPN(n9134), .CDN(n9149), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(n1143), .CPN(n9131), .CDN(n9153), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(n1241), .CPN(n9130), .CDN(n9151), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(n1243), .CPN(n9136), .CDN(n9149), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(n1245), .CPN(n9130), .CDN(n9151), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(n1247), .CPN(n9134), .CDN(n9152), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(n1249), .CPN(n9136), .CDN(n9154), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(n1251), .CPN(SerClock), .CDN(n9152), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(n1253), .CPN(n9136), .CDN(n9147), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(n1255), .CPN(n9134), .CDN(n9150), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(n1353), .CPN(n9146), .CDN(n9150), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(n1355), .CPN(n9132), .CDN(n9150), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(n1357), .CPN(n9136), .CDN(n9150), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(n1359), .CPN(SerClock), .CDN(n9150), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(n1361), .CPN(n9130), .CDN(n9154), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(n1363), .CPN(n9131), .CDN(n9152), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[0]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(n1365), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(n1367), .CPN(n9130), .CDN(n9148), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(n1464), .CPN(n9130), .CDN(n9149), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(n1561), .CPN(n9135), .CDN(n9148), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(n1658), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(n1661), .CPN(n9145), .CDN(n9147), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(n1665), .CPN(n9131), .CDN(n9148), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(n1762), .CPN(n9132), .CDN(n9149), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(n1860), .CPN(n9133), .CDN(n9150), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(n1862), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(n1865), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(n1868), .CPN(n9146), .CDN(n9147), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(n1871), .CPN(n9145), .CDN(n9147), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(n1875), .CPN(n9132), .CDN(n9147), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(n1972), .CPN(n9133), .CDN(n9149), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(n2069), .CPN(SerClock), .CDN(n9150), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(n2166), .CPN(n9135), .CDN(n9150), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(n2263), .CPN(n9131), .CDN(n9149), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(n2360), .CPN(SerClock), .CDN(n9150), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(n2457), .CPN(n9133), .CDN(n9148), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(n2554), .CPN(n9134), .CDN(n9148), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(n2556), .E(SerValid), .CP(n9137), .CDN(n9153), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n2557), .CPN(n9134), .CDN(n9147), .Q(
        Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n2691), .CPN(n9146), .CDN(n9153), .Q(
        Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n2827), .CPN(n9133), .CDN(n9149), .Q(
        Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n2963), .CPN(n9132), .CDN(n9151), .Q(
        Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n3099), .CPN(n9146), .CDN(n9149), .Q(
        Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n3235), .CPN(n9144), .CDN(n9154), .Q(
        Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n3371), .CPN(n9144), .CDN(n9153), .Q(
        Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n3507), .CPN(n9144), .CDN(n9147), .Q(
        Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n3643), .CPN(n9144), .CDN(n9153), .Q(
        Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n3779), .CPN(n9144), .CDN(n9153), .Q(
        Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n3915), .CPN(n9144), .CDN(n9151), .Q(
        Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n4051), .CPN(n9144), .CDN(n9151), .Q(
        Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n4188), .CPN(n9144), .CDN(n9154), .Q(
        Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n4324), .CPN(n9144), .CDN(n9148), .Q(
        Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n4460), .CPN(n9143), .CDN(n9152), .Q(
        Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n4596), .CPN(n9143), .CDN(n9153), .Q(
        Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n4732), .CPN(n9143), .CDN(n9152), .Q(
        Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n4868), .CPN(n9143), .CDN(n9153), .Q(
        Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n5004), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n5141), .CPN(n9143), .CDN(n9154), .Q(
        Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n5277), .CPN(n9143), .CDN(n9151), .Q(
        Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n5413), .CPN(n9143), .CDN(n9148), .Q(
        Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n5549), .CPN(n9143), .CDN(n9153), .Q(
        Decoder[9]) );
  DFNCND1 \Decoder_reg[8]  ( .D(n5685), .CPN(n9142), .CDN(n9151), .Q(
        Decoder[8]) );
  DFNCND1 \Decoder_reg[7]  ( .D(n5821), .CPN(n9142), .CDN(n9151), .Q(
        Decoder[7]) );
  DFNCND1 \Decoder_reg[6]  ( .D(n5958), .CPN(n9142), .CDN(n9152), .Q(
        Decoder[6]) );
  DFNCND1 \Decoder_reg[5]  ( .D(n6094), .CPN(n9142), .CDN(n9150), .Q(
        Decoder[5]) );
  DFNCND1 \Decoder_reg[4]  ( .D(n6231), .CPN(n9142), .CDN(n9150), .Q(
        Decoder[4]) );
  DFNCND1 \Decoder_reg[3]  ( .D(n6368), .CPN(n9142), .CDN(n9151), .Q(
        Decoder[3]) );
  DFNCND1 \Decoder_reg[2]  ( .D(n6505), .CPN(n9142), .CDN(n9149), .Q(
        Decoder[2]) );
  DFNCND1 \Decoder_reg[1]  ( .D(n6642), .CPN(n9142), .CDN(n9153), .Q(
        Decoder[1]) );
  DFNCND1 \Decoder_reg[0]  ( .D(n6779), .CPN(n9142), .CDN(n9148), .Q(
        Decoder[0]) );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n6916), .CPN(n9138), .CDN(n9153), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(n6918), .E(SerValid), .CP(n9137), .CDN(n9153), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n6920), .CPN(n9138), .CDN(n9150), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(n6922), .E(SerValid), .CP(n9137), .CDN(n9148), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(n6924), .E(SerValid), .CP(n9137), .CDN(n9147), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(n6926), .E(SerValid), .CP(n9137), .CDN(n9149), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n6928), .CPN(n9141), .CDN(n9151), .Q(ParOut[2]), .QN(n9229) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n6932), .CPN(n9141), .CDN(n9153), .Q(ParOut[1]), .QN(n9228) );
  EDFCNQD1 ParClkr_reg ( .D(n6936), .E(n6938), .CP(n9137), .CDN(n9151), .Q(
        ParClk) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n6940), .CPN(n9141), .CDN(n9154), .Q(ParOut[0]), .QN(n9227) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n6944), .CPN(n9141), .CDN(n9152), .Q(ParOut[5]), .QN(n9232) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n6948), .CPN(n9140), .CDN(n9150), .Q(
        ParOut[12]), .QN(n9239) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n6952), .CPN(n9139), .CDN(n9153), .Q(
        ParOut[19]), .QN(n9246) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n6956), .CPN(n9141), .CDN(n9151), .Q(ParOut[6]), .QN(n9233) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n6960), .CPN(n9140), .CDN(n9150), .Q(ParOut[9]), .QN(n9236) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n6964), .CPN(n9140), .CDN(n9151), .Q(
        ParOut[13]), .QN(n9240) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n6968), .CPN(n9139), .CDN(n9152), .Q(
        ParOut[16]), .QN(n9243) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n6972), .CPN(n9139), .CDN(n9154), .Q(
        ParOut[20]), .QN(n9247) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n6976), .CPN(n9139), .CDN(n9152), .Q(
        ParOut[23]), .QN(n9250) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n6980), .CPN(n9139), .CDN(n9151), .Q(
        ParOut[24]), .QN(n9251) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n6984), .CPN(n9138), .CDN(n9151), .Q(
        ParOut[27]), .QN(n9254) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n6988), .CPN(n9138), .CDN(n9154), .Q(
        ParOut[28]), .QN(n9255) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n6992), .CPN(n9138), .CDN(n9151), .Q(
        ParOut[31]), .QN(n9258) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n6996), .CPN(n9141), .CDN(n9154), .Q(ParOut[3]), .QN(n9230) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n7000), .CPN(n9141), .CDN(n9154), .Q(ParOut[4]), .QN(n9231) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n7004), .CPN(n9140), .CDN(n9147), .Q(
        ParOut[10]), .QN(n9237) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n7008), .CPN(n9140), .CDN(n9153), .Q(
        ParOut[11]), .QN(n9238) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n7012), .CPN(n9139), .CDN(n9149), .Q(
        ParOut[17]), .QN(n9244) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n7016), .CPN(n9139), .CDN(n9149), .Q(
        ParOut[18]), .QN(n9245) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n7020), .CPN(n9140), .CDN(n9152), .Q(ParOut[7]), .QN(n9234) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n7024), .CPN(n9140), .CDN(n9152), .Q(ParOut[8]), .QN(n9235) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n7028), .CPN(n9140), .CDN(n9148), .Q(
        ParOut[14]), .QN(n9241) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n7032), .CPN(n9140), .CDN(n9147), .Q(
        ParOut[15]), .QN(n9242) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n7036), .CPN(n9139), .CDN(n9154), .Q(
        ParOut[21]), .QN(n9248) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n7040), .CPN(n9139), .CDN(n9152), .Q(
        ParOut[22]), .QN(n9249) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n7044), .CPN(n9138), .CDN(n9152), .Q(
        ParOut[25]), .QN(n9252) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n7048), .CPN(n9138), .CDN(n9151), .Q(
        ParOut[26]), .QN(n9253) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n7052), .CPN(n9138), .CDN(n9152), .Q(
        ParOut[29]), .QN(n9256) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n7056), .CPN(n9138), .CDN(n9153), .Q(
        ParOut[30]), .QN(n9257) );
  DFNCND1 ParValidr_reg ( .D(n7060), .CPN(n9137), .CDN(n9152), .Q(ParValid), 
        .QN(n9259) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n9141), .CDN(n9154), .Q(n9261), .QN(
        n9284) );
  DFNCND1 UnLoad_reg ( .D(n9018), .CPN(n9141), .CDN(n9154), .Q(n1), .QN(n9156)
         );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n9019), .CPN(n9137), .CDN(n9154), .QN(
        n9155) );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n9022), .CPN(n9137), .CDN(n9154), .QN(
        n9157) );
  IOA22D0 U3 ( .B1(n9128), .B2(n9258), .A1(n1), .A2(Decoder[31]), .ZN(n9221)
         );
  CKAN2D0 U4 ( .A1(N30), .A2(n9284), .Z(N38) );
  INVD0 U5 ( .I(ParValidTimer[0]), .ZN(n9282) );
  BUFFD0 U6 ( .I(n2826), .Z(n4) );
  CKBD0 U7 ( .CLK(FrameSR[62]), .C(n5) );
  BUFFD0 U8 ( .I(n8992), .Z(n30) );
  CKBD0 U9 ( .CLK(FrameSR[21]), .C(n31) );
  CKBD0 U10 ( .CLK(n31), .C(n64) );
  BUFFD0 U11 ( .I(n64), .Z(n65) );
  CKBD0 U12 ( .CLK(n65), .C(n66) );
  CKBD0 U13 ( .CLK(n66), .C(n67) );
  CKBD0 U14 ( .CLK(n67), .C(n68) );
  CKBD0 U15 ( .CLK(n68), .C(n69) );
  CKBD0 U16 ( .CLK(n69), .C(n70) );
  CKBD0 U17 ( .CLK(n70), .C(n71) );
  CKBD0 U18 ( .CLK(n71), .C(n72) );
  CKBD0 U19 ( .CLK(n72), .C(n73) );
  CKBD0 U20 ( .CLK(n73), .C(n74) );
  CKBD0 U21 ( .CLK(n74), .C(n75) );
  BUFFD0 U22 ( .I(n75), .Z(n76) );
  CKBD0 U23 ( .CLK(n76), .C(n77) );
  CKBD0 U24 ( .CLK(n77), .C(n78) );
  CKBD0 U25 ( .CLK(n78), .C(n79) );
  CKBD0 U26 ( .CLK(n79), .C(n80) );
  CKBD0 U27 ( .CLK(n80), .C(n81) );
  CKBD0 U28 ( .CLK(n81), .C(n82) );
  CKBD0 U30 ( .CLK(n82), .C(n83) );
  CKBD0 U31 ( .CLK(n83), .C(n84) );
  CKBD0 U32 ( .CLK(n84), .C(n85) );
  BUFFD0 U33 ( .I(n85), .Z(n86) );
  CKBD0 U34 ( .CLK(n86), .C(n87) );
  CKBD0 U35 ( .CLK(n87), .C(n88) );
  CKBD0 U37 ( .CLK(n88), .C(n89) );
  CKBD0 U38 ( .CLK(n89), .C(n90) );
  CKBD0 U39 ( .CLK(n90), .C(n91) );
  CKBD0 U40 ( .CLK(n91), .C(n92) );
  CKBD0 U41 ( .CLK(n92), .C(n93) );
  CKBD0 U42 ( .CLK(n93), .C(n94) );
  CKBD0 U43 ( .CLK(n94), .C(n95) );
  CKBD0 U44 ( .CLK(n95), .C(n165) );
  BUFFD0 U45 ( .I(n165), .Z(n166) );
  CKBD0 U46 ( .CLK(n166), .C(n167) );
  CKBD0 U47 ( .CLK(n167), .C(n168) );
  CKBD0 U48 ( .CLK(n168), .C(n169) );
  CKBD0 U49 ( .CLK(n169), .C(n170) );
  CKBD0 U50 ( .CLK(n170), .C(n171) );
  CKBD0 U51 ( .CLK(n171), .C(n172) );
  CKBD0 U52 ( .CLK(n172), .C(n173) );
  CKBD0 U53 ( .CLK(n173), .C(n174) );
  CKBD0 U54 ( .CLK(n174), .C(n175) );
  CKBD0 U55 ( .CLK(n175), .C(n176) );
  BUFFD0 U56 ( .I(n176), .Z(n177) );
  CKBD0 U57 ( .CLK(n177), .C(n178) );
  CKBD0 U58 ( .CLK(n178), .C(n179) );
  CKBD0 U59 ( .CLK(n179), .C(n180) );
  CKBD0 U60 ( .CLK(n180), .C(n181) );
  CKBD0 U61 ( .CLK(n181), .C(n182) );
  CKBD0 U62 ( .CLK(n182), .C(n183) );
  CKBD0 U63 ( .CLK(n183), .C(n184) );
  CKBD0 U64 ( .CLK(n184), .C(n185) );
  CKBD0 U65 ( .CLK(n185), .C(n186) );
  CKBD0 U66 ( .CLK(n186), .C(n187) );
  BUFFD0 U67 ( .I(n187), .Z(n188) );
  CKBD0 U68 ( .CLK(n188), .C(n189) );
  CKBD0 U69 ( .CLK(n189), .C(n190) );
  CKBD0 U70 ( .CLK(n190), .C(n191) );
  CKBD0 U71 ( .CLK(n191), .C(n192) );
  CKBD0 U72 ( .CLK(n192), .C(n193) );
  CKBD0 U73 ( .CLK(n193), .C(n194) );
  CKBD0 U74 ( .CLK(n194), .C(n195) );
  CKBD0 U75 ( .CLK(n195), .C(n196) );
  CKBD0 U76 ( .CLK(n196), .C(n197) );
  CKBD0 U77 ( .CLK(n197), .C(n198) );
  BUFFD0 U78 ( .I(n198), .Z(n199) );
  CKBD0 U79 ( .CLK(n199), .C(n200) );
  CKBD0 U80 ( .CLK(n200), .C(n201) );
  CKBD0 U81 ( .CLK(n201), .C(n202) );
  CKBD0 U82 ( .CLK(n202), .C(n203) );
  CKBD0 U83 ( .CLK(n203), .C(n204) );
  CKBD0 U84 ( .CLK(n204), .C(n205) );
  CKBD0 U85 ( .CLK(n205), .C(n206) );
  CKBD0 U86 ( .CLK(n206), .C(n207) );
  CKBD0 U87 ( .CLK(n207), .C(n208) );
  CKBD0 U88 ( .CLK(n208), .C(n209) );
  BUFFD0 U89 ( .I(n209), .Z(n210) );
  CKBD0 U90 ( .CLK(n210), .C(n211) );
  CKBD0 U91 ( .CLK(n211), .C(n212) );
  CKBD0 U93 ( .CLK(n212), .C(n213) );
  CKBD0 U95 ( .CLK(n213), .C(n214) );
  CKBD0 U97 ( .CLK(n214), .C(n215) );
  CKBD0 U98 ( .CLK(n215), .C(n216) );
  CKBD0 U100 ( .CLK(n216), .C(n217) );
  CKBD0 U102 ( .CLK(n217), .C(n218) );
  CKBD0 U103 ( .CLK(n218), .C(n219) );
  CKBD0 U104 ( .CLK(n219), .C(n220) );
  BUFFD0 U105 ( .I(n220), .Z(n221) );
  CKBD0 U106 ( .CLK(n221), .C(n222) );
  CKBD0 U107 ( .CLK(n222), .C(n223) );
  CKBD0 U108 ( .CLK(n223), .C(n224) );
  CKBD0 U109 ( .CLK(n224), .C(n225) );
  CKBD0 U110 ( .CLK(n225), .C(n226) );
  CKBD0 U111 ( .CLK(n226), .C(n227) );
  BUFFD0 U112 ( .I(n8973), .Z(n228) );
  CKBD0 U113 ( .CLK(FrameSR[22]), .C(n229) );
  BUFFD0 U114 ( .I(n229), .Z(n233) );
  CKBD0 U115 ( .CLK(n233), .C(n234) );
  CKBD0 U116 ( .CLK(n234), .C(n235) );
  CKBD0 U117 ( .CLK(n235), .C(n236) );
  CKBD0 U118 ( .CLK(n236), .C(n237) );
  CKBD0 U119 ( .CLK(n237), .C(n238) );
  CKBD0 U120 ( .CLK(n238), .C(n239) );
  CKBD0 U121 ( .CLK(n239), .C(n240) );
  CKBD0 U122 ( .CLK(n240), .C(n241) );
  CKBD0 U123 ( .CLK(n241), .C(n242) );
  CKBD0 U124 ( .CLK(n242), .C(n243) );
  BUFFD0 U125 ( .I(n243), .Z(n244) );
  CKBD0 U126 ( .CLK(n244), .C(n245) );
  CKBD0 U127 ( .CLK(n245), .C(n246) );
  CKBD0 U128 ( .CLK(n246), .C(n247) );
  CKBD0 U129 ( .CLK(n247), .C(n248) );
  CKBD0 U130 ( .CLK(n248), .C(n249) );
  CKBD0 U131 ( .CLK(n249), .C(n250) );
  CKBD0 U132 ( .CLK(n250), .C(n251) );
  CKBD0 U133 ( .CLK(n251), .C(n252) );
  CKBD0 U134 ( .CLK(n252), .C(n253) );
  CKBD0 U135 ( .CLK(n253), .C(n254) );
  BUFFD0 U136 ( .I(n254), .Z(n255) );
  CKBD0 U137 ( .CLK(n255), .C(n256) );
  CKBD0 U138 ( .CLK(n256), .C(n257) );
  CKBD0 U139 ( .CLK(n257), .C(n258) );
  CKBD0 U140 ( .CLK(n258), .C(n259) );
  CKBD0 U141 ( .CLK(n259), .C(n260) );
  CKBD0 U142 ( .CLK(n260), .C(n261) );
  CKBD0 U143 ( .CLK(n261), .C(n262) );
  CKBD0 U144 ( .CLK(n262), .C(n263) );
  CKBD0 U145 ( .CLK(n263), .C(n264) );
  CKBD0 U146 ( .CLK(n264), .C(n265) );
  BUFFD0 U147 ( .I(n265), .Z(n266) );
  CKBD0 U148 ( .CLK(n266), .C(n267) );
  CKBD0 U149 ( .CLK(n267), .C(n268) );
  CKBD0 U150 ( .CLK(n268), .C(n269) );
  CKBD0 U151 ( .CLK(n269), .C(n270) );
  CKBD0 U152 ( .CLK(n270), .C(n271) );
  CKBD0 U153 ( .CLK(n271), .C(n272) );
  CKBD0 U154 ( .CLK(n272), .C(n273) );
  CKBD0 U155 ( .CLK(n273), .C(n274) );
  CKBD0 U156 ( .CLK(n274), .C(n275) );
  BUFFD0 U157 ( .I(n275), .Z(n276) );
  CKBD0 U158 ( .CLK(n276), .C(n277) );
  CKBD0 U159 ( .CLK(n277), .C(n278) );
  CKBD0 U160 ( .CLK(n278), .C(n279) );
  CKBD0 U161 ( .CLK(n279), .C(n280) );
  CKBD0 U162 ( .CLK(n280), .C(n281) );
  CKBD0 U163 ( .CLK(n281), .C(n282) );
  CKBD0 U164 ( .CLK(n282), .C(n283) );
  CKBD0 U165 ( .CLK(n283), .C(n284) );
  CKBD0 U166 ( .CLK(n284), .C(n285) );
  CKBD0 U167 ( .CLK(n285), .C(n286) );
  BUFFD0 U168 ( .I(n286), .Z(n287) );
  CKBD0 U169 ( .CLK(n287), .C(n288) );
  CKBD0 U170 ( .CLK(n288), .C(n289) );
  CKBD0 U171 ( .CLK(n289), .C(n290) );
  CKBD0 U172 ( .CLK(n290), .C(n291) );
  CKBD0 U173 ( .CLK(n291), .C(n292) );
  CKBD0 U174 ( .CLK(n292), .C(n293) );
  CKBD0 U175 ( .CLK(n293), .C(n294) );
  CKBD0 U176 ( .CLK(n294), .C(n295) );
  CKBD0 U177 ( .CLK(n295), .C(n296) );
  CKBD0 U178 ( .CLK(n296), .C(n297) );
  BUFFD0 U179 ( .I(n297), .Z(n298) );
  CKBD0 U180 ( .CLK(n298), .C(n299) );
  CKBD0 U181 ( .CLK(n299), .C(n300) );
  CKBD0 U182 ( .CLK(n300), .C(n301) );
  CKBD0 U183 ( .CLK(n301), .C(n302) );
  CKBD0 U184 ( .CLK(n302), .C(n303) );
  CKBD0 U185 ( .CLK(n303), .C(n304) );
  CKBD0 U186 ( .CLK(n304), .C(n305) );
  CKBD0 U187 ( .CLK(n305), .C(n306) );
  CKBD0 U188 ( .CLK(n306), .C(n307) );
  CKBD0 U189 ( .CLK(n307), .C(n308) );
  BUFFD0 U190 ( .I(n308), .Z(n309) );
  CKBD0 U191 ( .CLK(n309), .C(n310) );
  CKBD0 U192 ( .CLK(n310), .C(n311) );
  CKBD0 U193 ( .CLK(n311), .C(n312) );
  CKBD0 U194 ( .CLK(n312), .C(n313) );
  CKBD0 U195 ( .CLK(n313), .C(n314) );
  CKBD0 U196 ( .CLK(n314), .C(n315) );
  CKBD0 U197 ( .CLK(n315), .C(n316) );
  CKBD0 U198 ( .CLK(n316), .C(n317) );
  CKBD0 U199 ( .CLK(n317), .C(n318) );
  CKBD0 U200 ( .CLK(n318), .C(n319) );
  BUFFD0 U201 ( .I(n319), .Z(n320) );
  CKBD0 U202 ( .CLK(n320), .C(n321) );
  CKBD0 U203 ( .CLK(n321), .C(n322) );
  CKBD0 U204 ( .CLK(n322), .C(n323) );
  CKBD0 U205 ( .CLK(n323), .C(n324) );
  CKBD0 U206 ( .CLK(n324), .C(n325) );
  CKBD0 U207 ( .CLK(n325), .C(n326) );
  CKBD0 U208 ( .CLK(n326), .C(n327) );
  CKBD0 U209 ( .CLK(n327), .C(n328) );
  BUFFD0 U210 ( .I(n8979), .Z(n329) );
  CKBD0 U211 ( .CLK(FrameSR[36]), .C(n330) );
  CKBD0 U212 ( .CLK(n330), .C(n331) );
  CKBD0 U213 ( .CLK(n331), .C(n332) );
  CKBD0 U214 ( .CLK(n332), .C(n333) );
  CKBD0 U215 ( .CLK(n333), .C(n334) );
  CKBD0 U216 ( .CLK(n334), .C(n335) );
  CKBD0 U217 ( .CLK(n335), .C(n336) );
  CKBD0 U218 ( .CLK(n336), .C(n337) );
  CKBD0 U219 ( .CLK(n337), .C(n338) );
  CKBD0 U220 ( .CLK(n338), .C(n339) );
  BUFFD0 U221 ( .I(n339), .Z(n340) );
  CKBD0 U222 ( .CLK(n340), .C(n341) );
  CKBD0 U223 ( .CLK(n341), .C(n342) );
  CKBD0 U224 ( .CLK(n342), .C(n343) );
  CKBD0 U225 ( .CLK(n343), .C(n344) );
  CKBD0 U226 ( .CLK(n344), .C(n345) );
  CKBD0 U227 ( .CLK(n345), .C(n346) );
  CKBD0 U228 ( .CLK(n346), .C(n347) );
  CKBD0 U229 ( .CLK(n347), .C(n348) );
  CKBD0 U230 ( .CLK(n348), .C(n349) );
  CKBD0 U231 ( .CLK(n349), .C(n350) );
  BUFFD0 U232 ( .I(n350), .Z(n351) );
  CKBD0 U233 ( .CLK(n351), .C(n352) );
  CKBD0 U234 ( .CLK(n352), .C(n353) );
  CKBD0 U235 ( .CLK(n353), .C(n354) );
  CKBD0 U236 ( .CLK(n354), .C(n355) );
  CKBD0 U237 ( .CLK(n355), .C(n356) );
  CKBD0 U238 ( .CLK(n356), .C(n357) );
  CKBD0 U239 ( .CLK(n357), .C(n358) );
  CKBD0 U240 ( .CLK(n358), .C(n359) );
  CKBD0 U241 ( .CLK(n359), .C(n360) );
  CKBD0 U242 ( .CLK(n360), .C(n361) );
  BUFFD0 U243 ( .I(n361), .Z(n362) );
  CKBD0 U244 ( .CLK(n362), .C(n363) );
  CKBD0 U245 ( .CLK(n363), .C(n364) );
  CKBD0 U246 ( .CLK(n364), .C(n365) );
  CKBD0 U247 ( .CLK(n365), .C(n366) );
  CKBD0 U248 ( .CLK(n366), .C(n367) );
  CKBD0 U249 ( .CLK(n367), .C(n368) );
  CKBD0 U250 ( .CLK(n368), .C(n369) );
  CKBD0 U251 ( .CLK(n369), .C(n370) );
  CKBD0 U252 ( .CLK(n370), .C(n371) );
  BUFFD0 U253 ( .I(n371), .Z(n372) );
  CKBD0 U254 ( .CLK(n372), .C(n373) );
  CKBD0 U255 ( .CLK(n373), .C(n374) );
  CKBD0 U256 ( .CLK(n374), .C(n375) );
  CKBD0 U257 ( .CLK(n375), .C(n376) );
  CKBD0 U258 ( .CLK(n376), .C(n377) );
  CKBD0 U259 ( .CLK(n377), .C(n378) );
  CKBD0 U260 ( .CLK(n378), .C(n379) );
  CKBD0 U261 ( .CLK(n379), .C(n380) );
  CKBD0 U262 ( .CLK(n380), .C(n381) );
  CKBD0 U263 ( .CLK(n381), .C(n382) );
  BUFFD0 U264 ( .I(n382), .Z(n383) );
  CKBD0 U265 ( .CLK(n383), .C(n384) );
  CKBD0 U266 ( .CLK(n384), .C(n385) );
  CKBD0 U267 ( .CLK(n385), .C(n386) );
  CKBD0 U268 ( .CLK(n386), .C(n387) );
  CKBD0 U269 ( .CLK(n387), .C(n388) );
  CKBD0 U270 ( .CLK(n388), .C(n389) );
  CKBD0 U271 ( .CLK(n389), .C(n390) );
  CKBD0 U272 ( .CLK(n390), .C(n391) );
  CKBD0 U273 ( .CLK(n391), .C(n392) );
  CKBD0 U274 ( .CLK(n392), .C(n393) );
  BUFFD0 U275 ( .I(n393), .Z(n394) );
  CKBD0 U276 ( .CLK(n394), .C(n395) );
  CKBD0 U277 ( .CLK(n395), .C(n396) );
  CKBD0 U278 ( .CLK(n396), .C(n397) );
  CKBD0 U279 ( .CLK(n397), .C(n398) );
  CKBD0 U280 ( .CLK(n398), .C(n399) );
  CKBD0 U281 ( .CLK(n399), .C(n400) );
  CKBD0 U282 ( .CLK(n400), .C(n401) );
  CKBD0 U283 ( .CLK(n401), .C(n402) );
  CKBD0 U284 ( .CLK(n402), .C(n403) );
  CKBD0 U285 ( .CLK(n403), .C(n404) );
  BUFFD0 U286 ( .I(n404), .Z(n405) );
  CKBD0 U287 ( .CLK(n405), .C(n406) );
  CKBD0 U288 ( .CLK(n406), .C(n407) );
  CKBD0 U289 ( .CLK(n407), .C(n408) );
  CKBD0 U290 ( .CLK(n408), .C(n409) );
  CKBD0 U291 ( .CLK(n409), .C(n410) );
  CKBD0 U292 ( .CLK(n410), .C(n411) );
  CKBD0 U293 ( .CLK(n411), .C(n412) );
  CKBD0 U294 ( .CLK(n412), .C(n413) );
  CKBD0 U295 ( .CLK(n413), .C(n414) );
  CKBD0 U296 ( .CLK(n414), .C(n415) );
  BUFFD0 U297 ( .I(n415), .Z(n416) );
  CKBD0 U298 ( .CLK(n416), .C(n417) );
  CKBD0 U299 ( .CLK(n417), .C(n418) );
  CKBD0 U300 ( .CLK(n418), .C(n419) );
  CKBD0 U301 ( .CLK(n419), .C(n420) );
  CKBD0 U302 ( .CLK(n420), .C(n421) );
  CKBD0 U303 ( .CLK(n421), .C(n422) );
  CKBD0 U304 ( .CLK(n422), .C(n423) );
  CKBD0 U305 ( .CLK(n423), .C(n424) );
  CKBD0 U306 ( .CLK(n424), .C(n425) );
  BUFFD0 U307 ( .I(n8974), .Z(n426) );
  CKBD0 U308 ( .CLK(FrameSR[37]), .C(n427) );
  BUFFD0 U309 ( .I(n427), .Z(n428) );
  CKBD0 U310 ( .CLK(n428), .C(n429) );
  CKBD0 U311 ( .CLK(n429), .C(n430) );
  CKBD0 U312 ( .CLK(n430), .C(n431) );
  CKBD0 U313 ( .CLK(n431), .C(n432) );
  CKBD0 U314 ( .CLK(n432), .C(n433) );
  CKBD0 U315 ( .CLK(n433), .C(n434) );
  CKBD0 U316 ( .CLK(n434), .C(n435) );
  CKBD0 U317 ( .CLK(n435), .C(n436) );
  CKBD0 U318 ( .CLK(n436), .C(n437) );
  CKBD0 U319 ( .CLK(n437), .C(n438) );
  BUFFD0 U320 ( .I(n438), .Z(n439) );
  CKBD0 U321 ( .CLK(n439), .C(n440) );
  CKBD0 U322 ( .CLK(n440), .C(n441) );
  CKBD0 U323 ( .CLK(n441), .C(n442) );
  CKBD0 U324 ( .CLK(n442), .C(n443) );
  CKBD0 U325 ( .CLK(n443), .C(n444) );
  CKBD0 U326 ( .CLK(n444), .C(n445) );
  CKBD0 U327 ( .CLK(n445), .C(n446) );
  CKBD0 U328 ( .CLK(n446), .C(n447) );
  CKBD0 U329 ( .CLK(n447), .C(n448) );
  CKBD0 U330 ( .CLK(n448), .C(n449) );
  BUFFD0 U331 ( .I(n449), .Z(n450) );
  CKBD0 U332 ( .CLK(n450), .C(n451) );
  CKBD0 U333 ( .CLK(n451), .C(n452) );
  CKBD0 U334 ( .CLK(n452), .C(n453) );
  CKBD0 U335 ( .CLK(n453), .C(n454) );
  CKBD0 U336 ( .CLK(n454), .C(n455) );
  CKBD0 U337 ( .CLK(n455), .C(n456) );
  CKBD0 U338 ( .CLK(n456), .C(n457) );
  CKBD0 U339 ( .CLK(n457), .C(n458) );
  CKBD0 U340 ( .CLK(n458), .C(n459) );
  CKBD0 U341 ( .CLK(n459), .C(n460) );
  BUFFD0 U342 ( .I(n460), .Z(n461) );
  CKBD0 U343 ( .CLK(n461), .C(n462) );
  CKBD0 U344 ( .CLK(n462), .C(n463) );
  CKBD0 U345 ( .CLK(n463), .C(n464) );
  CKBD0 U346 ( .CLK(n464), .C(n465) );
  CKBD0 U347 ( .CLK(n465), .C(n466) );
  CKBD0 U348 ( .CLK(n466), .C(n467) );
  CKBD0 U349 ( .CLK(n467), .C(n468) );
  CKBD0 U350 ( .CLK(n468), .C(n469) );
  CKBD0 U351 ( .CLK(n469), .C(n470) );
  BUFFD0 U352 ( .I(n470), .Z(n471) );
  CKBD0 U353 ( .CLK(n471), .C(n472) );
  CKBD0 U354 ( .CLK(n472), .C(n473) );
  CKBD0 U355 ( .CLK(n473), .C(n474) );
  CKBD0 U356 ( .CLK(n474), .C(n475) );
  CKBD0 U357 ( .CLK(n475), .C(n476) );
  CKBD0 U358 ( .CLK(n476), .C(n477) );
  CKBD0 U359 ( .CLK(n477), .C(n478) );
  CKBD0 U360 ( .CLK(n478), .C(n479) );
  CKBD0 U361 ( .CLK(n479), .C(n480) );
  CKBD0 U362 ( .CLK(n480), .C(n481) );
  BUFFD0 U363 ( .I(n481), .Z(n482) );
  CKBD0 U364 ( .CLK(n482), .C(n483) );
  CKBD0 U365 ( .CLK(n483), .C(n484) );
  CKBD0 U366 ( .CLK(n484), .C(n485) );
  CKBD0 U367 ( .CLK(n485), .C(n486) );
  CKBD0 U368 ( .CLK(n486), .C(n487) );
  CKBD0 U369 ( .CLK(n487), .C(n488) );
  CKBD0 U370 ( .CLK(n488), .C(n489) );
  CKBD0 U371 ( .CLK(n489), .C(n490) );
  CKBD0 U372 ( .CLK(n490), .C(n491) );
  CKBD0 U373 ( .CLK(n491), .C(n492) );
  BUFFD0 U374 ( .I(n492), .Z(n493) );
  CKBD0 U375 ( .CLK(n493), .C(n494) );
  CKBD0 U376 ( .CLK(n494), .C(n495) );
  CKBD0 U377 ( .CLK(n495), .C(n496) );
  CKBD0 U378 ( .CLK(n496), .C(n497) );
  CKBD0 U379 ( .CLK(n497), .C(n498) );
  CKBD0 U380 ( .CLK(n498), .C(n499) );
  CKBD0 U381 ( .CLK(n499), .C(n500) );
  CKBD0 U382 ( .CLK(n500), .C(n501) );
  CKBD0 U383 ( .CLK(n501), .C(n502) );
  CKBD0 U384 ( .CLK(n502), .C(n503) );
  BUFFD0 U385 ( .I(n503), .Z(n504) );
  CKBD0 U386 ( .CLK(n504), .C(n505) );
  CKBD0 U387 ( .CLK(n505), .C(n506) );
  CKBD0 U388 ( .CLK(n506), .C(n507) );
  CKBD0 U389 ( .CLK(n507), .C(n508) );
  CKBD0 U390 ( .CLK(n508), .C(n509) );
  CKBD0 U391 ( .CLK(n509), .C(n510) );
  CKBD0 U392 ( .CLK(n510), .C(n511) );
  CKBD0 U393 ( .CLK(n511), .C(n512) );
  CKBD0 U394 ( .CLK(n512), .C(n513) );
  CKBD0 U395 ( .CLK(n513), .C(n514) );
  BUFFD0 U396 ( .I(n514), .Z(n515) );
  CKBD0 U397 ( .CLK(n515), .C(n516) );
  CKBD0 U398 ( .CLK(n516), .C(n517) );
  CKBD0 U399 ( .CLK(n517), .C(n518) );
  CKBD0 U400 ( .CLK(n518), .C(n519) );
  CKBD0 U401 ( .CLK(n519), .C(n520) );
  CKBD0 U402 ( .CLK(n520), .C(n521) );
  CKBD0 U403 ( .CLK(n521), .C(n522) );
  CKBD0 U404 ( .CLK(n522), .C(n523) );
  BUFFD0 U405 ( .I(n8978), .Z(n524) );
  CKBD0 U406 ( .CLK(FrameSR[52]), .C(n525) );
  CKBD0 U407 ( .CLK(n525), .C(n526) );
  CKBD0 U408 ( .CLK(n526), .C(n527) );
  CKBD0 U409 ( .CLK(n527), .C(n528) );
  CKBD0 U410 ( .CLK(n528), .C(n529) );
  CKBD0 U411 ( .CLK(n529), .C(n530) );
  CKBD0 U412 ( .CLK(n530), .C(n531) );
  CKBD0 U413 ( .CLK(n531), .C(n532) );
  CKBD0 U414 ( .CLK(n532), .C(n533) );
  CKBD0 U415 ( .CLK(n533), .C(n534) );
  BUFFD0 U416 ( .I(n534), .Z(n535) );
  CKBD0 U417 ( .CLK(n535), .C(n536) );
  CKBD0 U418 ( .CLK(n536), .C(n537) );
  CKBD0 U419 ( .CLK(n537), .C(n538) );
  CKBD0 U420 ( .CLK(n538), .C(n539) );
  CKBD0 U421 ( .CLK(n539), .C(n540) );
  CKBD0 U422 ( .CLK(n540), .C(n541) );
  CKBD0 U423 ( .CLK(n541), .C(n542) );
  CKBD0 U424 ( .CLK(n542), .C(n543) );
  CKBD0 U425 ( .CLK(n543), .C(n544) );
  CKBD0 U426 ( .CLK(n544), .C(n545) );
  BUFFD0 U427 ( .I(n545), .Z(n546) );
  CKBD0 U428 ( .CLK(n546), .C(n547) );
  CKBD0 U429 ( .CLK(n547), .C(n548) );
  CKBD0 U430 ( .CLK(n548), .C(n549) );
  CKBD0 U431 ( .CLK(n549), .C(n550) );
  CKBD0 U432 ( .CLK(n550), .C(n551) );
  CKBD0 U433 ( .CLK(n551), .C(n552) );
  CKBD0 U434 ( .CLK(n552), .C(n553) );
  CKBD0 U435 ( .CLK(n553), .C(n554) );
  CKBD0 U436 ( .CLK(n554), .C(n555) );
  CKBD0 U437 ( .CLK(n555), .C(n556) );
  BUFFD0 U438 ( .I(n556), .Z(n557) );
  CKBD0 U439 ( .CLK(n557), .C(n558) );
  CKBD0 U440 ( .CLK(n558), .C(n559) );
  CKBD0 U441 ( .CLK(n559), .C(n560) );
  CKBD0 U442 ( .CLK(n560), .C(n561) );
  CKBD0 U443 ( .CLK(n561), .C(n562) );
  CKBD0 U444 ( .CLK(n562), .C(n563) );
  CKBD0 U445 ( .CLK(n563), .C(n564) );
  CKBD0 U446 ( .CLK(n564), .C(n565) );
  CKBD0 U447 ( .CLK(n565), .C(n566) );
  CKBD0 U448 ( .CLK(n566), .C(n567) );
  BUFFD0 U449 ( .I(n567), .Z(n568) );
  CKBD0 U450 ( .CLK(n568), .C(n569) );
  CKBD0 U451 ( .CLK(n569), .C(n570) );
  CKBD0 U452 ( .CLK(n570), .C(n571) );
  CKBD0 U453 ( .CLK(n571), .C(n572) );
  CKBD0 U454 ( .CLK(n572), .C(n573) );
  CKBD0 U455 ( .CLK(n573), .C(n574) );
  CKBD0 U456 ( .CLK(n574), .C(n575) );
  CKBD0 U457 ( .CLK(n575), .C(n576) );
  CKBD0 U458 ( .CLK(n576), .C(n577) );
  CKBD0 U459 ( .CLK(n577), .C(n578) );
  BUFFD0 U460 ( .I(n578), .Z(n579) );
  CKBD0 U461 ( .CLK(n579), .C(n580) );
  CKBD0 U462 ( .CLK(n580), .C(n581) );
  CKBD0 U463 ( .CLK(n581), .C(n582) );
  CKBD0 U464 ( .CLK(n582), .C(n583) );
  CKBD0 U465 ( .CLK(n583), .C(n584) );
  CKBD0 U466 ( .CLK(n584), .C(n585) );
  CKBD0 U467 ( .CLK(n585), .C(n586) );
  CKBD0 U468 ( .CLK(n586), .C(n587) );
  CKBD0 U469 ( .CLK(n587), .C(n588) );
  CKBD0 U470 ( .CLK(n588), .C(n589) );
  BUFFD0 U471 ( .I(n589), .Z(n590) );
  CKBD0 U472 ( .CLK(n590), .C(n591) );
  CKBD0 U473 ( .CLK(n591), .C(n592) );
  CKBD0 U474 ( .CLK(n592), .C(n593) );
  CKBD0 U475 ( .CLK(n593), .C(n594) );
  CKBD0 U476 ( .CLK(n594), .C(n595) );
  CKBD0 U477 ( .CLK(n595), .C(n596) );
  CKBD0 U478 ( .CLK(n596), .C(n597) );
  CKBD0 U479 ( .CLK(n597), .C(n598) );
  CKBD0 U480 ( .CLK(n598), .C(n599) );
  BUFFD0 U481 ( .I(n599), .Z(n600) );
  CKBD0 U482 ( .CLK(n600), .C(n601) );
  CKBD0 U483 ( .CLK(n601), .C(n602) );
  CKBD0 U484 ( .CLK(n602), .C(n603) );
  CKBD0 U485 ( .CLK(n603), .C(n604) );
  CKBD0 U486 ( .CLK(n604), .C(n605) );
  CKBD0 U487 ( .CLK(n605), .C(n606) );
  CKBD0 U488 ( .CLK(n606), .C(n607) );
  CKBD0 U489 ( .CLK(n607), .C(n608) );
  CKBD0 U490 ( .CLK(n608), .C(n609) );
  CKBD0 U491 ( .CLK(n609), .C(n610) );
  BUFFD0 U492 ( .I(n610), .Z(n611) );
  CKBD0 U493 ( .CLK(n611), .C(n612) );
  CKBD0 U494 ( .CLK(n612), .C(n613) );
  CKBD0 U495 ( .CLK(n613), .C(n614) );
  CKBD0 U496 ( .CLK(n614), .C(n615) );
  CKBD0 U497 ( .CLK(n615), .C(n616) );
  CKBD0 U498 ( .CLK(n616), .C(n617) );
  CKBD0 U499 ( .CLK(n617), .C(n618) );
  CKBD0 U500 ( .CLK(n618), .C(n619) );
  CKBD0 U501 ( .CLK(n619), .C(n620) );
  BUFFD0 U502 ( .I(n8972), .Z(n621) );
  CKBD0 U503 ( .CLK(FrameSR[53]), .C(n622) );
  BUFFD0 U504 ( .I(n622), .Z(n623) );
  CKBD0 U505 ( .CLK(n623), .C(n624) );
  CKBD0 U506 ( .CLK(n624), .C(n625) );
  CKBD0 U507 ( .CLK(n625), .C(n626) );
  CKBD0 U508 ( .CLK(n626), .C(n627) );
  CKBD0 U509 ( .CLK(n627), .C(n628) );
  CKBD0 U510 ( .CLK(n628), .C(n629) );
  CKBD0 U511 ( .CLK(n629), .C(n630) );
  CKBD0 U512 ( .CLK(n630), .C(n631) );
  CKBD0 U513 ( .CLK(n631), .C(n632) );
  CKBD0 U514 ( .CLK(n632), .C(n633) );
  BUFFD0 U515 ( .I(n633), .Z(n634) );
  CKBD0 U516 ( .CLK(n634), .C(n635) );
  CKBD0 U517 ( .CLK(n635), .C(n636) );
  CKBD0 U518 ( .CLK(n636), .C(n637) );
  CKBD0 U519 ( .CLK(n637), .C(n638) );
  CKBD0 U520 ( .CLK(n638), .C(n639) );
  CKBD0 U521 ( .CLK(n639), .C(n640) );
  CKBD0 U522 ( .CLK(n640), .C(n641) );
  CKBD0 U523 ( .CLK(n641), .C(n642) );
  CKBD0 U524 ( .CLK(n642), .C(n643) );
  CKBD0 U525 ( .CLK(n643), .C(n644) );
  BUFFD0 U526 ( .I(n644), .Z(n645) );
  CKBD0 U527 ( .CLK(n645), .C(n646) );
  CKBD0 U528 ( .CLK(n646), .C(n647) );
  CKBD0 U529 ( .CLK(n647), .C(n648) );
  CKBD0 U530 ( .CLK(n648), .C(n649) );
  CKBD0 U531 ( .CLK(n649), .C(n650) );
  CKBD0 U532 ( .CLK(n650), .C(n651) );
  CKBD0 U533 ( .CLK(n651), .C(n652) );
  CKBD0 U534 ( .CLK(n652), .C(n653) );
  CKBD0 U535 ( .CLK(n653), .C(n654) );
  CKBD0 U536 ( .CLK(n654), .C(n655) );
  BUFFD0 U537 ( .I(n655), .Z(n656) );
  CKBD0 U538 ( .CLK(n656), .C(n657) );
  CKBD0 U539 ( .CLK(n657), .C(n658) );
  CKBD0 U540 ( .CLK(n658), .C(n659) );
  CKBD0 U541 ( .CLK(n659), .C(n660) );
  CKBD0 U542 ( .CLK(n660), .C(n661) );
  CKBD0 U543 ( .CLK(n661), .C(n662) );
  CKBD0 U544 ( .CLK(n662), .C(n663) );
  CKBD0 U545 ( .CLK(n663), .C(n664) );
  CKBD0 U546 ( .CLK(n664), .C(n665) );
  BUFFD0 U547 ( .I(n665), .Z(n666) );
  CKBD0 U548 ( .CLK(n666), .C(n667) );
  CKBD0 U549 ( .CLK(n667), .C(n668) );
  CKBD0 U550 ( .CLK(n668), .C(n669) );
  CKBD0 U551 ( .CLK(n669), .C(n670) );
  CKBD0 U552 ( .CLK(n670), .C(n671) );
  CKBD0 U553 ( .CLK(n671), .C(n672) );
  CKBD0 U554 ( .CLK(n672), .C(n673) );
  CKBD0 U555 ( .CLK(n673), .C(n674) );
  CKBD0 U556 ( .CLK(n674), .C(n675) );
  CKBD0 U557 ( .CLK(n675), .C(n676) );
  BUFFD0 U558 ( .I(n676), .Z(n677) );
  CKBD0 U559 ( .CLK(n677), .C(n678) );
  CKBD0 U560 ( .CLK(n678), .C(n679) );
  CKBD0 U561 ( .CLK(n679), .C(n680) );
  CKBD0 U562 ( .CLK(n680), .C(n681) );
  CKBD0 U563 ( .CLK(n681), .C(n682) );
  CKBD0 U564 ( .CLK(n682), .C(n683) );
  CKBD0 U565 ( .CLK(n683), .C(n684) );
  CKBD0 U566 ( .CLK(n684), .C(n685) );
  CKBD0 U567 ( .CLK(n685), .C(n686) );
  CKBD0 U568 ( .CLK(n686), .C(n687) );
  BUFFD0 U569 ( .I(n687), .Z(n688) );
  CKBD0 U570 ( .CLK(n688), .C(n689) );
  CKBD0 U571 ( .CLK(n689), .C(n690) );
  CKBD0 U572 ( .CLK(n690), .C(n691) );
  CKBD0 U573 ( .CLK(n691), .C(n692) );
  CKBD0 U574 ( .CLK(n692), .C(n693) );
  CKBD0 U575 ( .CLK(n693), .C(n694) );
  CKBD0 U576 ( .CLK(n694), .C(n695) );
  CKBD0 U577 ( .CLK(n695), .C(n696) );
  CKBD0 U578 ( .CLK(n696), .C(n697) );
  CKBD0 U579 ( .CLK(n697), .C(n698) );
  BUFFD0 U580 ( .I(n698), .Z(n699) );
  CKBD0 U581 ( .CLK(n699), .C(n700) );
  CKBD0 U582 ( .CLK(n700), .C(n701) );
  CKBD0 U583 ( .CLK(n701), .C(n702) );
  CKBD0 U584 ( .CLK(n702), .C(n703) );
  CKBD0 U585 ( .CLK(n703), .C(n704) );
  CKBD0 U586 ( .CLK(n704), .C(n705) );
  CKBD0 U587 ( .CLK(n705), .C(n706) );
  CKBD0 U588 ( .CLK(n706), .C(n707) );
  CKBD0 U589 ( .CLK(n707), .C(n708) );
  CKBD0 U590 ( .CLK(n708), .C(n709) );
  BUFFD0 U591 ( .I(n709), .Z(n710) );
  CKBD0 U592 ( .CLK(n710), .C(n711) );
  CKBD0 U593 ( .CLK(n711), .C(n712) );
  CKBD0 U594 ( .CLK(n712), .C(n713) );
  CKBD0 U595 ( .CLK(n713), .C(n714) );
  CKBD0 U596 ( .CLK(n714), .C(n715) );
  CKBD0 U597 ( .CLK(n715), .C(n716) );
  CKBD0 U598 ( .CLK(n716), .C(n717) );
  CKBD0 U599 ( .CLK(n717), .C(n718) );
  BUFFD0 U600 ( .I(n4867), .Z(n719) );
  CKBD0 U601 ( .CLK(FrameSR[31]), .C(n720) );
  BUFFD0 U602 ( .I(n8966), .Z(n721) );
  CKBD0 U603 ( .CLK(FrameSR[38]), .C(n722) );
  BUFFD0 U604 ( .I(n722), .Z(n723) );
  CKBD0 U605 ( .CLK(n723), .C(n724) );
  CKBD0 U606 ( .CLK(n724), .C(n725) );
  CKBD0 U607 ( .CLK(n725), .C(n726) );
  CKBD0 U608 ( .CLK(n726), .C(n727) );
  CKBD0 U609 ( .CLK(n727), .C(n728) );
  CKBD0 U610 ( .CLK(n728), .C(n729) );
  CKBD0 U611 ( .CLK(n729), .C(n730) );
  CKBD0 U612 ( .CLK(n730), .C(n731) );
  CKBD0 U613 ( .CLK(n731), .C(n732) );
  CKBD0 U614 ( .CLK(n732), .C(n733) );
  BUFFD0 U615 ( .I(n733), .Z(n734) );
  CKBD0 U616 ( .CLK(n734), .C(n735) );
  CKBD0 U617 ( .CLK(n735), .C(n736) );
  CKBD0 U618 ( .CLK(n736), .C(n737) );
  CKBD0 U619 ( .CLK(n737), .C(n738) );
  CKBD0 U620 ( .CLK(n738), .C(n739) );
  CKBD0 U621 ( .CLK(n739), .C(n740) );
  CKBD0 U622 ( .CLK(n740), .C(n741) );
  CKBD0 U623 ( .CLK(n741), .C(n742) );
  CKBD0 U624 ( .CLK(n742), .C(n743) );
  CKBD0 U625 ( .CLK(n743), .C(n744) );
  BUFFD0 U626 ( .I(n744), .Z(n745) );
  CKBD0 U627 ( .CLK(n745), .C(n746) );
  CKBD0 U628 ( .CLK(n746), .C(n747) );
  CKBD0 U629 ( .CLK(n747), .C(n748) );
  CKBD0 U630 ( .CLK(n748), .C(n749) );
  CKBD0 U631 ( .CLK(n749), .C(n750) );
  CKBD0 U632 ( .CLK(n750), .C(n751) );
  CKBD0 U633 ( .CLK(n751), .C(n752) );
  CKBD0 U634 ( .CLK(n752), .C(n753) );
  CKBD0 U635 ( .CLK(n753), .C(n754) );
  CKBD0 U636 ( .CLK(n754), .C(n755) );
  BUFFD0 U637 ( .I(n755), .Z(n756) );
  CKBD0 U638 ( .CLK(n756), .C(n757) );
  CKBD0 U639 ( .CLK(n757), .C(n758) );
  CKBD0 U640 ( .CLK(n758), .C(n759) );
  CKBD0 U641 ( .CLK(n759), .C(n760) );
  CKBD0 U642 ( .CLK(n760), .C(n761) );
  CKBD0 U643 ( .CLK(n761), .C(n762) );
  CKBD0 U644 ( .CLK(n762), .C(n763) );
  CKBD0 U645 ( .CLK(n763), .C(n764) );
  CKBD0 U646 ( .CLK(n764), .C(n765) );
  BUFFD0 U647 ( .I(n765), .Z(n766) );
  CKBD0 U648 ( .CLK(n766), .C(n767) );
  CKBD0 U649 ( .CLK(n767), .C(n768) );
  CKBD0 U650 ( .CLK(n768), .C(n769) );
  CKBD0 U651 ( .CLK(n769), .C(n770) );
  CKBD0 U652 ( .CLK(n770), .C(n771) );
  CKBD0 U653 ( .CLK(n771), .C(n772) );
  CKBD0 U654 ( .CLK(n772), .C(n773) );
  CKBD0 U655 ( .CLK(n773), .C(n774) );
  CKBD0 U656 ( .CLK(n774), .C(n775) );
  CKBD0 U657 ( .CLK(n775), .C(n776) );
  BUFFD0 U658 ( .I(n776), .Z(n777) );
  CKBD0 U659 ( .CLK(n777), .C(n778) );
  CKBD0 U660 ( .CLK(n778), .C(n779) );
  CKBD0 U661 ( .CLK(n779), .C(n780) );
  CKBD0 U662 ( .CLK(n780), .C(n781) );
  CKBD0 U663 ( .CLK(n781), .C(n782) );
  CKBD0 U664 ( .CLK(n782), .C(n783) );
  CKBD0 U665 ( .CLK(n783), .C(n784) );
  CKBD0 U666 ( .CLK(n784), .C(n785) );
  CKBD0 U667 ( .CLK(n785), .C(n786) );
  CKBD0 U668 ( .CLK(n786), .C(n787) );
  BUFFD0 U669 ( .I(n787), .Z(n788) );
  CKBD0 U670 ( .CLK(n788), .C(n789) );
  CKBD0 U671 ( .CLK(n789), .C(n790) );
  CKBD0 U672 ( .CLK(n790), .C(n791) );
  CKBD0 U673 ( .CLK(n791), .C(n792) );
  CKBD0 U674 ( .CLK(n792), .C(n793) );
  CKBD0 U675 ( .CLK(n793), .C(n794) );
  CKBD0 U676 ( .CLK(n794), .C(n795) );
  CKBD0 U677 ( .CLK(n795), .C(n796) );
  CKBD0 U678 ( .CLK(n796), .C(n797) );
  CKBD0 U679 ( .CLK(n797), .C(n798) );
  BUFFD0 U680 ( .I(n798), .Z(n799) );
  CKBD0 U681 ( .CLK(n799), .C(n800) );
  CKBD0 U682 ( .CLK(n800), .C(n801) );
  CKBD0 U683 ( .CLK(n801), .C(n802) );
  CKBD0 U684 ( .CLK(n802), .C(n803) );
  CKBD0 U685 ( .CLK(n803), .C(n804) );
  CKBD0 U686 ( .CLK(n804), .C(n805) );
  CKBD0 U687 ( .CLK(n805), .C(n806) );
  CKBD0 U688 ( .CLK(n806), .C(n807) );
  CKBD0 U689 ( .CLK(n807), .C(n808) );
  CKBD0 U690 ( .CLK(n808), .C(n809) );
  BUFFD0 U691 ( .I(n809), .Z(n810) );
  CKBD0 U692 ( .CLK(n810), .C(n811) );
  CKBD0 U693 ( .CLK(n811), .C(n812) );
  CKBD0 U694 ( .CLK(n812), .C(n813) );
  CKBD0 U695 ( .CLK(n813), .C(n814) );
  CKBD0 U696 ( .CLK(n814), .C(n815) );
  CKBD0 U697 ( .CLK(n815), .C(n816) );
  CKBD0 U698 ( .CLK(n816), .C(n817) );
  CKBD0 U699 ( .CLK(n817), .C(n818) );
  BUFFD0 U700 ( .I(n8963), .Z(n819) );
  CKBD0 U701 ( .CLK(FrameSR[54]), .C(n820) );
  BUFFD0 U702 ( .I(n820), .Z(n821) );
  CKBD0 U703 ( .CLK(n821), .C(n822) );
  CKBD0 U704 ( .CLK(n822), .C(n823) );
  CKBD0 U705 ( .CLK(n823), .C(n824) );
  CKBD0 U706 ( .CLK(n824), .C(n825) );
  CKBD0 U707 ( .CLK(n825), .C(n826) );
  CKBD0 U708 ( .CLK(n826), .C(n827) );
  CKBD0 U709 ( .CLK(n827), .C(n828) );
  CKBD0 U710 ( .CLK(n828), .C(n829) );
  CKBD0 U711 ( .CLK(n829), .C(n830) );
  CKBD0 U712 ( .CLK(n830), .C(n831) );
  BUFFD0 U713 ( .I(n831), .Z(n832) );
  CKBD0 U714 ( .CLK(n832), .C(n833) );
  CKBD0 U715 ( .CLK(n833), .C(n834) );
  CKBD0 U716 ( .CLK(n834), .C(n835) );
  CKBD0 U717 ( .CLK(n835), .C(n836) );
  CKBD0 U718 ( .CLK(n836), .C(n837) );
  CKBD0 U719 ( .CLK(n837), .C(n838) );
  CKBD0 U720 ( .CLK(n838), .C(n839) );
  CKBD0 U721 ( .CLK(n839), .C(n840) );
  CKBD0 U722 ( .CLK(n840), .C(n841) );
  CKBD0 U723 ( .CLK(n841), .C(n842) );
  BUFFD0 U724 ( .I(n842), .Z(n843) );
  CKBD0 U725 ( .CLK(n843), .C(n844) );
  CKBD0 U726 ( .CLK(n844), .C(n845) );
  CKBD0 U727 ( .CLK(n845), .C(n846) );
  CKBD0 U728 ( .CLK(n846), .C(n847) );
  CKBD0 U729 ( .CLK(n847), .C(n848) );
  CKBD0 U730 ( .CLK(n848), .C(n849) );
  CKBD0 U731 ( .CLK(n849), .C(n850) );
  CKBD0 U732 ( .CLK(n850), .C(n851) );
  CKBD0 U733 ( .CLK(n851), .C(n852) );
  CKBD0 U734 ( .CLK(n852), .C(n853) );
  BUFFD0 U735 ( .I(n853), .Z(n854) );
  CKBD0 U736 ( .CLK(n854), .C(n855) );
  CKBD0 U737 ( .CLK(n855), .C(n856) );
  CKBD0 U738 ( .CLK(n856), .C(n857) );
  CKBD0 U739 ( .CLK(n857), .C(n858) );
  CKBD0 U740 ( .CLK(n858), .C(n859) );
  CKBD0 U741 ( .CLK(n859), .C(n860) );
  CKBD0 U742 ( .CLK(n860), .C(n861) );
  CKBD0 U743 ( .CLK(n861), .C(n862) );
  CKBD0 U744 ( .CLK(n862), .C(n863) );
  BUFFD0 U745 ( .I(n863), .Z(n864) );
  CKBD0 U746 ( .CLK(n864), .C(n865) );
  CKBD0 U747 ( .CLK(n865), .C(n866) );
  CKBD0 U748 ( .CLK(n866), .C(n867) );
  CKBD0 U749 ( .CLK(n867), .C(n868) );
  CKBD0 U750 ( .CLK(n868), .C(n869) );
  CKBD0 U751 ( .CLK(n869), .C(n870) );
  CKBD0 U752 ( .CLK(n870), .C(n871) );
  CKBD0 U753 ( .CLK(n871), .C(n872) );
  CKBD0 U754 ( .CLK(n872), .C(n873) );
  CKBD0 U755 ( .CLK(n873), .C(n874) );
  BUFFD0 U756 ( .I(n874), .Z(n875) );
  CKBD0 U757 ( .CLK(n875), .C(n876) );
  CKBD0 U758 ( .CLK(n876), .C(n877) );
  CKBD0 U759 ( .CLK(n877), .C(n878) );
  CKBD0 U760 ( .CLK(n878), .C(n879) );
  CKBD0 U761 ( .CLK(n879), .C(n880) );
  CKBD0 U762 ( .CLK(n880), .C(n881) );
  CKBD0 U763 ( .CLK(n881), .C(n882) );
  CKBD0 U764 ( .CLK(n882), .C(n883) );
  CKBD0 U765 ( .CLK(n883), .C(n884) );
  CKBD0 U766 ( .CLK(n884), .C(n885) );
  BUFFD0 U767 ( .I(n885), .Z(n886) );
  CKBD0 U768 ( .CLK(n886), .C(n887) );
  CKBD0 U769 ( .CLK(n887), .C(n888) );
  CKBD0 U770 ( .CLK(n888), .C(n889) );
  CKBD0 U771 ( .CLK(n889), .C(n890) );
  CKBD0 U772 ( .CLK(n890), .C(n891) );
  CKBD0 U773 ( .CLK(n891), .C(n892) );
  CKBD0 U774 ( .CLK(n892), .C(n893) );
  CKBD0 U775 ( .CLK(n893), .C(n894) );
  CKBD0 U776 ( .CLK(n894), .C(n895) );
  CKBD0 U777 ( .CLK(n895), .C(n896) );
  BUFFD0 U778 ( .I(n896), .Z(n897) );
  CKBD0 U779 ( .CLK(n897), .C(n898) );
  CKBD0 U780 ( .CLK(n898), .C(n899) );
  CKBD0 U781 ( .CLK(n899), .C(n900) );
  CKBD0 U782 ( .CLK(n900), .C(n901) );
  CKBD0 U783 ( .CLK(n901), .C(n902) );
  CKBD0 U784 ( .CLK(n902), .C(n903) );
  CKBD0 U785 ( .CLK(n903), .C(n904) );
  CKBD0 U786 ( .CLK(n904), .C(n905) );
  CKBD0 U787 ( .CLK(n905), .C(n906) );
  CKBD0 U788 ( .CLK(n906), .C(n907) );
  BUFFD0 U789 ( .I(n907), .Z(n908) );
  CKBD0 U790 ( .CLK(n908), .C(n909) );
  CKBD0 U791 ( .CLK(n909), .C(n910) );
  CKBD0 U792 ( .CLK(n910), .C(n911) );
  CKBD0 U793 ( .CLK(n911), .C(n912) );
  CKBD0 U794 ( .CLK(n912), .C(n913) );
  CKBD0 U795 ( .CLK(n913), .C(n914) );
  CKBD0 U796 ( .CLK(n914), .C(n915) );
  CKBD0 U797 ( .CLK(n915), .C(n916) );
  BUFFD0 U798 ( .I(n9017), .Z(n917) );
  CKBD0 U799 ( .CLK(FrameSR[7]), .C(n918) );
  BUFFD0 U800 ( .I(n918), .Z(n919) );
  BUFFD0 U801 ( .I(n6915), .Z(n920) );
  CKBD0 U802 ( .CLK(FrameSR[8]), .C(n921) );
  BUFFD0 U803 ( .I(n6778), .Z(n922) );
  CKBD0 U804 ( .CLK(FrameSR[9]), .C(n923) );
  BUFFD0 U805 ( .I(n6641), .Z(n924) );
  CKBD0 U806 ( .CLK(FrameSR[10]), .C(n925) );
  BUFFD0 U807 ( .I(n6504), .Z(n926) );
  CKBD0 U808 ( .CLK(FrameSR[11]), .C(n927) );
  BUFFD0 U809 ( .I(n6367), .Z(n928) );
  CKBD0 U810 ( .CLK(FrameSR[12]), .C(n929) );
  BUFFD0 U811 ( .I(n6230), .Z(n930) );
  CKBD0 U812 ( .CLK(FrameSR[13]), .C(n931) );
  BUFFD0 U813 ( .I(n6093), .Z(n932) );
  CKBD0 U814 ( .CLK(FrameSR[14]), .C(n933) );
  BUFFD0 U815 ( .I(n9008), .Z(n934) );
  CKBD0 U816 ( .CLK(FrameSR[18]), .C(n935) );
  CKBD0 U817 ( .CLK(n935), .C(n936) );
  BUFFD0 U818 ( .I(n936), .Z(n937) );
  CKBD0 U819 ( .CLK(n937), .C(n938) );
  CKBD0 U820 ( .CLK(n938), .C(n939) );
  CKBD0 U821 ( .CLK(n939), .C(n940) );
  CKBD0 U822 ( .CLK(n940), .C(n941) );
  CKBD0 U823 ( .CLK(n941), .C(n942) );
  CKBD0 U824 ( .CLK(n942), .C(n943) );
  CKBD0 U825 ( .CLK(n943), .C(n944) );
  CKBD0 U826 ( .CLK(n944), .C(n945) );
  CKBD0 U827 ( .CLK(n945), .C(n946) );
  CKBD0 U828 ( .CLK(n946), .C(n947) );
  BUFFD0 U829 ( .I(n947), .Z(n948) );
  CKBD0 U830 ( .CLK(n948), .C(n949) );
  CKBD0 U831 ( .CLK(n949), .C(n950) );
  CKBD0 U832 ( .CLK(n950), .C(n951) );
  CKBD0 U833 ( .CLK(n951), .C(n952) );
  CKBD0 U834 ( .CLK(n952), .C(n953) );
  CKBD0 U835 ( .CLK(n953), .C(n954) );
  CKBD0 U836 ( .CLK(n954), .C(n955) );
  CKBD0 U837 ( .CLK(n955), .C(n956) );
  CKBD0 U838 ( .CLK(n956), .C(n957) );
  BUFFD0 U839 ( .I(n957), .Z(n958) );
  CKBD0 U840 ( .CLK(n958), .C(n959) );
  CKBD0 U841 ( .CLK(n959), .C(n960) );
  CKBD0 U842 ( .CLK(n960), .C(n961) );
  CKBD0 U843 ( .CLK(n961), .C(n962) );
  CKBD0 U844 ( .CLK(n962), .C(n963) );
  CKBD0 U845 ( .CLK(n963), .C(n964) );
  CKBD0 U846 ( .CLK(n964), .C(n965) );
  CKBD0 U847 ( .CLK(n965), .C(n966) );
  CKBD0 U848 ( .CLK(n966), .C(n967) );
  CKBD0 U849 ( .CLK(n967), .C(n968) );
  BUFFD0 U850 ( .I(n968), .Z(n969) );
  CKBD0 U851 ( .CLK(n969), .C(n970) );
  CKBD0 U852 ( .CLK(n970), .C(n971) );
  CKBD0 U853 ( .CLK(n971), .C(n972) );
  CKBD0 U854 ( .CLK(n972), .C(n973) );
  CKBD0 U855 ( .CLK(n973), .C(n974) );
  CKBD0 U856 ( .CLK(n974), .C(n975) );
  CKBD0 U857 ( .CLK(n975), .C(n976) );
  CKBD0 U858 ( .CLK(n976), .C(n977) );
  CKBD0 U859 ( .CLK(n977), .C(n978) );
  CKBD0 U860 ( .CLK(n978), .C(n979) );
  BUFFD0 U861 ( .I(n979), .Z(n980) );
  CKBD0 U862 ( .CLK(n980), .C(n981) );
  CKBD0 U863 ( .CLK(n981), .C(n982) );
  CKBD0 U864 ( .CLK(n982), .C(n983) );
  CKBD0 U865 ( .CLK(n983), .C(n984) );
  CKBD0 U866 ( .CLK(n984), .C(n985) );
  CKBD0 U867 ( .CLK(n985), .C(n986) );
  CKBD0 U868 ( .CLK(n986), .C(n987) );
  CKBD0 U869 ( .CLK(n987), .C(n988) );
  CKBD0 U870 ( .CLK(n988), .C(n989) );
  CKBD0 U871 ( .CLK(n989), .C(n990) );
  BUFFD0 U872 ( .I(n990), .Z(n991) );
  CKBD0 U873 ( .CLK(n991), .C(n992) );
  CKBD0 U874 ( .CLK(n992), .C(n993) );
  CKBD0 U875 ( .CLK(n993), .C(n994) );
  CKBD0 U876 ( .CLK(n994), .C(n995) );
  CKBD0 U877 ( .CLK(n995), .C(n996) );
  CKBD0 U878 ( .CLK(n996), .C(n997) );
  CKBD0 U879 ( .CLK(n997), .C(n998) );
  CKBD0 U880 ( .CLK(n998), .C(n999) );
  CKBD0 U881 ( .CLK(n999), .C(n1000) );
  CKBD0 U882 ( .CLK(n1000), .C(n1001) );
  BUFFD0 U883 ( .I(n1001), .Z(n1002) );
  CKBD0 U884 ( .CLK(n1002), .C(n1003) );
  CKBD0 U885 ( .CLK(n1003), .C(n1004) );
  CKBD0 U886 ( .CLK(n1004), .C(n1005) );
  CKBD0 U887 ( .CLK(n1005), .C(n1006) );
  CKBD0 U888 ( .CLK(n1006), .C(n1007) );
  CKBD0 U889 ( .CLK(n1007), .C(n1008) );
  CKBD0 U890 ( .CLK(n1008), .C(n1009) );
  CKBD0 U891 ( .CLK(n1009), .C(n1010) );
  CKBD0 U892 ( .CLK(n1010), .C(n1011) );
  CKBD0 U893 ( .CLK(n1011), .C(n1012) );
  BUFFD0 U894 ( .I(n1012), .Z(n1013) );
  CKBD0 U895 ( .CLK(n1013), .C(n1014) );
  CKBD0 U896 ( .CLK(n1014), .C(n1015) );
  CKBD0 U897 ( .CLK(n1015), .C(n1016) );
  CKBD0 U898 ( .CLK(n1016), .C(n1017) );
  CKBD0 U899 ( .CLK(n1017), .C(n1018) );
  CKBD0 U900 ( .CLK(n1018), .C(n1019) );
  CKBD0 U901 ( .CLK(n1019), .C(n1020) );
  CKBD0 U902 ( .CLK(n1020), .C(n1021) );
  CKBD0 U903 ( .CLK(n1021), .C(n1022) );
  CKBD0 U904 ( .CLK(n1022), .C(n1023) );
  BUFFD0 U905 ( .I(n1023), .Z(n1024) );
  CKBD0 U906 ( .CLK(n1024), .C(n1025) );
  CKBD0 U907 ( .CLK(n1025), .C(n1026) );
  CKBD0 U908 ( .CLK(n1026), .C(n1027) );
  CKBD0 U909 ( .CLK(n1027), .C(n1028) );
  CKBD0 U910 ( .CLK(n1028), .C(n1029) );
  CKBD0 U911 ( .CLK(n1029), .C(n1030) );
  BUFFD0 U912 ( .I(n8970), .Z(n1031) );
  CKBD0 U913 ( .CLK(FrameSR[23]), .C(n1032) );
  BUFFD0 U914 ( .I(n1032), .Z(n1033) );
  CKBD0 U915 ( .CLK(n1033), .C(n1034) );
  CKBD0 U916 ( .CLK(n1034), .C(n1035) );
  CKBD0 U917 ( .CLK(n1035), .C(n1036) );
  CKBD0 U918 ( .CLK(n1036), .C(n1037) );
  CKBD0 U919 ( .CLK(n1037), .C(n1038) );
  CKBD0 U920 ( .CLK(n1038), .C(n1039) );
  CKBD0 U921 ( .CLK(n1039), .C(n1040) );
  CKBD0 U922 ( .CLK(n1040), .C(n1041) );
  CKBD0 U923 ( .CLK(n1041), .C(n1042) );
  CKBD0 U924 ( .CLK(n1042), .C(n1043) );
  BUFFD0 U925 ( .I(n1043), .Z(n1044) );
  CKBD0 U926 ( .CLK(n1044), .C(n1045) );
  CKBD0 U927 ( .CLK(n1045), .C(n1046) );
  CKBD0 U928 ( .CLK(n1046), .C(n1047) );
  CKBD0 U929 ( .CLK(n1047), .C(n1048) );
  CKBD0 U930 ( .CLK(n1048), .C(n1049) );
  CKBD0 U931 ( .CLK(n1049), .C(n1050) );
  CKBD0 U932 ( .CLK(n1050), .C(n1051) );
  CKBD0 U933 ( .CLK(n1051), .C(n1052) );
  CKBD0 U934 ( .CLK(n1052), .C(n1053) );
  CKBD0 U935 ( .CLK(n1053), .C(n1054) );
  BUFFD0 U936 ( .I(n1054), .Z(n1055) );
  CKBD0 U937 ( .CLK(n1055), .C(n1056) );
  CKBD0 U938 ( .CLK(n1056), .C(n1057) );
  CKBD0 U939 ( .CLK(n1057), .C(n1058) );
  CKBD0 U940 ( .CLK(n1058), .C(n1059) );
  CKBD0 U941 ( .CLK(n1059), .C(n1060) );
  CKBD0 U942 ( .CLK(n1060), .C(n1061) );
  CKBD0 U943 ( .CLK(n1061), .C(n1062) );
  CKBD0 U944 ( .CLK(n1062), .C(n1063) );
  CKBD0 U945 ( .CLK(n1063), .C(n1064) );
  CKBD0 U946 ( .CLK(n1064), .C(n1065) );
  BUFFD0 U947 ( .I(n1065), .Z(n1066) );
  CKBD0 U948 ( .CLK(n1066), .C(n1067) );
  CKBD0 U949 ( .CLK(n1067), .C(n1068) );
  CKBD0 U950 ( .CLK(n1068), .C(n1069) );
  CKBD0 U951 ( .CLK(n1069), .C(n1070) );
  CKBD0 U952 ( .CLK(n1070), .C(n1071) );
  CKBD0 U953 ( .CLK(n1071), .C(n1072) );
  CKBD0 U954 ( .CLK(n1072), .C(n1073) );
  CKBD0 U955 ( .CLK(n1073), .C(n1074) );
  CKBD0 U956 ( .CLK(n1074), .C(n1075) );
  BUFFD0 U957 ( .I(n1075), .Z(n1076) );
  CKBD0 U958 ( .CLK(n1076), .C(n1077) );
  CKBD0 U959 ( .CLK(n1077), .C(n1078) );
  CKBD0 U960 ( .CLK(n1078), .C(n1079) );
  CKBD0 U961 ( .CLK(n1079), .C(n1080) );
  CKBD0 U962 ( .CLK(n1080), .C(n1081) );
  CKBD0 U963 ( .CLK(n1081), .C(n1082) );
  CKBD0 U964 ( .CLK(n1082), .C(n1083) );
  CKBD0 U965 ( .CLK(n1083), .C(n1084) );
  CKBD0 U966 ( .CLK(n1084), .C(n1085) );
  CKBD0 U967 ( .CLK(n1085), .C(n1086) );
  BUFFD0 U968 ( .I(n1086), .Z(n1087) );
  CKBD0 U969 ( .CLK(n1087), .C(n1088) );
  CKBD0 U970 ( .CLK(n1088), .C(n1089) );
  CKBD0 U971 ( .CLK(n1089), .C(n1090) );
  CKBD0 U972 ( .CLK(n1090), .C(n1091) );
  CKBD0 U973 ( .CLK(n1091), .C(n1092) );
  CKBD0 U974 ( .CLK(n1092), .C(n1093) );
  CKBD0 U975 ( .CLK(n1093), .C(n1094) );
  CKBD0 U976 ( .CLK(n1094), .C(n1095) );
  CKBD0 U977 ( .CLK(n1095), .C(n1096) );
  CKBD0 U978 ( .CLK(n1096), .C(n1097) );
  BUFFD0 U979 ( .I(n1097), .Z(n1098) );
  CKBD0 U980 ( .CLK(n1098), .C(n1099) );
  CKBD0 U981 ( .CLK(n1099), .C(n1100) );
  CKBD0 U982 ( .CLK(n1100), .C(n1101) );
  CKBD0 U983 ( .CLK(n1101), .C(n1102) );
  CKBD0 U984 ( .CLK(n1102), .C(n1103) );
  CKBD0 U985 ( .CLK(n1103), .C(n1104) );
  CKBD0 U986 ( .CLK(n1104), .C(n1105) );
  CKBD0 U987 ( .CLK(n1105), .C(n1106) );
  CKBD0 U988 ( .CLK(n1106), .C(n1107) );
  CKBD0 U989 ( .CLK(n1107), .C(n1108) );
  BUFFD0 U990 ( .I(n1108), .Z(n1109) );
  CKBD0 U991 ( .CLK(n1109), .C(n1110) );
  CKBD0 U992 ( .CLK(n1110), .C(n1111) );
  CKBD0 U993 ( .CLK(n1111), .C(n1112) );
  CKBD0 U994 ( .CLK(n1112), .C(n1113) );
  CKBD0 U995 ( .CLK(n1113), .C(n1114) );
  CKBD0 U996 ( .CLK(n1114), .C(n1115) );
  CKBD0 U997 ( .CLK(n1115), .C(n1116) );
  CKBD0 U998 ( .CLK(n1116), .C(n1117) );
  CKBD0 U999 ( .CLK(n1117), .C(n1118) );
  CKBD0 U1000 ( .CLK(n1118), .C(n1119) );
  BUFFD0 U1001 ( .I(n1119), .Z(n1120) );
  CKBD0 U1002 ( .CLK(n1120), .C(n1121) );
  CKBD0 U1003 ( .CLK(n1121), .C(n1122) );
  CKBD0 U1004 ( .CLK(n1122), .C(n1123) );
  CKBD0 U1005 ( .CLK(n1123), .C(n1124) );
  CKBD0 U1006 ( .CLK(n1124), .C(n1125) );
  CKBD0 U1007 ( .CLK(n1125), .C(n1126) );
  CKBD0 U1008 ( .CLK(n1126), .C(n1127) );
  CKBD0 U1009 ( .CLK(n1127), .C(n1128) );
  BUFFD0 U1010 ( .I(n5820), .Z(n1129) );
  CKBD0 U1011 ( .CLK(FrameSR[24]), .C(n1130) );
  BUFFD0 U1012 ( .I(n5684), .Z(n1131) );
  CKBD0 U1013 ( .CLK(FrameSR[25]), .C(n1132) );
  BUFFD0 U1014 ( .I(n5548), .Z(n1133) );
  CKBD0 U1015 ( .CLK(FrameSR[26]), .C(n1134) );
  BUFFD0 U1016 ( .I(n5412), .Z(n1135) );
  CKBD0 U1017 ( .CLK(FrameSR[27]), .C(n1136) );
  BUFFD0 U1018 ( .I(n5276), .Z(n1137) );
  CKBD0 U1019 ( .CLK(FrameSR[28]), .C(n1138) );
  BUFFD0 U1020 ( .I(n5139), .Z(n1139) );
  CKBD0 U1021 ( .CLK(FrameSR[29]), .C(n1140) );
  BUFFD0 U1022 ( .I(n5003), .Z(n1141) );
  CKBD0 U1023 ( .CLK(FrameSR[30]), .C(n1142) );
  BUFFD0 U1024 ( .I(n8962), .Z(n1143) );
  CKBD0 U1025 ( .CLK(FrameSR[39]), .C(n1144) );
  BUFFD0 U1026 ( .I(n1144), .Z(n1145) );
  CKBD0 U1027 ( .CLK(n1145), .C(n1146) );
  CKBD0 U1028 ( .CLK(n1146), .C(n1147) );
  CKBD0 U1029 ( .CLK(n1147), .C(n1148) );
  CKBD0 U1030 ( .CLK(n1148), .C(n1149) );
  CKBD0 U1031 ( .CLK(n1149), .C(n1150) );
  CKBD0 U1032 ( .CLK(n1150), .C(n1151) );
  CKBD0 U1033 ( .CLK(n1151), .C(n1152) );
  CKBD0 U1034 ( .CLK(n1152), .C(n1153) );
  CKBD0 U1035 ( .CLK(n1153), .C(n1154) );
  BUFFD0 U1036 ( .I(n1154), .Z(n1155) );
  CKBD0 U1037 ( .CLK(n1155), .C(n1156) );
  CKBD0 U1038 ( .CLK(n1156), .C(n1157) );
  CKBD0 U1039 ( .CLK(n1157), .C(n1158) );
  CKBD0 U1040 ( .CLK(n1158), .C(n1159) );
  CKBD0 U1041 ( .CLK(n1159), .C(n1160) );
  CKBD0 U1042 ( .CLK(n1160), .C(n1161) );
  CKBD0 U1043 ( .CLK(n1161), .C(n1162) );
  CKBD0 U1044 ( .CLK(n1162), .C(n1163) );
  CKBD0 U1045 ( .CLK(n1163), .C(n1164) );
  CKBD0 U1046 ( .CLK(n1164), .C(n1165) );
  BUFFD0 U1047 ( .I(n1165), .Z(n1166) );
  CKBD0 U1048 ( .CLK(n1166), .C(n1167) );
  CKBD0 U1049 ( .CLK(n1167), .C(n1168) );
  CKBD0 U1050 ( .CLK(n1168), .C(n1169) );
  CKBD0 U1051 ( .CLK(n1169), .C(n1170) );
  CKBD0 U1052 ( .CLK(n1170), .C(n1171) );
  CKBD0 U1053 ( .CLK(n1171), .C(n1172) );
  CKBD0 U1054 ( .CLK(n1172), .C(n1173) );
  CKBD0 U1055 ( .CLK(n1173), .C(n1174) );
  CKBD0 U1056 ( .CLK(n1174), .C(n1175) );
  CKBD0 U1057 ( .CLK(n1175), .C(n1176) );
  BUFFD0 U1058 ( .I(n1176), .Z(n1177) );
  CKBD0 U1059 ( .CLK(n1177), .C(n1178) );
  CKBD0 U1060 ( .CLK(n1178), .C(n1179) );
  CKBD0 U1061 ( .CLK(n1179), .C(n1180) );
  CKBD0 U1062 ( .CLK(n1180), .C(n1181) );
  CKBD0 U1063 ( .CLK(n1181), .C(n1182) );
  CKBD0 U1064 ( .CLK(n1182), .C(n1183) );
  CKBD0 U1065 ( .CLK(n1183), .C(n1184) );
  CKBD0 U1066 ( .CLK(n1184), .C(n1185) );
  CKBD0 U1067 ( .CLK(n1185), .C(n1186) );
  CKBD0 U1068 ( .CLK(n1186), .C(n1187) );
  BUFFD0 U1069 ( .I(n1187), .Z(n1188) );
  CKBD0 U1070 ( .CLK(n1188), .C(n1189) );
  CKBD0 U1071 ( .CLK(n1189), .C(n1190) );
  CKBD0 U1072 ( .CLK(n1190), .C(n1191) );
  CKBD0 U1073 ( .CLK(n1191), .C(n1192) );
  CKBD0 U1074 ( .CLK(n1192), .C(n1193) );
  CKBD0 U1075 ( .CLK(n1193), .C(n1194) );
  CKBD0 U1076 ( .CLK(n1194), .C(n1195) );
  CKBD0 U1077 ( .CLK(n1195), .C(n1196) );
  CKBD0 U1078 ( .CLK(n1196), .C(n1197) );
  CKBD0 U1079 ( .CLK(n1197), .C(n1198) );
  BUFFD0 U1080 ( .I(n1198), .Z(n1199) );
  CKBD0 U1081 ( .CLK(n1199), .C(n1200) );
  CKBD0 U1082 ( .CLK(n1200), .C(n1201) );
  CKBD0 U1083 ( .CLK(n1201), .C(n1202) );
  CKBD0 U1084 ( .CLK(n1202), .C(n1203) );
  CKBD0 U1085 ( .CLK(n1203), .C(n1204) );
  CKBD0 U1086 ( .CLK(n1204), .C(n1205) );
  CKBD0 U1087 ( .CLK(n1205), .C(n1206) );
  CKBD0 U1088 ( .CLK(n1206), .C(n1207) );
  CKBD0 U1089 ( .CLK(n1207), .C(n1208) );
  CKBD0 U1090 ( .CLK(n1208), .C(n1209) );
  BUFFD0 U1091 ( .I(n1209), .Z(n1210) );
  CKBD0 U1092 ( .CLK(n1210), .C(n1211) );
  CKBD0 U1093 ( .CLK(n1211), .C(n1212) );
  CKBD0 U1094 ( .CLK(n1212), .C(n1213) );
  CKBD0 U1095 ( .CLK(n1213), .C(n1214) );
  CKBD0 U1096 ( .CLK(n1214), .C(n1215) );
  CKBD0 U1097 ( .CLK(n1215), .C(n1216) );
  CKBD0 U1098 ( .CLK(n1216), .C(n1217) );
  CKBD0 U1099 ( .CLK(n1217), .C(n1218) );
  CKBD0 U1100 ( .CLK(n1218), .C(n1219) );
  CKBD0 U1101 ( .CLK(n1219), .C(n1220) );
  BUFFD0 U1102 ( .I(n1220), .Z(n1221) );
  CKBD0 U1103 ( .CLK(n1221), .C(n1222) );
  CKBD0 U1104 ( .CLK(n1222), .C(n1223) );
  CKBD0 U1105 ( .CLK(n1223), .C(n1224) );
  CKBD0 U1106 ( .CLK(n1224), .C(n1225) );
  CKBD0 U1107 ( .CLK(n1225), .C(n1226) );
  CKBD0 U1108 ( .CLK(n1226), .C(n1227) );
  CKBD0 U1109 ( .CLK(n1227), .C(n1228) );
  CKBD0 U1110 ( .CLK(n1228), .C(n1229) );
  CKBD0 U1111 ( .CLK(n1229), .C(n1230) );
  BUFFD0 U1112 ( .I(n1230), .Z(n1231) );
  CKBD0 U1113 ( .CLK(n1231), .C(n1232) );
  CKBD0 U1114 ( .CLK(n1232), .C(n1233) );
  CKBD0 U1115 ( .CLK(n1233), .C(n1234) );
  CKBD0 U1116 ( .CLK(n1234), .C(n1235) );
  CKBD0 U1117 ( .CLK(n1235), .C(n1236) );
  CKBD0 U1118 ( .CLK(n1236), .C(n1237) );
  CKBD0 U1119 ( .CLK(n1237), .C(n1238) );
  CKBD0 U1120 ( .CLK(n1238), .C(n1239) );
  CKBD0 U1121 ( .CLK(n1239), .C(n1240) );
  BUFFD0 U1122 ( .I(n4731), .Z(n1241) );
  CKBD0 U1123 ( .CLK(FrameSR[40]), .C(n1242) );
  BUFFD0 U1124 ( .I(n4595), .Z(n1243) );
  CKBD0 U1125 ( .CLK(FrameSR[41]), .C(n1244) );
  BUFFD0 U1126 ( .I(n4459), .Z(n1245) );
  CKBD0 U1127 ( .CLK(FrameSR[42]), .C(n1246) );
  BUFFD0 U1128 ( .I(n4323), .Z(n1247) );
  CKBD0 U1129 ( .CLK(FrameSR[43]), .C(n1248) );
  BUFFD0 U1130 ( .I(n4186), .Z(n1249) );
  CKBD0 U1131 ( .CLK(FrameSR[44]), .C(n1250) );
  BUFFD0 U1132 ( .I(n4050), .Z(n1251) );
  CKBD0 U1133 ( .CLK(FrameSR[45]), .C(n1252) );
  BUFFD0 U1134 ( .I(n3914), .Z(n1253) );
  CKBD0 U1135 ( .CLK(FrameSR[46]), .C(n1254) );
  BUFFD0 U1136 ( .I(n8960), .Z(n1255) );
  CKBD0 U1137 ( .CLK(FrameSR[55]), .C(n1256) );
  BUFFD0 U1138 ( .I(n1256), .Z(n1257) );
  CKBD0 U1139 ( .CLK(n1257), .C(n1258) );
  CKBD0 U1140 ( .CLK(n1258), .C(n1259) );
  CKBD0 U1141 ( .CLK(n1259), .C(n1260) );
  CKBD0 U1142 ( .CLK(n1260), .C(n1261) );
  CKBD0 U1143 ( .CLK(n1261), .C(n1262) );
  CKBD0 U1144 ( .CLK(n1262), .C(n1263) );
  CKBD0 U1145 ( .CLK(n1263), .C(n1264) );
  CKBD0 U1146 ( .CLK(n1264), .C(n1265) );
  CKBD0 U1147 ( .CLK(n1265), .C(n1266) );
  BUFFD0 U1148 ( .I(n1266), .Z(n1267) );
  CKBD0 U1149 ( .CLK(n1267), .C(n1268) );
  CKBD0 U1150 ( .CLK(n1268), .C(n1269) );
  CKBD0 U1151 ( .CLK(n1269), .C(n1270) );
  CKBD0 U1152 ( .CLK(n1270), .C(n1271) );
  CKBD0 U1153 ( .CLK(n1271), .C(n1272) );
  CKBD0 U1154 ( .CLK(n1272), .C(n1273) );
  CKBD0 U1155 ( .CLK(n1273), .C(n1274) );
  CKBD0 U1156 ( .CLK(n1274), .C(n1275) );
  CKBD0 U1157 ( .CLK(n1275), .C(n1276) );
  CKBD0 U1158 ( .CLK(n1276), .C(n1277) );
  BUFFD0 U1159 ( .I(n1277), .Z(n1278) );
  CKBD0 U1160 ( .CLK(n1278), .C(n1279) );
  CKBD0 U1161 ( .CLK(n1279), .C(n1280) );
  CKBD0 U1162 ( .CLK(n1280), .C(n1281) );
  CKBD0 U1163 ( .CLK(n1281), .C(n1282) );
  CKBD0 U1164 ( .CLK(n1282), .C(n1283) );
  CKBD0 U1165 ( .CLK(n1283), .C(n1284) );
  CKBD0 U1166 ( .CLK(n1284), .C(n1285) );
  CKBD0 U1167 ( .CLK(n1285), .C(n1286) );
  CKBD0 U1168 ( .CLK(n1286), .C(n1287) );
  CKBD0 U1169 ( .CLK(n1287), .C(n1288) );
  BUFFD0 U1170 ( .I(n1288), .Z(n1289) );
  CKBD0 U1171 ( .CLK(n1289), .C(n1290) );
  CKBD0 U1172 ( .CLK(n1290), .C(n1291) );
  CKBD0 U1173 ( .CLK(n1291), .C(n1292) );
  CKBD0 U1174 ( .CLK(n1292), .C(n1293) );
  CKBD0 U1175 ( .CLK(n1293), .C(n1294) );
  CKBD0 U1176 ( .CLK(n1294), .C(n1295) );
  CKBD0 U1177 ( .CLK(n1295), .C(n1296) );
  CKBD0 U1178 ( .CLK(n1296), .C(n1297) );
  CKBD0 U1179 ( .CLK(n1297), .C(n1298) );
  CKBD0 U1180 ( .CLK(n1298), .C(n1299) );
  BUFFD0 U1181 ( .I(n1299), .Z(n1300) );
  CKBD0 U1182 ( .CLK(n1300), .C(n1301) );
  CKBD0 U1183 ( .CLK(n1301), .C(n1302) );
  CKBD0 U1184 ( .CLK(n1302), .C(n1303) );
  CKBD0 U1185 ( .CLK(n1303), .C(n1304) );
  CKBD0 U1186 ( .CLK(n1304), .C(n1305) );
  CKBD0 U1187 ( .CLK(n1305), .C(n1306) );
  CKBD0 U1188 ( .CLK(n1306), .C(n1307) );
  CKBD0 U1189 ( .CLK(n1307), .C(n1308) );
  CKBD0 U1190 ( .CLK(n1308), .C(n1309) );
  CKBD0 U1191 ( .CLK(n1309), .C(n1310) );
  BUFFD0 U1192 ( .I(n1310), .Z(n1311) );
  CKBD0 U1193 ( .CLK(n1311), .C(n1312) );
  CKBD0 U1194 ( .CLK(n1312), .C(n1313) );
  CKBD0 U1195 ( .CLK(n1313), .C(n1314) );
  CKBD0 U1196 ( .CLK(n1314), .C(n1315) );
  CKBD0 U1197 ( .CLK(n1315), .C(n1316) );
  CKBD0 U1198 ( .CLK(n1316), .C(n1317) );
  CKBD0 U1199 ( .CLK(n1317), .C(n1318) );
  CKBD0 U1200 ( .CLK(n1318), .C(n1319) );
  CKBD0 U1201 ( .CLK(n1319), .C(n1320) );
  CKBD0 U1202 ( .CLK(n1320), .C(n1321) );
  BUFFD0 U1203 ( .I(n1321), .Z(n1322) );
  CKBD0 U1204 ( .CLK(n1322), .C(n1323) );
  CKBD0 U1205 ( .CLK(n1323), .C(n1324) );
  CKBD0 U1206 ( .CLK(n1324), .C(n1325) );
  CKBD0 U1207 ( .CLK(n1325), .C(n1326) );
  CKBD0 U1208 ( .CLK(n1326), .C(n1327) );
  CKBD0 U1209 ( .CLK(n1327), .C(n1328) );
  CKBD0 U1210 ( .CLK(n1328), .C(n1329) );
  CKBD0 U1211 ( .CLK(n1329), .C(n1330) );
  CKBD0 U1212 ( .CLK(n1330), .C(n1331) );
  CKBD0 U1213 ( .CLK(n1331), .C(n1332) );
  BUFFD0 U1214 ( .I(n1332), .Z(n1333) );
  CKBD0 U1215 ( .CLK(n1333), .C(n1334) );
  CKBD0 U1216 ( .CLK(n1334), .C(n1335) );
  CKBD0 U1217 ( .CLK(n1335), .C(n1336) );
  CKBD0 U1218 ( .CLK(n1336), .C(n1337) );
  CKBD0 U1219 ( .CLK(n1337), .C(n1338) );
  CKBD0 U1220 ( .CLK(n1338), .C(n1339) );
  CKBD0 U1221 ( .CLK(n1339), .C(n1340) );
  CKBD0 U1222 ( .CLK(n1340), .C(n1341) );
  CKBD0 U1223 ( .CLK(n1341), .C(n1342) );
  BUFFD0 U1224 ( .I(n1342), .Z(n1343) );
  CKBD0 U1225 ( .CLK(n1343), .C(n1344) );
  CKBD0 U1226 ( .CLK(n1344), .C(n1345) );
  CKBD0 U1227 ( .CLK(n1345), .C(n1346) );
  CKBD0 U1228 ( .CLK(n1346), .C(n1347) );
  CKBD0 U1229 ( .CLK(n1347), .C(n1348) );
  CKBD0 U1230 ( .CLK(n1348), .C(n1349) );
  CKBD0 U1231 ( .CLK(n1349), .C(n1350) );
  CKBD0 U1232 ( .CLK(n1350), .C(n1351) );
  CKBD0 U1233 ( .CLK(n1351), .C(n1352) );
  BUFFD0 U1234 ( .I(n3642), .Z(n1353) );
  CKBD0 U1235 ( .CLK(FrameSR[56]), .C(n1354) );
  BUFFD0 U1236 ( .I(n3506), .Z(n1355) );
  CKBD0 U1237 ( .CLK(FrameSR[57]), .C(n1356) );
  BUFFD0 U1238 ( .I(n3370), .Z(n1357) );
  CKBD0 U1239 ( .CLK(FrameSR[58]), .C(n1358) );
  BUFFD0 U1240 ( .I(n3234), .Z(n1359) );
  CKBD0 U1241 ( .CLK(FrameSR[59]), .C(n1360) );
  BUFFD0 U1242 ( .I(n3098), .Z(n1361) );
  CKBD0 U1243 ( .CLK(FrameSR[60]), .C(n1362) );
  BUFFD0 U1244 ( .I(n2962), .Z(n1363) );
  CKBD0 U1245 ( .CLK(FrameSR[61]), .C(n1364) );
  BUFFD0 U1246 ( .I(n9016), .Z(n1365) );
  CKBD0 U1247 ( .CLK(FrameSR[3]), .C(n1366) );
  BUFFD0 U1248 ( .I(n8982), .Z(n1367) );
  CKBD0 U1249 ( .CLK(FrameSR[19]), .C(n1368) );
  CKBD0 U1250 ( .CLK(n1368), .C(n1369) );
  BUFFD0 U1251 ( .I(n1369), .Z(n1370) );
  CKBD0 U1252 ( .CLK(n1370), .C(n1371) );
  CKBD0 U1253 ( .CLK(n1371), .C(n1372) );
  CKBD0 U1254 ( .CLK(n1372), .C(n1373) );
  CKBD0 U1255 ( .CLK(n1373), .C(n1374) );
  CKBD0 U1256 ( .CLK(n1374), .C(n1375) );
  CKBD0 U1257 ( .CLK(n1375), .C(n1376) );
  CKBD0 U1258 ( .CLK(n1376), .C(n1377) );
  CKBD0 U1259 ( .CLK(n1377), .C(n1378) );
  CKBD0 U1260 ( .CLK(n1378), .C(n1379) );
  CKBD0 U1261 ( .CLK(n1379), .C(n1380) );
  BUFFD0 U1262 ( .I(n1380), .Z(n1381) );
  CKBD0 U1263 ( .CLK(n1381), .C(n1382) );
  CKBD0 U1264 ( .CLK(n1382), .C(n1383) );
  CKBD0 U1265 ( .CLK(n1383), .C(n1384) );
  CKBD0 U1266 ( .CLK(n1384), .C(n1385) );
  CKBD0 U1267 ( .CLK(n1385), .C(n1386) );
  CKBD0 U1268 ( .CLK(n1386), .C(n1387) );
  CKBD0 U1269 ( .CLK(n1387), .C(n1388) );
  CKBD0 U1270 ( .CLK(n1388), .C(n1389) );
  CKBD0 U1271 ( .CLK(n1389), .C(n1390) );
  CKBD0 U1272 ( .CLK(n1390), .C(n1391) );
  BUFFD0 U1273 ( .I(n1391), .Z(n1392) );
  CKBD0 U1274 ( .CLK(n1392), .C(n1393) );
  CKBD0 U1275 ( .CLK(n1393), .C(n1394) );
  CKBD0 U1276 ( .CLK(n1394), .C(n1395) );
  CKBD0 U1277 ( .CLK(n1395), .C(n1396) );
  CKBD0 U1278 ( .CLK(n1396), .C(n1397) );
  CKBD0 U1279 ( .CLK(n1397), .C(n1398) );
  CKBD0 U1280 ( .CLK(n1398), .C(n1399) );
  CKBD0 U1281 ( .CLK(n1399), .C(n1400) );
  CKBD0 U1282 ( .CLK(n1400), .C(n1401) );
  CKBD0 U1283 ( .CLK(n1401), .C(n1402) );
  BUFFD0 U1284 ( .I(n1402), .Z(n1403) );
  CKBD0 U1285 ( .CLK(n1403), .C(n1404) );
  CKBD0 U1286 ( .CLK(n1404), .C(n1405) );
  CKBD0 U1287 ( .CLK(n1405), .C(n1406) );
  CKBD0 U1288 ( .CLK(n1406), .C(n1407) );
  CKBD0 U1289 ( .CLK(n1407), .C(n1408) );
  CKBD0 U1290 ( .CLK(n1408), .C(n1409) );
  CKBD0 U1291 ( .CLK(n1409), .C(n1410) );
  CKBD0 U1292 ( .CLK(n1410), .C(n1411) );
  CKBD0 U1293 ( .CLK(n1411), .C(n1412) );
  CKBD0 U1294 ( .CLK(n1412), .C(n1413) );
  BUFFD0 U1295 ( .I(n1413), .Z(n1414) );
  CKBD0 U1296 ( .CLK(n1414), .C(n1415) );
  CKBD0 U1297 ( .CLK(n1415), .C(n1416) );
  CKBD0 U1298 ( .CLK(n1416), .C(n1417) );
  CKBD0 U1299 ( .CLK(n1417), .C(n1418) );
  CKBD0 U1300 ( .CLK(n1418), .C(n1419) );
  CKBD0 U1301 ( .CLK(n1419), .C(n1420) );
  CKBD0 U1302 ( .CLK(n1420), .C(n1421) );
  CKBD0 U1303 ( .CLK(n1421), .C(n1422) );
  CKBD0 U1304 ( .CLK(n1422), .C(n1423) );
  CKBD0 U1305 ( .CLK(n1423), .C(n1424) );
  BUFFD0 U1306 ( .I(n1424), .Z(n1425) );
  CKBD0 U1307 ( .CLK(n1425), .C(n1426) );
  CKBD0 U1308 ( .CLK(n1426), .C(n1427) );
  CKBD0 U1309 ( .CLK(n1427), .C(n1428) );
  CKBD0 U1310 ( .CLK(n1428), .C(n1429) );
  CKBD0 U1311 ( .CLK(n1429), .C(n1430) );
  CKBD0 U1312 ( .CLK(n1430), .C(n1431) );
  CKBD0 U1313 ( .CLK(n1431), .C(n1432) );
  CKBD0 U1314 ( .CLK(n1432), .C(n1433) );
  CKBD0 U1315 ( .CLK(n1433), .C(n1434) );
  CKBD0 U1316 ( .CLK(n1434), .C(n1435) );
  BUFFD0 U1317 ( .I(n1435), .Z(n1436) );
  CKBD0 U1318 ( .CLK(n1436), .C(n1437) );
  CKBD0 U1319 ( .CLK(n1437), .C(n1438) );
  CKBD0 U1320 ( .CLK(n1438), .C(n1439) );
  CKBD0 U1321 ( .CLK(n1439), .C(n1440) );
  CKBD0 U1322 ( .CLK(n1440), .C(n1441) );
  CKBD0 U1323 ( .CLK(n1441), .C(n1442) );
  CKBD0 U1324 ( .CLK(n1442), .C(n1443) );
  CKBD0 U1325 ( .CLK(n1443), .C(n1444) );
  CKBD0 U1326 ( .CLK(n1444), .C(n1445) );
  BUFFD0 U1327 ( .I(n1445), .Z(n1446) );
  CKBD0 U1328 ( .CLK(n1446), .C(n1447) );
  CKBD0 U1329 ( .CLK(n1447), .C(n1448) );
  CKBD0 U1330 ( .CLK(n1448), .C(n1449) );
  CKBD0 U1331 ( .CLK(n1449), .C(n1450) );
  CKBD0 U1332 ( .CLK(n1450), .C(n1451) );
  CKBD0 U1333 ( .CLK(n1451), .C(n1452) );
  CKBD0 U1334 ( .CLK(n1452), .C(n1453) );
  CKBD0 U1335 ( .CLK(n1453), .C(n1454) );
  CKBD0 U1336 ( .CLK(n1454), .C(n1455) );
  CKBD0 U1337 ( .CLK(n1455), .C(n1456) );
  BUFFD0 U1338 ( .I(n1456), .Z(n1457) );
  CKBD0 U1339 ( .CLK(n1457), .C(n1458) );
  CKBD0 U1340 ( .CLK(n1458), .C(n1459) );
  CKBD0 U1341 ( .CLK(n1459), .C(n1460) );
  CKBD0 U1342 ( .CLK(n1460), .C(n1461) );
  CKBD0 U1343 ( .CLK(n1461), .C(n1462) );
  CKBD0 U1344 ( .CLK(n1462), .C(n1463) );
  BUFFD0 U1345 ( .I(n8997), .Z(n1464) );
  CKBD0 U1346 ( .CLK(FrameSR[33]), .C(n1465) );
  CKBD0 U1347 ( .CLK(n1465), .C(n1466) );
  BUFFD0 U1348 ( .I(n1466), .Z(n1467) );
  CKBD0 U1349 ( .CLK(n1467), .C(n1468) );
  CKBD0 U1350 ( .CLK(n1468), .C(n1469) );
  CKBD0 U1351 ( .CLK(n1469), .C(n1470) );
  CKBD0 U1352 ( .CLK(n1470), .C(n1471) );
  CKBD0 U1353 ( .CLK(n1471), .C(n1472) );
  CKBD0 U1354 ( .CLK(n1472), .C(n1473) );
  CKBD0 U1355 ( .CLK(n1473), .C(n1474) );
  CKBD0 U1356 ( .CLK(n1474), .C(n1475) );
  CKBD0 U1357 ( .CLK(n1475), .C(n1476) );
  CKBD0 U1358 ( .CLK(n1476), .C(n1477) );
  BUFFD0 U1359 ( .I(n1477), .Z(n1478) );
  CKBD0 U1360 ( .CLK(n1478), .C(n1479) );
  CKBD0 U1361 ( .CLK(n1479), .C(n1480) );
  CKBD0 U1362 ( .CLK(n1480), .C(n1481) );
  CKBD0 U1363 ( .CLK(n1481), .C(n1482) );
  CKBD0 U1364 ( .CLK(n1482), .C(n1483) );
  CKBD0 U1365 ( .CLK(n1483), .C(n1484) );
  CKBD0 U1366 ( .CLK(n1484), .C(n1485) );
  CKBD0 U1367 ( .CLK(n1485), .C(n1486) );
  CKBD0 U1368 ( .CLK(n1486), .C(n1487) );
  BUFFD0 U1369 ( .I(n1487), .Z(n1488) );
  CKBD0 U1370 ( .CLK(n1488), .C(n1489) );
  CKBD0 U1371 ( .CLK(n1489), .C(n1490) );
  CKBD0 U1372 ( .CLK(n1490), .C(n1491) );
  CKBD0 U1373 ( .CLK(n1491), .C(n1492) );
  CKBD0 U1374 ( .CLK(n1492), .C(n1493) );
  CKBD0 U1375 ( .CLK(n1493), .C(n1494) );
  CKBD0 U1376 ( .CLK(n1494), .C(n1495) );
  CKBD0 U1377 ( .CLK(n1495), .C(n1496) );
  CKBD0 U1378 ( .CLK(n1496), .C(n1497) );
  CKBD0 U1379 ( .CLK(n1497), .C(n1498) );
  BUFFD0 U1380 ( .I(n1498), .Z(n1499) );
  CKBD0 U1381 ( .CLK(n1499), .C(n1500) );
  CKBD0 U1382 ( .CLK(n1500), .C(n1501) );
  CKBD0 U1383 ( .CLK(n1501), .C(n1502) );
  CKBD0 U1384 ( .CLK(n1502), .C(n1503) );
  CKBD0 U1385 ( .CLK(n1503), .C(n1504) );
  CKBD0 U1386 ( .CLK(n1504), .C(n1505) );
  CKBD0 U1387 ( .CLK(n1505), .C(n1506) );
  CKBD0 U1388 ( .CLK(n1506), .C(n1507) );
  CKBD0 U1389 ( .CLK(n1507), .C(n1508) );
  CKBD0 U1390 ( .CLK(n1508), .C(n1509) );
  BUFFD0 U1391 ( .I(n1509), .Z(n1510) );
  CKBD0 U1392 ( .CLK(n1510), .C(n1511) );
  CKBD0 U1393 ( .CLK(n1511), .C(n1512) );
  CKBD0 U1394 ( .CLK(n1512), .C(n1513) );
  CKBD0 U1395 ( .CLK(n1513), .C(n1514) );
  CKBD0 U1396 ( .CLK(n1514), .C(n1515) );
  CKBD0 U1397 ( .CLK(n1515), .C(n1516) );
  CKBD0 U1398 ( .CLK(n1516), .C(n1517) );
  CKBD0 U1399 ( .CLK(n1517), .C(n1518) );
  CKBD0 U1400 ( .CLK(n1518), .C(n1519) );
  CKBD0 U1401 ( .CLK(n1519), .C(n1520) );
  BUFFD0 U1402 ( .I(n1520), .Z(n1521) );
  CKBD0 U1403 ( .CLK(n1521), .C(n1522) );
  CKBD0 U1404 ( .CLK(n1522), .C(n1523) );
  CKBD0 U1405 ( .CLK(n1523), .C(n1524) );
  CKBD0 U1406 ( .CLK(n1524), .C(n1525) );
  CKBD0 U1407 ( .CLK(n1525), .C(n1526) );
  CKBD0 U1408 ( .CLK(n1526), .C(n1527) );
  CKBD0 U1409 ( .CLK(n1527), .C(n1528) );
  CKBD0 U1410 ( .CLK(n1528), .C(n1529) );
  CKBD0 U1411 ( .CLK(n1529), .C(n1530) );
  CKBD0 U1412 ( .CLK(n1530), .C(n1531) );
  BUFFD0 U1413 ( .I(n1531), .Z(n1532) );
  CKBD0 U1414 ( .CLK(n1532), .C(n1533) );
  CKBD0 U1415 ( .CLK(n1533), .C(n1534) );
  CKBD0 U1416 ( .CLK(n1534), .C(n1535) );
  CKBD0 U1417 ( .CLK(n1535), .C(n1536) );
  CKBD0 U1418 ( .CLK(n1536), .C(n1537) );
  CKBD0 U1419 ( .CLK(n1537), .C(n1538) );
  CKBD0 U1420 ( .CLK(n1538), .C(n1539) );
  CKBD0 U1421 ( .CLK(n1539), .C(n1540) );
  CKBD0 U1422 ( .CLK(n1540), .C(n1541) );
  CKBD0 U1423 ( .CLK(n1541), .C(n1542) );
  BUFFD0 U1424 ( .I(n1542), .Z(n1543) );
  CKBD0 U1425 ( .CLK(n1543), .C(n1544) );
  CKBD0 U1426 ( .CLK(n1544), .C(n1545) );
  CKBD0 U1427 ( .CLK(n1545), .C(n1546) );
  CKBD0 U1428 ( .CLK(n1546), .C(n1547) );
  CKBD0 U1429 ( .CLK(n1547), .C(n1548) );
  CKBD0 U1430 ( .CLK(n1548), .C(n1549) );
  CKBD0 U1431 ( .CLK(n1549), .C(n1550) );
  CKBD0 U1432 ( .CLK(n1550), .C(n1551) );
  CKBD0 U1433 ( .CLK(n1551), .C(n1552) );
  CKBD0 U1434 ( .CLK(n1552), .C(n1553) );
  BUFFD0 U1435 ( .I(n1553), .Z(n1554) );
  CKBD0 U1436 ( .CLK(n1554), .C(n1555) );
  CKBD0 U1437 ( .CLK(n1555), .C(n1556) );
  CKBD0 U1438 ( .CLK(n1556), .C(n1557) );
  CKBD0 U1439 ( .CLK(n1557), .C(n1558) );
  CKBD0 U1440 ( .CLK(n1558), .C(n1559) );
  CKBD0 U1441 ( .CLK(n1559), .C(n1560) );
  BUFFD0 U1442 ( .I(n8996), .Z(n1561) );
  CKBD0 U1443 ( .CLK(FrameSR[48]), .C(n1562) );
  CKBD0 U1444 ( .CLK(n1562), .C(n1563) );
  BUFFD0 U1445 ( .I(n1563), .Z(n1564) );
  CKBD0 U1446 ( .CLK(n1564), .C(n1565) );
  CKBD0 U1447 ( .CLK(n1565), .C(n1566) );
  CKBD0 U1448 ( .CLK(n1566), .C(n1567) );
  CKBD0 U1449 ( .CLK(n1567), .C(n1568) );
  CKBD0 U1450 ( .CLK(n1568), .C(n1569) );
  CKBD0 U1451 ( .CLK(n1569), .C(n1570) );
  CKBD0 U1452 ( .CLK(n1570), .C(n1571) );
  CKBD0 U1453 ( .CLK(n1571), .C(n1572) );
  CKBD0 U1454 ( .CLK(n1572), .C(n1573) );
  CKBD0 U1455 ( .CLK(n1573), .C(n1574) );
  BUFFD0 U1456 ( .I(n1574), .Z(n1575) );
  CKBD0 U1457 ( .CLK(n1575), .C(n1576) );
  CKBD0 U1458 ( .CLK(n1576), .C(n1577) );
  CKBD0 U1459 ( .CLK(n1577), .C(n1578) );
  CKBD0 U1460 ( .CLK(n1578), .C(n1579) );
  CKBD0 U1461 ( .CLK(n1579), .C(n1580) );
  CKBD0 U1462 ( .CLK(n1580), .C(n1581) );
  CKBD0 U1463 ( .CLK(n1581), .C(n1582) );
  CKBD0 U1464 ( .CLK(n1582), .C(n1583) );
  CKBD0 U1465 ( .CLK(n1583), .C(n1584) );
  BUFFD0 U1466 ( .I(n1584), .Z(n1585) );
  CKBD0 U1467 ( .CLK(n1585), .C(n1586) );
  CKBD0 U1468 ( .CLK(n1586), .C(n1587) );
  CKBD0 U1469 ( .CLK(n1587), .C(n1588) );
  CKBD0 U1470 ( .CLK(n1588), .C(n1589) );
  CKBD0 U1471 ( .CLK(n1589), .C(n1590) );
  CKBD0 U1472 ( .CLK(n1590), .C(n1591) );
  CKBD0 U1473 ( .CLK(n1591), .C(n1592) );
  CKBD0 U1474 ( .CLK(n1592), .C(n1593) );
  CKBD0 U1475 ( .CLK(n1593), .C(n1594) );
  CKBD0 U1476 ( .CLK(n1594), .C(n1595) );
  BUFFD0 U1477 ( .I(n1595), .Z(n1596) );
  CKBD0 U1478 ( .CLK(n1596), .C(n1597) );
  CKBD0 U1479 ( .CLK(n1597), .C(n1598) );
  CKBD0 U1480 ( .CLK(n1598), .C(n1599) );
  CKBD0 U1481 ( .CLK(n1599), .C(n1600) );
  CKBD0 U1482 ( .CLK(n1600), .C(n1601) );
  CKBD0 U1483 ( .CLK(n1601), .C(n1602) );
  CKBD0 U1484 ( .CLK(n1602), .C(n1603) );
  CKBD0 U1485 ( .CLK(n1603), .C(n1604) );
  CKBD0 U1486 ( .CLK(n1604), .C(n1605) );
  CKBD0 U1487 ( .CLK(n1605), .C(n1606) );
  BUFFD0 U1488 ( .I(n1606), .Z(n1607) );
  CKBD0 U1489 ( .CLK(n1607), .C(n1608) );
  CKBD0 U1490 ( .CLK(n1608), .C(n1609) );
  CKBD0 U1491 ( .CLK(n1609), .C(n1610) );
  CKBD0 U1492 ( .CLK(n1610), .C(n1611) );
  CKBD0 U1493 ( .CLK(n1611), .C(n1612) );
  CKBD0 U1494 ( .CLK(n1612), .C(n1613) );
  CKBD0 U1495 ( .CLK(n1613), .C(n1614) );
  CKBD0 U1496 ( .CLK(n1614), .C(n1615) );
  CKBD0 U1497 ( .CLK(n1615), .C(n1616) );
  CKBD0 U1498 ( .CLK(n1616), .C(n1617) );
  BUFFD0 U1499 ( .I(n1617), .Z(n1618) );
  CKBD0 U1500 ( .CLK(n1618), .C(n1619) );
  CKBD0 U1501 ( .CLK(n1619), .C(n1620) );
  CKBD0 U1502 ( .CLK(n1620), .C(n1621) );
  CKBD0 U1503 ( .CLK(n1621), .C(n1622) );
  CKBD0 U1504 ( .CLK(n1622), .C(n1623) );
  CKBD0 U1505 ( .CLK(n1623), .C(n1624) );
  CKBD0 U1506 ( .CLK(n1624), .C(n1625) );
  CKBD0 U1507 ( .CLK(n1625), .C(n1626) );
  CKBD0 U1508 ( .CLK(n1626), .C(n1627) );
  CKBD0 U1509 ( .CLK(n1627), .C(n1628) );
  BUFFD0 U1510 ( .I(n1628), .Z(n1629) );
  CKBD0 U1511 ( .CLK(n1629), .C(n1630) );
  CKBD0 U1512 ( .CLK(n1630), .C(n1631) );
  CKBD0 U1513 ( .CLK(n1631), .C(n1632) );
  CKBD0 U1514 ( .CLK(n1632), .C(n1633) );
  CKBD0 U1515 ( .CLK(n1633), .C(n1634) );
  CKBD0 U1516 ( .CLK(n1634), .C(n1635) );
  CKBD0 U1517 ( .CLK(n1635), .C(n1636) );
  CKBD0 U1518 ( .CLK(n1636), .C(n1637) );
  CKBD0 U1519 ( .CLK(n1637), .C(n1638) );
  CKBD0 U1520 ( .CLK(n1638), .C(n1639) );
  BUFFD0 U1521 ( .I(n1639), .Z(n1640) );
  CKBD0 U1522 ( .CLK(n1640), .C(n1641) );
  CKBD0 U1523 ( .CLK(n1641), .C(n1642) );
  CKBD0 U1524 ( .CLK(n1642), .C(n1643) );
  CKBD0 U1525 ( .CLK(n1643), .C(n1644) );
  CKBD0 U1526 ( .CLK(n1644), .C(n1645) );
  CKBD0 U1527 ( .CLK(n1645), .C(n1646) );
  CKBD0 U1528 ( .CLK(n1646), .C(n1647) );
  CKBD0 U1529 ( .CLK(n1647), .C(n1648) );
  CKBD0 U1530 ( .CLK(n1648), .C(n1649) );
  CKBD0 U1531 ( .CLK(n1649), .C(n1650) );
  BUFFD0 U1532 ( .I(n1650), .Z(n1651) );
  CKBD0 U1533 ( .CLK(n1651), .C(n1652) );
  CKBD0 U1534 ( .CLK(n1652), .C(n1653) );
  CKBD0 U1535 ( .CLK(n1653), .C(n1654) );
  CKBD0 U1536 ( .CLK(n1654), .C(n1655) );
  CKBD0 U1537 ( .CLK(n1655), .C(n1656) );
  CKBD0 U1538 ( .CLK(n1656), .C(n1657) );
  BUFFD0 U1539 ( .I(n9010), .Z(n1658) );
  CKBD0 U1540 ( .CLK(FrameSR[1]), .C(n1659) );
  CKBD0 U1541 ( .CLK(n1659), .C(n1660) );
  BUFFD0 U1542 ( .I(n9012), .Z(n1661) );
  CKBD0 U1543 ( .CLK(FrameSR[5]), .C(n1662) );
  CKBD0 U1544 ( .CLK(n1662), .C(n1663) );
  BUFFD0 U1545 ( .I(n1663), .Z(n1664) );
  BUFFD0 U1546 ( .I(n9009), .Z(n1665) );
  CKBD0 U1547 ( .CLK(FrameSR[17]), .C(n1666) );
  BUFFD0 U1548 ( .I(n1666), .Z(n1667) );
  CKBD0 U1549 ( .CLK(n1667), .C(n1668) );
  CKBD0 U1550 ( .CLK(n1668), .C(n1669) );
  CKBD0 U1551 ( .CLK(n1669), .C(n1670) );
  CKBD0 U1552 ( .CLK(n1670), .C(n1671) );
  CKBD0 U1553 ( .CLK(n1671), .C(n1672) );
  CKBD0 U1554 ( .CLK(n1672), .C(n1673) );
  CKBD0 U1555 ( .CLK(n1673), .C(n1674) );
  CKBD0 U1556 ( .CLK(n1674), .C(n1675) );
  CKBD0 U1557 ( .CLK(n1675), .C(n1676) );
  CKBD0 U1558 ( .CLK(n1676), .C(n1677) );
  BUFFD0 U1559 ( .I(n1677), .Z(n1678) );
  CKBD0 U1560 ( .CLK(n1678), .C(n1679) );
  CKBD0 U1561 ( .CLK(n1679), .C(n1680) );
  CKBD0 U1562 ( .CLK(n1680), .C(n1681) );
  CKBD0 U1563 ( .CLK(n1681), .C(n1682) );
  CKBD0 U1564 ( .CLK(n1682), .C(n1683) );
  CKBD0 U1565 ( .CLK(n1683), .C(n1684) );
  CKBD0 U1566 ( .CLK(n1684), .C(n1685) );
  CKBD0 U1567 ( .CLK(n1685), .C(n1686) );
  CKBD0 U1568 ( .CLK(n1686), .C(n1687) );
  CKBD0 U1569 ( .CLK(n1687), .C(n1688) );
  BUFFD0 U1570 ( .I(n1688), .Z(n1689) );
  CKBD0 U1571 ( .CLK(n1689), .C(n1690) );
  CKBD0 U1572 ( .CLK(n1690), .C(n1691) );
  CKBD0 U1573 ( .CLK(n1691), .C(n1692) );
  CKBD0 U1574 ( .CLK(n1692), .C(n1693) );
  CKBD0 U1575 ( .CLK(n1693), .C(n1694) );
  CKBD0 U1576 ( .CLK(n1694), .C(n1695) );
  CKBD0 U1577 ( .CLK(n1695), .C(n1696) );
  CKBD0 U1578 ( .CLK(n1696), .C(n1697) );
  CKBD0 U1579 ( .CLK(n1697), .C(n1698) );
  CKBD0 U1580 ( .CLK(n1698), .C(n1699) );
  BUFFD0 U1581 ( .I(n1699), .Z(n1700) );
  CKBD0 U1582 ( .CLK(n1700), .C(n1701) );
  CKBD0 U1583 ( .CLK(n1701), .C(n1702) );
  CKBD0 U1584 ( .CLK(n1702), .C(n1703) );
  CKBD0 U1585 ( .CLK(n1703), .C(n1704) );
  CKBD0 U1586 ( .CLK(n1704), .C(n1705) );
  CKBD0 U1587 ( .CLK(n1705), .C(n1706) );
  CKBD0 U1588 ( .CLK(n1706), .C(n1707) );
  CKBD0 U1589 ( .CLK(n1707), .C(n1708) );
  CKBD0 U1590 ( .CLK(n1708), .C(n1709) );
  CKBD0 U1591 ( .CLK(n1709), .C(n1710) );
  BUFFD0 U1592 ( .I(n1710), .Z(n1711) );
  CKBD0 U1593 ( .CLK(n1711), .C(n1712) );
  CKBD0 U1594 ( .CLK(n1712), .C(n1713) );
  CKBD0 U1595 ( .CLK(n1713), .C(n1714) );
  CKBD0 U1596 ( .CLK(n1714), .C(n1715) );
  CKBD0 U1597 ( .CLK(n1715), .C(n1716) );
  CKBD0 U1598 ( .CLK(n1716), .C(n1717) );
  CKBD0 U1599 ( .CLK(n1717), .C(n1718) );
  CKBD0 U1600 ( .CLK(n1718), .C(n1719) );
  CKBD0 U1601 ( .CLK(n1719), .C(n1720) );
  CKBD0 U1602 ( .CLK(n1720), .C(n1721) );
  BUFFD0 U1603 ( .I(n1721), .Z(n1722) );
  CKBD0 U1604 ( .CLK(n1722), .C(n1723) );
  CKBD0 U1605 ( .CLK(n1723), .C(n1724) );
  CKBD0 U1606 ( .CLK(n1724), .C(n1725) );
  CKBD0 U1607 ( .CLK(n1725), .C(n1726) );
  CKBD0 U1608 ( .CLK(n1726), .C(n1727) );
  CKBD0 U1609 ( .CLK(n1727), .C(n1728) );
  CKBD0 U1610 ( .CLK(n1728), .C(n1729) );
  CKBD0 U1611 ( .CLK(n1729), .C(n1730) );
  CKBD0 U1612 ( .CLK(n1730), .C(n1731) );
  BUFFD0 U1613 ( .I(n1731), .Z(n1732) );
  CKBD0 U1614 ( .CLK(n1732), .C(n1733) );
  CKBD0 U1615 ( .CLK(n1733), .C(n1734) );
  CKBD0 U1616 ( .CLK(n1734), .C(n1735) );
  CKBD0 U1617 ( .CLK(n1735), .C(n1736) );
  CKBD0 U1618 ( .CLK(n1736), .C(n1737) );
  CKBD0 U1619 ( .CLK(n1737), .C(n1738) );
  CKBD0 U1620 ( .CLK(n1738), .C(n1739) );
  CKBD0 U1621 ( .CLK(n1739), .C(n1740) );
  CKBD0 U1622 ( .CLK(n1740), .C(n1741) );
  CKBD0 U1623 ( .CLK(n1741), .C(n1742) );
  BUFFD0 U1624 ( .I(n1742), .Z(n1743) );
  CKBD0 U1625 ( .CLK(n1743), .C(n1744) );
  CKBD0 U1626 ( .CLK(n1744), .C(n1745) );
  CKBD0 U1627 ( .CLK(n1745), .C(n1746) );
  CKBD0 U1628 ( .CLK(n1746), .C(n1747) );
  CKBD0 U1629 ( .CLK(n1747), .C(n1748) );
  CKBD0 U1630 ( .CLK(n1748), .C(n1749) );
  CKBD0 U1631 ( .CLK(n1749), .C(n1750) );
  CKBD0 U1632 ( .CLK(n1750), .C(n1751) );
  CKBD0 U1633 ( .CLK(n1751), .C(n1752) );
  CKBD0 U1634 ( .CLK(n1752), .C(n1753) );
  BUFFD0 U1635 ( .I(n1753), .Z(n1754) );
  CKBD0 U1636 ( .CLK(n1754), .C(n1755) );
  CKBD0 U1637 ( .CLK(n1755), .C(n1756) );
  CKBD0 U1638 ( .CLK(n1756), .C(n1757) );
  CKBD0 U1639 ( .CLK(n1757), .C(n1758) );
  CKBD0 U1640 ( .CLK(n1758), .C(n1759) );
  CKBD0 U1641 ( .CLK(n1759), .C(n1760) );
  CKBD0 U1642 ( .CLK(n1760), .C(n1761) );
  BUFFD0 U1643 ( .I(n8964), .Z(n1762) );
  CKBD0 U1644 ( .CLK(FrameSR[32]), .C(n1763) );
  BUFFD0 U1645 ( .I(n1763), .Z(n1764) );
  CKBD0 U1646 ( .CLK(n1764), .C(n1765) );
  CKBD0 U1647 ( .CLK(n1765), .C(n1766) );
  CKBD0 U1648 ( .CLK(n1766), .C(n1767) );
  CKBD0 U1649 ( .CLK(n1767), .C(n1768) );
  CKBD0 U1650 ( .CLK(n1768), .C(n1769) );
  CKBD0 U1651 ( .CLK(n1769), .C(n1770) );
  CKBD0 U1652 ( .CLK(n1770), .C(n1771) );
  CKBD0 U1653 ( .CLK(n1771), .C(n1772) );
  CKBD0 U1654 ( .CLK(n1772), .C(n1773) );
  BUFFD0 U1655 ( .I(n1773), .Z(n1774) );
  CKBD0 U1656 ( .CLK(n1774), .C(n1775) );
  CKBD0 U1657 ( .CLK(n1775), .C(n1776) );
  CKBD0 U1658 ( .CLK(n1776), .C(n1777) );
  CKBD0 U1659 ( .CLK(n1777), .C(n1778) );
  CKBD0 U1660 ( .CLK(n1778), .C(n1779) );
  CKBD0 U1661 ( .CLK(n1779), .C(n1780) );
  CKBD0 U1662 ( .CLK(n1780), .C(n1781) );
  CKBD0 U1663 ( .CLK(n1781), .C(n1782) );
  CKBD0 U1664 ( .CLK(n1782), .C(n1783) );
  CKBD0 U1665 ( .CLK(n1783), .C(n1784) );
  BUFFD0 U1666 ( .I(n1784), .Z(n1785) );
  CKBD0 U1667 ( .CLK(n1785), .C(n1786) );
  CKBD0 U1668 ( .CLK(n1786), .C(n1787) );
  CKBD0 U1669 ( .CLK(n1787), .C(n1788) );
  CKBD0 U1670 ( .CLK(n1788), .C(n1789) );
  CKBD0 U1671 ( .CLK(n1789), .C(n1790) );
  CKBD0 U1672 ( .CLK(n1790), .C(n1791) );
  CKBD0 U1673 ( .CLK(n1791), .C(n1792) );
  CKBD0 U1674 ( .CLK(n1792), .C(n1793) );
  CKBD0 U1675 ( .CLK(n1793), .C(n1794) );
  CKBD0 U1676 ( .CLK(n1794), .C(n1795) );
  BUFFD0 U1677 ( .I(n1795), .Z(n1796) );
  CKBD0 U1678 ( .CLK(n1796), .C(n1797) );
  CKBD0 U1679 ( .CLK(n1797), .C(n1798) );
  CKBD0 U1680 ( .CLK(n1798), .C(n1799) );
  CKBD0 U1681 ( .CLK(n1799), .C(n1800) );
  CKBD0 U1682 ( .CLK(n1800), .C(n1801) );
  CKBD0 U1683 ( .CLK(n1801), .C(n1802) );
  CKBD0 U1684 ( .CLK(n1802), .C(n1803) );
  CKBD0 U1685 ( .CLK(n1803), .C(n1804) );
  CKBD0 U1686 ( .CLK(n1804), .C(n1805) );
  CKBD0 U1687 ( .CLK(n1805), .C(n1806) );
  BUFFD0 U1688 ( .I(n1806), .Z(n1807) );
  CKBD0 U1689 ( .CLK(n1807), .C(n1808) );
  CKBD0 U1690 ( .CLK(n1808), .C(n1809) );
  CKBD0 U1691 ( .CLK(n1809), .C(n1810) );
  CKBD0 U1692 ( .CLK(n1810), .C(n1811) );
  CKBD0 U1693 ( .CLK(n1811), .C(n1812) );
  CKBD0 U1694 ( .CLK(n1812), .C(n1813) );
  CKBD0 U1695 ( .CLK(n1813), .C(n1814) );
  CKBD0 U1696 ( .CLK(n1814), .C(n1815) );
  CKBD0 U1697 ( .CLK(n1815), .C(n1816) );
  CKBD0 U1698 ( .CLK(n1816), .C(n1817) );
  BUFFD0 U1699 ( .I(n1817), .Z(n1818) );
  CKBD0 U1700 ( .CLK(n1818), .C(n1819) );
  CKBD0 U1701 ( .CLK(n1819), .C(n1820) );
  CKBD0 U1702 ( .CLK(n1820), .C(n1821) );
  CKBD0 U1703 ( .CLK(n1821), .C(n1822) );
  CKBD0 U1704 ( .CLK(n1822), .C(n1823) );
  CKBD0 U1705 ( .CLK(n1823), .C(n1824) );
  CKBD0 U1706 ( .CLK(n1824), .C(n1825) );
  CKBD0 U1707 ( .CLK(n1825), .C(n1826) );
  CKBD0 U1708 ( .CLK(n1826), .C(n1827) );
  CKBD0 U1709 ( .CLK(n1827), .C(n1828) );
  BUFFD0 U1710 ( .I(n1828), .Z(n1829) );
  CKBD0 U1711 ( .CLK(n1829), .C(n1830) );
  CKBD0 U1712 ( .CLK(n1830), .C(n1831) );
  CKBD0 U1713 ( .CLK(n1831), .C(n1832) );
  CKBD0 U1714 ( .CLK(n1832), .C(n1833) );
  CKBD0 U1715 ( .CLK(n1833), .C(n1834) );
  CKBD0 U1716 ( .CLK(n1834), .C(n1835) );
  CKBD0 U1717 ( .CLK(n1835), .C(n1836) );
  CKBD0 U1718 ( .CLK(n1836), .C(n1837) );
  CKBD0 U1719 ( .CLK(n1837), .C(n1838) );
  CKBD0 U1720 ( .CLK(n1838), .C(n1839) );
  BUFFD0 U1721 ( .I(n1839), .Z(n1840) );
  CKBD0 U1722 ( .CLK(n1840), .C(n1841) );
  CKBD0 U1723 ( .CLK(n1841), .C(n1842) );
  CKBD0 U1724 ( .CLK(n1842), .C(n1843) );
  CKBD0 U1725 ( .CLK(n1843), .C(n1844) );
  CKBD0 U1726 ( .CLK(n1844), .C(n1845) );
  CKBD0 U1727 ( .CLK(n1845), .C(n1846) );
  CKBD0 U1728 ( .CLK(n1846), .C(n1847) );
  CKBD0 U1729 ( .CLK(n1847), .C(n1848) );
  CKBD0 U1730 ( .CLK(n1848), .C(n1849) );
  BUFFD0 U1731 ( .I(n1849), .Z(n1850) );
  CKBD0 U1732 ( .CLK(n1850), .C(n1851) );
  CKBD0 U1733 ( .CLK(n1851), .C(n1852) );
  CKBD0 U1734 ( .CLK(n1852), .C(n1853) );
  CKBD0 U1735 ( .CLK(n1853), .C(n1854) );
  CKBD0 U1736 ( .CLK(n1854), .C(n1855) );
  CKBD0 U1737 ( .CLK(n1855), .C(n1856) );
  CKBD0 U1738 ( .CLK(n1856), .C(n1857) );
  CKBD0 U1739 ( .CLK(n1857), .C(n1858) );
  CKBD0 U1740 ( .CLK(n1858), .C(n1859) );
  BUFFD0 U1741 ( .I(n3778), .Z(n1860) );
  CKBD0 U1742 ( .CLK(FrameSR[47]), .C(n1861) );
  BUFFD0 U1743 ( .I(n9007), .Z(n1862) );
  CKBD0 U1744 ( .CLK(FrameSR[0]), .C(n1863) );
  CKBD0 U1745 ( .CLK(n1863), .C(n1864) );
  BUFFD0 U1746 ( .I(n9014), .Z(n1865) );
  CKBD0 U1747 ( .CLK(FrameSR[2]), .C(n1866) );
  CKBD0 U1748 ( .CLK(n1866), .C(n1867) );
  BUFFD0 U1749 ( .I(n9011), .Z(n1868) );
  CKBD0 U1750 ( .CLK(FrameSR[4]), .C(n1869) );
  CKBD0 U1751 ( .CLK(n1869), .C(n1870) );
  BUFFD0 U1752 ( .I(n9015), .Z(n1871) );
  CKBD0 U1753 ( .CLK(FrameSR[6]), .C(n1872) );
  CKBD0 U1754 ( .CLK(n1872), .C(n1873) );
  BUFFD0 U1755 ( .I(n1873), .Z(n1874) );
  BUFFD0 U1756 ( .I(n8989), .Z(n1875) );
  CKBD0 U1757 ( .CLK(FrameSR[20]), .C(n1876) );
  CKBD0 U1758 ( .CLK(n1876), .C(n1877) );
  BUFFD0 U1759 ( .I(n1877), .Z(n1878) );
  CKBD0 U1760 ( .CLK(n1878), .C(n1879) );
  CKBD0 U1761 ( .CLK(n1879), .C(n1880) );
  CKBD0 U1762 ( .CLK(n1880), .C(n1881) );
  CKBD0 U1763 ( .CLK(n1881), .C(n1882) );
  CKBD0 U1764 ( .CLK(n1882), .C(n1883) );
  CKBD0 U1765 ( .CLK(n1883), .C(n1884) );
  CKBD0 U1766 ( .CLK(n1884), .C(n1885) );
  CKBD0 U1767 ( .CLK(n1885), .C(n1886) );
  CKBD0 U1768 ( .CLK(n1886), .C(n1887) );
  CKBD0 U1769 ( .CLK(n1887), .C(n1888) );
  BUFFD0 U1770 ( .I(n1888), .Z(n1889) );
  CKBD0 U1771 ( .CLK(n1889), .C(n1890) );
  CKBD0 U1772 ( .CLK(n1890), .C(n1891) );
  CKBD0 U1773 ( .CLK(n1891), .C(n1892) );
  CKBD0 U1774 ( .CLK(n1892), .C(n1893) );
  CKBD0 U1775 ( .CLK(n1893), .C(n1894) );
  CKBD0 U1776 ( .CLK(n1894), .C(n1895) );
  CKBD0 U1777 ( .CLK(n1895), .C(n1896) );
  CKBD0 U1778 ( .CLK(n1896), .C(n1897) );
  CKBD0 U1779 ( .CLK(n1897), .C(n1898) );
  BUFFD0 U1780 ( .I(n1898), .Z(n1899) );
  CKBD0 U1781 ( .CLK(n1899), .C(n1900) );
  CKBD0 U1782 ( .CLK(n1900), .C(n1901) );
  CKBD0 U1783 ( .CLK(n1901), .C(n1902) );
  CKBD0 U1784 ( .CLK(n1902), .C(n1903) );
  CKBD0 U1785 ( .CLK(n1903), .C(n1904) );
  CKBD0 U1786 ( .CLK(n1904), .C(n1905) );
  CKBD0 U1787 ( .CLK(n1905), .C(n1906) );
  CKBD0 U1788 ( .CLK(n1906), .C(n1907) );
  CKBD0 U1789 ( .CLK(n1907), .C(n1908) );
  CKBD0 U1790 ( .CLK(n1908), .C(n1909) );
  BUFFD0 U1791 ( .I(n1909), .Z(n1910) );
  CKBD0 U1792 ( .CLK(n1910), .C(n1911) );
  CKBD0 U1793 ( .CLK(n1911), .C(n1912) );
  CKBD0 U1794 ( .CLK(n1912), .C(n1913) );
  CKBD0 U1795 ( .CLK(n1913), .C(n1914) );
  CKBD0 U1796 ( .CLK(n1914), .C(n1915) );
  CKBD0 U1797 ( .CLK(n1915), .C(n1916) );
  CKBD0 U1798 ( .CLK(n1916), .C(n1917) );
  CKBD0 U1799 ( .CLK(n1917), .C(n1918) );
  CKBD0 U1800 ( .CLK(n1918), .C(n1919) );
  CKBD0 U1801 ( .CLK(n1919), .C(n1920) );
  BUFFD0 U1802 ( .I(n1920), .Z(n1921) );
  CKBD0 U1803 ( .CLK(n1921), .C(n1922) );
  CKBD0 U1804 ( .CLK(n1922), .C(n1923) );
  CKBD0 U1805 ( .CLK(n1923), .C(n1924) );
  CKBD0 U1806 ( .CLK(n1924), .C(n1925) );
  CKBD0 U1807 ( .CLK(n1925), .C(n1926) );
  CKBD0 U1808 ( .CLK(n1926), .C(n1927) );
  CKBD0 U1809 ( .CLK(n1927), .C(n1928) );
  CKBD0 U1810 ( .CLK(n1928), .C(n1929) );
  CKBD0 U1811 ( .CLK(n1929), .C(n1930) );
  CKBD0 U1812 ( .CLK(n1930), .C(n1931) );
  BUFFD0 U1813 ( .I(n1931), .Z(n1932) );
  CKBD0 U1814 ( .CLK(n1932), .C(n1933) );
  CKBD0 U1815 ( .CLK(n1933), .C(n1934) );
  CKBD0 U1816 ( .CLK(n1934), .C(n1935) );
  CKBD0 U1817 ( .CLK(n1935), .C(n1936) );
  CKBD0 U1818 ( .CLK(n1936), .C(n1937) );
  CKBD0 U1819 ( .CLK(n1937), .C(n1938) );
  CKBD0 U1820 ( .CLK(n1938), .C(n1939) );
  CKBD0 U1821 ( .CLK(n1939), .C(n1940) );
  CKBD0 U1822 ( .CLK(n1940), .C(n1941) );
  CKBD0 U1823 ( .CLK(n1941), .C(n1942) );
  BUFFD0 U1824 ( .I(n1942), .Z(n1943) );
  CKBD0 U1825 ( .CLK(n1943), .C(n1944) );
  CKBD0 U1826 ( .CLK(n1944), .C(n1945) );
  CKBD0 U1827 ( .CLK(n1945), .C(n1946) );
  CKBD0 U1828 ( .CLK(n1946), .C(n1947) );
  CKBD0 U1829 ( .CLK(n1947), .C(n1948) );
  CKBD0 U1830 ( .CLK(n1948), .C(n1949) );
  CKBD0 U1831 ( .CLK(n1949), .C(n1950) );
  CKBD0 U1832 ( .CLK(n1950), .C(n1951) );
  CKBD0 U1833 ( .CLK(n1951), .C(n1952) );
  CKBD0 U1834 ( .CLK(n1952), .C(n1953) );
  BUFFD0 U1835 ( .I(n1953), .Z(n1954) );
  CKBD0 U1836 ( .CLK(n1954), .C(n1955) );
  CKBD0 U1837 ( .CLK(n1955), .C(n1956) );
  CKBD0 U1838 ( .CLK(n1956), .C(n1957) );
  CKBD0 U1839 ( .CLK(n1957), .C(n1958) );
  CKBD0 U1840 ( .CLK(n1958), .C(n1959) );
  CKBD0 U1841 ( .CLK(n1959), .C(n1960) );
  CKBD0 U1842 ( .CLK(n1960), .C(n1961) );
  CKBD0 U1843 ( .CLK(n1961), .C(n1962) );
  CKBD0 U1844 ( .CLK(n1962), .C(n1963) );
  CKBD0 U1845 ( .CLK(n1963), .C(n1964) );
  BUFFD0 U1846 ( .I(n1964), .Z(n1965) );
  CKBD0 U1847 ( .CLK(n1965), .C(n1966) );
  CKBD0 U1848 ( .CLK(n1966), .C(n1967) );
  CKBD0 U1849 ( .CLK(n1967), .C(n1968) );
  CKBD0 U1850 ( .CLK(n1968), .C(n1969) );
  CKBD0 U1851 ( .CLK(n1969), .C(n1970) );
  CKBD0 U1852 ( .CLK(n1970), .C(n1971) );
  BUFFD0 U1853 ( .I(n8990), .Z(n1972) );
  CKBD0 U1854 ( .CLK(FrameSR[34]), .C(n1973) );
  CKBD0 U1855 ( .CLK(n1973), .C(n1974) );
  BUFFD0 U1856 ( .I(n1974), .Z(n1975) );
  CKBD0 U1857 ( .CLK(n1975), .C(n1976) );
  CKBD0 U1858 ( .CLK(n1976), .C(n1977) );
  CKBD0 U1859 ( .CLK(n1977), .C(n1978) );
  CKBD0 U1860 ( .CLK(n1978), .C(n1979) );
  CKBD0 U1861 ( .CLK(n1979), .C(n1980) );
  CKBD0 U1862 ( .CLK(n1980), .C(n1981) );
  CKBD0 U1863 ( .CLK(n1981), .C(n1982) );
  CKBD0 U1864 ( .CLK(n1982), .C(n1983) );
  CKBD0 U1865 ( .CLK(n1983), .C(n1984) );
  CKBD0 U1866 ( .CLK(n1984), .C(n1985) );
  BUFFD0 U1867 ( .I(n1985), .Z(n1986) );
  CKBD0 U1868 ( .CLK(n1986), .C(n1987) );
  CKBD0 U1869 ( .CLK(n1987), .C(n1988) );
  CKBD0 U1870 ( .CLK(n1988), .C(n1989) );
  CKBD0 U1871 ( .CLK(n1989), .C(n1990) );
  CKBD0 U1872 ( .CLK(n1990), .C(n1991) );
  CKBD0 U1873 ( .CLK(n1991), .C(n1992) );
  CKBD0 U1874 ( .CLK(n1992), .C(n1993) );
  CKBD0 U1875 ( .CLK(n1993), .C(n1994) );
  CKBD0 U1876 ( .CLK(n1994), .C(n1995) );
  BUFFD0 U1877 ( .I(n1995), .Z(n1996) );
  CKBD0 U1878 ( .CLK(n1996), .C(n1997) );
  CKBD0 U1879 ( .CLK(n1997), .C(n1998) );
  CKBD0 U1880 ( .CLK(n1998), .C(n1999) );
  CKBD0 U1881 ( .CLK(n1999), .C(n2000) );
  CKBD0 U1882 ( .CLK(n2000), .C(n2001) );
  CKBD0 U1883 ( .CLK(n2001), .C(n2002) );
  CKBD0 U1884 ( .CLK(n2002), .C(n2003) );
  CKBD0 U1885 ( .CLK(n2003), .C(n2004) );
  CKBD0 U1886 ( .CLK(n2004), .C(n2005) );
  CKBD0 U1887 ( .CLK(n2005), .C(n2006) );
  BUFFD0 U1888 ( .I(n2006), .Z(n2007) );
  CKBD0 U1889 ( .CLK(n2007), .C(n2008) );
  CKBD0 U1890 ( .CLK(n2008), .C(n2009) );
  CKBD0 U1891 ( .CLK(n2009), .C(n2010) );
  CKBD0 U1892 ( .CLK(n2010), .C(n2011) );
  CKBD0 U1893 ( .CLK(n2011), .C(n2012) );
  CKBD0 U1894 ( .CLK(n2012), .C(n2013) );
  CKBD0 U1895 ( .CLK(n2013), .C(n2014) );
  CKBD0 U1896 ( .CLK(n2014), .C(n2015) );
  CKBD0 U1897 ( .CLK(n2015), .C(n2016) );
  CKBD0 U1898 ( .CLK(n2016), .C(n2017) );
  BUFFD0 U1899 ( .I(n2017), .Z(n2018) );
  CKBD0 U1900 ( .CLK(n2018), .C(n2019) );
  CKBD0 U1901 ( .CLK(n2019), .C(n2020) );
  CKBD0 U1902 ( .CLK(n2020), .C(n2021) );
  CKBD0 U1903 ( .CLK(n2021), .C(n2022) );
  CKBD0 U1904 ( .CLK(n2022), .C(n2023) );
  CKBD0 U1905 ( .CLK(n2023), .C(n2024) );
  CKBD0 U1906 ( .CLK(n2024), .C(n2025) );
  CKBD0 U1907 ( .CLK(n2025), .C(n2026) );
  CKBD0 U1908 ( .CLK(n2026), .C(n2027) );
  CKBD0 U1909 ( .CLK(n2027), .C(n2028) );
  BUFFD0 U1910 ( .I(n2028), .Z(n2029) );
  CKBD0 U1911 ( .CLK(n2029), .C(n2030) );
  CKBD0 U1912 ( .CLK(n2030), .C(n2031) );
  CKBD0 U1913 ( .CLK(n2031), .C(n2032) );
  CKBD0 U1914 ( .CLK(n2032), .C(n2033) );
  CKBD0 U1915 ( .CLK(n2033), .C(n2034) );
  CKBD0 U1916 ( .CLK(n2034), .C(n2035) );
  CKBD0 U1917 ( .CLK(n2035), .C(n2036) );
  CKBD0 U1918 ( .CLK(n2036), .C(n2037) );
  CKBD0 U1919 ( .CLK(n2037), .C(n2038) );
  CKBD0 U1920 ( .CLK(n2038), .C(n2039) );
  BUFFD0 U1921 ( .I(n2039), .Z(n2040) );
  CKBD0 U1922 ( .CLK(n2040), .C(n2041) );
  CKBD0 U1923 ( .CLK(n2041), .C(n2042) );
  CKBD0 U1924 ( .CLK(n2042), .C(n2043) );
  CKBD0 U1925 ( .CLK(n2043), .C(n2044) );
  CKBD0 U1926 ( .CLK(n2044), .C(n2045) );
  CKBD0 U1927 ( .CLK(n2045), .C(n2046) );
  CKBD0 U1928 ( .CLK(n2046), .C(n2047) );
  CKBD0 U1929 ( .CLK(n2047), .C(n2048) );
  CKBD0 U1930 ( .CLK(n2048), .C(n2049) );
  CKBD0 U1931 ( .CLK(n2049), .C(n2050) );
  BUFFD0 U1932 ( .I(n2050), .Z(n2051) );
  CKBD0 U1933 ( .CLK(n2051), .C(n2052) );
  CKBD0 U1934 ( .CLK(n2052), .C(n2053) );
  CKBD0 U1935 ( .CLK(n2053), .C(n2054) );
  CKBD0 U1936 ( .CLK(n2054), .C(n2055) );
  CKBD0 U1937 ( .CLK(n2055), .C(n2056) );
  CKBD0 U1938 ( .CLK(n2056), .C(n2057) );
  CKBD0 U1939 ( .CLK(n2057), .C(n2058) );
  CKBD0 U1940 ( .CLK(n2058), .C(n2059) );
  CKBD0 U1941 ( .CLK(n2059), .C(n2060) );
  CKBD0 U1942 ( .CLK(n2060), .C(n2061) );
  BUFFD0 U1943 ( .I(n2061), .Z(n2062) );
  CKBD0 U1944 ( .CLK(n2062), .C(n2063) );
  CKBD0 U1945 ( .CLK(n2063), .C(n2064) );
  CKBD0 U1946 ( .CLK(n2064), .C(n2065) );
  CKBD0 U1947 ( .CLK(n2065), .C(n2066) );
  CKBD0 U1948 ( .CLK(n2066), .C(n2067) );
  CKBD0 U1949 ( .CLK(n2067), .C(n2068) );
  BUFFD0 U1950 ( .I(n8988), .Z(n2069) );
  CKBD0 U1951 ( .CLK(FrameSR[49]), .C(n2070) );
  CKBD0 U1952 ( .CLK(n2070), .C(n2071) );
  BUFFD0 U1953 ( .I(n2071), .Z(n2072) );
  CKBD0 U1954 ( .CLK(n2072), .C(n2073) );
  CKBD0 U1955 ( .CLK(n2073), .C(n2074) );
  CKBD0 U1956 ( .CLK(n2074), .C(n2075) );
  CKBD0 U1957 ( .CLK(n2075), .C(n2076) );
  CKBD0 U1958 ( .CLK(n2076), .C(n2077) );
  CKBD0 U1959 ( .CLK(n2077), .C(n2078) );
  CKBD0 U1960 ( .CLK(n2078), .C(n2079) );
  CKBD0 U1961 ( .CLK(n2079), .C(n2080) );
  CKBD0 U1962 ( .CLK(n2080), .C(n2081) );
  CKBD0 U1963 ( .CLK(n2081), .C(n2082) );
  BUFFD0 U1964 ( .I(n2082), .Z(n2083) );
  CKBD0 U1965 ( .CLK(n2083), .C(n2084) );
  CKBD0 U1966 ( .CLK(n2084), .C(n2085) );
  CKBD0 U1967 ( .CLK(n2085), .C(n2086) );
  CKBD0 U1968 ( .CLK(n2086), .C(n2087) );
  CKBD0 U1969 ( .CLK(n2087), .C(n2088) );
  CKBD0 U1970 ( .CLK(n2088), .C(n2089) );
  CKBD0 U1971 ( .CLK(n2089), .C(n2090) );
  CKBD0 U1972 ( .CLK(n2090), .C(n2091) );
  CKBD0 U1973 ( .CLK(n2091), .C(n2092) );
  BUFFD0 U1974 ( .I(n2092), .Z(n2093) );
  CKBD0 U1975 ( .CLK(n2093), .C(n2094) );
  CKBD0 U1976 ( .CLK(n2094), .C(n2095) );
  CKBD0 U1977 ( .CLK(n2095), .C(n2096) );
  CKBD0 U1978 ( .CLK(n2096), .C(n2097) );
  CKBD0 U1979 ( .CLK(n2097), .C(n2098) );
  CKBD0 U1980 ( .CLK(n2098), .C(n2099) );
  CKBD0 U1981 ( .CLK(n2099), .C(n2100) );
  CKBD0 U1982 ( .CLK(n2100), .C(n2101) );
  CKBD0 U1983 ( .CLK(n2101), .C(n2102) );
  CKBD0 U1984 ( .CLK(n2102), .C(n2103) );
  BUFFD0 U1985 ( .I(n2103), .Z(n2104) );
  CKBD0 U1986 ( .CLK(n2104), .C(n2105) );
  CKBD0 U1987 ( .CLK(n2105), .C(n2106) );
  CKBD0 U1988 ( .CLK(n2106), .C(n2107) );
  CKBD0 U1989 ( .CLK(n2107), .C(n2108) );
  CKBD0 U1990 ( .CLK(n2108), .C(n2109) );
  CKBD0 U1991 ( .CLK(n2109), .C(n2110) );
  CKBD0 U1992 ( .CLK(n2110), .C(n2111) );
  CKBD0 U1993 ( .CLK(n2111), .C(n2112) );
  CKBD0 U1994 ( .CLK(n2112), .C(n2113) );
  CKBD0 U1995 ( .CLK(n2113), .C(n2114) );
  BUFFD0 U1996 ( .I(n2114), .Z(n2115) );
  CKBD0 U1997 ( .CLK(n2115), .C(n2116) );
  CKBD0 U1998 ( .CLK(n2116), .C(n2117) );
  CKBD0 U1999 ( .CLK(n2117), .C(n2118) );
  CKBD0 U2000 ( .CLK(n2118), .C(n2119) );
  CKBD0 U2001 ( .CLK(n2119), .C(n2120) );
  CKBD0 U2002 ( .CLK(n2120), .C(n2121) );
  CKBD0 U2003 ( .CLK(n2121), .C(n2122) );
  CKBD0 U2004 ( .CLK(n2122), .C(n2123) );
  CKBD0 U2005 ( .CLK(n2123), .C(n2124) );
  CKBD0 U2006 ( .CLK(n2124), .C(n2125) );
  BUFFD0 U2007 ( .I(n2125), .Z(n2126) );
  CKBD0 U2008 ( .CLK(n2126), .C(n2127) );
  CKBD0 U2009 ( .CLK(n2127), .C(n2128) );
  CKBD0 U2010 ( .CLK(n2128), .C(n2129) );
  CKBD0 U2011 ( .CLK(n2129), .C(n2130) );
  CKBD0 U2012 ( .CLK(n2130), .C(n2131) );
  CKBD0 U2013 ( .CLK(n2131), .C(n2132) );
  CKBD0 U2014 ( .CLK(n2132), .C(n2133) );
  CKBD0 U2015 ( .CLK(n2133), .C(n2134) );
  CKBD0 U2016 ( .CLK(n2134), .C(n2135) );
  CKBD0 U2017 ( .CLK(n2135), .C(n2136) );
  BUFFD0 U2018 ( .I(n2136), .Z(n2137) );
  CKBD0 U2019 ( .CLK(n2137), .C(n2138) );
  CKBD0 U2020 ( .CLK(n2138), .C(n2139) );
  CKBD0 U2021 ( .CLK(n2139), .C(n2140) );
  CKBD0 U2022 ( .CLK(n2140), .C(n2141) );
  CKBD0 U2023 ( .CLK(n2141), .C(n2142) );
  CKBD0 U2024 ( .CLK(n2142), .C(n2143) );
  CKBD0 U2025 ( .CLK(n2143), .C(n2144) );
  CKBD0 U2026 ( .CLK(n2144), .C(n2145) );
  CKBD0 U2027 ( .CLK(n2145), .C(n2146) );
  CKBD0 U2028 ( .CLK(n2146), .C(n2147) );
  BUFFD0 U2029 ( .I(n2147), .Z(n2148) );
  CKBD0 U2030 ( .CLK(n2148), .C(n2149) );
  CKBD0 U2031 ( .CLK(n2149), .C(n2150) );
  CKBD0 U2032 ( .CLK(n2150), .C(n2151) );
  CKBD0 U2033 ( .CLK(n2151), .C(n2152) );
  CKBD0 U2034 ( .CLK(n2152), .C(n2153) );
  CKBD0 U2035 ( .CLK(n2153), .C(n2154) );
  CKBD0 U2036 ( .CLK(n2154), .C(n2155) );
  CKBD0 U2037 ( .CLK(n2155), .C(n2156) );
  CKBD0 U2038 ( .CLK(n2156), .C(n2157) );
  CKBD0 U2039 ( .CLK(n2157), .C(n2158) );
  BUFFD0 U2040 ( .I(n2158), .Z(n2159) );
  CKBD0 U2041 ( .CLK(n2159), .C(n2160) );
  CKBD0 U2042 ( .CLK(n2160), .C(n2161) );
  CKBD0 U2043 ( .CLK(n2161), .C(n2162) );
  CKBD0 U2044 ( .CLK(n2162), .C(n2163) );
  CKBD0 U2045 ( .CLK(n2163), .C(n2164) );
  CKBD0 U2046 ( .CLK(n2164), .C(n2165) );
  BUFFD0 U2047 ( .I(n8991), .Z(n2166) );
  CKBD0 U2048 ( .CLK(FrameSR[50]), .C(n2167) );
  CKBD0 U2049 ( .CLK(n2167), .C(n2168) );
  BUFFD0 U2050 ( .I(n2168), .Z(n2169) );
  CKBD0 U2051 ( .CLK(n2169), .C(n2170) );
  CKBD0 U2052 ( .CLK(n2170), .C(n2171) );
  CKBD0 U2053 ( .CLK(n2171), .C(n2172) );
  CKBD0 U2054 ( .CLK(n2172), .C(n2173) );
  CKBD0 U2055 ( .CLK(n2173), .C(n2174) );
  CKBD0 U2056 ( .CLK(n2174), .C(n2175) );
  CKBD0 U2057 ( .CLK(n2175), .C(n2176) );
  CKBD0 U2058 ( .CLK(n2176), .C(n2177) );
  CKBD0 U2059 ( .CLK(n2177), .C(n2178) );
  CKBD0 U2060 ( .CLK(n2178), .C(n2179) );
  BUFFD0 U2061 ( .I(n2179), .Z(n2180) );
  CKBD0 U2062 ( .CLK(n2180), .C(n2181) );
  CKBD0 U2063 ( .CLK(n2181), .C(n2182) );
  CKBD0 U2064 ( .CLK(n2182), .C(n2183) );
  CKBD0 U2065 ( .CLK(n2183), .C(n2184) );
  CKBD0 U2066 ( .CLK(n2184), .C(n2185) );
  CKBD0 U2067 ( .CLK(n2185), .C(n2186) );
  CKBD0 U2068 ( .CLK(n2186), .C(n2187) );
  CKBD0 U2069 ( .CLK(n2187), .C(n2188) );
  CKBD0 U2070 ( .CLK(n2188), .C(n2189) );
  BUFFD0 U2071 ( .I(n2189), .Z(n2190) );
  CKBD0 U2072 ( .CLK(n2190), .C(n2191) );
  CKBD0 U2073 ( .CLK(n2191), .C(n2192) );
  CKBD0 U2074 ( .CLK(n2192), .C(n2193) );
  CKBD0 U2075 ( .CLK(n2193), .C(n2194) );
  CKBD0 U2076 ( .CLK(n2194), .C(n2195) );
  CKBD0 U2077 ( .CLK(n2195), .C(n2196) );
  CKBD0 U2078 ( .CLK(n2196), .C(n2197) );
  CKBD0 U2079 ( .CLK(n2197), .C(n2198) );
  CKBD0 U2080 ( .CLK(n2198), .C(n2199) );
  CKBD0 U2081 ( .CLK(n2199), .C(n2200) );
  BUFFD0 U2082 ( .I(n2200), .Z(n2201) );
  CKBD0 U2083 ( .CLK(n2201), .C(n2202) );
  CKBD0 U2084 ( .CLK(n2202), .C(n2203) );
  CKBD0 U2085 ( .CLK(n2203), .C(n2204) );
  CKBD0 U2086 ( .CLK(n2204), .C(n2205) );
  CKBD0 U2087 ( .CLK(n2205), .C(n2206) );
  CKBD0 U2088 ( .CLK(n2206), .C(n2207) );
  CKBD0 U2089 ( .CLK(n2207), .C(n2208) );
  CKBD0 U2090 ( .CLK(n2208), .C(n2209) );
  CKBD0 U2091 ( .CLK(n2209), .C(n2210) );
  CKBD0 U2092 ( .CLK(n2210), .C(n2211) );
  BUFFD0 U2093 ( .I(n2211), .Z(n2212) );
  CKBD0 U2094 ( .CLK(n2212), .C(n2213) );
  CKBD0 U2095 ( .CLK(n2213), .C(n2214) );
  CKBD0 U2096 ( .CLK(n2214), .C(n2215) );
  CKBD0 U2097 ( .CLK(n2215), .C(n2216) );
  CKBD0 U2098 ( .CLK(n2216), .C(n2217) );
  CKBD0 U2099 ( .CLK(n2217), .C(n2218) );
  CKBD0 U2100 ( .CLK(n2218), .C(n2219) );
  CKBD0 U2101 ( .CLK(n2219), .C(n2220) );
  CKBD0 U2102 ( .CLK(n2220), .C(n2221) );
  CKBD0 U2103 ( .CLK(n2221), .C(n2222) );
  BUFFD0 U2104 ( .I(n2222), .Z(n2223) );
  CKBD0 U2105 ( .CLK(n2223), .C(n2224) );
  CKBD0 U2106 ( .CLK(n2224), .C(n2225) );
  CKBD0 U2107 ( .CLK(n2225), .C(n2226) );
  CKBD0 U2108 ( .CLK(n2226), .C(n2227) );
  CKBD0 U2109 ( .CLK(n2227), .C(n2228) );
  CKBD0 U2110 ( .CLK(n2228), .C(n2229) );
  CKBD0 U2111 ( .CLK(n2229), .C(n2230) );
  CKBD0 U2112 ( .CLK(n2230), .C(n2231) );
  CKBD0 U2113 ( .CLK(n2231), .C(n2232) );
  CKBD0 U2114 ( .CLK(n2232), .C(n2233) );
  BUFFD0 U2115 ( .I(n2233), .Z(n2234) );
  CKBD0 U2116 ( .CLK(n2234), .C(n2235) );
  CKBD0 U2117 ( .CLK(n2235), .C(n2236) );
  CKBD0 U2118 ( .CLK(n2236), .C(n2237) );
  CKBD0 U2119 ( .CLK(n2237), .C(n2238) );
  CKBD0 U2120 ( .CLK(n2238), .C(n2239) );
  CKBD0 U2121 ( .CLK(n2239), .C(n2240) );
  CKBD0 U2122 ( .CLK(n2240), .C(n2241) );
  CKBD0 U2123 ( .CLK(n2241), .C(n2242) );
  CKBD0 U2124 ( .CLK(n2242), .C(n2243) );
  CKBD0 U2125 ( .CLK(n2243), .C(n2244) );
  BUFFD0 U2126 ( .I(n2244), .Z(n2245) );
  CKBD0 U2127 ( .CLK(n2245), .C(n2246) );
  CKBD0 U2128 ( .CLK(n2246), .C(n2247) );
  CKBD0 U2129 ( .CLK(n2247), .C(n2248) );
  CKBD0 U2130 ( .CLK(n2248), .C(n2249) );
  CKBD0 U2131 ( .CLK(n2249), .C(n2250) );
  CKBD0 U2132 ( .CLK(n2250), .C(n2251) );
  CKBD0 U2133 ( .CLK(n2251), .C(n2252) );
  CKBD0 U2134 ( .CLK(n2252), .C(n2253) );
  CKBD0 U2135 ( .CLK(n2253), .C(n2254) );
  CKBD0 U2136 ( .CLK(n2254), .C(n2255) );
  BUFFD0 U2137 ( .I(n2255), .Z(n2256) );
  CKBD0 U2138 ( .CLK(n2256), .C(n2257) );
  CKBD0 U2139 ( .CLK(n2257), .C(n2258) );
  CKBD0 U2140 ( .CLK(n2258), .C(n2259) );
  CKBD0 U2141 ( .CLK(n2259), .C(n2260) );
  CKBD0 U2142 ( .CLK(n2260), .C(n2261) );
  CKBD0 U2143 ( .CLK(n2261), .C(n2262) );
  BUFFD0 U2144 ( .I(n8993), .Z(n2263) );
  CKBD0 U2145 ( .CLK(FrameSR[35]), .C(n2264) );
  CKBD0 U2146 ( .CLK(n2264), .C(n2265) );
  BUFFD0 U2147 ( .I(n2265), .Z(n2266) );
  CKBD0 U2148 ( .CLK(n2266), .C(n2267) );
  CKBD0 U2149 ( .CLK(n2267), .C(n2268) );
  CKBD0 U2150 ( .CLK(n2268), .C(n2269) );
  CKBD0 U2151 ( .CLK(n2269), .C(n2270) );
  CKBD0 U2152 ( .CLK(n2270), .C(n2271) );
  CKBD0 U2153 ( .CLK(n2271), .C(n2272) );
  CKBD0 U2154 ( .CLK(n2272), .C(n2273) );
  CKBD0 U2155 ( .CLK(n2273), .C(n2274) );
  CKBD0 U2156 ( .CLK(n2274), .C(n2275) );
  CKBD0 U2157 ( .CLK(n2275), .C(n2276) );
  BUFFD0 U2158 ( .I(n2276), .Z(n2277) );
  CKBD0 U2159 ( .CLK(n2277), .C(n2278) );
  CKBD0 U2160 ( .CLK(n2278), .C(n2279) );
  CKBD0 U2161 ( .CLK(n2279), .C(n2280) );
  CKBD0 U2162 ( .CLK(n2280), .C(n2281) );
  CKBD0 U2163 ( .CLK(n2281), .C(n2282) );
  CKBD0 U2164 ( .CLK(n2282), .C(n2283) );
  CKBD0 U2165 ( .CLK(n2283), .C(n2284) );
  CKBD0 U2166 ( .CLK(n2284), .C(n2285) );
  CKBD0 U2167 ( .CLK(n2285), .C(n2286) );
  BUFFD0 U2168 ( .I(n2286), .Z(n2287) );
  CKBD0 U2169 ( .CLK(n2287), .C(n2288) );
  CKBD0 U2170 ( .CLK(n2288), .C(n2289) );
  CKBD0 U2171 ( .CLK(n2289), .C(n2290) );
  CKBD0 U2172 ( .CLK(n2290), .C(n2291) );
  CKBD0 U2173 ( .CLK(n2291), .C(n2292) );
  CKBD0 U2174 ( .CLK(n2292), .C(n2293) );
  CKBD0 U2175 ( .CLK(n2293), .C(n2294) );
  CKBD0 U2176 ( .CLK(n2294), .C(n2295) );
  CKBD0 U2177 ( .CLK(n2295), .C(n2296) );
  CKBD0 U2178 ( .CLK(n2296), .C(n2297) );
  BUFFD0 U2179 ( .I(n2297), .Z(n2298) );
  CKBD0 U2180 ( .CLK(n2298), .C(n2299) );
  CKBD0 U2181 ( .CLK(n2299), .C(n2300) );
  CKBD0 U2182 ( .CLK(n2300), .C(n2301) );
  CKBD0 U2183 ( .CLK(n2301), .C(n2302) );
  CKBD0 U2184 ( .CLK(n2302), .C(n2303) );
  CKBD0 U2185 ( .CLK(n2303), .C(n2304) );
  CKBD0 U2186 ( .CLK(n2304), .C(n2305) );
  CKBD0 U2187 ( .CLK(n2305), .C(n2306) );
  CKBD0 U2188 ( .CLK(n2306), .C(n2307) );
  CKBD0 U2189 ( .CLK(n2307), .C(n2308) );
  BUFFD0 U2190 ( .I(n2308), .Z(n2309) );
  CKBD0 U2191 ( .CLK(n2309), .C(n2310) );
  CKBD0 U2192 ( .CLK(n2310), .C(n2311) );
  CKBD0 U2193 ( .CLK(n2311), .C(n2312) );
  CKBD0 U2194 ( .CLK(n2312), .C(n2313) );
  CKBD0 U2195 ( .CLK(n2313), .C(n2314) );
  CKBD0 U2196 ( .CLK(n2314), .C(n2315) );
  CKBD0 U2197 ( .CLK(n2315), .C(n2316) );
  CKBD0 U2198 ( .CLK(n2316), .C(n2317) );
  CKBD0 U2199 ( .CLK(n2317), .C(n2318) );
  CKBD0 U2200 ( .CLK(n2318), .C(n2319) );
  BUFFD0 U2201 ( .I(n2319), .Z(n2320) );
  CKBD0 U2202 ( .CLK(n2320), .C(n2321) );
  CKBD0 U2203 ( .CLK(n2321), .C(n2322) );
  CKBD0 U2204 ( .CLK(n2322), .C(n2323) );
  CKBD0 U2205 ( .CLK(n2323), .C(n2324) );
  CKBD0 U2206 ( .CLK(n2324), .C(n2325) );
  CKBD0 U2207 ( .CLK(n2325), .C(n2326) );
  CKBD0 U2208 ( .CLK(n2326), .C(n2327) );
  CKBD0 U2209 ( .CLK(n2327), .C(n2328) );
  CKBD0 U2210 ( .CLK(n2328), .C(n2329) );
  CKBD0 U2211 ( .CLK(n2329), .C(n2330) );
  BUFFD0 U2212 ( .I(n2330), .Z(n2331) );
  CKBD0 U2213 ( .CLK(n2331), .C(n2332) );
  CKBD0 U2214 ( .CLK(n2332), .C(n2333) );
  CKBD0 U2215 ( .CLK(n2333), .C(n2334) );
  CKBD0 U2216 ( .CLK(n2334), .C(n2335) );
  CKBD0 U2217 ( .CLK(n2335), .C(n2336) );
  CKBD0 U2218 ( .CLK(n2336), .C(n2337) );
  CKBD0 U2219 ( .CLK(n2337), .C(n2338) );
  CKBD0 U2220 ( .CLK(n2338), .C(n2339) );
  CKBD0 U2221 ( .CLK(n2339), .C(n2340) );
  CKBD0 U2222 ( .CLK(n2340), .C(n2341) );
  BUFFD0 U2223 ( .I(n2341), .Z(n2342) );
  CKBD0 U2224 ( .CLK(n2342), .C(n2343) );
  CKBD0 U2225 ( .CLK(n2343), .C(n2344) );
  CKBD0 U2226 ( .CLK(n2344), .C(n2345) );
  CKBD0 U2227 ( .CLK(n2345), .C(n2346) );
  CKBD0 U2228 ( .CLK(n2346), .C(n2347) );
  CKBD0 U2229 ( .CLK(n2347), .C(n2348) );
  CKBD0 U2230 ( .CLK(n2348), .C(n2349) );
  CKBD0 U2231 ( .CLK(n2349), .C(n2350) );
  CKBD0 U2232 ( .CLK(n2350), .C(n2351) );
  CKBD0 U2233 ( .CLK(n2351), .C(n2352) );
  BUFFD0 U2234 ( .I(n2352), .Z(n2353) );
  CKBD0 U2235 ( .CLK(n2353), .C(n2354) );
  CKBD0 U2236 ( .CLK(n2354), .C(n2355) );
  CKBD0 U2237 ( .CLK(n2355), .C(n2356) );
  CKBD0 U2238 ( .CLK(n2356), .C(n2357) );
  CKBD0 U2239 ( .CLK(n2357), .C(n2358) );
  CKBD0 U2240 ( .CLK(n2358), .C(n2359) );
  BUFFD0 U2241 ( .I(n8980), .Z(n2360) );
  CKBD0 U2242 ( .CLK(FrameSR[51]), .C(n2361) );
  CKBD0 U2243 ( .CLK(n2361), .C(n2362) );
  CKBD0 U2244 ( .CLK(n2362), .C(n2363) );
  CKBD0 U2245 ( .CLK(n2363), .C(n2364) );
  CKBD0 U2246 ( .CLK(n2364), .C(n2365) );
  CKBD0 U2247 ( .CLK(n2365), .C(n2366) );
  CKBD0 U2248 ( .CLK(n2366), .C(n2367) );
  CKBD0 U2249 ( .CLK(n2367), .C(n2368) );
  CKBD0 U2250 ( .CLK(n2368), .C(n2369) );
  CKBD0 U2251 ( .CLK(n2369), .C(n2370) );
  BUFFD0 U2252 ( .I(n2370), .Z(n2371) );
  CKBD0 U2253 ( .CLK(n2371), .C(n2372) );
  CKBD0 U2254 ( .CLK(n2372), .C(n2373) );
  CKBD0 U2255 ( .CLK(n2373), .C(n2374) );
  CKBD0 U2256 ( .CLK(n2374), .C(n2375) );
  CKBD0 U2257 ( .CLK(n2375), .C(n2376) );
  CKBD0 U2258 ( .CLK(n2376), .C(n2377) );
  CKBD0 U2259 ( .CLK(n2377), .C(n2378) );
  CKBD0 U2260 ( .CLK(n2378), .C(n2379) );
  CKBD0 U2261 ( .CLK(n2379), .C(n2380) );
  BUFFD0 U2262 ( .I(n2380), .Z(n2381) );
  CKBD0 U2263 ( .CLK(n2381), .C(n2382) );
  CKBD0 U2264 ( .CLK(n2382), .C(n2383) );
  CKBD0 U2265 ( .CLK(n2383), .C(n2384) );
  CKBD0 U2266 ( .CLK(n2384), .C(n2385) );
  CKBD0 U2267 ( .CLK(n2385), .C(n2386) );
  CKBD0 U2268 ( .CLK(n2386), .C(n2387) );
  CKBD0 U2269 ( .CLK(n2387), .C(n2388) );
  CKBD0 U2270 ( .CLK(n2388), .C(n2389) );
  CKBD0 U2271 ( .CLK(n2389), .C(n2390) );
  CKBD0 U2272 ( .CLK(n2390), .C(n2391) );
  BUFFD0 U2273 ( .I(n2391), .Z(n2392) );
  CKBD0 U2274 ( .CLK(n2392), .C(n2393) );
  CKBD0 U2275 ( .CLK(n2393), .C(n2394) );
  CKBD0 U2276 ( .CLK(n2394), .C(n2395) );
  CKBD0 U2277 ( .CLK(n2395), .C(n2396) );
  CKBD0 U2278 ( .CLK(n2396), .C(n2397) );
  CKBD0 U2279 ( .CLK(n2397), .C(n2398) );
  CKBD0 U2280 ( .CLK(n2398), .C(n2399) );
  CKBD0 U2281 ( .CLK(n2399), .C(n2400) );
  CKBD0 U2282 ( .CLK(n2400), .C(n2401) );
  CKBD0 U2283 ( .CLK(n2401), .C(n2402) );
  BUFFD0 U2284 ( .I(n2402), .Z(n2403) );
  CKBD0 U2285 ( .CLK(n2403), .C(n2404) );
  CKBD0 U2286 ( .CLK(n2404), .C(n2405) );
  CKBD0 U2287 ( .CLK(n2405), .C(n2406) );
  CKBD0 U2288 ( .CLK(n2406), .C(n2407) );
  CKBD0 U2289 ( .CLK(n2407), .C(n2408) );
  CKBD0 U2290 ( .CLK(n2408), .C(n2409) );
  CKBD0 U2291 ( .CLK(n2409), .C(n2410) );
  CKBD0 U2292 ( .CLK(n2410), .C(n2411) );
  CKBD0 U2293 ( .CLK(n2411), .C(n2412) );
  CKBD0 U2294 ( .CLK(n2412), .C(n2413) );
  BUFFD0 U2295 ( .I(n2413), .Z(n2414) );
  CKBD0 U2296 ( .CLK(n2414), .C(n2415) );
  CKBD0 U2297 ( .CLK(n2415), .C(n2416) );
  CKBD0 U2298 ( .CLK(n2416), .C(n2417) );
  CKBD0 U2299 ( .CLK(n2417), .C(n2418) );
  CKBD0 U2300 ( .CLK(n2418), .C(n2419) );
  CKBD0 U2301 ( .CLK(n2419), .C(n2420) );
  CKBD0 U2302 ( .CLK(n2420), .C(n2421) );
  CKBD0 U2303 ( .CLK(n2421), .C(n2422) );
  CKBD0 U2304 ( .CLK(n2422), .C(n2423) );
  CKBD0 U2305 ( .CLK(n2423), .C(n2424) );
  BUFFD0 U2306 ( .I(n2424), .Z(n2425) );
  CKBD0 U2307 ( .CLK(n2425), .C(n2426) );
  CKBD0 U2308 ( .CLK(n2426), .C(n2427) );
  CKBD0 U2309 ( .CLK(n2427), .C(n2428) );
  CKBD0 U2310 ( .CLK(n2428), .C(n2429) );
  CKBD0 U2311 ( .CLK(n2429), .C(n2430) );
  CKBD0 U2312 ( .CLK(n2430), .C(n2431) );
  CKBD0 U2313 ( .CLK(n2431), .C(n2432) );
  CKBD0 U2314 ( .CLK(n2432), .C(n2433) );
  CKBD0 U2315 ( .CLK(n2433), .C(n2434) );
  CKBD0 U2316 ( .CLK(n2434), .C(n2435) );
  BUFFD0 U2317 ( .I(n2435), .Z(n2436) );
  CKBD0 U2318 ( .CLK(n2436), .C(n2437) );
  CKBD0 U2319 ( .CLK(n2437), .C(n2438) );
  CKBD0 U2320 ( .CLK(n2438), .C(n2439) );
  CKBD0 U2321 ( .CLK(n2439), .C(n2440) );
  CKBD0 U2322 ( .CLK(n2440), .C(n2441) );
  CKBD0 U2323 ( .CLK(n2441), .C(n2442) );
  CKBD0 U2324 ( .CLK(n2442), .C(n2443) );
  CKBD0 U2325 ( .CLK(n2443), .C(n2444) );
  CKBD0 U2326 ( .CLK(n2444), .C(n2445) );
  BUFFD0 U2327 ( .I(n2445), .Z(n2446) );
  CKBD0 U2328 ( .CLK(n2446), .C(n2447) );
  CKBD0 U2329 ( .CLK(n2447), .C(n2448) );
  CKBD0 U2330 ( .CLK(n2448), .C(n2449) );
  CKBD0 U2331 ( .CLK(n2449), .C(n2450) );
  CKBD0 U2332 ( .CLK(n2450), .C(n2451) );
  CKBD0 U2333 ( .CLK(n2451), .C(n2452) );
  CKBD0 U2334 ( .CLK(n2452), .C(n2453) );
  CKBD0 U2335 ( .CLK(n2453), .C(n2454) );
  CKBD0 U2336 ( .CLK(n2454), .C(n2455) );
  BUFFD0 U2337 ( .I(n2455), .Z(n2456) );
  BUFFD0 U2338 ( .I(n9013), .Z(n2457) );
  CKBD0 U2339 ( .CLK(FrameSR[16]), .C(n2458) );
  BUFFD0 U2340 ( .I(n2458), .Z(n2459) );
  CKBD0 U2341 ( .CLK(n2459), .C(n2460) );
  CKBD0 U2342 ( .CLK(n2460), .C(n2461) );
  CKBD0 U2343 ( .CLK(n2461), .C(n2462) );
  CKBD0 U2344 ( .CLK(n2462), .C(n2463) );
  CKBD0 U2345 ( .CLK(n2463), .C(n2464) );
  CKBD0 U2346 ( .CLK(n2464), .C(n2465) );
  CKBD0 U2347 ( .CLK(n2465), .C(n2466) );
  CKBD0 U2348 ( .CLK(n2466), .C(n2467) );
  CKBD0 U2349 ( .CLK(n2467), .C(n2468) );
  CKBD0 U2350 ( .CLK(n2468), .C(n2469) );
  BUFFD0 U2351 ( .I(n2469), .Z(n2470) );
  CKBD0 U2352 ( .CLK(n2470), .C(n2471) );
  CKBD0 U2353 ( .CLK(n2471), .C(n2472) );
  CKBD0 U2354 ( .CLK(n2472), .C(n2473) );
  CKBD0 U2355 ( .CLK(n2473), .C(n2474) );
  CKBD0 U2356 ( .CLK(n2474), .C(n2475) );
  CKBD0 U2357 ( .CLK(n2475), .C(n2476) );
  CKBD0 U2358 ( .CLK(n2476), .C(n2477) );
  CKBD0 U2359 ( .CLK(n2477), .C(n2478) );
  CKBD0 U2360 ( .CLK(n2478), .C(n2479) );
  CKBD0 U2361 ( .CLK(n2479), .C(n2480) );
  BUFFD0 U2362 ( .I(n2480), .Z(n2481) );
  CKBD0 U2363 ( .CLK(n2481), .C(n2482) );
  CKBD0 U2364 ( .CLK(n2482), .C(n2483) );
  CKBD0 U2365 ( .CLK(n2483), .C(n2484) );
  CKBD0 U2366 ( .CLK(n2484), .C(n2485) );
  CKBD0 U2367 ( .CLK(n2485), .C(n2486) );
  CKBD0 U2368 ( .CLK(n2486), .C(n2487) );
  CKBD0 U2369 ( .CLK(n2487), .C(n2488) );
  CKBD0 U2370 ( .CLK(n2488), .C(n2489) );
  CKBD0 U2371 ( .CLK(n2489), .C(n2490) );
  CKBD0 U2372 ( .CLK(n2490), .C(n2491) );
  BUFFD0 U2373 ( .I(n2491), .Z(n2492) );
  CKBD0 U2374 ( .CLK(n2492), .C(n2493) );
  CKBD0 U2375 ( .CLK(n2493), .C(n2494) );
  CKBD0 U2376 ( .CLK(n2494), .C(n2495) );
  CKBD0 U2377 ( .CLK(n2495), .C(n2496) );
  CKBD0 U2378 ( .CLK(n2496), .C(n2497) );
  CKBD0 U2379 ( .CLK(n2497), .C(n2498) );
  CKBD0 U2380 ( .CLK(n2498), .C(n2499) );
  CKBD0 U2381 ( .CLK(n2499), .C(n2500) );
  CKBD0 U2382 ( .CLK(n2500), .C(n2501) );
  BUFFD0 U2383 ( .I(n2501), .Z(n2502) );
  CKBD0 U2384 ( .CLK(n2502), .C(n2503) );
  CKBD0 U2385 ( .CLK(n2503), .C(n2504) );
  CKBD0 U2386 ( .CLK(n2504), .C(n2505) );
  CKBD0 U2387 ( .CLK(n2505), .C(n2506) );
  CKBD0 U2388 ( .CLK(n2506), .C(n2507) );
  CKBD0 U2389 ( .CLK(n2507), .C(n2508) );
  CKBD0 U2390 ( .CLK(n2508), .C(n2509) );
  CKBD0 U2391 ( .CLK(n2509), .C(n2510) );
  CKBD0 U2392 ( .CLK(n2510), .C(n2511) );
  CKBD0 U2393 ( .CLK(n2511), .C(n2512) );
  BUFFD0 U2394 ( .I(n2512), .Z(n2513) );
  CKBD0 U2395 ( .CLK(n2513), .C(n2514) );
  CKBD0 U2396 ( .CLK(n2514), .C(n2515) );
  CKBD0 U2397 ( .CLK(n2515), .C(n2516) );
  CKBD0 U2398 ( .CLK(n2516), .C(n2517) );
  CKBD0 U2399 ( .CLK(n2517), .C(n2518) );
  CKBD0 U2400 ( .CLK(n2518), .C(n2519) );
  CKBD0 U2401 ( .CLK(n2519), .C(n2520) );
  CKBD0 U2402 ( .CLK(n2520), .C(n2521) );
  CKBD0 U2403 ( .CLK(n2521), .C(n2522) );
  CKBD0 U2404 ( .CLK(n2522), .C(n2523) );
  BUFFD0 U2405 ( .I(n2523), .Z(n2524) );
  CKBD0 U2406 ( .CLK(n2524), .C(n2525) );
  CKBD0 U2407 ( .CLK(n2525), .C(n2526) );
  CKBD0 U2408 ( .CLK(n2526), .C(n2527) );
  CKBD0 U2409 ( .CLK(n2527), .C(n2528) );
  CKBD0 U2410 ( .CLK(n2528), .C(n2529) );
  CKBD0 U2411 ( .CLK(n2529), .C(n2530) );
  CKBD0 U2412 ( .CLK(n2530), .C(n2531) );
  CKBD0 U2413 ( .CLK(n2531), .C(n2532) );
  CKBD0 U2414 ( .CLK(n2532), .C(n2533) );
  CKBD0 U2415 ( .CLK(n2533), .C(n2534) );
  BUFFD0 U2416 ( .I(n2534), .Z(n2535) );
  CKBD0 U2417 ( .CLK(n2535), .C(n2536) );
  CKBD0 U2418 ( .CLK(n2536), .C(n2537) );
  CKBD0 U2419 ( .CLK(n2537), .C(n2538) );
  CKBD0 U2420 ( .CLK(n2538), .C(n2539) );
  CKBD0 U2421 ( .CLK(n2539), .C(n2540) );
  CKBD0 U2422 ( .CLK(n2540), .C(n2541) );
  CKBD0 U2423 ( .CLK(n2541), .C(n2542) );
  CKBD0 U2424 ( .CLK(n2542), .C(n2543) );
  CKBD0 U2425 ( .CLK(n2543), .C(n2544) );
  CKBD0 U2426 ( .CLK(n2544), .C(n2545) );
  BUFFD0 U2427 ( .I(n2545), .Z(n2546) );
  CKBD0 U2428 ( .CLK(n2546), .C(n2547) );
  CKBD0 U2429 ( .CLK(n2547), .C(n2548) );
  CKBD0 U2430 ( .CLK(n2548), .C(n2549) );
  CKBD0 U2431 ( .CLK(n2549), .C(n2550) );
  CKBD0 U2432 ( .CLK(n2550), .C(n2551) );
  CKBD0 U2433 ( .CLK(n2551), .C(n2552) );
  CKBD0 U2434 ( .CLK(n2552), .C(n2553) );
  BUFFD0 U2435 ( .I(n5956), .Z(n2554) );
  CKBD0 U2436 ( .CLK(FrameSR[15]), .C(n2555) );
  BUFFD0 U2437 ( .I(N42), .Z(n2556) );
  BUFFD0 U2438 ( .I(n2688), .Z(n2557) );
  CKBD0 U2439 ( .CLK(FrameSR[63]), .C(n2558) );
  CKBD0 U2440 ( .CLK(n2558), .C(n2559) );
  CKBD0 U2441 ( .CLK(n2559), .C(n2560) );
  CKBD0 U2442 ( .CLK(n2560), .C(n2561) );
  CKBD0 U2443 ( .CLK(n2561), .C(n2562) );
  CKBD0 U2444 ( .CLK(n2562), .C(n2563) );
  CKBD0 U2445 ( .CLK(n2563), .C(n2564) );
  CKBD0 U2446 ( .CLK(n2564), .C(n2565) );
  CKBD0 U2447 ( .CLK(n2565), .C(n2566) );
  CKBD0 U2448 ( .CLK(n2566), .C(n2567) );
  BUFFD0 U2449 ( .I(n2567), .Z(n2568) );
  CKBD0 U2450 ( .CLK(n2568), .C(n2569) );
  CKBD0 U2451 ( .CLK(n2569), .C(n2570) );
  CKBD0 U2452 ( .CLK(n2570), .C(n2571) );
  CKBD0 U2453 ( .CLK(n2571), .C(n2572) );
  CKBD0 U2454 ( .CLK(n2572), .C(n2573) );
  CKBD0 U2455 ( .CLK(n2573), .C(n2574) );
  CKBD0 U2456 ( .CLK(n2574), .C(n2575) );
  CKBD0 U2457 ( .CLK(n2575), .C(n2576) );
  CKBD0 U2458 ( .CLK(n2576), .C(n2577) );
  CKBD0 U2459 ( .CLK(n2577), .C(n2578) );
  BUFFD0 U2460 ( .I(n2578), .Z(n2579) );
  CKBD0 U2461 ( .CLK(n2579), .C(n2580) );
  CKBD0 U2462 ( .CLK(n2580), .C(n2581) );
  CKBD0 U2463 ( .CLK(n2581), .C(n2582) );
  CKBD0 U2464 ( .CLK(n2582), .C(n2583) );
  CKBD0 U2465 ( .CLK(n2583), .C(n2584) );
  CKBD0 U2466 ( .CLK(n2584), .C(n2585) );
  CKBD0 U2467 ( .CLK(n2585), .C(n2586) );
  CKBD0 U2468 ( .CLK(n2586), .C(n2587) );
  CKBD0 U2469 ( .CLK(n2587), .C(n2588) );
  CKBD0 U2470 ( .CLK(n2588), .C(n2589) );
  BUFFD0 U2471 ( .I(n2589), .Z(n2590) );
  CKBD0 U2472 ( .CLK(n2590), .C(n2591) );
  CKBD0 U2473 ( .CLK(n2591), .C(n2592) );
  CKBD0 U2474 ( .CLK(n2592), .C(n2593) );
  CKBD0 U2475 ( .CLK(n2593), .C(n2594) );
  CKBD0 U2476 ( .CLK(n2594), .C(n2595) );
  CKBD0 U2477 ( .CLK(n2595), .C(n2596) );
  CKBD0 U2478 ( .CLK(n2596), .C(n2597) );
  CKBD0 U2479 ( .CLK(n2597), .C(n2598) );
  CKBD0 U2480 ( .CLK(n2598), .C(n2599) );
  CKBD0 U2481 ( .CLK(n2599), .C(n2600) );
  BUFFD0 U2482 ( .I(n2600), .Z(n2601) );
  CKBD0 U2483 ( .CLK(n2601), .C(n2602) );
  CKBD0 U2484 ( .CLK(n2602), .C(n2603) );
  CKBD0 U2485 ( .CLK(n2603), .C(n2604) );
  CKBD0 U2486 ( .CLK(n2604), .C(n2605) );
  CKBD0 U2487 ( .CLK(n2605), .C(n2606) );
  CKBD0 U2488 ( .CLK(n2606), .C(n2607) );
  CKBD0 U2489 ( .CLK(n2607), .C(n2608) );
  CKBD0 U2490 ( .CLK(n2608), .C(n2609) );
  CKBD0 U2491 ( .CLK(n2609), .C(n2610) );
  CKBD0 U2492 ( .CLK(n2610), .C(n2611) );
  BUFFD0 U2493 ( .I(n2611), .Z(n2612) );
  CKBD0 U2494 ( .CLK(n2612), .C(n2613) );
  CKBD0 U2495 ( .CLK(n2613), .C(n2614) );
  CKBD0 U2496 ( .CLK(n2614), .C(n2615) );
  CKBD0 U2497 ( .CLK(n2615), .C(n2616) );
  CKBD0 U2498 ( .CLK(n2616), .C(n2617) );
  CKBD0 U2499 ( .CLK(n2617), .C(n2618) );
  CKBD0 U2500 ( .CLK(n2618), .C(n2619) );
  CKBD0 U2501 ( .CLK(n2619), .C(n2620) );
  CKBD0 U2502 ( .CLK(n2620), .C(n2621) );
  CKBD0 U2503 ( .CLK(n2621), .C(n2622) );
  BUFFD0 U2504 ( .I(n2622), .Z(n2623) );
  CKBD0 U2505 ( .CLK(n2623), .C(n2624) );
  CKBD0 U2506 ( .CLK(n2624), .C(n2625) );
  CKBD0 U2507 ( .CLK(n2625), .C(n2626) );
  CKBD0 U2508 ( .CLK(n2626), .C(n2627) );
  CKBD0 U2509 ( .CLK(n2627), .C(n2628) );
  CKBD0 U2510 ( .CLK(n2628), .C(n2629) );
  CKBD0 U2511 ( .CLK(n2629), .C(n2630) );
  CKBD0 U2512 ( .CLK(n2630), .C(n2631) );
  CKBD0 U2513 ( .CLK(n2631), .C(n2632) );
  BUFFD0 U2514 ( .I(n2632), .Z(n2633) );
  CKBD0 U2515 ( .CLK(n2633), .C(n2634) );
  CKBD0 U2516 ( .CLK(n2634), .C(n2635) );
  CKBD0 U2517 ( .CLK(n2635), .C(n2636) );
  CKBD0 U2518 ( .CLK(n2636), .C(n2637) );
  CKBD0 U2519 ( .CLK(n2637), .C(n2638) );
  CKBD0 U2520 ( .CLK(n2638), .C(n2639) );
  CKBD0 U2521 ( .CLK(n2639), .C(n2640) );
  CKBD0 U2522 ( .CLK(n2640), .C(n2641) );
  CKBD0 U2523 ( .CLK(n2641), .C(n2642) );
  CKBD0 U2524 ( .CLK(n2642), .C(n2643) );
  BUFFD0 U2525 ( .I(n2643), .Z(n2644) );
  CKBD0 U2526 ( .CLK(n2644), .C(n2645) );
  CKBD0 U2527 ( .CLK(n2645), .C(n2646) );
  CKBD0 U2528 ( .CLK(n2646), .C(n2647) );
  CKBD0 U2529 ( .CLK(n2647), .C(n2648) );
  CKBD0 U2530 ( .CLK(n2648), .C(n2649) );
  CKBD0 U2531 ( .CLK(n2649), .C(n2650) );
  CKBD0 U2532 ( .CLK(n2650), .C(n2651) );
  CKBD0 U2533 ( .CLK(n2651), .C(n2652) );
  CKBD0 U2534 ( .CLK(n2652), .C(n2653) );
  CKBD0 U2535 ( .CLK(n2653), .C(n2654) );
  BUFFD0 U2536 ( .I(n2654), .Z(n2655) );
  CKBD0 U2537 ( .CLK(n2655), .C(n2656) );
  CKBD0 U2538 ( .CLK(n2656), .C(n2657) );
  CKBD0 U2539 ( .CLK(n2657), .C(n2658) );
  CKBD0 U2540 ( .CLK(n2658), .C(n2659) );
  BUFFD0 U2541 ( .I(n2659), .Z(n2660) );
  CKBD0 U2542 ( .CLK(n2660), .C(n2661) );
  BUFFD0 U2543 ( .I(n2661), .Z(n2662) );
  CKBD0 U2544 ( .CLK(n2662), .C(n2663) );
  BUFFD0 U2545 ( .I(n2663), .Z(n2664) );
  CKBD0 U2546 ( .CLK(n2664), .C(n2665) );
  BUFFD0 U2547 ( .I(n2665), .Z(n2666) );
  CKBD0 U2548 ( .CLK(n2666), .C(n2667) );
  BUFFD0 U2549 ( .I(n2667), .Z(n2668) );
  CKBD0 U2550 ( .CLK(n2668), .C(n2669) );
  BUFFD0 U2551 ( .I(n2669), .Z(n2670) );
  CKBD0 U2552 ( .CLK(n2670), .C(n2671) );
  BUFFD0 U2553 ( .I(n2671), .Z(n2672) );
  CKBD0 U2554 ( .CLK(n2672), .C(n2673) );
  BUFFD0 U2555 ( .I(n2673), .Z(n2674) );
  CKBD0 U2556 ( .CLK(n2674), .C(n2675) );
  BUFFD0 U2557 ( .I(n2675), .Z(n2676) );
  CKBD0 U2558 ( .CLK(n2676), .C(n2677) );
  BUFFD0 U2559 ( .I(n2677), .Z(n2678) );
  CKBD0 U2560 ( .CLK(n2678), .C(n2679) );
  BUFFD0 U2561 ( .I(n2679), .Z(n2680) );
  CKBD0 U2562 ( .CLK(n2680), .C(n2681) );
  BUFFD0 U2563 ( .I(n2681), .Z(n2682) );
  CKBD0 U2564 ( .CLK(n2682), .C(n2683) );
  BUFFD0 U2565 ( .I(n2683), .Z(n2684) );
  CKBD0 U2566 ( .CLK(n2684), .C(n2685) );
  BUFFD0 U2567 ( .I(n2685), .Z(n2686) );
  CKBD0 U2568 ( .CLK(n2686), .C(n2687) );
  BUFFD0 U2569 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2570 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2571 ( .I(n9158), .Z(n2690) );
  BUFFD0 U2572 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2573 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2574 ( .I(n9159), .Z(n2693) );
  CKBD0 U2575 ( .CLK(n5), .C(n2694) );
  CKBD0 U2576 ( .CLK(n2694), .C(n2695) );
  CKBD0 U2577 ( .CLK(n2695), .C(n2696) );
  BUFFD0 U2578 ( .I(n2696), .Z(n2697) );
  CKBD0 U2579 ( .CLK(n2697), .C(n2698) );
  CKBD0 U2580 ( .CLK(n2698), .C(n2699) );
  CKBD0 U2581 ( .CLK(n2699), .C(n2700) );
  CKBD0 U2582 ( .CLK(n2700), .C(n2701) );
  CKBD0 U2583 ( .CLK(n2701), .C(n2702) );
  CKBD0 U2584 ( .CLK(n2702), .C(n2703) );
  CKBD0 U2585 ( .CLK(n2703), .C(n2704) );
  CKBD0 U2586 ( .CLK(n2704), .C(n2705) );
  CKBD0 U2587 ( .CLK(n2705), .C(n2706) );
  CKBD0 U2588 ( .CLK(n2706), .C(n2707) );
  BUFFD0 U2589 ( .I(n2707), .Z(n2708) );
  CKBD0 U2590 ( .CLK(n2708), .C(n2709) );
  CKBD0 U2591 ( .CLK(n2709), .C(n2710) );
  CKBD0 U2592 ( .CLK(n2710), .C(n2711) );
  CKBD0 U2593 ( .CLK(n2711), .C(n2712) );
  CKBD0 U2594 ( .CLK(n2712), .C(n2713) );
  CKBD0 U2595 ( .CLK(n2713), .C(n2714) );
  CKBD0 U2596 ( .CLK(n2714), .C(n2715) );
  CKBD0 U2597 ( .CLK(n2715), .C(n2716) );
  CKBD0 U2598 ( .CLK(n2716), .C(n2717) );
  BUFFD0 U2599 ( .I(n2717), .Z(n2718) );
  CKBD0 U2600 ( .CLK(n2718), .C(n2719) );
  CKBD0 U2601 ( .CLK(n2719), .C(n2720) );
  CKBD0 U2602 ( .CLK(n2720), .C(n2721) );
  CKBD0 U2603 ( .CLK(n2721), .C(n2722) );
  CKBD0 U2604 ( .CLK(n2722), .C(n2723) );
  CKBD0 U2605 ( .CLK(n2723), .C(n2724) );
  CKBD0 U2606 ( .CLK(n2724), .C(n2725) );
  CKBD0 U2607 ( .CLK(n2725), .C(n2726) );
  CKBD0 U2608 ( .CLK(n2726), .C(n2727) );
  CKBD0 U2609 ( .CLK(n2727), .C(n2728) );
  BUFFD0 U2610 ( .I(n2728), .Z(n2729) );
  CKBD0 U2611 ( .CLK(n2729), .C(n2730) );
  CKBD0 U2612 ( .CLK(n2730), .C(n2731) );
  CKBD0 U2613 ( .CLK(n2731), .C(n2732) );
  CKBD0 U2614 ( .CLK(n2732), .C(n2733) );
  CKBD0 U2615 ( .CLK(n2733), .C(n2734) );
  CKBD0 U2616 ( .CLK(n2734), .C(n2735) );
  CKBD0 U2617 ( .CLK(n2735), .C(n2736) );
  CKBD0 U2618 ( .CLK(n2736), .C(n2737) );
  CKBD0 U2619 ( .CLK(n2737), .C(n2738) );
  CKBD0 U2620 ( .CLK(n2738), .C(n2739) );
  BUFFD0 U2621 ( .I(n2739), .Z(n2740) );
  CKBD0 U2622 ( .CLK(n2740), .C(n2741) );
  CKBD0 U2623 ( .CLK(n2741), .C(n2742) );
  CKBD0 U2624 ( .CLK(n2742), .C(n2743) );
  CKBD0 U2625 ( .CLK(n2743), .C(n2744) );
  CKBD0 U2626 ( .CLK(n2744), .C(n2745) );
  CKBD0 U2627 ( .CLK(n2745), .C(n2746) );
  CKBD0 U2628 ( .CLK(n2746), .C(n2747) );
  CKBD0 U2629 ( .CLK(n2747), .C(n2748) );
  CKBD0 U2630 ( .CLK(n2748), .C(n2749) );
  CKBD0 U2631 ( .CLK(n2749), .C(n2750) );
  BUFFD0 U2632 ( .I(n2750), .Z(n2751) );
  CKBD0 U2633 ( .CLK(n2751), .C(n2752) );
  CKBD0 U2634 ( .CLK(n2752), .C(n2753) );
  CKBD0 U2635 ( .CLK(n2753), .C(n2754) );
  CKBD0 U2636 ( .CLK(n2754), .C(n2755) );
  CKBD0 U2637 ( .CLK(n2755), .C(n2756) );
  CKBD0 U2638 ( .CLK(n2756), .C(n2757) );
  CKBD0 U2639 ( .CLK(n2757), .C(n2758) );
  CKBD0 U2640 ( .CLK(n2758), .C(n2759) );
  CKBD0 U2641 ( .CLK(n2759), .C(n2760) );
  CKBD0 U2642 ( .CLK(n2760), .C(n2761) );
  BUFFD0 U2643 ( .I(n2761), .Z(n2762) );
  CKBD0 U2644 ( .CLK(n2762), .C(n2763) );
  CKBD0 U2645 ( .CLK(n2763), .C(n2764) );
  CKBD0 U2646 ( .CLK(n2764), .C(n2765) );
  CKBD0 U2647 ( .CLK(n2765), .C(n2766) );
  CKBD0 U2648 ( .CLK(n2766), .C(n2767) );
  CKBD0 U2649 ( .CLK(n2767), .C(n2768) );
  CKBD0 U2650 ( .CLK(n2768), .C(n2769) );
  CKBD0 U2651 ( .CLK(n2769), .C(n2770) );
  CKBD0 U2652 ( .CLK(n2770), .C(n2771) );
  CKBD0 U2653 ( .CLK(n2771), .C(n2772) );
  BUFFD0 U2654 ( .I(n2772), .Z(n2773) );
  CKBD0 U2655 ( .CLK(n2773), .C(n2774) );
  CKBD0 U2656 ( .CLK(n2774), .C(n2775) );
  CKBD0 U2657 ( .CLK(n2775), .C(n2776) );
  CKBD0 U2658 ( .CLK(n2776), .C(n2777) );
  CKBD0 U2659 ( .CLK(n2777), .C(n2778) );
  CKBD0 U2660 ( .CLK(n2778), .C(n2779) );
  CKBD0 U2661 ( .CLK(n2779), .C(n2780) );
  CKBD0 U2662 ( .CLK(n2780), .C(n2781) );
  CKBD0 U2663 ( .CLK(n2781), .C(n2782) );
  BUFFD0 U2664 ( .I(n2782), .Z(n2783) );
  CKBD0 U2665 ( .CLK(n2783), .C(n2784) );
  CKBD0 U2666 ( .CLK(n2784), .C(n2785) );
  CKBD0 U2667 ( .CLK(n2785), .C(n2786) );
  CKBD0 U2668 ( .CLK(n2786), .C(n2787) );
  CKBD0 U2669 ( .CLK(n2787), .C(n2788) );
  CKBD0 U2670 ( .CLK(n2788), .C(n2789) );
  CKBD0 U2671 ( .CLK(n2789), .C(n2790) );
  CKBD0 U2672 ( .CLK(n2790), .C(n2791) );
  CKBD0 U2673 ( .CLK(n2791), .C(n2792) );
  CKBD0 U2674 ( .CLK(n2792), .C(n2793) );
  BUFFD0 U2675 ( .I(n2793), .Z(n2794) );
  CKBD0 U2676 ( .CLK(n2794), .C(n2795) );
  CKBD0 U2677 ( .CLK(n2795), .C(n2796) );
  CKBD0 U2678 ( .CLK(n2796), .C(n2797) );
  CKBD0 U2679 ( .CLK(n2797), .C(n2798) );
  CKBD0 U2680 ( .CLK(n2798), .C(n2799) );
  CKBD0 U2681 ( .CLK(n2799), .C(n2800) );
  CKBD0 U2682 ( .CLK(n2800), .C(n2801) );
  CKBD0 U2683 ( .CLK(n2801), .C(n2802) );
  CKBD0 U2684 ( .CLK(n2802), .C(n2803) );
  CKBD0 U2685 ( .CLK(n2803), .C(n2804) );
  BUFFD0 U2686 ( .I(n2804), .Z(n2805) );
  CKBD0 U2687 ( .CLK(n2805), .C(n2806) );
  CKBD0 U2688 ( .CLK(n2806), .C(n2807) );
  CKBD0 U2689 ( .CLK(n2807), .C(n2808) );
  CKBD0 U2690 ( .CLK(n2808), .C(n2809) );
  CKBD0 U2691 ( .CLK(n2809), .C(n2810) );
  CKBD0 U2692 ( .CLK(n2810), .C(n2811) );
  BUFFD0 U2693 ( .I(n2811), .Z(n2812) );
  CKBD0 U2694 ( .CLK(n2812), .C(n2813) );
  BUFFD0 U2695 ( .I(n2813), .Z(n2814) );
  CKBD0 U2696 ( .CLK(n2814), .C(n2815) );
  BUFFD0 U2697 ( .I(n2815), .Z(n2816) );
  CKBD0 U2698 ( .CLK(n2816), .C(n2817) );
  BUFFD0 U2699 ( .I(n2817), .Z(n2818) );
  CKBD0 U2700 ( .CLK(n2818), .C(n2819) );
  BUFFD0 U2701 ( .I(n2819), .Z(n2820) );
  CKBD0 U2702 ( .CLK(n2820), .C(n2821) );
  BUFFD0 U2703 ( .I(n2821), .Z(n2822) );
  CKBD0 U2704 ( .CLK(n2822), .C(n2823) );
  BUFFD0 U2705 ( .I(n2823), .Z(n2824) );
  CKBD0 U2706 ( .CLK(n2824), .C(n2825) );
  BUFFD0 U2707 ( .I(n2825), .Z(n2826) );
  BUFFD0 U2708 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2709 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2710 ( .I(n9160), .Z(n2829) );
  CKBD0 U2711 ( .CLK(n1364), .C(n2830) );
  CKBD0 U2712 ( .CLK(n2830), .C(n2831) );
  CKBD0 U2713 ( .CLK(n2831), .C(n2832) );
  BUFFD0 U2714 ( .I(n2832), .Z(n2833) );
  CKBD0 U2715 ( .CLK(n2833), .C(n2834) );
  CKBD0 U2716 ( .CLK(n2834), .C(n2835) );
  CKBD0 U2717 ( .CLK(n2835), .C(n2836) );
  CKBD0 U2718 ( .CLK(n2836), .C(n2837) );
  CKBD0 U2719 ( .CLK(n2837), .C(n2838) );
  CKBD0 U2720 ( .CLK(n2838), .C(n2839) );
  CKBD0 U2721 ( .CLK(n2839), .C(n2840) );
  CKBD0 U2722 ( .CLK(n2840), .C(n2841) );
  CKBD0 U2723 ( .CLK(n2841), .C(n2842) );
  CKBD0 U2724 ( .CLK(n2842), .C(n2843) );
  BUFFD0 U2725 ( .I(n2843), .Z(n2844) );
  CKBD0 U2726 ( .CLK(n2844), .C(n2845) );
  CKBD0 U2727 ( .CLK(n2845), .C(n2846) );
  CKBD0 U2728 ( .CLK(n2846), .C(n2847) );
  CKBD0 U2729 ( .CLK(n2847), .C(n2848) );
  CKBD0 U2730 ( .CLK(n2848), .C(n2849) );
  CKBD0 U2731 ( .CLK(n2849), .C(n2850) );
  CKBD0 U2732 ( .CLK(n2850), .C(n2851) );
  CKBD0 U2733 ( .CLK(n2851), .C(n2852) );
  CKBD0 U2734 ( .CLK(n2852), .C(n2853) );
  BUFFD0 U2735 ( .I(n2853), .Z(n2854) );
  CKBD0 U2736 ( .CLK(n2854), .C(n2855) );
  CKBD0 U2737 ( .CLK(n2855), .C(n2856) );
  CKBD0 U2738 ( .CLK(n2856), .C(n2857) );
  CKBD0 U2739 ( .CLK(n2857), .C(n2858) );
  CKBD0 U2740 ( .CLK(n2858), .C(n2859) );
  CKBD0 U2741 ( .CLK(n2859), .C(n2860) );
  CKBD0 U2742 ( .CLK(n2860), .C(n2861) );
  CKBD0 U2743 ( .CLK(n2861), .C(n2862) );
  CKBD0 U2744 ( .CLK(n2862), .C(n2863) );
  CKBD0 U2745 ( .CLK(n2863), .C(n2864) );
  BUFFD0 U2746 ( .I(n2864), .Z(n2865) );
  CKBD0 U2747 ( .CLK(n2865), .C(n2866) );
  CKBD0 U2748 ( .CLK(n2866), .C(n2867) );
  CKBD0 U2749 ( .CLK(n2867), .C(n2868) );
  CKBD0 U2750 ( .CLK(n2868), .C(n2869) );
  CKBD0 U2751 ( .CLK(n2869), .C(n2870) );
  CKBD0 U2752 ( .CLK(n2870), .C(n2871) );
  CKBD0 U2753 ( .CLK(n2871), .C(n2872) );
  CKBD0 U2754 ( .CLK(n2872), .C(n2873) );
  CKBD0 U2755 ( .CLK(n2873), .C(n2874) );
  CKBD0 U2756 ( .CLK(n2874), .C(n2875) );
  BUFFD0 U2757 ( .I(n2875), .Z(n2876) );
  CKBD0 U2758 ( .CLK(n2876), .C(n2877) );
  CKBD0 U2759 ( .CLK(n2877), .C(n2878) );
  CKBD0 U2760 ( .CLK(n2878), .C(n2879) );
  CKBD0 U2761 ( .CLK(n2879), .C(n2880) );
  CKBD0 U2762 ( .CLK(n2880), .C(n2881) );
  CKBD0 U2763 ( .CLK(n2881), .C(n2882) );
  CKBD0 U2764 ( .CLK(n2882), .C(n2883) );
  CKBD0 U2765 ( .CLK(n2883), .C(n2884) );
  CKBD0 U2766 ( .CLK(n2884), .C(n2885) );
  CKBD0 U2767 ( .CLK(n2885), .C(n2886) );
  BUFFD0 U2768 ( .I(n2886), .Z(n2887) );
  CKBD0 U2769 ( .CLK(n2887), .C(n2888) );
  CKBD0 U2770 ( .CLK(n2888), .C(n2889) );
  CKBD0 U2771 ( .CLK(n2889), .C(n2890) );
  CKBD0 U2772 ( .CLK(n2890), .C(n2891) );
  CKBD0 U2773 ( .CLK(n2891), .C(n2892) );
  CKBD0 U2774 ( .CLK(n2892), .C(n2893) );
  CKBD0 U2775 ( .CLK(n2893), .C(n2894) );
  CKBD0 U2776 ( .CLK(n2894), .C(n2895) );
  CKBD0 U2777 ( .CLK(n2895), .C(n2896) );
  CKBD0 U2778 ( .CLK(n2896), .C(n2897) );
  BUFFD0 U2779 ( .I(n2897), .Z(n2898) );
  CKBD0 U2780 ( .CLK(n2898), .C(n2899) );
  CKBD0 U2781 ( .CLK(n2899), .C(n2900) );
  CKBD0 U2782 ( .CLK(n2900), .C(n2901) );
  CKBD0 U2783 ( .CLK(n2901), .C(n2902) );
  CKBD0 U2784 ( .CLK(n2902), .C(n2903) );
  CKBD0 U2785 ( .CLK(n2903), .C(n2904) );
  CKBD0 U2786 ( .CLK(n2904), .C(n2905) );
  CKBD0 U2787 ( .CLK(n2905), .C(n2906) );
  CKBD0 U2788 ( .CLK(n2906), .C(n2907) );
  CKBD0 U2789 ( .CLK(n2907), .C(n2908) );
  BUFFD0 U2790 ( .I(n2908), .Z(n2909) );
  CKBD0 U2791 ( .CLK(n2909), .C(n2910) );
  CKBD0 U2792 ( .CLK(n2910), .C(n2911) );
  CKBD0 U2793 ( .CLK(n2911), .C(n2912) );
  CKBD0 U2794 ( .CLK(n2912), .C(n2913) );
  CKBD0 U2795 ( .CLK(n2913), .C(n2914) );
  CKBD0 U2796 ( .CLK(n2914), .C(n2915) );
  CKBD0 U2797 ( .CLK(n2915), .C(n2916) );
  CKBD0 U2798 ( .CLK(n2916), .C(n2917) );
  CKBD0 U2799 ( .CLK(n2917), .C(n2918) );
  CKBD0 U2800 ( .CLK(n2918), .C(n2919) );
  BUFFD0 U2801 ( .I(n2919), .Z(n2920) );
  CKBD0 U2802 ( .CLK(n2920), .C(n2921) );
  CKBD0 U2803 ( .CLK(n2921), .C(n2922) );
  CKBD0 U2804 ( .CLK(n2922), .C(n2923) );
  CKBD0 U2805 ( .CLK(n2923), .C(n2924) );
  CKBD0 U2806 ( .CLK(n2924), .C(n2925) );
  CKBD0 U2807 ( .CLK(n2925), .C(n2926) );
  CKBD0 U2808 ( .CLK(n2926), .C(n2927) );
  CKBD0 U2809 ( .CLK(n2927), .C(n2928) );
  CKBD0 U2810 ( .CLK(n2928), .C(n2929) );
  BUFFD0 U2811 ( .I(n2929), .Z(n2930) );
  CKBD0 U2812 ( .CLK(n2930), .C(n2931) );
  CKBD0 U2813 ( .CLK(n2931), .C(n2932) );
  CKBD0 U2814 ( .CLK(n2932), .C(n2933) );
  CKBD0 U2815 ( .CLK(n2933), .C(n2934) );
  CKBD0 U2816 ( .CLK(n2934), .C(n2935) );
  CKBD0 U2817 ( .CLK(n2935), .C(n2936) );
  CKBD0 U2818 ( .CLK(n2936), .C(n2937) );
  CKBD0 U2819 ( .CLK(n2937), .C(n2938) );
  CKBD0 U2820 ( .CLK(n2938), .C(n2939) );
  CKBD0 U2821 ( .CLK(n2939), .C(n2940) );
  BUFFD0 U2822 ( .I(n2940), .Z(n2941) );
  CKBD0 U2823 ( .CLK(n2941), .C(n2942) );
  CKBD0 U2824 ( .CLK(n2942), .C(n2943) );
  CKBD0 U2825 ( .CLK(n2943), .C(n2944) );
  CKBD0 U2826 ( .CLK(n2944), .C(n2945) );
  CKBD0 U2827 ( .CLK(n2945), .C(n2946) );
  CKBD0 U2828 ( .CLK(n2946), .C(n2947) );
  BUFFD0 U2829 ( .I(n2947), .Z(n2948) );
  CKBD0 U2830 ( .CLK(n2948), .C(n2949) );
  BUFFD0 U2831 ( .I(n2949), .Z(n2950) );
  CKBD0 U2832 ( .CLK(n2950), .C(n2951) );
  BUFFD0 U2833 ( .I(n2951), .Z(n2952) );
  CKBD0 U2834 ( .CLK(n2952), .C(n2953) );
  BUFFD0 U2835 ( .I(n2953), .Z(n2954) );
  CKBD0 U2836 ( .CLK(n2954), .C(n2955) );
  BUFFD0 U2837 ( .I(n2955), .Z(n2956) );
  CKBD0 U2838 ( .CLK(n2956), .C(n2957) );
  BUFFD0 U2839 ( .I(n2957), .Z(n2958) );
  CKBD0 U2840 ( .CLK(n2958), .C(n2959) );
  BUFFD0 U2841 ( .I(n2959), .Z(n2960) );
  CKBD0 U2842 ( .CLK(n2960), .C(n2961) );
  BUFFD0 U2843 ( .I(n2961), .Z(n2962) );
  BUFFD0 U2844 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2845 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2846 ( .I(n9161), .Z(n2965) );
  CKBD0 U2847 ( .CLK(n1362), .C(n2966) );
  CKBD0 U2848 ( .CLK(n2966), .C(n2967) );
  CKBD0 U2849 ( .CLK(n2967), .C(n2968) );
  BUFFD0 U2850 ( .I(n2968), .Z(n2969) );
  CKBD0 U2851 ( .CLK(n2969), .C(n2970) );
  CKBD0 U2852 ( .CLK(n2970), .C(n2971) );
  CKBD0 U2853 ( .CLK(n2971), .C(n2972) );
  CKBD0 U2854 ( .CLK(n2972), .C(n2973) );
  CKBD0 U2855 ( .CLK(n2973), .C(n2974) );
  CKBD0 U2856 ( .CLK(n2974), .C(n2975) );
  CKBD0 U2857 ( .CLK(n2975), .C(n2976) );
  CKBD0 U2858 ( .CLK(n2976), .C(n2977) );
  CKBD0 U2859 ( .CLK(n2977), .C(n2978) );
  CKBD0 U2860 ( .CLK(n2978), .C(n2979) );
  BUFFD0 U2861 ( .I(n2979), .Z(n2980) );
  CKBD0 U2862 ( .CLK(n2980), .C(n2981) );
  CKBD0 U2863 ( .CLK(n2981), .C(n2982) );
  CKBD0 U2864 ( .CLK(n2982), .C(n2983) );
  CKBD0 U2865 ( .CLK(n2983), .C(n2984) );
  CKBD0 U2866 ( .CLK(n2984), .C(n2985) );
  CKBD0 U2867 ( .CLK(n2985), .C(n2986) );
  CKBD0 U2868 ( .CLK(n2986), .C(n2987) );
  CKBD0 U2869 ( .CLK(n2987), .C(n2988) );
  CKBD0 U2870 ( .CLK(n2988), .C(n2989) );
  BUFFD0 U2871 ( .I(n2989), .Z(n2990) );
  CKBD0 U2872 ( .CLK(n2990), .C(n2991) );
  CKBD0 U2873 ( .CLK(n2991), .C(n2992) );
  CKBD0 U2874 ( .CLK(n2992), .C(n2993) );
  CKBD0 U2875 ( .CLK(n2993), .C(n2994) );
  CKBD0 U2876 ( .CLK(n2994), .C(n2995) );
  CKBD0 U2877 ( .CLK(n2995), .C(n2996) );
  CKBD0 U2878 ( .CLK(n2996), .C(n2997) );
  CKBD0 U2879 ( .CLK(n2997), .C(n2998) );
  CKBD0 U2880 ( .CLK(n2998), .C(n2999) );
  CKBD0 U2881 ( .CLK(n2999), .C(n3000) );
  BUFFD0 U2882 ( .I(n3000), .Z(n3001) );
  CKBD0 U2883 ( .CLK(n3001), .C(n3002) );
  CKBD0 U2884 ( .CLK(n3002), .C(n3003) );
  CKBD0 U2885 ( .CLK(n3003), .C(n3004) );
  CKBD0 U2886 ( .CLK(n3004), .C(n3005) );
  CKBD0 U2887 ( .CLK(n3005), .C(n3006) );
  CKBD0 U2888 ( .CLK(n3006), .C(n3007) );
  CKBD0 U2889 ( .CLK(n3007), .C(n3008) );
  CKBD0 U2890 ( .CLK(n3008), .C(n3009) );
  CKBD0 U2891 ( .CLK(n3009), .C(n3010) );
  CKBD0 U2892 ( .CLK(n3010), .C(n3011) );
  BUFFD0 U2893 ( .I(n3011), .Z(n3012) );
  CKBD0 U2894 ( .CLK(n3012), .C(n3013) );
  CKBD0 U2895 ( .CLK(n3013), .C(n3014) );
  CKBD0 U2896 ( .CLK(n3014), .C(n3015) );
  CKBD0 U2897 ( .CLK(n3015), .C(n3016) );
  CKBD0 U2898 ( .CLK(n3016), .C(n3017) );
  CKBD0 U2899 ( .CLK(n3017), .C(n3018) );
  CKBD0 U2900 ( .CLK(n3018), .C(n3019) );
  CKBD0 U2901 ( .CLK(n3019), .C(n3020) );
  CKBD0 U2902 ( .CLK(n3020), .C(n3021) );
  CKBD0 U2903 ( .CLK(n3021), .C(n3022) );
  BUFFD0 U2904 ( .I(n3022), .Z(n3023) );
  CKBD0 U2905 ( .CLK(n3023), .C(n3024) );
  CKBD0 U2906 ( .CLK(n3024), .C(n3025) );
  CKBD0 U2907 ( .CLK(n3025), .C(n3026) );
  CKBD0 U2908 ( .CLK(n3026), .C(n3027) );
  CKBD0 U2909 ( .CLK(n3027), .C(n3028) );
  CKBD0 U2910 ( .CLK(n3028), .C(n3029) );
  CKBD0 U2911 ( .CLK(n3029), .C(n3030) );
  CKBD0 U2912 ( .CLK(n3030), .C(n3031) );
  CKBD0 U2913 ( .CLK(n3031), .C(n3032) );
  CKBD0 U2914 ( .CLK(n3032), .C(n3033) );
  BUFFD0 U2915 ( .I(n3033), .Z(n3034) );
  CKBD0 U2916 ( .CLK(n3034), .C(n3035) );
  CKBD0 U2917 ( .CLK(n3035), .C(n3036) );
  CKBD0 U2918 ( .CLK(n3036), .C(n3037) );
  CKBD0 U2919 ( .CLK(n3037), .C(n3038) );
  CKBD0 U2920 ( .CLK(n3038), .C(n3039) );
  CKBD0 U2921 ( .CLK(n3039), .C(n3040) );
  CKBD0 U2922 ( .CLK(n3040), .C(n3041) );
  CKBD0 U2923 ( .CLK(n3041), .C(n3042) );
  CKBD0 U2924 ( .CLK(n3042), .C(n3043) );
  CKBD0 U2925 ( .CLK(n3043), .C(n3044) );
  BUFFD0 U2926 ( .I(n3044), .Z(n3045) );
  CKBD0 U2927 ( .CLK(n3045), .C(n3046) );
  CKBD0 U2928 ( .CLK(n3046), .C(n3047) );
  CKBD0 U2929 ( .CLK(n3047), .C(n3048) );
  CKBD0 U2930 ( .CLK(n3048), .C(n3049) );
  CKBD0 U2931 ( .CLK(n3049), .C(n3050) );
  CKBD0 U2932 ( .CLK(n3050), .C(n3051) );
  CKBD0 U2933 ( .CLK(n3051), .C(n3052) );
  CKBD0 U2934 ( .CLK(n3052), .C(n3053) );
  CKBD0 U2935 ( .CLK(n3053), .C(n3054) );
  CKBD0 U2936 ( .CLK(n3054), .C(n3055) );
  BUFFD0 U2937 ( .I(n3055), .Z(n3056) );
  CKBD0 U2938 ( .CLK(n3056), .C(n3057) );
  CKBD0 U2939 ( .CLK(n3057), .C(n3058) );
  CKBD0 U2940 ( .CLK(n3058), .C(n3059) );
  CKBD0 U2941 ( .CLK(n3059), .C(n3060) );
  CKBD0 U2942 ( .CLK(n3060), .C(n3061) );
  CKBD0 U2943 ( .CLK(n3061), .C(n3062) );
  CKBD0 U2944 ( .CLK(n3062), .C(n3063) );
  CKBD0 U2945 ( .CLK(n3063), .C(n3064) );
  CKBD0 U2946 ( .CLK(n3064), .C(n3065) );
  BUFFD0 U2947 ( .I(n3065), .Z(n3066) );
  CKBD0 U2948 ( .CLK(n3066), .C(n3067) );
  CKBD0 U2949 ( .CLK(n3067), .C(n3068) );
  CKBD0 U2950 ( .CLK(n3068), .C(n3069) );
  CKBD0 U2951 ( .CLK(n3069), .C(n3070) );
  CKBD0 U2952 ( .CLK(n3070), .C(n3071) );
  CKBD0 U2953 ( .CLK(n3071), .C(n3072) );
  CKBD0 U2954 ( .CLK(n3072), .C(n3073) );
  CKBD0 U2955 ( .CLK(n3073), .C(n3074) );
  CKBD0 U2956 ( .CLK(n3074), .C(n3075) );
  CKBD0 U2957 ( .CLK(n3075), .C(n3076) );
  BUFFD0 U2958 ( .I(n3076), .Z(n3077) );
  CKBD0 U2959 ( .CLK(n3077), .C(n3078) );
  CKBD0 U2960 ( .CLK(n3078), .C(n3079) );
  CKBD0 U2961 ( .CLK(n3079), .C(n3080) );
  CKBD0 U2962 ( .CLK(n3080), .C(n3081) );
  CKBD0 U2963 ( .CLK(n3081), .C(n3082) );
  CKBD0 U2964 ( .CLK(n3082), .C(n3083) );
  BUFFD0 U2965 ( .I(n3083), .Z(n3084) );
  CKBD0 U2966 ( .CLK(n3084), .C(n3085) );
  BUFFD0 U2967 ( .I(n3085), .Z(n3086) );
  CKBD0 U2968 ( .CLK(n3086), .C(n3087) );
  BUFFD0 U2969 ( .I(n3087), .Z(n3088) );
  CKBD0 U2970 ( .CLK(n3088), .C(n3089) );
  BUFFD0 U2971 ( .I(n3089), .Z(n3090) );
  CKBD0 U2972 ( .CLK(n3090), .C(n3091) );
  BUFFD0 U2973 ( .I(n3091), .Z(n3092) );
  CKBD0 U2974 ( .CLK(n3092), .C(n3093) );
  BUFFD0 U2975 ( .I(n3093), .Z(n3094) );
  CKBD0 U2976 ( .CLK(n3094), .C(n3095) );
  BUFFD0 U2977 ( .I(n3095), .Z(n3096) );
  CKBD0 U2978 ( .CLK(n3096), .C(n3097) );
  BUFFD0 U2979 ( .I(n3097), .Z(n3098) );
  BUFFD0 U2980 ( .I(n3100), .Z(n3099) );
  BUFFD0 U2981 ( .I(n3101), .Z(n3100) );
  BUFFD0 U2982 ( .I(n9162), .Z(n3101) );
  CKBD0 U2983 ( .CLK(n1360), .C(n3102) );
  CKBD0 U2984 ( .CLK(n3102), .C(n3103) );
  CKBD0 U2985 ( .CLK(n3103), .C(n3104) );
  BUFFD0 U2986 ( .I(n3104), .Z(n3105) );
  CKBD0 U2987 ( .CLK(n3105), .C(n3106) );
  CKBD0 U2988 ( .CLK(n3106), .C(n3107) );
  CKBD0 U2989 ( .CLK(n3107), .C(n3108) );
  CKBD0 U2990 ( .CLK(n3108), .C(n3109) );
  CKBD0 U2991 ( .CLK(n3109), .C(n3110) );
  CKBD0 U2992 ( .CLK(n3110), .C(n3111) );
  CKBD0 U2993 ( .CLK(n3111), .C(n3112) );
  CKBD0 U2994 ( .CLK(n3112), .C(n3113) );
  CKBD0 U2995 ( .CLK(n3113), .C(n3114) );
  CKBD0 U2996 ( .CLK(n3114), .C(n3115) );
  BUFFD0 U2997 ( .I(n3115), .Z(n3116) );
  CKBD0 U2998 ( .CLK(n3116), .C(n3117) );
  CKBD0 U2999 ( .CLK(n3117), .C(n3118) );
  CKBD0 U3000 ( .CLK(n3118), .C(n3119) );
  CKBD0 U3001 ( .CLK(n3119), .C(n3120) );
  CKBD0 U3002 ( .CLK(n3120), .C(n3121) );
  CKBD0 U3003 ( .CLK(n3121), .C(n3122) );
  CKBD0 U3004 ( .CLK(n3122), .C(n3123) );
  CKBD0 U3005 ( .CLK(n3123), .C(n3124) );
  CKBD0 U3006 ( .CLK(n3124), .C(n3125) );
  BUFFD0 U3007 ( .I(n3125), .Z(n3126) );
  CKBD0 U3008 ( .CLK(n3126), .C(n3127) );
  CKBD0 U3009 ( .CLK(n3127), .C(n3128) );
  CKBD0 U3010 ( .CLK(n3128), .C(n3129) );
  CKBD0 U3011 ( .CLK(n3129), .C(n3130) );
  CKBD0 U3012 ( .CLK(n3130), .C(n3131) );
  CKBD0 U3013 ( .CLK(n3131), .C(n3132) );
  CKBD0 U3014 ( .CLK(n3132), .C(n3133) );
  CKBD0 U3015 ( .CLK(n3133), .C(n3134) );
  CKBD0 U3016 ( .CLK(n3134), .C(n3135) );
  CKBD0 U3017 ( .CLK(n3135), .C(n3136) );
  BUFFD0 U3018 ( .I(n3136), .Z(n3137) );
  CKBD0 U3019 ( .CLK(n3137), .C(n3138) );
  CKBD0 U3020 ( .CLK(n3138), .C(n3139) );
  CKBD0 U3021 ( .CLK(n3139), .C(n3140) );
  CKBD0 U3022 ( .CLK(n3140), .C(n3141) );
  CKBD0 U3023 ( .CLK(n3141), .C(n3142) );
  CKBD0 U3024 ( .CLK(n3142), .C(n3143) );
  CKBD0 U3025 ( .CLK(n3143), .C(n3144) );
  CKBD0 U3026 ( .CLK(n3144), .C(n3145) );
  CKBD0 U3027 ( .CLK(n3145), .C(n3146) );
  CKBD0 U3028 ( .CLK(n3146), .C(n3147) );
  BUFFD0 U3029 ( .I(n3147), .Z(n3148) );
  CKBD0 U3030 ( .CLK(n3148), .C(n3149) );
  CKBD0 U3031 ( .CLK(n3149), .C(n3150) );
  CKBD0 U3032 ( .CLK(n3150), .C(n3151) );
  CKBD0 U3033 ( .CLK(n3151), .C(n3152) );
  CKBD0 U3034 ( .CLK(n3152), .C(n3153) );
  CKBD0 U3035 ( .CLK(n3153), .C(n3154) );
  CKBD0 U3036 ( .CLK(n3154), .C(n3155) );
  CKBD0 U3037 ( .CLK(n3155), .C(n3156) );
  CKBD0 U3038 ( .CLK(n3156), .C(n3157) );
  CKBD0 U3039 ( .CLK(n3157), .C(n3158) );
  BUFFD0 U3040 ( .I(n3158), .Z(n3159) );
  CKBD0 U3041 ( .CLK(n3159), .C(n3160) );
  CKBD0 U3042 ( .CLK(n3160), .C(n3161) );
  CKBD0 U3043 ( .CLK(n3161), .C(n3162) );
  CKBD0 U3044 ( .CLK(n3162), .C(n3163) );
  CKBD0 U3045 ( .CLK(n3163), .C(n3164) );
  CKBD0 U3046 ( .CLK(n3164), .C(n3165) );
  CKBD0 U3047 ( .CLK(n3165), .C(n3166) );
  CKBD0 U3048 ( .CLK(n3166), .C(n3167) );
  CKBD0 U3049 ( .CLK(n3167), .C(n3168) );
  CKBD0 U3050 ( .CLK(n3168), .C(n3169) );
  BUFFD0 U3051 ( .I(n3169), .Z(n3170) );
  CKBD0 U3052 ( .CLK(n3170), .C(n3171) );
  CKBD0 U3053 ( .CLK(n3171), .C(n3172) );
  CKBD0 U3054 ( .CLK(n3172), .C(n3173) );
  CKBD0 U3055 ( .CLK(n3173), .C(n3174) );
  CKBD0 U3056 ( .CLK(n3174), .C(n3175) );
  CKBD0 U3057 ( .CLK(n3175), .C(n3176) );
  CKBD0 U3058 ( .CLK(n3176), .C(n3177) );
  CKBD0 U3059 ( .CLK(n3177), .C(n3178) );
  CKBD0 U3060 ( .CLK(n3178), .C(n3179) );
  CKBD0 U3061 ( .CLK(n3179), .C(n3180) );
  BUFFD0 U3062 ( .I(n3180), .Z(n3181) );
  CKBD0 U3063 ( .CLK(n3181), .C(n3182) );
  CKBD0 U3064 ( .CLK(n3182), .C(n3183) );
  CKBD0 U3065 ( .CLK(n3183), .C(n3184) );
  CKBD0 U3066 ( .CLK(n3184), .C(n3185) );
  CKBD0 U3067 ( .CLK(n3185), .C(n3186) );
  CKBD0 U3068 ( .CLK(n3186), .C(n3187) );
  CKBD0 U3069 ( .CLK(n3187), .C(n3188) );
  CKBD0 U3070 ( .CLK(n3188), .C(n3189) );
  CKBD0 U3071 ( .CLK(n3189), .C(n3190) );
  BUFFD0 U3072 ( .I(n3190), .Z(n3191) );
  CKBD0 U3073 ( .CLK(n3191), .C(n3192) );
  CKBD0 U3074 ( .CLK(n3192), .C(n3193) );
  CKBD0 U3075 ( .CLK(n3193), .C(n3194) );
  CKBD0 U3076 ( .CLK(n3194), .C(n3195) );
  CKBD0 U3077 ( .CLK(n3195), .C(n3196) );
  CKBD0 U3078 ( .CLK(n3196), .C(n3197) );
  CKBD0 U3079 ( .CLK(n3197), .C(n3198) );
  CKBD0 U3080 ( .CLK(n3198), .C(n3199) );
  CKBD0 U3081 ( .CLK(n3199), .C(n3200) );
  CKBD0 U3082 ( .CLK(n3200), .C(n3201) );
  BUFFD0 U3083 ( .I(n3201), .Z(n3202) );
  CKBD0 U3084 ( .CLK(n3202), .C(n3203) );
  CKBD0 U3085 ( .CLK(n3203), .C(n3204) );
  CKBD0 U3086 ( .CLK(n3204), .C(n3205) );
  CKBD0 U3087 ( .CLK(n3205), .C(n3206) );
  CKBD0 U3088 ( .CLK(n3206), .C(n3207) );
  CKBD0 U3089 ( .CLK(n3207), .C(n3208) );
  CKBD0 U3090 ( .CLK(n3208), .C(n3209) );
  CKBD0 U3091 ( .CLK(n3209), .C(n3210) );
  CKBD0 U3092 ( .CLK(n3210), .C(n3211) );
  CKBD0 U3093 ( .CLK(n3211), .C(n3212) );
  BUFFD0 U3094 ( .I(n3212), .Z(n3213) );
  CKBD0 U3095 ( .CLK(n3213), .C(n3214) );
  CKBD0 U3096 ( .CLK(n3214), .C(n3215) );
  CKBD0 U3097 ( .CLK(n3215), .C(n3216) );
  CKBD0 U3098 ( .CLK(n3216), .C(n3217) );
  CKBD0 U3099 ( .CLK(n3217), .C(n3218) );
  CKBD0 U3100 ( .CLK(n3218), .C(n3219) );
  BUFFD0 U3101 ( .I(n3219), .Z(n3220) );
  CKBD0 U3102 ( .CLK(n3220), .C(n3221) );
  BUFFD0 U3103 ( .I(n3221), .Z(n3222) );
  CKBD0 U3104 ( .CLK(n3222), .C(n3223) );
  BUFFD0 U3105 ( .I(n3223), .Z(n3224) );
  CKBD0 U3106 ( .CLK(n3224), .C(n3225) );
  BUFFD0 U3107 ( .I(n3225), .Z(n3226) );
  CKBD0 U3108 ( .CLK(n3226), .C(n3227) );
  BUFFD0 U3109 ( .I(n3227), .Z(n3228) );
  CKBD0 U3110 ( .CLK(n3228), .C(n3229) );
  BUFFD0 U3111 ( .I(n3229), .Z(n3230) );
  CKBD0 U3112 ( .CLK(n3230), .C(n3231) );
  BUFFD0 U3113 ( .I(n3231), .Z(n3232) );
  CKBD0 U3114 ( .CLK(n3232), .C(n3233) );
  BUFFD0 U3115 ( .I(n3233), .Z(n3234) );
  BUFFD0 U3116 ( .I(n3236), .Z(n3235) );
  BUFFD0 U3117 ( .I(n3237), .Z(n3236) );
  BUFFD0 U3118 ( .I(n9163), .Z(n3237) );
  CKBD0 U3119 ( .CLK(n1358), .C(n3238) );
  CKBD0 U3120 ( .CLK(n3238), .C(n3239) );
  CKBD0 U3121 ( .CLK(n3239), .C(n3240) );
  BUFFD0 U3122 ( .I(n3240), .Z(n3241) );
  CKBD0 U3123 ( .CLK(n3241), .C(n3242) );
  CKBD0 U3124 ( .CLK(n3242), .C(n3243) );
  CKBD0 U3125 ( .CLK(n3243), .C(n3244) );
  CKBD0 U3126 ( .CLK(n3244), .C(n3245) );
  CKBD0 U3127 ( .CLK(n3245), .C(n3246) );
  CKBD0 U3128 ( .CLK(n3246), .C(n3247) );
  CKBD0 U3129 ( .CLK(n3247), .C(n3248) );
  CKBD0 U3130 ( .CLK(n3248), .C(n3249) );
  CKBD0 U3131 ( .CLK(n3249), .C(n3250) );
  CKBD0 U3132 ( .CLK(n3250), .C(n3251) );
  BUFFD0 U3133 ( .I(n3251), .Z(n3252) );
  CKBD0 U3134 ( .CLK(n3252), .C(n3253) );
  CKBD0 U3135 ( .CLK(n3253), .C(n3254) );
  CKBD0 U3136 ( .CLK(n3254), .C(n3255) );
  CKBD0 U3137 ( .CLK(n3255), .C(n3256) );
  CKBD0 U3138 ( .CLK(n3256), .C(n3257) );
  CKBD0 U3139 ( .CLK(n3257), .C(n3258) );
  CKBD0 U3140 ( .CLK(n3258), .C(n3259) );
  CKBD0 U3141 ( .CLK(n3259), .C(n3260) );
  CKBD0 U3142 ( .CLK(n3260), .C(n3261) );
  BUFFD0 U3143 ( .I(n3261), .Z(n3262) );
  CKBD0 U3144 ( .CLK(n3262), .C(n3263) );
  CKBD0 U3145 ( .CLK(n3263), .C(n3264) );
  CKBD0 U3146 ( .CLK(n3264), .C(n3265) );
  CKBD0 U3147 ( .CLK(n3265), .C(n3266) );
  CKBD0 U3148 ( .CLK(n3266), .C(n3267) );
  CKBD0 U3149 ( .CLK(n3267), .C(n3268) );
  CKBD0 U3150 ( .CLK(n3268), .C(n3269) );
  CKBD0 U3151 ( .CLK(n3269), .C(n3270) );
  CKBD0 U3152 ( .CLK(n3270), .C(n3271) );
  CKBD0 U3153 ( .CLK(n3271), .C(n3272) );
  BUFFD0 U3154 ( .I(n3272), .Z(n3273) );
  CKBD0 U3155 ( .CLK(n3273), .C(n3274) );
  CKBD0 U3156 ( .CLK(n3274), .C(n3275) );
  CKBD0 U3157 ( .CLK(n3275), .C(n3276) );
  CKBD0 U3158 ( .CLK(n3276), .C(n3277) );
  CKBD0 U3159 ( .CLK(n3277), .C(n3278) );
  CKBD0 U3160 ( .CLK(n3278), .C(n3279) );
  CKBD0 U3161 ( .CLK(n3279), .C(n3280) );
  CKBD0 U3162 ( .CLK(n3280), .C(n3281) );
  CKBD0 U3163 ( .CLK(n3281), .C(n3282) );
  CKBD0 U3164 ( .CLK(n3282), .C(n3283) );
  BUFFD0 U3165 ( .I(n3283), .Z(n3284) );
  CKBD0 U3166 ( .CLK(n3284), .C(n3285) );
  CKBD0 U3167 ( .CLK(n3285), .C(n3286) );
  CKBD0 U3168 ( .CLK(n3286), .C(n3287) );
  CKBD0 U3169 ( .CLK(n3287), .C(n3288) );
  CKBD0 U3170 ( .CLK(n3288), .C(n3289) );
  CKBD0 U3171 ( .CLK(n3289), .C(n3290) );
  CKBD0 U3172 ( .CLK(n3290), .C(n3291) );
  CKBD0 U3173 ( .CLK(n3291), .C(n3292) );
  CKBD0 U3174 ( .CLK(n3292), .C(n3293) );
  CKBD0 U3175 ( .CLK(n3293), .C(n3294) );
  BUFFD0 U3176 ( .I(n3294), .Z(n3295) );
  CKBD0 U3177 ( .CLK(n3295), .C(n3296) );
  CKBD0 U3178 ( .CLK(n3296), .C(n3297) );
  CKBD0 U3179 ( .CLK(n3297), .C(n3298) );
  CKBD0 U3180 ( .CLK(n3298), .C(n3299) );
  CKBD0 U3181 ( .CLK(n3299), .C(n3300) );
  CKBD0 U3182 ( .CLK(n3300), .C(n3301) );
  CKBD0 U3183 ( .CLK(n3301), .C(n3302) );
  CKBD0 U3184 ( .CLK(n3302), .C(n3303) );
  CKBD0 U3185 ( .CLK(n3303), .C(n3304) );
  CKBD0 U3186 ( .CLK(n3304), .C(n3305) );
  BUFFD0 U3187 ( .I(n3305), .Z(n3306) );
  CKBD0 U3188 ( .CLK(n3306), .C(n3307) );
  CKBD0 U3189 ( .CLK(n3307), .C(n3308) );
  CKBD0 U3190 ( .CLK(n3308), .C(n3309) );
  CKBD0 U3191 ( .CLK(n3309), .C(n3310) );
  CKBD0 U3192 ( .CLK(n3310), .C(n3311) );
  CKBD0 U3193 ( .CLK(n3311), .C(n3312) );
  CKBD0 U3194 ( .CLK(n3312), .C(n3313) );
  CKBD0 U3195 ( .CLK(n3313), .C(n3314) );
  CKBD0 U3196 ( .CLK(n3314), .C(n3315) );
  CKBD0 U3197 ( .CLK(n3315), .C(n3316) );
  BUFFD0 U3198 ( .I(n3316), .Z(n3317) );
  CKBD0 U3199 ( .CLK(n3317), .C(n3318) );
  CKBD0 U3200 ( .CLK(n3318), .C(n3319) );
  CKBD0 U3201 ( .CLK(n3319), .C(n3320) );
  CKBD0 U3202 ( .CLK(n3320), .C(n3321) );
  CKBD0 U3203 ( .CLK(n3321), .C(n3322) );
  CKBD0 U3204 ( .CLK(n3322), .C(n3323) );
  CKBD0 U3205 ( .CLK(n3323), .C(n3324) );
  CKBD0 U3206 ( .CLK(n3324), .C(n3325) );
  CKBD0 U3207 ( .CLK(n3325), .C(n3326) );
  BUFFD0 U3208 ( .I(n3326), .Z(n3327) );
  CKBD0 U3209 ( .CLK(n3327), .C(n3328) );
  CKBD0 U3210 ( .CLK(n3328), .C(n3329) );
  CKBD0 U3211 ( .CLK(n3329), .C(n3330) );
  CKBD0 U3212 ( .CLK(n3330), .C(n3331) );
  CKBD0 U3213 ( .CLK(n3331), .C(n3332) );
  CKBD0 U3214 ( .CLK(n3332), .C(n3333) );
  CKBD0 U3215 ( .CLK(n3333), .C(n3334) );
  CKBD0 U3216 ( .CLK(n3334), .C(n3335) );
  CKBD0 U3217 ( .CLK(n3335), .C(n3336) );
  CKBD0 U3218 ( .CLK(n3336), .C(n3337) );
  BUFFD0 U3219 ( .I(n3337), .Z(n3338) );
  CKBD0 U3220 ( .CLK(n3338), .C(n3339) );
  CKBD0 U3221 ( .CLK(n3339), .C(n3340) );
  CKBD0 U3222 ( .CLK(n3340), .C(n3341) );
  CKBD0 U3223 ( .CLK(n3341), .C(n3342) );
  CKBD0 U3224 ( .CLK(n3342), .C(n3343) );
  CKBD0 U3225 ( .CLK(n3343), .C(n3344) );
  CKBD0 U3226 ( .CLK(n3344), .C(n3345) );
  CKBD0 U3227 ( .CLK(n3345), .C(n3346) );
  CKBD0 U3228 ( .CLK(n3346), .C(n3347) );
  CKBD0 U3229 ( .CLK(n3347), .C(n3348) );
  BUFFD0 U3230 ( .I(n3348), .Z(n3349) );
  CKBD0 U3231 ( .CLK(n3349), .C(n3350) );
  CKBD0 U3232 ( .CLK(n3350), .C(n3351) );
  CKBD0 U3233 ( .CLK(n3351), .C(n3352) );
  CKBD0 U3234 ( .CLK(n3352), .C(n3353) );
  CKBD0 U3235 ( .CLK(n3353), .C(n3354) );
  CKBD0 U3236 ( .CLK(n3354), .C(n3355) );
  BUFFD0 U3237 ( .I(n3355), .Z(n3356) );
  CKBD0 U3238 ( .CLK(n3356), .C(n3357) );
  BUFFD0 U3239 ( .I(n3357), .Z(n3358) );
  CKBD0 U3240 ( .CLK(n3358), .C(n3359) );
  BUFFD0 U3241 ( .I(n3359), .Z(n3360) );
  CKBD0 U3242 ( .CLK(n3360), .C(n3361) );
  BUFFD0 U3243 ( .I(n3361), .Z(n3362) );
  CKBD0 U3244 ( .CLK(n3362), .C(n3363) );
  BUFFD0 U3245 ( .I(n3363), .Z(n3364) );
  CKBD0 U3246 ( .CLK(n3364), .C(n3365) );
  BUFFD0 U3247 ( .I(n3365), .Z(n3366) );
  CKBD0 U3248 ( .CLK(n3366), .C(n3367) );
  BUFFD0 U3249 ( .I(n3367), .Z(n3368) );
  CKBD0 U3250 ( .CLK(n3368), .C(n3369) );
  BUFFD0 U3251 ( .I(n3369), .Z(n3370) );
  BUFFD0 U3252 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3253 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3254 ( .I(n9164), .Z(n3373) );
  CKBD0 U3255 ( .CLK(n1356), .C(n3374) );
  CKBD0 U3256 ( .CLK(n3374), .C(n3375) );
  CKBD0 U3257 ( .CLK(n3375), .C(n3376) );
  BUFFD0 U3258 ( .I(n3376), .Z(n3377) );
  CKBD0 U3259 ( .CLK(n3377), .C(n3378) );
  CKBD0 U3260 ( .CLK(n3378), .C(n3379) );
  CKBD0 U3261 ( .CLK(n3379), .C(n3380) );
  CKBD0 U3262 ( .CLK(n3380), .C(n3381) );
  CKBD0 U3263 ( .CLK(n3381), .C(n3382) );
  CKBD0 U3264 ( .CLK(n3382), .C(n3383) );
  CKBD0 U3265 ( .CLK(n3383), .C(n3384) );
  CKBD0 U3266 ( .CLK(n3384), .C(n3385) );
  CKBD0 U3267 ( .CLK(n3385), .C(n3386) );
  CKBD0 U3268 ( .CLK(n3386), .C(n3387) );
  BUFFD0 U3269 ( .I(n3387), .Z(n3388) );
  CKBD0 U3270 ( .CLK(n3388), .C(n3389) );
  CKBD0 U3271 ( .CLK(n3389), .C(n3390) );
  CKBD0 U3272 ( .CLK(n3390), .C(n3391) );
  CKBD0 U3273 ( .CLK(n3391), .C(n3392) );
  CKBD0 U3274 ( .CLK(n3392), .C(n3393) );
  CKBD0 U3275 ( .CLK(n3393), .C(n3394) );
  CKBD0 U3276 ( .CLK(n3394), .C(n3395) );
  CKBD0 U3277 ( .CLK(n3395), .C(n3396) );
  CKBD0 U3278 ( .CLK(n3396), .C(n3397) );
  BUFFD0 U3279 ( .I(n3397), .Z(n3398) );
  CKBD0 U3280 ( .CLK(n3398), .C(n3399) );
  CKBD0 U3281 ( .CLK(n3399), .C(n3400) );
  CKBD0 U3282 ( .CLK(n3400), .C(n3401) );
  CKBD0 U3283 ( .CLK(n3401), .C(n3402) );
  CKBD0 U3284 ( .CLK(n3402), .C(n3403) );
  CKBD0 U3285 ( .CLK(n3403), .C(n3404) );
  CKBD0 U3286 ( .CLK(n3404), .C(n3405) );
  CKBD0 U3287 ( .CLK(n3405), .C(n3406) );
  CKBD0 U3288 ( .CLK(n3406), .C(n3407) );
  CKBD0 U3289 ( .CLK(n3407), .C(n3408) );
  BUFFD0 U3290 ( .I(n3408), .Z(n3409) );
  CKBD0 U3291 ( .CLK(n3409), .C(n3410) );
  CKBD0 U3292 ( .CLK(n3410), .C(n3411) );
  CKBD0 U3293 ( .CLK(n3411), .C(n3412) );
  CKBD0 U3294 ( .CLK(n3412), .C(n3413) );
  CKBD0 U3295 ( .CLK(n3413), .C(n3414) );
  CKBD0 U3296 ( .CLK(n3414), .C(n3415) );
  CKBD0 U3297 ( .CLK(n3415), .C(n3416) );
  CKBD0 U3298 ( .CLK(n3416), .C(n3417) );
  CKBD0 U3299 ( .CLK(n3417), .C(n3418) );
  CKBD0 U3300 ( .CLK(n3418), .C(n3419) );
  BUFFD0 U3301 ( .I(n3419), .Z(n3420) );
  CKBD0 U3302 ( .CLK(n3420), .C(n3421) );
  CKBD0 U3303 ( .CLK(n3421), .C(n3422) );
  CKBD0 U3304 ( .CLK(n3422), .C(n3423) );
  CKBD0 U3305 ( .CLK(n3423), .C(n3424) );
  CKBD0 U3306 ( .CLK(n3424), .C(n3425) );
  CKBD0 U3307 ( .CLK(n3425), .C(n3426) );
  CKBD0 U3308 ( .CLK(n3426), .C(n3427) );
  CKBD0 U3309 ( .CLK(n3427), .C(n3428) );
  CKBD0 U3310 ( .CLK(n3428), .C(n3429) );
  CKBD0 U3311 ( .CLK(n3429), .C(n3430) );
  BUFFD0 U3312 ( .I(n3430), .Z(n3431) );
  CKBD0 U3313 ( .CLK(n3431), .C(n3432) );
  CKBD0 U3314 ( .CLK(n3432), .C(n3433) );
  CKBD0 U3315 ( .CLK(n3433), .C(n3434) );
  CKBD0 U3316 ( .CLK(n3434), .C(n3435) );
  CKBD0 U3317 ( .CLK(n3435), .C(n3436) );
  CKBD0 U3318 ( .CLK(n3436), .C(n3437) );
  CKBD0 U3319 ( .CLK(n3437), .C(n3438) );
  CKBD0 U3320 ( .CLK(n3438), .C(n3439) );
  CKBD0 U3321 ( .CLK(n3439), .C(n3440) );
  CKBD0 U3322 ( .CLK(n3440), .C(n3441) );
  BUFFD0 U3323 ( .I(n3441), .Z(n3442) );
  CKBD0 U3324 ( .CLK(n3442), .C(n3443) );
  CKBD0 U3325 ( .CLK(n3443), .C(n3444) );
  CKBD0 U3326 ( .CLK(n3444), .C(n3445) );
  CKBD0 U3327 ( .CLK(n3445), .C(n3446) );
  CKBD0 U3328 ( .CLK(n3446), .C(n3447) );
  CKBD0 U3329 ( .CLK(n3447), .C(n3448) );
  CKBD0 U3330 ( .CLK(n3448), .C(n3449) );
  CKBD0 U3331 ( .CLK(n3449), .C(n3450) );
  CKBD0 U3332 ( .CLK(n3450), .C(n3451) );
  CKBD0 U3333 ( .CLK(n3451), .C(n3452) );
  BUFFD0 U3334 ( .I(n3452), .Z(n3453) );
  CKBD0 U3335 ( .CLK(n3453), .C(n3454) );
  CKBD0 U3336 ( .CLK(n3454), .C(n3455) );
  CKBD0 U3337 ( .CLK(n3455), .C(n3456) );
  CKBD0 U3338 ( .CLK(n3456), .C(n3457) );
  CKBD0 U3339 ( .CLK(n3457), .C(n3458) );
  CKBD0 U3340 ( .CLK(n3458), .C(n3459) );
  CKBD0 U3341 ( .CLK(n3459), .C(n3460) );
  CKBD0 U3342 ( .CLK(n3460), .C(n3461) );
  CKBD0 U3343 ( .CLK(n3461), .C(n3462) );
  CKBD0 U3344 ( .CLK(n3462), .C(n3463) );
  BUFFD0 U3345 ( .I(n3463), .Z(n3464) );
  CKBD0 U3346 ( .CLK(n3464), .C(n3465) );
  CKBD0 U3347 ( .CLK(n3465), .C(n3466) );
  CKBD0 U3348 ( .CLK(n3466), .C(n3467) );
  CKBD0 U3349 ( .CLK(n3467), .C(n3468) );
  CKBD0 U3350 ( .CLK(n3468), .C(n3469) );
  CKBD0 U3351 ( .CLK(n3469), .C(n3470) );
  CKBD0 U3352 ( .CLK(n3470), .C(n3471) );
  CKBD0 U3353 ( .CLK(n3471), .C(n3472) );
  CKBD0 U3354 ( .CLK(n3472), .C(n3473) );
  BUFFD0 U3355 ( .I(n3473), .Z(n3474) );
  CKBD0 U3356 ( .CLK(n3474), .C(n3475) );
  CKBD0 U3357 ( .CLK(n3475), .C(n3476) );
  CKBD0 U3358 ( .CLK(n3476), .C(n3477) );
  CKBD0 U3359 ( .CLK(n3477), .C(n3478) );
  CKBD0 U3360 ( .CLK(n3478), .C(n3479) );
  CKBD0 U3361 ( .CLK(n3479), .C(n3480) );
  CKBD0 U3362 ( .CLK(n3480), .C(n3481) );
  CKBD0 U3363 ( .CLK(n3481), .C(n3482) );
  CKBD0 U3364 ( .CLK(n3482), .C(n3483) );
  CKBD0 U3365 ( .CLK(n3483), .C(n3484) );
  BUFFD0 U3366 ( .I(n3484), .Z(n3485) );
  CKBD0 U3367 ( .CLK(n3485), .C(n3486) );
  CKBD0 U3368 ( .CLK(n3486), .C(n3487) );
  CKBD0 U3369 ( .CLK(n3487), .C(n3488) );
  CKBD0 U3370 ( .CLK(n3488), .C(n3489) );
  CKBD0 U3371 ( .CLK(n3489), .C(n3490) );
  CKBD0 U3372 ( .CLK(n3490), .C(n3491) );
  BUFFD0 U3373 ( .I(n3491), .Z(n3492) );
  CKBD0 U3374 ( .CLK(n3492), .C(n3493) );
  BUFFD0 U3375 ( .I(n3493), .Z(n3494) );
  CKBD0 U3376 ( .CLK(n3494), .C(n3495) );
  BUFFD0 U3377 ( .I(n3495), .Z(n3496) );
  CKBD0 U3378 ( .CLK(n3496), .C(n3497) );
  BUFFD0 U3379 ( .I(n3497), .Z(n3498) );
  CKBD0 U3380 ( .CLK(n3498), .C(n3499) );
  BUFFD0 U3381 ( .I(n3499), .Z(n3500) );
  CKBD0 U3382 ( .CLK(n3500), .C(n3501) );
  BUFFD0 U3383 ( .I(n3501), .Z(n3502) );
  CKBD0 U3384 ( .CLK(n3502), .C(n3503) );
  BUFFD0 U3385 ( .I(n3503), .Z(n3504) );
  CKBD0 U3386 ( .CLK(n3504), .C(n3505) );
  BUFFD0 U3387 ( .I(n3505), .Z(n3506) );
  BUFFD0 U3388 ( .I(n3508), .Z(n3507) );
  BUFFD0 U3389 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3390 ( .I(n9165), .Z(n3509) );
  CKBD0 U3391 ( .CLK(n1354), .C(n3510) );
  CKBD0 U3392 ( .CLK(n3510), .C(n3511) );
  CKBD0 U3393 ( .CLK(n3511), .C(n3512) );
  BUFFD0 U3394 ( .I(n3512), .Z(n3513) );
  CKBD0 U3395 ( .CLK(n3513), .C(n3514) );
  CKBD0 U3396 ( .CLK(n3514), .C(n3515) );
  CKBD0 U3397 ( .CLK(n3515), .C(n3516) );
  CKBD0 U3398 ( .CLK(n3516), .C(n3517) );
  CKBD0 U3399 ( .CLK(n3517), .C(n3518) );
  CKBD0 U3400 ( .CLK(n3518), .C(n3519) );
  CKBD0 U3401 ( .CLK(n3519), .C(n3520) );
  CKBD0 U3402 ( .CLK(n3520), .C(n3521) );
  CKBD0 U3403 ( .CLK(n3521), .C(n3522) );
  CKBD0 U3404 ( .CLK(n3522), .C(n3523) );
  BUFFD0 U3405 ( .I(n3523), .Z(n3524) );
  CKBD0 U3406 ( .CLK(n3524), .C(n3525) );
  CKBD0 U3407 ( .CLK(n3525), .C(n3526) );
  CKBD0 U3408 ( .CLK(n3526), .C(n3527) );
  CKBD0 U3409 ( .CLK(n3527), .C(n3528) );
  CKBD0 U3410 ( .CLK(n3528), .C(n3529) );
  CKBD0 U3411 ( .CLK(n3529), .C(n3530) );
  CKBD0 U3412 ( .CLK(n3530), .C(n3531) );
  CKBD0 U3413 ( .CLK(n3531), .C(n3532) );
  CKBD0 U3414 ( .CLK(n3532), .C(n3533) );
  BUFFD0 U3415 ( .I(n3533), .Z(n3534) );
  CKBD0 U3416 ( .CLK(n3534), .C(n3535) );
  CKBD0 U3417 ( .CLK(n3535), .C(n3536) );
  CKBD0 U3418 ( .CLK(n3536), .C(n3537) );
  CKBD0 U3419 ( .CLK(n3537), .C(n3538) );
  CKBD0 U3420 ( .CLK(n3538), .C(n3539) );
  CKBD0 U3421 ( .CLK(n3539), .C(n3540) );
  CKBD0 U3422 ( .CLK(n3540), .C(n3541) );
  CKBD0 U3423 ( .CLK(n3541), .C(n3542) );
  CKBD0 U3424 ( .CLK(n3542), .C(n3543) );
  CKBD0 U3425 ( .CLK(n3543), .C(n3544) );
  BUFFD0 U3426 ( .I(n3544), .Z(n3545) );
  CKBD0 U3427 ( .CLK(n3545), .C(n3546) );
  CKBD0 U3428 ( .CLK(n3546), .C(n3547) );
  CKBD0 U3429 ( .CLK(n3547), .C(n3548) );
  CKBD0 U3430 ( .CLK(n3548), .C(n3549) );
  CKBD0 U3431 ( .CLK(n3549), .C(n3550) );
  CKBD0 U3432 ( .CLK(n3550), .C(n3551) );
  CKBD0 U3433 ( .CLK(n3551), .C(n3552) );
  CKBD0 U3434 ( .CLK(n3552), .C(n3553) );
  CKBD0 U3435 ( .CLK(n3553), .C(n3554) );
  CKBD0 U3436 ( .CLK(n3554), .C(n3555) );
  BUFFD0 U3437 ( .I(n3555), .Z(n3556) );
  CKBD0 U3438 ( .CLK(n3556), .C(n3557) );
  CKBD0 U3439 ( .CLK(n3557), .C(n3558) );
  CKBD0 U3440 ( .CLK(n3558), .C(n3559) );
  CKBD0 U3441 ( .CLK(n3559), .C(n3560) );
  CKBD0 U3442 ( .CLK(n3560), .C(n3561) );
  CKBD0 U3443 ( .CLK(n3561), .C(n3562) );
  CKBD0 U3444 ( .CLK(n3562), .C(n3563) );
  CKBD0 U3445 ( .CLK(n3563), .C(n3564) );
  CKBD0 U3446 ( .CLK(n3564), .C(n3565) );
  CKBD0 U3447 ( .CLK(n3565), .C(n3566) );
  BUFFD0 U3448 ( .I(n3566), .Z(n3567) );
  CKBD0 U3449 ( .CLK(n3567), .C(n3568) );
  CKBD0 U3450 ( .CLK(n3568), .C(n3569) );
  CKBD0 U3451 ( .CLK(n3569), .C(n3570) );
  CKBD0 U3452 ( .CLK(n3570), .C(n3571) );
  CKBD0 U3453 ( .CLK(n3571), .C(n3572) );
  CKBD0 U3454 ( .CLK(n3572), .C(n3573) );
  CKBD0 U3455 ( .CLK(n3573), .C(n3574) );
  CKBD0 U3456 ( .CLK(n3574), .C(n3575) );
  CKBD0 U3457 ( .CLK(n3575), .C(n3576) );
  CKBD0 U3458 ( .CLK(n3576), .C(n3577) );
  BUFFD0 U3459 ( .I(n3577), .Z(n3578) );
  CKBD0 U3460 ( .CLK(n3578), .C(n3579) );
  CKBD0 U3461 ( .CLK(n3579), .C(n3580) );
  CKBD0 U3462 ( .CLK(n3580), .C(n3581) );
  CKBD0 U3463 ( .CLK(n3581), .C(n3582) );
  CKBD0 U3464 ( .CLK(n3582), .C(n3583) );
  CKBD0 U3465 ( .CLK(n3583), .C(n3584) );
  CKBD0 U3466 ( .CLK(n3584), .C(n3585) );
  CKBD0 U3467 ( .CLK(n3585), .C(n3586) );
  CKBD0 U3468 ( .CLK(n3586), .C(n3587) );
  CKBD0 U3469 ( .CLK(n3587), .C(n3588) );
  BUFFD0 U3470 ( .I(n3588), .Z(n3589) );
  CKBD0 U3471 ( .CLK(n3589), .C(n3590) );
  CKBD0 U3472 ( .CLK(n3590), .C(n3591) );
  CKBD0 U3473 ( .CLK(n3591), .C(n3592) );
  CKBD0 U3474 ( .CLK(n3592), .C(n3593) );
  CKBD0 U3475 ( .CLK(n3593), .C(n3594) );
  CKBD0 U3476 ( .CLK(n3594), .C(n3595) );
  CKBD0 U3477 ( .CLK(n3595), .C(n3596) );
  CKBD0 U3478 ( .CLK(n3596), .C(n3597) );
  CKBD0 U3479 ( .CLK(n3597), .C(n3598) );
  CKBD0 U3480 ( .CLK(n3598), .C(n3599) );
  BUFFD0 U3481 ( .I(n3599), .Z(n3600) );
  CKBD0 U3482 ( .CLK(n3600), .C(n3601) );
  CKBD0 U3483 ( .CLK(n3601), .C(n3602) );
  CKBD0 U3484 ( .CLK(n3602), .C(n3603) );
  CKBD0 U3485 ( .CLK(n3603), .C(n3604) );
  CKBD0 U3486 ( .CLK(n3604), .C(n3605) );
  CKBD0 U3487 ( .CLK(n3605), .C(n3606) );
  CKBD0 U3488 ( .CLK(n3606), .C(n3607) );
  CKBD0 U3489 ( .CLK(n3607), .C(n3608) );
  CKBD0 U3490 ( .CLK(n3608), .C(n3609) );
  BUFFD0 U3491 ( .I(n3609), .Z(n3610) );
  CKBD0 U3492 ( .CLK(n3610), .C(n3611) );
  CKBD0 U3493 ( .CLK(n3611), .C(n3612) );
  CKBD0 U3494 ( .CLK(n3612), .C(n3613) );
  CKBD0 U3495 ( .CLK(n3613), .C(n3614) );
  CKBD0 U3496 ( .CLK(n3614), .C(n3615) );
  CKBD0 U3497 ( .CLK(n3615), .C(n3616) );
  CKBD0 U3498 ( .CLK(n3616), .C(n3617) );
  CKBD0 U3499 ( .CLK(n3617), .C(n3618) );
  CKBD0 U3500 ( .CLK(n3618), .C(n3619) );
  CKBD0 U3501 ( .CLK(n3619), .C(n3620) );
  BUFFD0 U3502 ( .I(n3620), .Z(n3621) );
  CKBD0 U3503 ( .CLK(n3621), .C(n3622) );
  CKBD0 U3504 ( .CLK(n3622), .C(n3623) );
  CKBD0 U3505 ( .CLK(n3623), .C(n3624) );
  CKBD0 U3506 ( .CLK(n3624), .C(n3625) );
  CKBD0 U3507 ( .CLK(n3625), .C(n3626) );
  CKBD0 U3508 ( .CLK(n3626), .C(n3627) );
  BUFFD0 U3509 ( .I(n3627), .Z(n3628) );
  CKBD0 U3510 ( .CLK(n3628), .C(n3629) );
  BUFFD0 U3511 ( .I(n3629), .Z(n3630) );
  CKBD0 U3512 ( .CLK(n3630), .C(n3631) );
  BUFFD0 U3513 ( .I(n3631), .Z(n3632) );
  CKBD0 U3514 ( .CLK(n3632), .C(n3633) );
  BUFFD0 U3515 ( .I(n3633), .Z(n3634) );
  CKBD0 U3516 ( .CLK(n3634), .C(n3635) );
  BUFFD0 U3517 ( .I(n3635), .Z(n3636) );
  CKBD0 U3518 ( .CLK(n3636), .C(n3637) );
  BUFFD0 U3519 ( .I(n3637), .Z(n3638) );
  CKBD0 U3520 ( .CLK(n3638), .C(n3639) );
  BUFFD0 U3521 ( .I(n3639), .Z(n3640) );
  CKBD0 U3522 ( .CLK(n3640), .C(n3641) );
  BUFFD0 U3523 ( .I(n3641), .Z(n3642) );
  BUFFD0 U3524 ( .I(n3644), .Z(n3643) );
  BUFFD0 U3525 ( .I(n3645), .Z(n3644) );
  BUFFD0 U3526 ( .I(n9166), .Z(n3645) );
  CKBD0 U3527 ( .CLK(n1861), .C(n3646) );
  CKBD0 U3528 ( .CLK(n3646), .C(n3647) );
  CKBD0 U3529 ( .CLK(n3647), .C(n3648) );
  BUFFD0 U3530 ( .I(n3648), .Z(n3649) );
  CKBD0 U3531 ( .CLK(n3649), .C(n3650) );
  CKBD0 U3532 ( .CLK(n3650), .C(n3651) );
  CKBD0 U3533 ( .CLK(n3651), .C(n3652) );
  CKBD0 U3534 ( .CLK(n3652), .C(n3653) );
  CKBD0 U3535 ( .CLK(n3653), .C(n3654) );
  CKBD0 U3536 ( .CLK(n3654), .C(n3655) );
  CKBD0 U3537 ( .CLK(n3655), .C(n3656) );
  CKBD0 U3538 ( .CLK(n3656), .C(n3657) );
  CKBD0 U3539 ( .CLK(n3657), .C(n3658) );
  CKBD0 U3540 ( .CLK(n3658), .C(n3659) );
  BUFFD0 U3541 ( .I(n3659), .Z(n3660) );
  CKBD0 U3542 ( .CLK(n3660), .C(n3661) );
  CKBD0 U3543 ( .CLK(n3661), .C(n3662) );
  CKBD0 U3544 ( .CLK(n3662), .C(n3663) );
  CKBD0 U3545 ( .CLK(n3663), .C(n3664) );
  CKBD0 U3546 ( .CLK(n3664), .C(n3665) );
  CKBD0 U3547 ( .CLK(n3665), .C(n3666) );
  CKBD0 U3548 ( .CLK(n3666), .C(n3667) );
  CKBD0 U3549 ( .CLK(n3667), .C(n3668) );
  CKBD0 U3550 ( .CLK(n3668), .C(n3669) );
  BUFFD0 U3551 ( .I(n3669), .Z(n3670) );
  CKBD0 U3552 ( .CLK(n3670), .C(n3671) );
  CKBD0 U3553 ( .CLK(n3671), .C(n3672) );
  CKBD0 U3554 ( .CLK(n3672), .C(n3673) );
  CKBD0 U3555 ( .CLK(n3673), .C(n3674) );
  CKBD0 U3556 ( .CLK(n3674), .C(n3675) );
  CKBD0 U3557 ( .CLK(n3675), .C(n3676) );
  CKBD0 U3558 ( .CLK(n3676), .C(n3677) );
  CKBD0 U3559 ( .CLK(n3677), .C(n3678) );
  CKBD0 U3560 ( .CLK(n3678), .C(n3679) );
  CKBD0 U3561 ( .CLK(n3679), .C(n3680) );
  BUFFD0 U3562 ( .I(n3680), .Z(n3681) );
  CKBD0 U3563 ( .CLK(n3681), .C(n3682) );
  CKBD0 U3564 ( .CLK(n3682), .C(n3683) );
  CKBD0 U3565 ( .CLK(n3683), .C(n3684) );
  CKBD0 U3566 ( .CLK(n3684), .C(n3685) );
  CKBD0 U3567 ( .CLK(n3685), .C(n3686) );
  CKBD0 U3568 ( .CLK(n3686), .C(n3687) );
  CKBD0 U3569 ( .CLK(n3687), .C(n3688) );
  CKBD0 U3570 ( .CLK(n3688), .C(n3689) );
  CKBD0 U3571 ( .CLK(n3689), .C(n3690) );
  CKBD0 U3572 ( .CLK(n3690), .C(n3691) );
  BUFFD0 U3573 ( .I(n3691), .Z(n3692) );
  CKBD0 U3574 ( .CLK(n3692), .C(n3693) );
  CKBD0 U3575 ( .CLK(n3693), .C(n3694) );
  CKBD0 U3576 ( .CLK(n3694), .C(n3695) );
  CKBD0 U3577 ( .CLK(n3695), .C(n3696) );
  CKBD0 U3578 ( .CLK(n3696), .C(n3697) );
  CKBD0 U3579 ( .CLK(n3697), .C(n3698) );
  CKBD0 U3580 ( .CLK(n3698), .C(n3699) );
  CKBD0 U3581 ( .CLK(n3699), .C(n3700) );
  CKBD0 U3582 ( .CLK(n3700), .C(n3701) );
  CKBD0 U3583 ( .CLK(n3701), .C(n3702) );
  BUFFD0 U3584 ( .I(n3702), .Z(n3703) );
  CKBD0 U3585 ( .CLK(n3703), .C(n3704) );
  CKBD0 U3586 ( .CLK(n3704), .C(n3705) );
  CKBD0 U3587 ( .CLK(n3705), .C(n3706) );
  CKBD0 U3588 ( .CLK(n3706), .C(n3707) );
  CKBD0 U3589 ( .CLK(n3707), .C(n3708) );
  CKBD0 U3590 ( .CLK(n3708), .C(n3709) );
  CKBD0 U3591 ( .CLK(n3709), .C(n3710) );
  CKBD0 U3592 ( .CLK(n3710), .C(n3711) );
  CKBD0 U3593 ( .CLK(n3711), .C(n3712) );
  CKBD0 U3594 ( .CLK(n3712), .C(n3713) );
  BUFFD0 U3595 ( .I(n3713), .Z(n3714) );
  CKBD0 U3596 ( .CLK(n3714), .C(n3715) );
  CKBD0 U3597 ( .CLK(n3715), .C(n3716) );
  CKBD0 U3598 ( .CLK(n3716), .C(n3717) );
  CKBD0 U3599 ( .CLK(n3717), .C(n3718) );
  CKBD0 U3600 ( .CLK(n3718), .C(n3719) );
  CKBD0 U3601 ( .CLK(n3719), .C(n3720) );
  CKBD0 U3602 ( .CLK(n3720), .C(n3721) );
  CKBD0 U3603 ( .CLK(n3721), .C(n3722) );
  CKBD0 U3604 ( .CLK(n3722), .C(n3723) );
  CKBD0 U3605 ( .CLK(n3723), .C(n3724) );
  BUFFD0 U3606 ( .I(n3724), .Z(n3725) );
  CKBD0 U3607 ( .CLK(n3725), .C(n3726) );
  CKBD0 U3608 ( .CLK(n3726), .C(n3727) );
  CKBD0 U3609 ( .CLK(n3727), .C(n3728) );
  CKBD0 U3610 ( .CLK(n3728), .C(n3729) );
  CKBD0 U3611 ( .CLK(n3729), .C(n3730) );
  CKBD0 U3612 ( .CLK(n3730), .C(n3731) );
  CKBD0 U3613 ( .CLK(n3731), .C(n3732) );
  CKBD0 U3614 ( .CLK(n3732), .C(n3733) );
  CKBD0 U3615 ( .CLK(n3733), .C(n3734) );
  BUFFD0 U3616 ( .I(n3734), .Z(n3735) );
  CKBD0 U3617 ( .CLK(n3735), .C(n3736) );
  CKBD0 U3618 ( .CLK(n3736), .C(n3737) );
  CKBD0 U3619 ( .CLK(n3737), .C(n3738) );
  CKBD0 U3620 ( .CLK(n3738), .C(n3739) );
  CKBD0 U3621 ( .CLK(n3739), .C(n3740) );
  CKBD0 U3622 ( .CLK(n3740), .C(n3741) );
  CKBD0 U3623 ( .CLK(n3741), .C(n3742) );
  CKBD0 U3624 ( .CLK(n3742), .C(n3743) );
  CKBD0 U3625 ( .CLK(n3743), .C(n3744) );
  CKBD0 U3626 ( .CLK(n3744), .C(n3745) );
  BUFFD0 U3627 ( .I(n3745), .Z(n3746) );
  CKBD0 U3628 ( .CLK(n3746), .C(n3747) );
  CKBD0 U3629 ( .CLK(n3747), .C(n3748) );
  CKBD0 U3630 ( .CLK(n3748), .C(n3749) );
  CKBD0 U3631 ( .CLK(n3749), .C(n3750) );
  CKBD0 U3632 ( .CLK(n3750), .C(n3751) );
  CKBD0 U3633 ( .CLK(n3751), .C(n3752) );
  CKBD0 U3634 ( .CLK(n3752), .C(n3753) );
  CKBD0 U3635 ( .CLK(n3753), .C(n3754) );
  CKBD0 U3636 ( .CLK(n3754), .C(n3755) );
  CKBD0 U3637 ( .CLK(n3755), .C(n3756) );
  BUFFD0 U3638 ( .I(n3756), .Z(n3757) );
  CKBD0 U3639 ( .CLK(n3757), .C(n3758) );
  CKBD0 U3640 ( .CLK(n3758), .C(n3759) );
  CKBD0 U3641 ( .CLK(n3759), .C(n3760) );
  CKBD0 U3642 ( .CLK(n3760), .C(n3761) );
  CKBD0 U3643 ( .CLK(n3761), .C(n3762) );
  CKBD0 U3644 ( .CLK(n3762), .C(n3763) );
  BUFFD0 U3645 ( .I(n3763), .Z(n3764) );
  CKBD0 U3646 ( .CLK(n3764), .C(n3765) );
  BUFFD0 U3647 ( .I(n3765), .Z(n3766) );
  CKBD0 U3648 ( .CLK(n3766), .C(n3767) );
  BUFFD0 U3649 ( .I(n3767), .Z(n3768) );
  CKBD0 U3650 ( .CLK(n3768), .C(n3769) );
  BUFFD0 U3651 ( .I(n3769), .Z(n3770) );
  CKBD0 U3652 ( .CLK(n3770), .C(n3771) );
  BUFFD0 U3653 ( .I(n3771), .Z(n3772) );
  CKBD0 U3654 ( .CLK(n3772), .C(n3773) );
  BUFFD0 U3655 ( .I(n3773), .Z(n3774) );
  CKBD0 U3656 ( .CLK(n3774), .C(n3775) );
  BUFFD0 U3657 ( .I(n3775), .Z(n3776) );
  CKBD0 U3658 ( .CLK(n3776), .C(n3777) );
  BUFFD0 U3659 ( .I(n3777), .Z(n3778) );
  BUFFD0 U3660 ( .I(n3780), .Z(n3779) );
  BUFFD0 U3661 ( .I(n3781), .Z(n3780) );
  BUFFD0 U3662 ( .I(n9167), .Z(n3781) );
  CKBD0 U3663 ( .CLK(n1254), .C(n3782) );
  CKBD0 U3664 ( .CLK(n3782), .C(n3783) );
  CKBD0 U3665 ( .CLK(n3783), .C(n3784) );
  BUFFD0 U3666 ( .I(n3784), .Z(n3785) );
  CKBD0 U3667 ( .CLK(n3785), .C(n3786) );
  CKBD0 U3668 ( .CLK(n3786), .C(n3787) );
  CKBD0 U3669 ( .CLK(n3787), .C(n3788) );
  CKBD0 U3670 ( .CLK(n3788), .C(n3789) );
  CKBD0 U3671 ( .CLK(n3789), .C(n3790) );
  CKBD0 U3672 ( .CLK(n3790), .C(n3791) );
  CKBD0 U3673 ( .CLK(n3791), .C(n3792) );
  CKBD0 U3674 ( .CLK(n3792), .C(n3793) );
  CKBD0 U3675 ( .CLK(n3793), .C(n3794) );
  CKBD0 U3676 ( .CLK(n3794), .C(n3795) );
  BUFFD0 U3677 ( .I(n3795), .Z(n3796) );
  CKBD0 U3678 ( .CLK(n3796), .C(n3797) );
  CKBD0 U3679 ( .CLK(n3797), .C(n3798) );
  CKBD0 U3680 ( .CLK(n3798), .C(n3799) );
  CKBD0 U3681 ( .CLK(n3799), .C(n3800) );
  CKBD0 U3682 ( .CLK(n3800), .C(n3801) );
  CKBD0 U3683 ( .CLK(n3801), .C(n3802) );
  CKBD0 U3684 ( .CLK(n3802), .C(n3803) );
  CKBD0 U3685 ( .CLK(n3803), .C(n3804) );
  CKBD0 U3686 ( .CLK(n3804), .C(n3805) );
  BUFFD0 U3687 ( .I(n3805), .Z(n3806) );
  CKBD0 U3688 ( .CLK(n3806), .C(n3807) );
  CKBD0 U3689 ( .CLK(n3807), .C(n3808) );
  CKBD0 U3690 ( .CLK(n3808), .C(n3809) );
  CKBD0 U3691 ( .CLK(n3809), .C(n3810) );
  CKBD0 U3692 ( .CLK(n3810), .C(n3811) );
  CKBD0 U3693 ( .CLK(n3811), .C(n3812) );
  CKBD0 U3694 ( .CLK(n3812), .C(n3813) );
  CKBD0 U3695 ( .CLK(n3813), .C(n3814) );
  CKBD0 U3696 ( .CLK(n3814), .C(n3815) );
  CKBD0 U3697 ( .CLK(n3815), .C(n3816) );
  BUFFD0 U3698 ( .I(n3816), .Z(n3817) );
  CKBD0 U3699 ( .CLK(n3817), .C(n3818) );
  CKBD0 U3700 ( .CLK(n3818), .C(n3819) );
  CKBD0 U3701 ( .CLK(n3819), .C(n3820) );
  CKBD0 U3702 ( .CLK(n3820), .C(n3821) );
  CKBD0 U3703 ( .CLK(n3821), .C(n3822) );
  CKBD0 U3704 ( .CLK(n3822), .C(n3823) );
  CKBD0 U3705 ( .CLK(n3823), .C(n3824) );
  CKBD0 U3706 ( .CLK(n3824), .C(n3825) );
  CKBD0 U3707 ( .CLK(n3825), .C(n3826) );
  CKBD0 U3708 ( .CLK(n3826), .C(n3827) );
  BUFFD0 U3709 ( .I(n3827), .Z(n3828) );
  CKBD0 U3710 ( .CLK(n3828), .C(n3829) );
  CKBD0 U3711 ( .CLK(n3829), .C(n3830) );
  CKBD0 U3712 ( .CLK(n3830), .C(n3831) );
  CKBD0 U3713 ( .CLK(n3831), .C(n3832) );
  CKBD0 U3714 ( .CLK(n3832), .C(n3833) );
  CKBD0 U3715 ( .CLK(n3833), .C(n3834) );
  CKBD0 U3716 ( .CLK(n3834), .C(n3835) );
  CKBD0 U3717 ( .CLK(n3835), .C(n3836) );
  CKBD0 U3718 ( .CLK(n3836), .C(n3837) );
  CKBD0 U3719 ( .CLK(n3837), .C(n3838) );
  BUFFD0 U3720 ( .I(n3838), .Z(n3839) );
  CKBD0 U3721 ( .CLK(n3839), .C(n3840) );
  CKBD0 U3722 ( .CLK(n3840), .C(n3841) );
  CKBD0 U3723 ( .CLK(n3841), .C(n3842) );
  CKBD0 U3724 ( .CLK(n3842), .C(n3843) );
  CKBD0 U3725 ( .CLK(n3843), .C(n3844) );
  CKBD0 U3726 ( .CLK(n3844), .C(n3845) );
  CKBD0 U3727 ( .CLK(n3845), .C(n3846) );
  CKBD0 U3728 ( .CLK(n3846), .C(n3847) );
  CKBD0 U3729 ( .CLK(n3847), .C(n3848) );
  CKBD0 U3730 ( .CLK(n3848), .C(n3849) );
  BUFFD0 U3731 ( .I(n3849), .Z(n3850) );
  CKBD0 U3732 ( .CLK(n3850), .C(n3851) );
  CKBD0 U3733 ( .CLK(n3851), .C(n3852) );
  CKBD0 U3734 ( .CLK(n3852), .C(n3853) );
  CKBD0 U3735 ( .CLK(n3853), .C(n3854) );
  CKBD0 U3736 ( .CLK(n3854), .C(n3855) );
  CKBD0 U3737 ( .CLK(n3855), .C(n3856) );
  CKBD0 U3738 ( .CLK(n3856), .C(n3857) );
  CKBD0 U3739 ( .CLK(n3857), .C(n3858) );
  CKBD0 U3740 ( .CLK(n3858), .C(n3859) );
  CKBD0 U3741 ( .CLK(n3859), .C(n3860) );
  BUFFD0 U3742 ( .I(n3860), .Z(n3861) );
  CKBD0 U3743 ( .CLK(n3861), .C(n3862) );
  CKBD0 U3744 ( .CLK(n3862), .C(n3863) );
  CKBD0 U3745 ( .CLK(n3863), .C(n3864) );
  CKBD0 U3746 ( .CLK(n3864), .C(n3865) );
  CKBD0 U3747 ( .CLK(n3865), .C(n3866) );
  CKBD0 U3748 ( .CLK(n3866), .C(n3867) );
  CKBD0 U3749 ( .CLK(n3867), .C(n3868) );
  CKBD0 U3750 ( .CLK(n3868), .C(n3869) );
  CKBD0 U3751 ( .CLK(n3869), .C(n3870) );
  BUFFD0 U3752 ( .I(n3870), .Z(n3871) );
  CKBD0 U3753 ( .CLK(n3871), .C(n3872) );
  CKBD0 U3754 ( .CLK(n3872), .C(n3873) );
  CKBD0 U3755 ( .CLK(n3873), .C(n3874) );
  CKBD0 U3756 ( .CLK(n3874), .C(n3875) );
  CKBD0 U3757 ( .CLK(n3875), .C(n3876) );
  CKBD0 U3758 ( .CLK(n3876), .C(n3877) );
  CKBD0 U3759 ( .CLK(n3877), .C(n3878) );
  CKBD0 U3760 ( .CLK(n3878), .C(n3879) );
  CKBD0 U3761 ( .CLK(n3879), .C(n3880) );
  CKBD0 U3762 ( .CLK(n3880), .C(n3881) );
  BUFFD0 U3763 ( .I(n3881), .Z(n3882) );
  CKBD0 U3764 ( .CLK(n3882), .C(n3883) );
  CKBD0 U3765 ( .CLK(n3883), .C(n3884) );
  CKBD0 U3766 ( .CLK(n3884), .C(n3885) );
  CKBD0 U3767 ( .CLK(n3885), .C(n3886) );
  CKBD0 U3768 ( .CLK(n3886), .C(n3887) );
  CKBD0 U3769 ( .CLK(n3887), .C(n3888) );
  CKBD0 U3770 ( .CLK(n3888), .C(n3889) );
  CKBD0 U3771 ( .CLK(n3889), .C(n3890) );
  CKBD0 U3772 ( .CLK(n3890), .C(n3891) );
  CKBD0 U3773 ( .CLK(n3891), .C(n3892) );
  BUFFD0 U3774 ( .I(n3892), .Z(n3893) );
  CKBD0 U3775 ( .CLK(n3893), .C(n3894) );
  CKBD0 U3776 ( .CLK(n3894), .C(n3895) );
  CKBD0 U3777 ( .CLK(n3895), .C(n3896) );
  CKBD0 U3778 ( .CLK(n3896), .C(n3897) );
  CKBD0 U3779 ( .CLK(n3897), .C(n3898) );
  CKBD0 U3780 ( .CLK(n3898), .C(n3899) );
  BUFFD0 U3781 ( .I(n3899), .Z(n3900) );
  CKBD0 U3782 ( .CLK(n3900), .C(n3901) );
  BUFFD0 U3783 ( .I(n3901), .Z(n3902) );
  CKBD0 U3784 ( .CLK(n3902), .C(n3903) );
  BUFFD0 U3785 ( .I(n3903), .Z(n3904) );
  CKBD0 U3786 ( .CLK(n3904), .C(n3905) );
  BUFFD0 U3787 ( .I(n3905), .Z(n3906) );
  CKBD0 U3788 ( .CLK(n3906), .C(n3907) );
  BUFFD0 U3789 ( .I(n3907), .Z(n3908) );
  CKBD0 U3790 ( .CLK(n3908), .C(n3909) );
  BUFFD0 U3791 ( .I(n3909), .Z(n3910) );
  CKBD0 U3792 ( .CLK(n3910), .C(n3911) );
  BUFFD0 U3793 ( .I(n3911), .Z(n3912) );
  CKBD0 U3794 ( .CLK(n3912), .C(n3913) );
  BUFFD0 U3795 ( .I(n3913), .Z(n3914) );
  BUFFD0 U3796 ( .I(n3916), .Z(n3915) );
  BUFFD0 U3797 ( .I(n3917), .Z(n3916) );
  BUFFD0 U3798 ( .I(n9168), .Z(n3917) );
  CKBD0 U3799 ( .CLK(n1252), .C(n3918) );
  CKBD0 U3800 ( .CLK(n3918), .C(n3919) );
  CKBD0 U3801 ( .CLK(n3919), .C(n3920) );
  BUFFD0 U3802 ( .I(n3920), .Z(n3921) );
  CKBD0 U3803 ( .CLK(n3921), .C(n3922) );
  CKBD0 U3804 ( .CLK(n3922), .C(n3923) );
  CKBD0 U3805 ( .CLK(n3923), .C(n3924) );
  CKBD0 U3806 ( .CLK(n3924), .C(n3925) );
  CKBD0 U3807 ( .CLK(n3925), .C(n3926) );
  CKBD0 U3808 ( .CLK(n3926), .C(n3927) );
  CKBD0 U3809 ( .CLK(n3927), .C(n3928) );
  CKBD0 U3810 ( .CLK(n3928), .C(n3929) );
  CKBD0 U3811 ( .CLK(n3929), .C(n3930) );
  CKBD0 U3812 ( .CLK(n3930), .C(n3931) );
  BUFFD0 U3813 ( .I(n3931), .Z(n3932) );
  CKBD0 U3814 ( .CLK(n3932), .C(n3933) );
  CKBD0 U3815 ( .CLK(n3933), .C(n3934) );
  CKBD0 U3816 ( .CLK(n3934), .C(n3935) );
  CKBD0 U3817 ( .CLK(n3935), .C(n3936) );
  CKBD0 U3818 ( .CLK(n3936), .C(n3937) );
  CKBD0 U3819 ( .CLK(n3937), .C(n3938) );
  CKBD0 U3820 ( .CLK(n3938), .C(n3939) );
  CKBD0 U3821 ( .CLK(n3939), .C(n3940) );
  CKBD0 U3822 ( .CLK(n3940), .C(n3941) );
  BUFFD0 U3823 ( .I(n3941), .Z(n3942) );
  CKBD0 U3824 ( .CLK(n3942), .C(n3943) );
  CKBD0 U3825 ( .CLK(n3943), .C(n3944) );
  CKBD0 U3826 ( .CLK(n3944), .C(n3945) );
  CKBD0 U3827 ( .CLK(n3945), .C(n3946) );
  CKBD0 U3828 ( .CLK(n3946), .C(n3947) );
  CKBD0 U3829 ( .CLK(n3947), .C(n3948) );
  CKBD0 U3830 ( .CLK(n3948), .C(n3949) );
  CKBD0 U3831 ( .CLK(n3949), .C(n3950) );
  CKBD0 U3832 ( .CLK(n3950), .C(n3951) );
  CKBD0 U3833 ( .CLK(n3951), .C(n3952) );
  BUFFD0 U3834 ( .I(n3952), .Z(n3953) );
  CKBD0 U3835 ( .CLK(n3953), .C(n3954) );
  CKBD0 U3836 ( .CLK(n3954), .C(n3955) );
  CKBD0 U3837 ( .CLK(n3955), .C(n3956) );
  CKBD0 U3838 ( .CLK(n3956), .C(n3957) );
  CKBD0 U3839 ( .CLK(n3957), .C(n3958) );
  CKBD0 U3840 ( .CLK(n3958), .C(n3959) );
  CKBD0 U3841 ( .CLK(n3959), .C(n3960) );
  CKBD0 U3842 ( .CLK(n3960), .C(n3961) );
  CKBD0 U3843 ( .CLK(n3961), .C(n3962) );
  CKBD0 U3844 ( .CLK(n3962), .C(n3963) );
  BUFFD0 U3845 ( .I(n3963), .Z(n3964) );
  CKBD0 U3846 ( .CLK(n3964), .C(n3965) );
  CKBD0 U3847 ( .CLK(n3965), .C(n3966) );
  CKBD0 U3848 ( .CLK(n3966), .C(n3967) );
  CKBD0 U3849 ( .CLK(n3967), .C(n3968) );
  CKBD0 U3850 ( .CLK(n3968), .C(n3969) );
  CKBD0 U3851 ( .CLK(n3969), .C(n3970) );
  CKBD0 U3852 ( .CLK(n3970), .C(n3971) );
  CKBD0 U3853 ( .CLK(n3971), .C(n3972) );
  CKBD0 U3854 ( .CLK(n3972), .C(n3973) );
  CKBD0 U3855 ( .CLK(n3973), .C(n3974) );
  BUFFD0 U3856 ( .I(n3974), .Z(n3975) );
  CKBD0 U3857 ( .CLK(n3975), .C(n3976) );
  CKBD0 U3858 ( .CLK(n3976), .C(n3977) );
  CKBD0 U3859 ( .CLK(n3977), .C(n3978) );
  CKBD0 U3860 ( .CLK(n3978), .C(n3979) );
  CKBD0 U3861 ( .CLK(n3979), .C(n3980) );
  CKBD0 U3862 ( .CLK(n3980), .C(n3981) );
  CKBD0 U3863 ( .CLK(n3981), .C(n3982) );
  CKBD0 U3864 ( .CLK(n3982), .C(n3983) );
  CKBD0 U3865 ( .CLK(n3983), .C(n3984) );
  CKBD0 U3866 ( .CLK(n3984), .C(n3985) );
  BUFFD0 U3867 ( .I(n3985), .Z(n3986) );
  CKBD0 U3868 ( .CLK(n3986), .C(n3987) );
  CKBD0 U3869 ( .CLK(n3987), .C(n3988) );
  CKBD0 U3870 ( .CLK(n3988), .C(n3989) );
  CKBD0 U3871 ( .CLK(n3989), .C(n3990) );
  CKBD0 U3872 ( .CLK(n3990), .C(n3991) );
  CKBD0 U3873 ( .CLK(n3991), .C(n3992) );
  CKBD0 U3874 ( .CLK(n3992), .C(n3993) );
  CKBD0 U3875 ( .CLK(n3993), .C(n3994) );
  CKBD0 U3876 ( .CLK(n3994), .C(n3995) );
  CKBD0 U3877 ( .CLK(n3995), .C(n3996) );
  BUFFD0 U3878 ( .I(n3996), .Z(n3997) );
  CKBD0 U3879 ( .CLK(n3997), .C(n3998) );
  CKBD0 U3880 ( .CLK(n3998), .C(n3999) );
  CKBD0 U3881 ( .CLK(n3999), .C(n4000) );
  CKBD0 U3882 ( .CLK(n4000), .C(n4001) );
  CKBD0 U3883 ( .CLK(n4001), .C(n4002) );
  CKBD0 U3884 ( .CLK(n4002), .C(n4003) );
  CKBD0 U3885 ( .CLK(n4003), .C(n4004) );
  CKBD0 U3886 ( .CLK(n4004), .C(n4005) );
  CKBD0 U3887 ( .CLK(n4005), .C(n4006) );
  BUFFD0 U3888 ( .I(n4006), .Z(n4007) );
  CKBD0 U3889 ( .CLK(n4007), .C(n4008) );
  CKBD0 U3890 ( .CLK(n4008), .C(n4009) );
  CKBD0 U3891 ( .CLK(n4009), .C(n4010) );
  CKBD0 U3892 ( .CLK(n4010), .C(n4011) );
  CKBD0 U3893 ( .CLK(n4011), .C(n4012) );
  CKBD0 U3894 ( .CLK(n4012), .C(n4013) );
  CKBD0 U3895 ( .CLK(n4013), .C(n4014) );
  CKBD0 U3896 ( .CLK(n4014), .C(n4015) );
  CKBD0 U3897 ( .CLK(n4015), .C(n4016) );
  CKBD0 U3898 ( .CLK(n4016), .C(n4017) );
  BUFFD0 U3899 ( .I(n4017), .Z(n4018) );
  CKBD0 U3900 ( .CLK(n4018), .C(n4019) );
  CKBD0 U3901 ( .CLK(n4019), .C(n4020) );
  CKBD0 U3902 ( .CLK(n4020), .C(n4021) );
  CKBD0 U3903 ( .CLK(n4021), .C(n4022) );
  CKBD0 U3904 ( .CLK(n4022), .C(n4023) );
  CKBD0 U3905 ( .CLK(n4023), .C(n4024) );
  CKBD0 U3906 ( .CLK(n4024), .C(n4025) );
  CKBD0 U3907 ( .CLK(n4025), .C(n4026) );
  CKBD0 U3908 ( .CLK(n4026), .C(n4027) );
  CKBD0 U3909 ( .CLK(n4027), .C(n4028) );
  BUFFD0 U3910 ( .I(n4028), .Z(n4029) );
  CKBD0 U3911 ( .CLK(n4029), .C(n4030) );
  CKBD0 U3912 ( .CLK(n4030), .C(n4031) );
  CKBD0 U3913 ( .CLK(n4031), .C(n4032) );
  CKBD0 U3914 ( .CLK(n4032), .C(n4033) );
  CKBD0 U3915 ( .CLK(n4033), .C(n4034) );
  CKBD0 U3916 ( .CLK(n4034), .C(n4035) );
  BUFFD0 U3917 ( .I(n4035), .Z(n4036) );
  CKBD0 U3918 ( .CLK(n4036), .C(n4037) );
  BUFFD0 U3919 ( .I(n4037), .Z(n4038) );
  CKBD0 U3920 ( .CLK(n4038), .C(n4039) );
  BUFFD0 U3921 ( .I(n4039), .Z(n4040) );
  CKBD0 U3922 ( .CLK(n4040), .C(n4041) );
  BUFFD0 U3923 ( .I(n4041), .Z(n4042) );
  CKBD0 U3924 ( .CLK(n4042), .C(n4043) );
  BUFFD0 U3925 ( .I(n4043), .Z(n4044) );
  CKBD0 U3926 ( .CLK(n4044), .C(n4045) );
  BUFFD0 U3927 ( .I(n4045), .Z(n4046) );
  CKBD0 U3928 ( .CLK(n4046), .C(n4047) );
  BUFFD0 U3929 ( .I(n4047), .Z(n4048) );
  CKBD0 U3930 ( .CLK(n4048), .C(n4049) );
  BUFFD0 U3931 ( .I(n4049), .Z(n4050) );
  BUFFD0 U3932 ( .I(n4052), .Z(n4051) );
  BUFFD0 U3933 ( .I(n4053), .Z(n4052) );
  BUFFD0 U3934 ( .I(n9169), .Z(n4053) );
  CKBD0 U3935 ( .CLK(n1250), .C(n4054) );
  CKBD0 U3936 ( .CLK(n4054), .C(n4055) );
  CKBD0 U3937 ( .CLK(n4055), .C(n4056) );
  BUFFD0 U3938 ( .I(n4056), .Z(n4057) );
  CKBD0 U3939 ( .CLK(n4057), .C(n4058) );
  CKBD0 U3940 ( .CLK(n4058), .C(n4059) );
  CKBD0 U3941 ( .CLK(n4059), .C(n4060) );
  CKBD0 U3942 ( .CLK(n4060), .C(n4061) );
  CKBD0 U3943 ( .CLK(n4061), .C(n4062) );
  CKBD0 U3944 ( .CLK(n4062), .C(n4063) );
  CKBD0 U3945 ( .CLK(n4063), .C(n4064) );
  CKBD0 U3946 ( .CLK(n4064), .C(n4065) );
  CKBD0 U3947 ( .CLK(n4065), .C(n4066) );
  CKBD0 U3948 ( .CLK(n4066), .C(n4067) );
  BUFFD0 U3949 ( .I(n4067), .Z(n4068) );
  CKBD0 U3950 ( .CLK(n4068), .C(n4069) );
  CKBD0 U3951 ( .CLK(n4069), .C(n4070) );
  CKBD0 U3952 ( .CLK(n4070), .C(n4071) );
  CKBD0 U3953 ( .CLK(n4071), .C(n4072) );
  CKBD0 U3954 ( .CLK(n4072), .C(n4073) );
  CKBD0 U3955 ( .CLK(n4073), .C(n4074) );
  CKBD0 U3956 ( .CLK(n4074), .C(n4075) );
  CKBD0 U3957 ( .CLK(n4075), .C(n4076) );
  CKBD0 U3958 ( .CLK(n4076), .C(n4077) );
  BUFFD0 U3959 ( .I(n4077), .Z(n4078) );
  CKBD0 U3960 ( .CLK(n4078), .C(n4079) );
  CKBD0 U3961 ( .CLK(n4079), .C(n4080) );
  CKBD0 U3962 ( .CLK(n4080), .C(n4081) );
  CKBD0 U3963 ( .CLK(n4081), .C(n4082) );
  CKBD0 U3964 ( .CLK(n4082), .C(n4083) );
  CKBD0 U3965 ( .CLK(n4083), .C(n4084) );
  CKBD0 U3966 ( .CLK(n4084), .C(n4085) );
  CKBD0 U3967 ( .CLK(n4085), .C(n4086) );
  CKBD0 U3968 ( .CLK(n4086), .C(n4087) );
  CKBD0 U3969 ( .CLK(n4087), .C(n4088) );
  BUFFD0 U3970 ( .I(n4088), .Z(n4089) );
  CKBD0 U3971 ( .CLK(n4089), .C(n4090) );
  CKBD0 U3972 ( .CLK(n4090), .C(n4091) );
  CKBD0 U3973 ( .CLK(n4091), .C(n4092) );
  CKBD0 U3974 ( .CLK(n4092), .C(n4093) );
  CKBD0 U3975 ( .CLK(n4093), .C(n4094) );
  CKBD0 U3976 ( .CLK(n4094), .C(n4095) );
  CKBD0 U3977 ( .CLK(n4095), .C(n4096) );
  CKBD0 U3978 ( .CLK(n4096), .C(n4097) );
  CKBD0 U3979 ( .CLK(n4097), .C(n4098) );
  CKBD0 U3980 ( .CLK(n4098), .C(n4099) );
  BUFFD0 U3981 ( .I(n4099), .Z(n4100) );
  CKBD0 U3982 ( .CLK(n4100), .C(n4101) );
  CKBD0 U3983 ( .CLK(n4101), .C(n4102) );
  CKBD0 U3984 ( .CLK(n4102), .C(n4103) );
  CKBD0 U3985 ( .CLK(n4103), .C(n4104) );
  CKBD0 U3986 ( .CLK(n4104), .C(n4105) );
  CKBD0 U3987 ( .CLK(n4105), .C(n4106) );
  CKBD0 U3988 ( .CLK(n4106), .C(n4107) );
  CKBD0 U3989 ( .CLK(n4107), .C(n4108) );
  CKBD0 U3990 ( .CLK(n4108), .C(n4109) );
  CKBD0 U3991 ( .CLK(n4109), .C(n4110) );
  BUFFD0 U3992 ( .I(n4110), .Z(n4111) );
  CKBD0 U3993 ( .CLK(n4111), .C(n4112) );
  CKBD0 U3994 ( .CLK(n4112), .C(n4113) );
  CKBD0 U3995 ( .CLK(n4113), .C(n4114) );
  CKBD0 U3996 ( .CLK(n4114), .C(n4115) );
  CKBD0 U3997 ( .CLK(n4115), .C(n4116) );
  CKBD0 U3998 ( .CLK(n4116), .C(n4117) );
  CKBD0 U3999 ( .CLK(n4117), .C(n4118) );
  CKBD0 U4000 ( .CLK(n4118), .C(n4119) );
  CKBD0 U4001 ( .CLK(n4119), .C(n4120) );
  CKBD0 U4002 ( .CLK(n4120), .C(n4121) );
  BUFFD0 U4003 ( .I(n4121), .Z(n4122) );
  CKBD0 U4004 ( .CLK(n4122), .C(n4123) );
  CKBD0 U4005 ( .CLK(n4123), .C(n4124) );
  CKBD0 U4006 ( .CLK(n4124), .C(n4125) );
  CKBD0 U4007 ( .CLK(n4125), .C(n4126) );
  CKBD0 U4008 ( .CLK(n4126), .C(n4127) );
  CKBD0 U4009 ( .CLK(n4127), .C(n4128) );
  CKBD0 U4010 ( .CLK(n4128), .C(n4129) );
  CKBD0 U4011 ( .CLK(n4129), .C(n4130) );
  CKBD0 U4012 ( .CLK(n4130), .C(n4131) );
  CKBD0 U4013 ( .CLK(n4131), .C(n4132) );
  BUFFD0 U4014 ( .I(n4132), .Z(n4133) );
  CKBD0 U4015 ( .CLK(n4133), .C(n4134) );
  CKBD0 U4016 ( .CLK(n4134), .C(n4135) );
  CKBD0 U4017 ( .CLK(n4135), .C(n4136) );
  CKBD0 U4018 ( .CLK(n4136), .C(n4137) );
  CKBD0 U4019 ( .CLK(n4137), .C(n4138) );
  CKBD0 U4020 ( .CLK(n4138), .C(n4139) );
  CKBD0 U4021 ( .CLK(n4139), .C(n4140) );
  CKBD0 U4022 ( .CLK(n4140), .C(n4141) );
  CKBD0 U4023 ( .CLK(n4141), .C(n4142) );
  CKBD0 U4024 ( .CLK(n4142), .C(n4143) );
  BUFFD0 U4025 ( .I(n4143), .Z(n4144) );
  CKBD0 U4026 ( .CLK(n4144), .C(n4145) );
  CKBD0 U4027 ( .CLK(n4145), .C(n4146) );
  CKBD0 U4028 ( .CLK(n4146), .C(n4147) );
  CKBD0 U4029 ( .CLK(n4147), .C(n4148) );
  CKBD0 U4030 ( .CLK(n4148), .C(n4149) );
  CKBD0 U4031 ( .CLK(n4149), .C(n4150) );
  CKBD0 U4032 ( .CLK(n4150), .C(n4151) );
  CKBD0 U4033 ( .CLK(n4151), .C(n4152) );
  CKBD0 U4034 ( .CLK(n4152), .C(n4153) );
  BUFFD0 U4035 ( .I(n4153), .Z(n4154) );
  CKBD0 U4036 ( .CLK(n4154), .C(n4155) );
  CKBD0 U4037 ( .CLK(n4155), .C(n4156) );
  CKBD0 U4038 ( .CLK(n4156), .C(n4157) );
  CKBD0 U4039 ( .CLK(n4157), .C(n4158) );
  CKBD0 U4040 ( .CLK(n4158), .C(n4159) );
  CKBD0 U4041 ( .CLK(n4159), .C(n4160) );
  CKBD0 U4042 ( .CLK(n4160), .C(n4161) );
  CKBD0 U4043 ( .CLK(n4161), .C(n4162) );
  CKBD0 U4044 ( .CLK(n4162), .C(n4163) );
  CKBD0 U4045 ( .CLK(n4163), .C(n4164) );
  BUFFD0 U4046 ( .I(n4164), .Z(n4165) );
  CKBD0 U4047 ( .CLK(n4165), .C(n4166) );
  CKBD0 U4048 ( .CLK(n4166), .C(n4167) );
  CKBD0 U4049 ( .CLK(n4167), .C(n4168) );
  CKBD0 U4050 ( .CLK(n4168), .C(n4169) );
  CKBD0 U4051 ( .CLK(n4169), .C(n4170) );
  CKBD0 U4052 ( .CLK(n4170), .C(n4171) );
  BUFFD0 U4053 ( .I(n4171), .Z(n4172) );
  CKBD0 U4054 ( .CLK(n4172), .C(n4173) );
  BUFFD0 U4055 ( .I(n4173), .Z(n4174) );
  CKBD0 U4056 ( .CLK(n4174), .C(n4175) );
  BUFFD0 U4057 ( .I(n4175), .Z(n4176) );
  CKBD0 U4058 ( .CLK(n4176), .C(n4177) );
  BUFFD0 U4059 ( .I(n4177), .Z(n4178) );
  CKBD0 U4060 ( .CLK(n4178), .C(n4179) );
  BUFFD0 U4061 ( .I(n4179), .Z(n4180) );
  CKBD0 U4062 ( .CLK(n4180), .C(n4181) );
  BUFFD0 U4063 ( .I(n4181), .Z(n4182) );
  CKBD0 U4064 ( .CLK(n4182), .C(n4183) );
  BUFFD0 U4065 ( .I(n4183), .Z(n4184) );
  CKBD0 U4066 ( .CLK(n4184), .C(n4185) );
  BUFFD0 U4067 ( .I(n4185), .Z(n4186) );
  BUFFD0 U4068 ( .I(Decoder[19]), .Z(n4187) );
  BUFFD0 U4069 ( .I(n4189), .Z(n4188) );
  BUFFD0 U4070 ( .I(n4190), .Z(n4189) );
  BUFFD0 U4071 ( .I(n9170), .Z(n4190) );
  CKBD0 U4072 ( .CLK(n1248), .C(n4191) );
  CKBD0 U4073 ( .CLK(n4191), .C(n4192) );
  CKBD0 U4074 ( .CLK(n4192), .C(n4193) );
  BUFFD0 U4075 ( .I(n4193), .Z(n4194) );
  CKBD0 U4076 ( .CLK(n4194), .C(n4195) );
  CKBD0 U4077 ( .CLK(n4195), .C(n4196) );
  CKBD0 U4078 ( .CLK(n4196), .C(n4197) );
  CKBD0 U4079 ( .CLK(n4197), .C(n4198) );
  CKBD0 U4080 ( .CLK(n4198), .C(n4199) );
  CKBD0 U4081 ( .CLK(n4199), .C(n4200) );
  CKBD0 U4082 ( .CLK(n4200), .C(n4201) );
  CKBD0 U4083 ( .CLK(n4201), .C(n4202) );
  CKBD0 U4084 ( .CLK(n4202), .C(n4203) );
  CKBD0 U4085 ( .CLK(n4203), .C(n4204) );
  BUFFD0 U4086 ( .I(n4204), .Z(n4205) );
  CKBD0 U4087 ( .CLK(n4205), .C(n4206) );
  CKBD0 U4088 ( .CLK(n4206), .C(n4207) );
  CKBD0 U4089 ( .CLK(n4207), .C(n4208) );
  CKBD0 U4090 ( .CLK(n4208), .C(n4209) );
  CKBD0 U4091 ( .CLK(n4209), .C(n4210) );
  CKBD0 U4092 ( .CLK(n4210), .C(n4211) );
  CKBD0 U4093 ( .CLK(n4211), .C(n4212) );
  CKBD0 U4094 ( .CLK(n4212), .C(n4213) );
  CKBD0 U4095 ( .CLK(n4213), .C(n4214) );
  BUFFD0 U4096 ( .I(n4214), .Z(n4215) );
  CKBD0 U4097 ( .CLK(n4215), .C(n4216) );
  CKBD0 U4098 ( .CLK(n4216), .C(n4217) );
  CKBD0 U4099 ( .CLK(n4217), .C(n4218) );
  CKBD0 U4100 ( .CLK(n4218), .C(n4219) );
  CKBD0 U4101 ( .CLK(n4219), .C(n4220) );
  CKBD0 U4102 ( .CLK(n4220), .C(n4221) );
  CKBD0 U4103 ( .CLK(n4221), .C(n4222) );
  CKBD0 U4104 ( .CLK(n4222), .C(n4223) );
  CKBD0 U4105 ( .CLK(n4223), .C(n4224) );
  CKBD0 U4106 ( .CLK(n4224), .C(n4225) );
  BUFFD0 U4107 ( .I(n4225), .Z(n4226) );
  CKBD0 U4108 ( .CLK(n4226), .C(n4227) );
  CKBD0 U4109 ( .CLK(n4227), .C(n4228) );
  CKBD0 U4110 ( .CLK(n4228), .C(n4229) );
  CKBD0 U4111 ( .CLK(n4229), .C(n4230) );
  CKBD0 U4112 ( .CLK(n4230), .C(n4231) );
  CKBD0 U4113 ( .CLK(n4231), .C(n4232) );
  CKBD0 U4114 ( .CLK(n4232), .C(n4233) );
  CKBD0 U4115 ( .CLK(n4233), .C(n4234) );
  CKBD0 U4116 ( .CLK(n4234), .C(n4235) );
  CKBD0 U4117 ( .CLK(n4235), .C(n4236) );
  BUFFD0 U4118 ( .I(n4236), .Z(n4237) );
  CKBD0 U4119 ( .CLK(n4237), .C(n4238) );
  CKBD0 U4120 ( .CLK(n4238), .C(n4239) );
  CKBD0 U4121 ( .CLK(n4239), .C(n4240) );
  CKBD0 U4122 ( .CLK(n4240), .C(n4241) );
  CKBD0 U4123 ( .CLK(n4241), .C(n4242) );
  CKBD0 U4124 ( .CLK(n4242), .C(n4243) );
  CKBD0 U4125 ( .CLK(n4243), .C(n4244) );
  CKBD0 U4126 ( .CLK(n4244), .C(n4245) );
  CKBD0 U4127 ( .CLK(n4245), .C(n4246) );
  CKBD0 U4128 ( .CLK(n4246), .C(n4247) );
  BUFFD0 U4129 ( .I(n4247), .Z(n4248) );
  CKBD0 U4130 ( .CLK(n4248), .C(n4249) );
  CKBD0 U4131 ( .CLK(n4249), .C(n4250) );
  CKBD0 U4132 ( .CLK(n4250), .C(n4251) );
  CKBD0 U4133 ( .CLK(n4251), .C(n4252) );
  CKBD0 U4134 ( .CLK(n4252), .C(n4253) );
  CKBD0 U4135 ( .CLK(n4253), .C(n4254) );
  CKBD0 U4136 ( .CLK(n4254), .C(n4255) );
  CKBD0 U4137 ( .CLK(n4255), .C(n4256) );
  CKBD0 U4138 ( .CLK(n4256), .C(n4257) );
  CKBD0 U4139 ( .CLK(n4257), .C(n4258) );
  BUFFD0 U4140 ( .I(n4258), .Z(n4259) );
  CKBD0 U4141 ( .CLK(n4259), .C(n4260) );
  CKBD0 U4142 ( .CLK(n4260), .C(n4261) );
  CKBD0 U4143 ( .CLK(n4261), .C(n4262) );
  CKBD0 U4144 ( .CLK(n4262), .C(n4263) );
  CKBD0 U4145 ( .CLK(n4263), .C(n4264) );
  CKBD0 U4146 ( .CLK(n4264), .C(n4265) );
  CKBD0 U4147 ( .CLK(n4265), .C(n4266) );
  CKBD0 U4148 ( .CLK(n4266), .C(n4267) );
  CKBD0 U4149 ( .CLK(n4267), .C(n4268) );
  CKBD0 U4150 ( .CLK(n4268), .C(n4269) );
  BUFFD0 U4151 ( .I(n4269), .Z(n4270) );
  CKBD0 U4152 ( .CLK(n4270), .C(n4271) );
  CKBD0 U4153 ( .CLK(n4271), .C(n4272) );
  CKBD0 U4154 ( .CLK(n4272), .C(n4273) );
  CKBD0 U4155 ( .CLK(n4273), .C(n4274) );
  CKBD0 U4156 ( .CLK(n4274), .C(n4275) );
  CKBD0 U4157 ( .CLK(n4275), .C(n4276) );
  CKBD0 U4158 ( .CLK(n4276), .C(n4277) );
  CKBD0 U4159 ( .CLK(n4277), .C(n4278) );
  CKBD0 U4160 ( .CLK(n4278), .C(n4279) );
  CKBD0 U4161 ( .CLK(n4279), .C(n4280) );
  BUFFD0 U4162 ( .I(n4280), .Z(n4281) );
  CKBD0 U4163 ( .CLK(n4281), .C(n4282) );
  CKBD0 U4164 ( .CLK(n4282), .C(n4283) );
  CKBD0 U4165 ( .CLK(n4283), .C(n4284) );
  CKBD0 U4166 ( .CLK(n4284), .C(n4285) );
  CKBD0 U4167 ( .CLK(n4285), .C(n4286) );
  CKBD0 U4168 ( .CLK(n4286), .C(n4287) );
  CKBD0 U4169 ( .CLK(n4287), .C(n4288) );
  CKBD0 U4170 ( .CLK(n4288), .C(n4289) );
  CKBD0 U4171 ( .CLK(n4289), .C(n4290) );
  BUFFD0 U4172 ( .I(n4290), .Z(n4291) );
  CKBD0 U4173 ( .CLK(n4291), .C(n4292) );
  CKBD0 U4174 ( .CLK(n4292), .C(n4293) );
  CKBD0 U4175 ( .CLK(n4293), .C(n4294) );
  CKBD0 U4176 ( .CLK(n4294), .C(n4295) );
  CKBD0 U4177 ( .CLK(n4295), .C(n4296) );
  CKBD0 U4178 ( .CLK(n4296), .C(n4297) );
  CKBD0 U4179 ( .CLK(n4297), .C(n4298) );
  CKBD0 U4180 ( .CLK(n4298), .C(n4299) );
  CKBD0 U4181 ( .CLK(n4299), .C(n4300) );
  CKBD0 U4182 ( .CLK(n4300), .C(n4301) );
  BUFFD0 U4183 ( .I(n4301), .Z(n4302) );
  CKBD0 U4184 ( .CLK(n4302), .C(n4303) );
  CKBD0 U4185 ( .CLK(n4303), .C(n4304) );
  CKBD0 U4186 ( .CLK(n4304), .C(n4305) );
  CKBD0 U4187 ( .CLK(n4305), .C(n4306) );
  CKBD0 U4188 ( .CLK(n4306), .C(n4307) );
  CKBD0 U4189 ( .CLK(n4307), .C(n4308) );
  BUFFD0 U4190 ( .I(n4308), .Z(n4309) );
  CKBD0 U4191 ( .CLK(n4309), .C(n4310) );
  BUFFD0 U4192 ( .I(n4310), .Z(n4311) );
  CKBD0 U4193 ( .CLK(n4311), .C(n4312) );
  BUFFD0 U4194 ( .I(n4312), .Z(n4313) );
  CKBD0 U4195 ( .CLK(n4313), .C(n4314) );
  BUFFD0 U4196 ( .I(n4314), .Z(n4315) );
  CKBD0 U4197 ( .CLK(n4315), .C(n4316) );
  BUFFD0 U4198 ( .I(n4316), .Z(n4317) );
  CKBD0 U4199 ( .CLK(n4317), .C(n4318) );
  BUFFD0 U4200 ( .I(n4318), .Z(n4319) );
  CKBD0 U4201 ( .CLK(n4319), .C(n4320) );
  BUFFD0 U4202 ( .I(n4320), .Z(n4321) );
  CKBD0 U4203 ( .CLK(n4321), .C(n4322) );
  BUFFD0 U4204 ( .I(n4322), .Z(n4323) );
  BUFFD0 U4205 ( .I(n4325), .Z(n4324) );
  BUFFD0 U4206 ( .I(n4326), .Z(n4325) );
  BUFFD0 U4207 ( .I(n9171), .Z(n4326) );
  CKBD0 U4208 ( .CLK(n1246), .C(n4327) );
  CKBD0 U4209 ( .CLK(n4327), .C(n4328) );
  CKBD0 U4210 ( .CLK(n4328), .C(n4329) );
  BUFFD0 U4211 ( .I(n4329), .Z(n4330) );
  CKBD0 U4212 ( .CLK(n4330), .C(n4331) );
  CKBD0 U4213 ( .CLK(n4331), .C(n4332) );
  CKBD0 U4214 ( .CLK(n4332), .C(n4333) );
  CKBD0 U4215 ( .CLK(n4333), .C(n4334) );
  CKBD0 U4216 ( .CLK(n4334), .C(n4335) );
  CKBD0 U4217 ( .CLK(n4335), .C(n4336) );
  CKBD0 U4218 ( .CLK(n4336), .C(n4337) );
  CKBD0 U4219 ( .CLK(n4337), .C(n4338) );
  CKBD0 U4220 ( .CLK(n4338), .C(n4339) );
  BUFFD0 U4221 ( .I(n4339), .Z(n4340) );
  CKBD0 U4222 ( .CLK(n4340), .C(n4341) );
  CKBD0 U4223 ( .CLK(n4341), .C(n4342) );
  CKBD0 U4224 ( .CLK(n4342), .C(n4343) );
  CKBD0 U4225 ( .CLK(n4343), .C(n4344) );
  CKBD0 U4226 ( .CLK(n4344), .C(n4345) );
  CKBD0 U4227 ( .CLK(n4345), .C(n4346) );
  CKBD0 U4228 ( .CLK(n4346), .C(n4347) );
  CKBD0 U4229 ( .CLK(n4347), .C(n4348) );
  CKBD0 U4230 ( .CLK(n4348), .C(n4349) );
  CKBD0 U4231 ( .CLK(n4349), .C(n4350) );
  BUFFD0 U4232 ( .I(n4350), .Z(n4351) );
  CKBD0 U4233 ( .CLK(n4351), .C(n4352) );
  CKBD0 U4234 ( .CLK(n4352), .C(n4353) );
  CKBD0 U4235 ( .CLK(n4353), .C(n4354) );
  CKBD0 U4236 ( .CLK(n4354), .C(n4355) );
  CKBD0 U4237 ( .CLK(n4355), .C(n4356) );
  CKBD0 U4238 ( .CLK(n4356), .C(n4357) );
  CKBD0 U4239 ( .CLK(n4357), .C(n4358) );
  CKBD0 U4240 ( .CLK(n4358), .C(n4359) );
  CKBD0 U4241 ( .CLK(n4359), .C(n4360) );
  CKBD0 U4242 ( .CLK(n4360), .C(n4361) );
  BUFFD0 U4243 ( .I(n4361), .Z(n4362) );
  CKBD0 U4244 ( .CLK(n4362), .C(n4363) );
  CKBD0 U4245 ( .CLK(n4363), .C(n4364) );
  CKBD0 U4246 ( .CLK(n4364), .C(n4365) );
  CKBD0 U4247 ( .CLK(n4365), .C(n4366) );
  CKBD0 U4248 ( .CLK(n4366), .C(n4367) );
  CKBD0 U4249 ( .CLK(n4367), .C(n4368) );
  CKBD0 U4250 ( .CLK(n4368), .C(n4369) );
  CKBD0 U4251 ( .CLK(n4369), .C(n4370) );
  CKBD0 U4252 ( .CLK(n4370), .C(n4371) );
  CKBD0 U4253 ( .CLK(n4371), .C(n4372) );
  BUFFD0 U4254 ( .I(n4372), .Z(n4373) );
  CKBD0 U4255 ( .CLK(n4373), .C(n4374) );
  CKBD0 U4256 ( .CLK(n4374), .C(n4375) );
  CKBD0 U4257 ( .CLK(n4375), .C(n4376) );
  CKBD0 U4258 ( .CLK(n4376), .C(n4377) );
  CKBD0 U4259 ( .CLK(n4377), .C(n4378) );
  CKBD0 U4260 ( .CLK(n4378), .C(n4379) );
  CKBD0 U4261 ( .CLK(n4379), .C(n4380) );
  CKBD0 U4262 ( .CLK(n4380), .C(n4381) );
  CKBD0 U4263 ( .CLK(n4381), .C(n4382) );
  CKBD0 U4264 ( .CLK(n4382), .C(n4383) );
  BUFFD0 U4265 ( .I(n4383), .Z(n4384) );
  CKBD0 U4266 ( .CLK(n4384), .C(n4385) );
  CKBD0 U4267 ( .CLK(n4385), .C(n4386) );
  CKBD0 U4268 ( .CLK(n4386), .C(n4387) );
  CKBD0 U4269 ( .CLK(n4387), .C(n4388) );
  CKBD0 U4270 ( .CLK(n4388), .C(n4389) );
  CKBD0 U4271 ( .CLK(n4389), .C(n4390) );
  CKBD0 U4272 ( .CLK(n4390), .C(n4391) );
  CKBD0 U4273 ( .CLK(n4391), .C(n4392) );
  CKBD0 U4274 ( .CLK(n4392), .C(n4393) );
  CKBD0 U4275 ( .CLK(n4393), .C(n4394) );
  BUFFD0 U4276 ( .I(n4394), .Z(n4395) );
  CKBD0 U4277 ( .CLK(n4395), .C(n4396) );
  CKBD0 U4278 ( .CLK(n4396), .C(n4397) );
  CKBD0 U4279 ( .CLK(n4397), .C(n4398) );
  CKBD0 U4280 ( .CLK(n4398), .C(n4399) );
  CKBD0 U4281 ( .CLK(n4399), .C(n4400) );
  CKBD0 U4282 ( .CLK(n4400), .C(n4401) );
  CKBD0 U4283 ( .CLK(n4401), .C(n4402) );
  CKBD0 U4284 ( .CLK(n4402), .C(n4403) );
  CKBD0 U4285 ( .CLK(n4403), .C(n4404) );
  CKBD0 U4286 ( .CLK(n4404), .C(n4405) );
  BUFFD0 U4287 ( .I(n4405), .Z(n4406) );
  CKBD0 U4288 ( .CLK(n4406), .C(n4407) );
  CKBD0 U4289 ( .CLK(n4407), .C(n4408) );
  CKBD0 U4290 ( .CLK(n4408), .C(n4409) );
  CKBD0 U4291 ( .CLK(n4409), .C(n4410) );
  CKBD0 U4292 ( .CLK(n4410), .C(n4411) );
  CKBD0 U4293 ( .CLK(n4411), .C(n4412) );
  CKBD0 U4294 ( .CLK(n4412), .C(n4413) );
  CKBD0 U4295 ( .CLK(n4413), .C(n4414) );
  CKBD0 U4296 ( .CLK(n4414), .C(n4415) );
  BUFFD0 U4297 ( .I(n4415), .Z(n4416) );
  CKBD0 U4298 ( .CLK(n4416), .C(n4417) );
  CKBD0 U4299 ( .CLK(n4417), .C(n4418) );
  CKBD0 U4300 ( .CLK(n4418), .C(n4419) );
  CKBD0 U4301 ( .CLK(n4419), .C(n4420) );
  CKBD0 U4302 ( .CLK(n4420), .C(n4421) );
  CKBD0 U4303 ( .CLK(n4421), .C(n4422) );
  CKBD0 U4304 ( .CLK(n4422), .C(n4423) );
  CKBD0 U4305 ( .CLK(n4423), .C(n4424) );
  CKBD0 U4306 ( .CLK(n4424), .C(n4425) );
  CKBD0 U4307 ( .CLK(n4425), .C(n4426) );
  BUFFD0 U4308 ( .I(n4426), .Z(n4427) );
  CKBD0 U4309 ( .CLK(n4427), .C(n4428) );
  CKBD0 U4310 ( .CLK(n4428), .C(n4429) );
  CKBD0 U4311 ( .CLK(n4429), .C(n4430) );
  CKBD0 U4312 ( .CLK(n4430), .C(n4431) );
  CKBD0 U4313 ( .CLK(n4431), .C(n4432) );
  CKBD0 U4314 ( .CLK(n4432), .C(n4433) );
  CKBD0 U4315 ( .CLK(n4433), .C(n4434) );
  CKBD0 U4316 ( .CLK(n4434), .C(n4435) );
  CKBD0 U4317 ( .CLK(n4435), .C(n4436) );
  CKBD0 U4318 ( .CLK(n4436), .C(n4437) );
  BUFFD0 U4319 ( .I(n4437), .Z(n4438) );
  CKBD0 U4320 ( .CLK(n4438), .C(n4439) );
  CKBD0 U4321 ( .CLK(n4439), .C(n4440) );
  CKBD0 U4322 ( .CLK(n4440), .C(n4441) );
  CKBD0 U4323 ( .CLK(n4441), .C(n4442) );
  CKBD0 U4324 ( .CLK(n4442), .C(n4443) );
  CKBD0 U4325 ( .CLK(n4443), .C(n4444) );
  BUFFD0 U4326 ( .I(n4444), .Z(n4445) );
  CKBD0 U4327 ( .CLK(n4445), .C(n4446) );
  BUFFD0 U4328 ( .I(n4446), .Z(n4447) );
  CKBD0 U4329 ( .CLK(n4447), .C(n4448) );
  BUFFD0 U4330 ( .I(n4448), .Z(n4449) );
  CKBD0 U4331 ( .CLK(n4449), .C(n4450) );
  BUFFD0 U4332 ( .I(n4450), .Z(n4451) );
  CKBD0 U4333 ( .CLK(n4451), .C(n4452) );
  BUFFD0 U4334 ( .I(n4452), .Z(n4453) );
  CKBD0 U4335 ( .CLK(n4453), .C(n4454) );
  BUFFD0 U4336 ( .I(n4454), .Z(n4455) );
  CKBD0 U4337 ( .CLK(n4455), .C(n4456) );
  BUFFD0 U4338 ( .I(n4456), .Z(n4457) );
  CKBD0 U4339 ( .CLK(n4457), .C(n4458) );
  BUFFD0 U4340 ( .I(n4458), .Z(n4459) );
  BUFFD0 U4341 ( .I(n4461), .Z(n4460) );
  BUFFD0 U4342 ( .I(n4462), .Z(n4461) );
  BUFFD0 U4343 ( .I(n9172), .Z(n4462) );
  CKBD0 U4344 ( .CLK(n1244), .C(n4463) );
  CKBD0 U4345 ( .CLK(n4463), .C(n4464) );
  CKBD0 U4346 ( .CLK(n4464), .C(n4465) );
  BUFFD0 U4347 ( .I(n4465), .Z(n4466) );
  CKBD0 U4348 ( .CLK(n4466), .C(n4467) );
  CKBD0 U4349 ( .CLK(n4467), .C(n4468) );
  CKBD0 U4350 ( .CLK(n4468), .C(n4469) );
  CKBD0 U4351 ( .CLK(n4469), .C(n4470) );
  CKBD0 U4352 ( .CLK(n4470), .C(n4471) );
  CKBD0 U4353 ( .CLK(n4471), .C(n4472) );
  CKBD0 U4354 ( .CLK(n4472), .C(n4473) );
  CKBD0 U4355 ( .CLK(n4473), .C(n4474) );
  CKBD0 U4356 ( .CLK(n4474), .C(n4475) );
  CKBD0 U4357 ( .CLK(n4475), .C(n4476) );
  BUFFD0 U4358 ( .I(n4476), .Z(n4477) );
  CKBD0 U4359 ( .CLK(n4477), .C(n4478) );
  CKBD0 U4360 ( .CLK(n4478), .C(n4479) );
  CKBD0 U4361 ( .CLK(n4479), .C(n4480) );
  CKBD0 U4362 ( .CLK(n4480), .C(n4481) );
  CKBD0 U4363 ( .CLK(n4481), .C(n4482) );
  CKBD0 U4364 ( .CLK(n4482), .C(n4483) );
  CKBD0 U4365 ( .CLK(n4483), .C(n4484) );
  CKBD0 U4366 ( .CLK(n4484), .C(n4485) );
  CKBD0 U4367 ( .CLK(n4485), .C(n4486) );
  BUFFD0 U4368 ( .I(n4486), .Z(n4487) );
  CKBD0 U4369 ( .CLK(n4487), .C(n4488) );
  CKBD0 U4370 ( .CLK(n4488), .C(n4489) );
  CKBD0 U4371 ( .CLK(n4489), .C(n4490) );
  CKBD0 U4372 ( .CLK(n4490), .C(n4491) );
  CKBD0 U4373 ( .CLK(n4491), .C(n4492) );
  CKBD0 U4374 ( .CLK(n4492), .C(n4493) );
  CKBD0 U4375 ( .CLK(n4493), .C(n4494) );
  CKBD0 U4376 ( .CLK(n4494), .C(n4495) );
  CKBD0 U4377 ( .CLK(n4495), .C(n4496) );
  CKBD0 U4378 ( .CLK(n4496), .C(n4497) );
  BUFFD0 U4379 ( .I(n4497), .Z(n4498) );
  CKBD0 U4380 ( .CLK(n4498), .C(n4499) );
  CKBD0 U4381 ( .CLK(n4499), .C(n4500) );
  CKBD0 U4382 ( .CLK(n4500), .C(n4501) );
  CKBD0 U4383 ( .CLK(n4501), .C(n4502) );
  CKBD0 U4384 ( .CLK(n4502), .C(n4503) );
  CKBD0 U4385 ( .CLK(n4503), .C(n4504) );
  CKBD0 U4386 ( .CLK(n4504), .C(n4505) );
  CKBD0 U4387 ( .CLK(n4505), .C(n4506) );
  CKBD0 U4388 ( .CLK(n4506), .C(n4507) );
  CKBD0 U4389 ( .CLK(n4507), .C(n4508) );
  BUFFD0 U4390 ( .I(n4508), .Z(n4509) );
  CKBD0 U4391 ( .CLK(n4509), .C(n4510) );
  CKBD0 U4392 ( .CLK(n4510), .C(n4511) );
  CKBD0 U4393 ( .CLK(n4511), .C(n4512) );
  CKBD0 U4394 ( .CLK(n4512), .C(n4513) );
  CKBD0 U4395 ( .CLK(n4513), .C(n4514) );
  CKBD0 U4396 ( .CLK(n4514), .C(n4515) );
  CKBD0 U4397 ( .CLK(n4515), .C(n4516) );
  CKBD0 U4398 ( .CLK(n4516), .C(n4517) );
  CKBD0 U4399 ( .CLK(n4517), .C(n4518) );
  CKBD0 U4400 ( .CLK(n4518), .C(n4519) );
  BUFFD0 U4401 ( .I(n4519), .Z(n4520) );
  CKBD0 U4402 ( .CLK(n4520), .C(n4521) );
  CKBD0 U4403 ( .CLK(n4521), .C(n4522) );
  CKBD0 U4404 ( .CLK(n4522), .C(n4523) );
  CKBD0 U4405 ( .CLK(n4523), .C(n4524) );
  CKBD0 U4406 ( .CLK(n4524), .C(n4525) );
  CKBD0 U4407 ( .CLK(n4525), .C(n4526) );
  CKBD0 U4408 ( .CLK(n4526), .C(n4527) );
  CKBD0 U4409 ( .CLK(n4527), .C(n4528) );
  CKBD0 U4410 ( .CLK(n4528), .C(n4529) );
  CKBD0 U4411 ( .CLK(n4529), .C(n4530) );
  BUFFD0 U4412 ( .I(n4530), .Z(n4531) );
  CKBD0 U4413 ( .CLK(n4531), .C(n4532) );
  CKBD0 U4414 ( .CLK(n4532), .C(n4533) );
  CKBD0 U4415 ( .CLK(n4533), .C(n4534) );
  CKBD0 U4416 ( .CLK(n4534), .C(n4535) );
  CKBD0 U4417 ( .CLK(n4535), .C(n4536) );
  CKBD0 U4418 ( .CLK(n4536), .C(n4537) );
  CKBD0 U4419 ( .CLK(n4537), .C(n4538) );
  CKBD0 U4420 ( .CLK(n4538), .C(n4539) );
  CKBD0 U4421 ( .CLK(n4539), .C(n4540) );
  CKBD0 U4422 ( .CLK(n4540), .C(n4541) );
  BUFFD0 U4423 ( .I(n4541), .Z(n4542) );
  CKBD0 U4424 ( .CLK(n4542), .C(n4543) );
  CKBD0 U4425 ( .CLK(n4543), .C(n4544) );
  CKBD0 U4426 ( .CLK(n4544), .C(n4545) );
  CKBD0 U4427 ( .CLK(n4545), .C(n4546) );
  CKBD0 U4428 ( .CLK(n4546), .C(n4547) );
  CKBD0 U4429 ( .CLK(n4547), .C(n4548) );
  CKBD0 U4430 ( .CLK(n4548), .C(n4549) );
  CKBD0 U4431 ( .CLK(n4549), .C(n4550) );
  CKBD0 U4432 ( .CLK(n4550), .C(n4551) );
  BUFFD0 U4433 ( .I(n4551), .Z(n4552) );
  CKBD0 U4434 ( .CLK(n4552), .C(n4553) );
  CKBD0 U4435 ( .CLK(n4553), .C(n4554) );
  CKBD0 U4436 ( .CLK(n4554), .C(n4555) );
  CKBD0 U4437 ( .CLK(n4555), .C(n4556) );
  CKBD0 U4438 ( .CLK(n4556), .C(n4557) );
  CKBD0 U4439 ( .CLK(n4557), .C(n4558) );
  CKBD0 U4440 ( .CLK(n4558), .C(n4559) );
  CKBD0 U4441 ( .CLK(n4559), .C(n4560) );
  CKBD0 U4442 ( .CLK(n4560), .C(n4561) );
  CKBD0 U4443 ( .CLK(n4561), .C(n4562) );
  BUFFD0 U4444 ( .I(n4562), .Z(n4563) );
  CKBD0 U4445 ( .CLK(n4563), .C(n4564) );
  CKBD0 U4446 ( .CLK(n4564), .C(n4565) );
  CKBD0 U4447 ( .CLK(n4565), .C(n4566) );
  CKBD0 U4448 ( .CLK(n4566), .C(n4567) );
  CKBD0 U4449 ( .CLK(n4567), .C(n4568) );
  CKBD0 U4450 ( .CLK(n4568), .C(n4569) );
  CKBD0 U4451 ( .CLK(n4569), .C(n4570) );
  CKBD0 U4452 ( .CLK(n4570), .C(n4571) );
  CKBD0 U4453 ( .CLK(n4571), .C(n4572) );
  CKBD0 U4454 ( .CLK(n4572), .C(n4573) );
  BUFFD0 U4455 ( .I(n4573), .Z(n4574) );
  CKBD0 U4456 ( .CLK(n4574), .C(n4575) );
  CKBD0 U4457 ( .CLK(n4575), .C(n4576) );
  CKBD0 U4458 ( .CLK(n4576), .C(n4577) );
  CKBD0 U4459 ( .CLK(n4577), .C(n4578) );
  CKBD0 U4460 ( .CLK(n4578), .C(n4579) );
  CKBD0 U4461 ( .CLK(n4579), .C(n4580) );
  BUFFD0 U4462 ( .I(n4580), .Z(n4581) );
  CKBD0 U4463 ( .CLK(n4581), .C(n4582) );
  BUFFD0 U4464 ( .I(n4582), .Z(n4583) );
  CKBD0 U4465 ( .CLK(n4583), .C(n4584) );
  BUFFD0 U4466 ( .I(n4584), .Z(n4585) );
  CKBD0 U4467 ( .CLK(n4585), .C(n4586) );
  BUFFD0 U4468 ( .I(n4586), .Z(n4587) );
  CKBD0 U4469 ( .CLK(n4587), .C(n4588) );
  BUFFD0 U4470 ( .I(n4588), .Z(n4589) );
  CKBD0 U4471 ( .CLK(n4589), .C(n4590) );
  BUFFD0 U4472 ( .I(n4590), .Z(n4591) );
  CKBD0 U4473 ( .CLK(n4591), .C(n4592) );
  BUFFD0 U4474 ( .I(n4592), .Z(n4593) );
  CKBD0 U4475 ( .CLK(n4593), .C(n4594) );
  BUFFD0 U4476 ( .I(n4594), .Z(n4595) );
  BUFFD0 U4477 ( .I(n4597), .Z(n4596) );
  BUFFD0 U4478 ( .I(n4598), .Z(n4597) );
  BUFFD0 U4479 ( .I(n9173), .Z(n4598) );
  CKBD0 U4480 ( .CLK(n1242), .C(n4599) );
  CKBD0 U4481 ( .CLK(n4599), .C(n4600) );
  CKBD0 U4482 ( .CLK(n4600), .C(n4601) );
  BUFFD0 U4483 ( .I(n4601), .Z(n4602) );
  CKBD0 U4484 ( .CLK(n4602), .C(n4603) );
  CKBD0 U4485 ( .CLK(n4603), .C(n4604) );
  CKBD0 U4486 ( .CLK(n4604), .C(n4605) );
  CKBD0 U4487 ( .CLK(n4605), .C(n4606) );
  CKBD0 U4488 ( .CLK(n4606), .C(n4607) );
  CKBD0 U4489 ( .CLK(n4607), .C(n4608) );
  CKBD0 U4490 ( .CLK(n4608), .C(n4609) );
  CKBD0 U4491 ( .CLK(n4609), .C(n4610) );
  CKBD0 U4492 ( .CLK(n4610), .C(n4611) );
  CKBD0 U4493 ( .CLK(n4611), .C(n4612) );
  BUFFD0 U4494 ( .I(n4612), .Z(n4613) );
  CKBD0 U4495 ( .CLK(n4613), .C(n4614) );
  CKBD0 U4496 ( .CLK(n4614), .C(n4615) );
  CKBD0 U4497 ( .CLK(n4615), .C(n4616) );
  CKBD0 U4498 ( .CLK(n4616), .C(n4617) );
  CKBD0 U4499 ( .CLK(n4617), .C(n4618) );
  CKBD0 U4500 ( .CLK(n4618), .C(n4619) );
  CKBD0 U4501 ( .CLK(n4619), .C(n4620) );
  CKBD0 U4502 ( .CLK(n4620), .C(n4621) );
  CKBD0 U4503 ( .CLK(n4621), .C(n4622) );
  BUFFD0 U4504 ( .I(n4622), .Z(n4623) );
  CKBD0 U4505 ( .CLK(n4623), .C(n4624) );
  CKBD0 U4506 ( .CLK(n4624), .C(n4625) );
  CKBD0 U4507 ( .CLK(n4625), .C(n4626) );
  CKBD0 U4508 ( .CLK(n4626), .C(n4627) );
  CKBD0 U4509 ( .CLK(n4627), .C(n4628) );
  CKBD0 U4510 ( .CLK(n4628), .C(n4629) );
  CKBD0 U4511 ( .CLK(n4629), .C(n4630) );
  CKBD0 U4512 ( .CLK(n4630), .C(n4631) );
  CKBD0 U4513 ( .CLK(n4631), .C(n4632) );
  CKBD0 U4514 ( .CLK(n4632), .C(n4633) );
  BUFFD0 U4515 ( .I(n4633), .Z(n4634) );
  CKBD0 U4516 ( .CLK(n4634), .C(n4635) );
  CKBD0 U4517 ( .CLK(n4635), .C(n4636) );
  CKBD0 U4518 ( .CLK(n4636), .C(n4637) );
  CKBD0 U4519 ( .CLK(n4637), .C(n4638) );
  CKBD0 U4520 ( .CLK(n4638), .C(n4639) );
  CKBD0 U4521 ( .CLK(n4639), .C(n4640) );
  CKBD0 U4522 ( .CLK(n4640), .C(n4641) );
  CKBD0 U4523 ( .CLK(n4641), .C(n4642) );
  CKBD0 U4524 ( .CLK(n4642), .C(n4643) );
  CKBD0 U4525 ( .CLK(n4643), .C(n4644) );
  BUFFD0 U4526 ( .I(n4644), .Z(n4645) );
  CKBD0 U4527 ( .CLK(n4645), .C(n4646) );
  CKBD0 U4528 ( .CLK(n4646), .C(n4647) );
  CKBD0 U4529 ( .CLK(n4647), .C(n4648) );
  CKBD0 U4530 ( .CLK(n4648), .C(n4649) );
  CKBD0 U4531 ( .CLK(n4649), .C(n4650) );
  CKBD0 U4532 ( .CLK(n4650), .C(n4651) );
  CKBD0 U4533 ( .CLK(n4651), .C(n4652) );
  CKBD0 U4534 ( .CLK(n4652), .C(n4653) );
  CKBD0 U4535 ( .CLK(n4653), .C(n4654) );
  CKBD0 U4536 ( .CLK(n4654), .C(n4655) );
  BUFFD0 U4537 ( .I(n4655), .Z(n4656) );
  CKBD0 U4538 ( .CLK(n4656), .C(n4657) );
  CKBD0 U4539 ( .CLK(n4657), .C(n4658) );
  CKBD0 U4540 ( .CLK(n4658), .C(n4659) );
  CKBD0 U4541 ( .CLK(n4659), .C(n4660) );
  CKBD0 U4542 ( .CLK(n4660), .C(n4661) );
  CKBD0 U4543 ( .CLK(n4661), .C(n4662) );
  CKBD0 U4544 ( .CLK(n4662), .C(n4663) );
  CKBD0 U4545 ( .CLK(n4663), .C(n4664) );
  CKBD0 U4546 ( .CLK(n4664), .C(n4665) );
  CKBD0 U4547 ( .CLK(n4665), .C(n4666) );
  BUFFD0 U4548 ( .I(n4666), .Z(n4667) );
  CKBD0 U4549 ( .CLK(n4667), .C(n4668) );
  CKBD0 U4550 ( .CLK(n4668), .C(n4669) );
  CKBD0 U4551 ( .CLK(n4669), .C(n4670) );
  CKBD0 U4552 ( .CLK(n4670), .C(n4671) );
  CKBD0 U4553 ( .CLK(n4671), .C(n4672) );
  CKBD0 U4554 ( .CLK(n4672), .C(n4673) );
  CKBD0 U4555 ( .CLK(n4673), .C(n4674) );
  CKBD0 U4556 ( .CLK(n4674), .C(n4675) );
  CKBD0 U4557 ( .CLK(n4675), .C(n4676) );
  CKBD0 U4558 ( .CLK(n4676), .C(n4677) );
  BUFFD0 U4559 ( .I(n4677), .Z(n4678) );
  CKBD0 U4560 ( .CLK(n4678), .C(n4679) );
  CKBD0 U4561 ( .CLK(n4679), .C(n4680) );
  CKBD0 U4562 ( .CLK(n4680), .C(n4681) );
  CKBD0 U4563 ( .CLK(n4681), .C(n4682) );
  CKBD0 U4564 ( .CLK(n4682), .C(n4683) );
  CKBD0 U4565 ( .CLK(n4683), .C(n4684) );
  CKBD0 U4566 ( .CLK(n4684), .C(n4685) );
  CKBD0 U4567 ( .CLK(n4685), .C(n4686) );
  CKBD0 U4568 ( .CLK(n4686), .C(n4687) );
  CKBD0 U4569 ( .CLK(n4687), .C(n4688) );
  BUFFD0 U4570 ( .I(n4688), .Z(n4689) );
  CKBD0 U4571 ( .CLK(n4689), .C(n4690) );
  CKBD0 U4572 ( .CLK(n4690), .C(n4691) );
  CKBD0 U4573 ( .CLK(n4691), .C(n4692) );
  CKBD0 U4574 ( .CLK(n4692), .C(n4693) );
  CKBD0 U4575 ( .CLK(n4693), .C(n4694) );
  CKBD0 U4576 ( .CLK(n4694), .C(n4695) );
  CKBD0 U4577 ( .CLK(n4695), .C(n4696) );
  CKBD0 U4578 ( .CLK(n4696), .C(n4697) );
  CKBD0 U4579 ( .CLK(n4697), .C(n4698) );
  BUFFD0 U4580 ( .I(n4698), .Z(n4699) );
  CKBD0 U4581 ( .CLK(n4699), .C(n4700) );
  CKBD0 U4582 ( .CLK(n4700), .C(n4701) );
  CKBD0 U4583 ( .CLK(n4701), .C(n4702) );
  CKBD0 U4584 ( .CLK(n4702), .C(n4703) );
  CKBD0 U4585 ( .CLK(n4703), .C(n4704) );
  CKBD0 U4586 ( .CLK(n4704), .C(n4705) );
  CKBD0 U4587 ( .CLK(n4705), .C(n4706) );
  CKBD0 U4588 ( .CLK(n4706), .C(n4707) );
  CKBD0 U4589 ( .CLK(n4707), .C(n4708) );
  CKBD0 U4590 ( .CLK(n4708), .C(n4709) );
  BUFFD0 U4591 ( .I(n4709), .Z(n4710) );
  CKBD0 U4592 ( .CLK(n4710), .C(n4711) );
  CKBD0 U4593 ( .CLK(n4711), .C(n4712) );
  CKBD0 U4594 ( .CLK(n4712), .C(n4713) );
  CKBD0 U4595 ( .CLK(n4713), .C(n4714) );
  CKBD0 U4596 ( .CLK(n4714), .C(n4715) );
  CKBD0 U4597 ( .CLK(n4715), .C(n4716) );
  BUFFD0 U4598 ( .I(n4716), .Z(n4717) );
  CKBD0 U4599 ( .CLK(n4717), .C(n4718) );
  BUFFD0 U4600 ( .I(n4718), .Z(n4719) );
  CKBD0 U4601 ( .CLK(n4719), .C(n4720) );
  BUFFD0 U4602 ( .I(n4720), .Z(n4721) );
  CKBD0 U4603 ( .CLK(n4721), .C(n4722) );
  BUFFD0 U4604 ( .I(n4722), .Z(n4723) );
  CKBD0 U4605 ( .CLK(n4723), .C(n4724) );
  BUFFD0 U4606 ( .I(n4724), .Z(n4725) );
  CKBD0 U4607 ( .CLK(n4725), .C(n4726) );
  BUFFD0 U4608 ( .I(n4726), .Z(n4727) );
  CKBD0 U4609 ( .CLK(n4727), .C(n4728) );
  BUFFD0 U4610 ( .I(n4728), .Z(n4729) );
  CKBD0 U4611 ( .CLK(n4729), .C(n4730) );
  BUFFD0 U4612 ( .I(n4730), .Z(n4731) );
  BUFFD0 U4613 ( .I(n4733), .Z(n4732) );
  BUFFD0 U4614 ( .I(n4734), .Z(n4733) );
  BUFFD0 U4615 ( .I(n9174), .Z(n4734) );
  CKBD0 U4616 ( .CLK(n720), .C(n4735) );
  CKBD0 U4617 ( .CLK(n4735), .C(n4736) );
  CKBD0 U4618 ( .CLK(n4736), .C(n4737) );
  BUFFD0 U4619 ( .I(n4737), .Z(n4738) );
  CKBD0 U4620 ( .CLK(n4738), .C(n4739) );
  CKBD0 U4621 ( .CLK(n4739), .C(n4740) );
  CKBD0 U4622 ( .CLK(n4740), .C(n4741) );
  CKBD0 U4623 ( .CLK(n4741), .C(n4742) );
  CKBD0 U4624 ( .CLK(n4742), .C(n4743) );
  CKBD0 U4625 ( .CLK(n4743), .C(n4744) );
  CKBD0 U4626 ( .CLK(n4744), .C(n4745) );
  CKBD0 U4627 ( .CLK(n4745), .C(n4746) );
  CKBD0 U4628 ( .CLK(n4746), .C(n4747) );
  CKBD0 U4629 ( .CLK(n4747), .C(n4748) );
  BUFFD0 U4630 ( .I(n4748), .Z(n4749) );
  CKBD0 U4631 ( .CLK(n4749), .C(n4750) );
  CKBD0 U4632 ( .CLK(n4750), .C(n4751) );
  CKBD0 U4633 ( .CLK(n4751), .C(n4752) );
  CKBD0 U4634 ( .CLK(n4752), .C(n4753) );
  CKBD0 U4635 ( .CLK(n4753), .C(n4754) );
  CKBD0 U4636 ( .CLK(n4754), .C(n4755) );
  CKBD0 U4637 ( .CLK(n4755), .C(n4756) );
  CKBD0 U4638 ( .CLK(n4756), .C(n4757) );
  CKBD0 U4639 ( .CLK(n4757), .C(n4758) );
  BUFFD0 U4640 ( .I(n4758), .Z(n4759) );
  CKBD0 U4641 ( .CLK(n4759), .C(n4760) );
  CKBD0 U4642 ( .CLK(n4760), .C(n4761) );
  CKBD0 U4643 ( .CLK(n4761), .C(n4762) );
  CKBD0 U4644 ( .CLK(n4762), .C(n4763) );
  CKBD0 U4645 ( .CLK(n4763), .C(n4764) );
  CKBD0 U4646 ( .CLK(n4764), .C(n4765) );
  CKBD0 U4647 ( .CLK(n4765), .C(n4766) );
  CKBD0 U4648 ( .CLK(n4766), .C(n4767) );
  CKBD0 U4649 ( .CLK(n4767), .C(n4768) );
  CKBD0 U4650 ( .CLK(n4768), .C(n4769) );
  BUFFD0 U4651 ( .I(n4769), .Z(n4770) );
  CKBD0 U4652 ( .CLK(n4770), .C(n4771) );
  CKBD0 U4653 ( .CLK(n4771), .C(n4772) );
  CKBD0 U4654 ( .CLK(n4772), .C(n4773) );
  CKBD0 U4655 ( .CLK(n4773), .C(n4774) );
  CKBD0 U4656 ( .CLK(n4774), .C(n4775) );
  CKBD0 U4657 ( .CLK(n4775), .C(n4776) );
  CKBD0 U4658 ( .CLK(n4776), .C(n4777) );
  CKBD0 U4659 ( .CLK(n4777), .C(n4778) );
  CKBD0 U4660 ( .CLK(n4778), .C(n4779) );
  CKBD0 U4661 ( .CLK(n4779), .C(n4780) );
  BUFFD0 U4662 ( .I(n4780), .Z(n4781) );
  CKBD0 U4663 ( .CLK(n4781), .C(n4782) );
  CKBD0 U4664 ( .CLK(n4782), .C(n4783) );
  CKBD0 U4665 ( .CLK(n4783), .C(n4784) );
  CKBD0 U4666 ( .CLK(n4784), .C(n4785) );
  CKBD0 U4667 ( .CLK(n4785), .C(n4786) );
  CKBD0 U4668 ( .CLK(n4786), .C(n4787) );
  CKBD0 U4669 ( .CLK(n4787), .C(n4788) );
  CKBD0 U4670 ( .CLK(n4788), .C(n4789) );
  CKBD0 U4671 ( .CLK(n4789), .C(n4790) );
  CKBD0 U4672 ( .CLK(n4790), .C(n4791) );
  BUFFD0 U4673 ( .I(n4791), .Z(n4792) );
  CKBD0 U4674 ( .CLK(n4792), .C(n4793) );
  CKBD0 U4675 ( .CLK(n4793), .C(n4794) );
  CKBD0 U4676 ( .CLK(n4794), .C(n4795) );
  CKBD0 U4677 ( .CLK(n4795), .C(n4796) );
  CKBD0 U4678 ( .CLK(n4796), .C(n4797) );
  CKBD0 U4679 ( .CLK(n4797), .C(n4798) );
  CKBD0 U4680 ( .CLK(n4798), .C(n4799) );
  CKBD0 U4681 ( .CLK(n4799), .C(n4800) );
  CKBD0 U4682 ( .CLK(n4800), .C(n4801) );
  CKBD0 U4683 ( .CLK(n4801), .C(n4802) );
  BUFFD0 U4684 ( .I(n4802), .Z(n4803) );
  CKBD0 U4685 ( .CLK(n4803), .C(n4804) );
  CKBD0 U4686 ( .CLK(n4804), .C(n4805) );
  CKBD0 U4687 ( .CLK(n4805), .C(n4806) );
  CKBD0 U4688 ( .CLK(n4806), .C(n4807) );
  CKBD0 U4689 ( .CLK(n4807), .C(n4808) );
  CKBD0 U4690 ( .CLK(n4808), .C(n4809) );
  CKBD0 U4691 ( .CLK(n4809), .C(n4810) );
  CKBD0 U4692 ( .CLK(n4810), .C(n4811) );
  CKBD0 U4693 ( .CLK(n4811), .C(n4812) );
  CKBD0 U4694 ( .CLK(n4812), .C(n4813) );
  BUFFD0 U4695 ( .I(n4813), .Z(n4814) );
  CKBD0 U4696 ( .CLK(n4814), .C(n4815) );
  CKBD0 U4697 ( .CLK(n4815), .C(n4816) );
  CKBD0 U4698 ( .CLK(n4816), .C(n4817) );
  CKBD0 U4699 ( .CLK(n4817), .C(n4818) );
  CKBD0 U4700 ( .CLK(n4818), .C(n4819) );
  CKBD0 U4701 ( .CLK(n4819), .C(n4820) );
  CKBD0 U4702 ( .CLK(n4820), .C(n4821) );
  CKBD0 U4703 ( .CLK(n4821), .C(n4822) );
  CKBD0 U4704 ( .CLK(n4822), .C(n4823) );
  CKBD0 U4705 ( .CLK(n4823), .C(n4824) );
  BUFFD0 U4706 ( .I(n4824), .Z(n4825) );
  CKBD0 U4707 ( .CLK(n4825), .C(n4826) );
  CKBD0 U4708 ( .CLK(n4826), .C(n4827) );
  CKBD0 U4709 ( .CLK(n4827), .C(n4828) );
  CKBD0 U4710 ( .CLK(n4828), .C(n4829) );
  CKBD0 U4711 ( .CLK(n4829), .C(n4830) );
  CKBD0 U4712 ( .CLK(n4830), .C(n4831) );
  CKBD0 U4713 ( .CLK(n4831), .C(n4832) );
  CKBD0 U4714 ( .CLK(n4832), .C(n4833) );
  CKBD0 U4715 ( .CLK(n4833), .C(n4834) );
  BUFFD0 U4716 ( .I(n4834), .Z(n4835) );
  CKBD0 U4717 ( .CLK(n4835), .C(n4836) );
  CKBD0 U4718 ( .CLK(n4836), .C(n4837) );
  CKBD0 U4719 ( .CLK(n4837), .C(n4838) );
  CKBD0 U4720 ( .CLK(n4838), .C(n4839) );
  CKBD0 U4721 ( .CLK(n4839), .C(n4840) );
  CKBD0 U4722 ( .CLK(n4840), .C(n4841) );
  CKBD0 U4723 ( .CLK(n4841), .C(n4842) );
  CKBD0 U4724 ( .CLK(n4842), .C(n4843) );
  CKBD0 U4725 ( .CLK(n4843), .C(n4844) );
  CKBD0 U4726 ( .CLK(n4844), .C(n4845) );
  BUFFD0 U4727 ( .I(n4845), .Z(n4846) );
  CKBD0 U4728 ( .CLK(n4846), .C(n4847) );
  CKBD0 U4729 ( .CLK(n4847), .C(n4848) );
  CKBD0 U4730 ( .CLK(n4848), .C(n4849) );
  CKBD0 U4731 ( .CLK(n4849), .C(n4850) );
  CKBD0 U4732 ( .CLK(n4850), .C(n4851) );
  CKBD0 U4733 ( .CLK(n4851), .C(n4852) );
  BUFFD0 U4734 ( .I(n4852), .Z(n4853) );
  CKBD0 U4735 ( .CLK(n4853), .C(n4854) );
  BUFFD0 U4736 ( .I(n4854), .Z(n4855) );
  CKBD0 U4737 ( .CLK(n4855), .C(n4856) );
  BUFFD0 U4738 ( .I(n4856), .Z(n4857) );
  CKBD0 U4739 ( .CLK(n4857), .C(n4858) );
  BUFFD0 U4740 ( .I(n4858), .Z(n4859) );
  CKBD0 U4741 ( .CLK(n4859), .C(n4860) );
  BUFFD0 U4742 ( .I(n4860), .Z(n4861) );
  CKBD0 U4743 ( .CLK(n4861), .C(n4862) );
  BUFFD0 U4744 ( .I(n4862), .Z(n4863) );
  CKBD0 U4745 ( .CLK(n4863), .C(n4864) );
  BUFFD0 U4746 ( .I(n4864), .Z(n4865) );
  CKBD0 U4747 ( .CLK(n4865), .C(n4866) );
  BUFFD0 U4748 ( .I(n4866), .Z(n4867) );
  BUFFD0 U4749 ( .I(n4869), .Z(n4868) );
  BUFFD0 U4750 ( .I(n4870), .Z(n4869) );
  BUFFD0 U4751 ( .I(n9175), .Z(n4870) );
  CKBD0 U4752 ( .CLK(n1142), .C(n4871) );
  CKBD0 U4753 ( .CLK(n4871), .C(n4872) );
  CKBD0 U4754 ( .CLK(n4872), .C(n4873) );
  BUFFD0 U4755 ( .I(n4873), .Z(n4874) );
  CKBD0 U4756 ( .CLK(n4874), .C(n4875) );
  CKBD0 U4757 ( .CLK(n4875), .C(n4876) );
  CKBD0 U4758 ( .CLK(n4876), .C(n4877) );
  CKBD0 U4759 ( .CLK(n4877), .C(n4878) );
  CKBD0 U4760 ( .CLK(n4878), .C(n4879) );
  CKBD0 U4761 ( .CLK(n4879), .C(n4880) );
  CKBD0 U4762 ( .CLK(n4880), .C(n4881) );
  CKBD0 U4763 ( .CLK(n4881), .C(n4882) );
  CKBD0 U4764 ( .CLK(n4882), .C(n4883) );
  BUFFD0 U4765 ( .I(n4883), .Z(n4884) );
  CKBD0 U4766 ( .CLK(n4884), .C(n4885) );
  CKBD0 U4767 ( .CLK(n4885), .C(n4886) );
  CKBD0 U4768 ( .CLK(n4886), .C(n4887) );
  CKBD0 U4769 ( .CLK(n4887), .C(n4888) );
  CKBD0 U4770 ( .CLK(n4888), .C(n4889) );
  CKBD0 U4771 ( .CLK(n4889), .C(n4890) );
  CKBD0 U4772 ( .CLK(n4890), .C(n4891) );
  CKBD0 U4773 ( .CLK(n4891), .C(n4892) );
  CKBD0 U4774 ( .CLK(n4892), .C(n4893) );
  CKBD0 U4775 ( .CLK(n4893), .C(n4894) );
  BUFFD0 U4776 ( .I(n4894), .Z(n4895) );
  CKBD0 U4777 ( .CLK(n4895), .C(n4896) );
  CKBD0 U4778 ( .CLK(n4896), .C(n4897) );
  CKBD0 U4779 ( .CLK(n4897), .C(n4898) );
  CKBD0 U4780 ( .CLK(n4898), .C(n4899) );
  CKBD0 U4781 ( .CLK(n4899), .C(n4900) );
  CKBD0 U4782 ( .CLK(n4900), .C(n4901) );
  CKBD0 U4783 ( .CLK(n4901), .C(n4902) );
  CKBD0 U4784 ( .CLK(n4902), .C(n4903) );
  CKBD0 U4785 ( .CLK(n4903), .C(n4904) );
  CKBD0 U4786 ( .CLK(n4904), .C(n4905) );
  BUFFD0 U4787 ( .I(n4905), .Z(n4906) );
  CKBD0 U4788 ( .CLK(n4906), .C(n4907) );
  CKBD0 U4789 ( .CLK(n4907), .C(n4908) );
  CKBD0 U4790 ( .CLK(n4908), .C(n4909) );
  CKBD0 U4791 ( .CLK(n4909), .C(n4910) );
  CKBD0 U4792 ( .CLK(n4910), .C(n4911) );
  CKBD0 U4793 ( .CLK(n4911), .C(n4912) );
  CKBD0 U4794 ( .CLK(n4912), .C(n4913) );
  CKBD0 U4795 ( .CLK(n4913), .C(n4914) );
  CKBD0 U4796 ( .CLK(n4914), .C(n4915) );
  CKBD0 U4797 ( .CLK(n4915), .C(n4916) );
  BUFFD0 U4798 ( .I(n4916), .Z(n4917) );
  CKBD0 U4799 ( .CLK(n4917), .C(n4918) );
  CKBD0 U4800 ( .CLK(n4918), .C(n4919) );
  CKBD0 U4801 ( .CLK(n4919), .C(n4920) );
  CKBD0 U4802 ( .CLK(n4920), .C(n4921) );
  CKBD0 U4803 ( .CLK(n4921), .C(n4922) );
  CKBD0 U4804 ( .CLK(n4922), .C(n4923) );
  CKBD0 U4805 ( .CLK(n4923), .C(n4924) );
  CKBD0 U4806 ( .CLK(n4924), .C(n4925) );
  CKBD0 U4807 ( .CLK(n4925), .C(n4926) );
  CKBD0 U4808 ( .CLK(n4926), .C(n4927) );
  BUFFD0 U4809 ( .I(n4927), .Z(n4928) );
  CKBD0 U4810 ( .CLK(n4928), .C(n4929) );
  CKBD0 U4811 ( .CLK(n4929), .C(n4930) );
  CKBD0 U4812 ( .CLK(n4930), .C(n4931) );
  CKBD0 U4813 ( .CLK(n4931), .C(n4932) );
  CKBD0 U4814 ( .CLK(n4932), .C(n4933) );
  CKBD0 U4815 ( .CLK(n4933), .C(n4934) );
  CKBD0 U4816 ( .CLK(n4934), .C(n4935) );
  CKBD0 U4817 ( .CLK(n4935), .C(n4936) );
  CKBD0 U4818 ( .CLK(n4936), .C(n4937) );
  CKBD0 U4819 ( .CLK(n4937), .C(n4938) );
  BUFFD0 U4820 ( .I(n4938), .Z(n4939) );
  CKBD0 U4821 ( .CLK(n4939), .C(n4940) );
  CKBD0 U4822 ( .CLK(n4940), .C(n4941) );
  CKBD0 U4823 ( .CLK(n4941), .C(n4942) );
  CKBD0 U4824 ( .CLK(n4942), .C(n4943) );
  CKBD0 U4825 ( .CLK(n4943), .C(n4944) );
  CKBD0 U4826 ( .CLK(n4944), .C(n4945) );
  CKBD0 U4827 ( .CLK(n4945), .C(n4946) );
  CKBD0 U4828 ( .CLK(n4946), .C(n4947) );
  CKBD0 U4829 ( .CLK(n4947), .C(n4948) );
  CKBD0 U4830 ( .CLK(n4948), .C(n4949) );
  BUFFD0 U4831 ( .I(n4949), .Z(n4950) );
  CKBD0 U4832 ( .CLK(n4950), .C(n4951) );
  CKBD0 U4833 ( .CLK(n4951), .C(n4952) );
  CKBD0 U4834 ( .CLK(n4952), .C(n4953) );
  CKBD0 U4835 ( .CLK(n4953), .C(n4954) );
  CKBD0 U4836 ( .CLK(n4954), .C(n4955) );
  CKBD0 U4837 ( .CLK(n4955), .C(n4956) );
  CKBD0 U4838 ( .CLK(n4956), .C(n4957) );
  CKBD0 U4839 ( .CLK(n4957), .C(n4958) );
  CKBD0 U4840 ( .CLK(n4958), .C(n4959) );
  BUFFD0 U4841 ( .I(n4959), .Z(n4960) );
  CKBD0 U4842 ( .CLK(n4960), .C(n4961) );
  CKBD0 U4843 ( .CLK(n4961), .C(n4962) );
  CKBD0 U4844 ( .CLK(n4962), .C(n4963) );
  CKBD0 U4845 ( .CLK(n4963), .C(n4964) );
  CKBD0 U4846 ( .CLK(n4964), .C(n4965) );
  CKBD0 U4847 ( .CLK(n4965), .C(n4966) );
  CKBD0 U4848 ( .CLK(n4966), .C(n4967) );
  CKBD0 U4849 ( .CLK(n4967), .C(n4968) );
  CKBD0 U4850 ( .CLK(n4968), .C(n4969) );
  CKBD0 U4851 ( .CLK(n4969), .C(n4970) );
  BUFFD0 U4852 ( .I(n4970), .Z(n4971) );
  CKBD0 U4853 ( .CLK(n4971), .C(n4972) );
  CKBD0 U4854 ( .CLK(n4972), .C(n4973) );
  CKBD0 U4855 ( .CLK(n4973), .C(n4974) );
  CKBD0 U4856 ( .CLK(n4974), .C(n4975) );
  CKBD0 U4857 ( .CLK(n4975), .C(n4976) );
  CKBD0 U4858 ( .CLK(n4976), .C(n4977) );
  CKBD0 U4859 ( .CLK(n4977), .C(n4978) );
  CKBD0 U4860 ( .CLK(n4978), .C(n4979) );
  CKBD0 U4861 ( .CLK(n4979), .C(n4980) );
  CKBD0 U4862 ( .CLK(n4980), .C(n4981) );
  BUFFD0 U4863 ( .I(n4981), .Z(n4982) );
  CKBD0 U4864 ( .CLK(n4982), .C(n4983) );
  CKBD0 U4865 ( .CLK(n4983), .C(n4984) );
  CKBD0 U4866 ( .CLK(n4984), .C(n4985) );
  CKBD0 U4867 ( .CLK(n4985), .C(n4986) );
  CKBD0 U4868 ( .CLK(n4986), .C(n4987) );
  CKBD0 U4869 ( .CLK(n4987), .C(n4988) );
  BUFFD0 U4870 ( .I(n4988), .Z(n4989) );
  CKBD0 U4871 ( .CLK(n4989), .C(n4990) );
  BUFFD0 U4872 ( .I(n4990), .Z(n4991) );
  CKBD0 U4873 ( .CLK(n4991), .C(n4992) );
  BUFFD0 U4874 ( .I(n4992), .Z(n4993) );
  CKBD0 U4875 ( .CLK(n4993), .C(n4994) );
  BUFFD0 U4876 ( .I(n4994), .Z(n4995) );
  CKBD0 U4877 ( .CLK(n4995), .C(n4996) );
  BUFFD0 U4878 ( .I(n4996), .Z(n4997) );
  CKBD0 U4879 ( .CLK(n4997), .C(n4998) );
  BUFFD0 U4880 ( .I(n4998), .Z(n4999) );
  CKBD0 U4881 ( .CLK(n4999), .C(n5000) );
  BUFFD0 U4882 ( .I(n5000), .Z(n5001) );
  CKBD0 U4883 ( .CLK(n5001), .C(n5002) );
  BUFFD0 U4884 ( .I(n5002), .Z(n5003) );
  BUFFD0 U4885 ( .I(n5005), .Z(n5004) );
  BUFFD0 U4886 ( .I(n5006), .Z(n5005) );
  BUFFD0 U4887 ( .I(n9176), .Z(n5006) );
  CKBD0 U4888 ( .CLK(n1140), .C(n5007) );
  CKBD0 U4889 ( .CLK(n5007), .C(n5008) );
  CKBD0 U4890 ( .CLK(n5008), .C(n5009) );
  BUFFD0 U4891 ( .I(n5009), .Z(n5010) );
  CKBD0 U4892 ( .CLK(n5010), .C(n5011) );
  CKBD0 U4893 ( .CLK(n5011), .C(n5012) );
  CKBD0 U4894 ( .CLK(n5012), .C(n5013) );
  CKBD0 U4895 ( .CLK(n5013), .C(n5014) );
  CKBD0 U4896 ( .CLK(n5014), .C(n5015) );
  CKBD0 U4897 ( .CLK(n5015), .C(n5016) );
  CKBD0 U4898 ( .CLK(n5016), .C(n5017) );
  CKBD0 U4899 ( .CLK(n5017), .C(n5018) );
  CKBD0 U4900 ( .CLK(n5018), .C(n5019) );
  CKBD0 U4901 ( .CLK(n5019), .C(n5020) );
  BUFFD0 U4902 ( .I(n5020), .Z(n5021) );
  CKBD0 U4903 ( .CLK(n5021), .C(n5022) );
  CKBD0 U4904 ( .CLK(n5022), .C(n5023) );
  CKBD0 U4905 ( .CLK(n5023), .C(n5024) );
  CKBD0 U4906 ( .CLK(n5024), .C(n5025) );
  CKBD0 U4907 ( .CLK(n5025), .C(n5026) );
  CKBD0 U4908 ( .CLK(n5026), .C(n5027) );
  CKBD0 U4909 ( .CLK(n5027), .C(n5028) );
  CKBD0 U4910 ( .CLK(n5028), .C(n5029) );
  CKBD0 U4911 ( .CLK(n5029), .C(n5030) );
  BUFFD0 U4912 ( .I(n5030), .Z(n5031) );
  CKBD0 U4913 ( .CLK(n5031), .C(n5032) );
  CKBD0 U4914 ( .CLK(n5032), .C(n5033) );
  CKBD0 U4915 ( .CLK(n5033), .C(n5034) );
  CKBD0 U4916 ( .CLK(n5034), .C(n5035) );
  CKBD0 U4917 ( .CLK(n5035), .C(n5036) );
  CKBD0 U4918 ( .CLK(n5036), .C(n5037) );
  CKBD0 U4919 ( .CLK(n5037), .C(n5038) );
  CKBD0 U4920 ( .CLK(n5038), .C(n5039) );
  CKBD0 U4921 ( .CLK(n5039), .C(n5040) );
  CKBD0 U4922 ( .CLK(n5040), .C(n5041) );
  BUFFD0 U4923 ( .I(n5041), .Z(n5042) );
  CKBD0 U4924 ( .CLK(n5042), .C(n5043) );
  CKBD0 U4925 ( .CLK(n5043), .C(n5044) );
  CKBD0 U4926 ( .CLK(n5044), .C(n5045) );
  CKBD0 U4927 ( .CLK(n5045), .C(n5046) );
  CKBD0 U4928 ( .CLK(n5046), .C(n5047) );
  CKBD0 U4929 ( .CLK(n5047), .C(n5048) );
  CKBD0 U4930 ( .CLK(n5048), .C(n5049) );
  CKBD0 U4931 ( .CLK(n5049), .C(n5050) );
  CKBD0 U4932 ( .CLK(n5050), .C(n5051) );
  CKBD0 U4933 ( .CLK(n5051), .C(n5052) );
  BUFFD0 U4934 ( .I(n5052), .Z(n5053) );
  CKBD0 U4935 ( .CLK(n5053), .C(n5054) );
  CKBD0 U4936 ( .CLK(n5054), .C(n5055) );
  CKBD0 U4937 ( .CLK(n5055), .C(n5056) );
  CKBD0 U4938 ( .CLK(n5056), .C(n5057) );
  CKBD0 U4939 ( .CLK(n5057), .C(n5058) );
  CKBD0 U4940 ( .CLK(n5058), .C(n5059) );
  CKBD0 U4941 ( .CLK(n5059), .C(n5060) );
  CKBD0 U4942 ( .CLK(n5060), .C(n5061) );
  CKBD0 U4943 ( .CLK(n5061), .C(n5062) );
  CKBD0 U4944 ( .CLK(n5062), .C(n5063) );
  BUFFD0 U4945 ( .I(n5063), .Z(n5064) );
  CKBD0 U4946 ( .CLK(n5064), .C(n5065) );
  CKBD0 U4947 ( .CLK(n5065), .C(n5066) );
  CKBD0 U4948 ( .CLK(n5066), .C(n5067) );
  CKBD0 U4949 ( .CLK(n5067), .C(n5068) );
  CKBD0 U4950 ( .CLK(n5068), .C(n5069) );
  CKBD0 U4951 ( .CLK(n5069), .C(n5070) );
  CKBD0 U4952 ( .CLK(n5070), .C(n5071) );
  CKBD0 U4953 ( .CLK(n5071), .C(n5072) );
  CKBD0 U4954 ( .CLK(n5072), .C(n5073) );
  CKBD0 U4955 ( .CLK(n5073), .C(n5074) );
  BUFFD0 U4956 ( .I(n5074), .Z(n5075) );
  CKBD0 U4957 ( .CLK(n5075), .C(n5076) );
  CKBD0 U4958 ( .CLK(n5076), .C(n5077) );
  CKBD0 U4959 ( .CLK(n5077), .C(n5078) );
  CKBD0 U4960 ( .CLK(n5078), .C(n5079) );
  CKBD0 U4961 ( .CLK(n5079), .C(n5080) );
  CKBD0 U4962 ( .CLK(n5080), .C(n5081) );
  CKBD0 U4963 ( .CLK(n5081), .C(n5082) );
  CKBD0 U4964 ( .CLK(n5082), .C(n5083) );
  CKBD0 U4965 ( .CLK(n5083), .C(n5084) );
  CKBD0 U4966 ( .CLK(n5084), .C(n5085) );
  BUFFD0 U4967 ( .I(n5085), .Z(n5086) );
  CKBD0 U4968 ( .CLK(n5086), .C(n5087) );
  CKBD0 U4969 ( .CLK(n5087), .C(n5088) );
  CKBD0 U4970 ( .CLK(n5088), .C(n5089) );
  CKBD0 U4971 ( .CLK(n5089), .C(n5090) );
  CKBD0 U4972 ( .CLK(n5090), .C(n5091) );
  CKBD0 U4973 ( .CLK(n5091), .C(n5092) );
  CKBD0 U4974 ( .CLK(n5092), .C(n5093) );
  CKBD0 U4975 ( .CLK(n5093), .C(n5094) );
  CKBD0 U4976 ( .CLK(n5094), .C(n5095) );
  BUFFD0 U4977 ( .I(n5095), .Z(n5096) );
  CKBD0 U4978 ( .CLK(n5096), .C(n5097) );
  CKBD0 U4979 ( .CLK(n5097), .C(n5098) );
  CKBD0 U4980 ( .CLK(n5098), .C(n5099) );
  CKBD0 U4981 ( .CLK(n5099), .C(n5100) );
  CKBD0 U4982 ( .CLK(n5100), .C(n5101) );
  CKBD0 U4983 ( .CLK(n5101), .C(n5102) );
  CKBD0 U4984 ( .CLK(n5102), .C(n5103) );
  CKBD0 U4985 ( .CLK(n5103), .C(n5104) );
  CKBD0 U4986 ( .CLK(n5104), .C(n5105) );
  CKBD0 U4987 ( .CLK(n5105), .C(n5106) );
  BUFFD0 U4988 ( .I(n5106), .Z(n5107) );
  CKBD0 U4989 ( .CLK(n5107), .C(n5108) );
  CKBD0 U4990 ( .CLK(n5108), .C(n5109) );
  CKBD0 U4991 ( .CLK(n5109), .C(n5110) );
  CKBD0 U4992 ( .CLK(n5110), .C(n5111) );
  CKBD0 U4993 ( .CLK(n5111), .C(n5112) );
  CKBD0 U4994 ( .CLK(n5112), .C(n5113) );
  CKBD0 U4995 ( .CLK(n5113), .C(n5114) );
  CKBD0 U4996 ( .CLK(n5114), .C(n5115) );
  CKBD0 U4997 ( .CLK(n5115), .C(n5116) );
  CKBD0 U4998 ( .CLK(n5116), .C(n5117) );
  BUFFD0 U4999 ( .I(n5117), .Z(n5118) );
  CKBD0 U5000 ( .CLK(n5118), .C(n5119) );
  CKBD0 U5001 ( .CLK(n5119), .C(n5120) );
  CKBD0 U5002 ( .CLK(n5120), .C(n5121) );
  CKBD0 U5003 ( .CLK(n5121), .C(n5122) );
  CKBD0 U5004 ( .CLK(n5122), .C(n5123) );
  CKBD0 U5005 ( .CLK(n5123), .C(n5124) );
  BUFFD0 U5006 ( .I(n5124), .Z(n5125) );
  CKBD0 U5007 ( .CLK(n5125), .C(n5126) );
  BUFFD0 U5008 ( .I(n5126), .Z(n5127) );
  CKBD0 U5009 ( .CLK(n5127), .C(n5128) );
  BUFFD0 U5010 ( .I(n5128), .Z(n5129) );
  CKBD0 U5011 ( .CLK(n5129), .C(n5130) );
  BUFFD0 U5012 ( .I(n5130), .Z(n5131) );
  CKBD0 U5013 ( .CLK(n5131), .C(n5132) );
  BUFFD0 U5014 ( .I(n5132), .Z(n5133) );
  CKBD0 U5015 ( .CLK(n5133), .C(n5134) );
  BUFFD0 U5016 ( .I(n5134), .Z(n5135) );
  CKBD0 U5017 ( .CLK(n5135), .C(n5136) );
  BUFFD0 U5018 ( .I(n5136), .Z(n5137) );
  CKBD0 U5019 ( .CLK(n5137), .C(n5138) );
  BUFFD0 U5020 ( .I(n5138), .Z(n5139) );
  BUFFD0 U5021 ( .I(Decoder[12]), .Z(n5140) );
  BUFFD0 U5022 ( .I(n5142), .Z(n5141) );
  BUFFD0 U5023 ( .I(n5143), .Z(n5142) );
  BUFFD0 U5024 ( .I(n9177), .Z(n5143) );
  CKBD0 U5025 ( .CLK(n1138), .C(n5144) );
  CKBD0 U5026 ( .CLK(n5144), .C(n5145) );
  CKBD0 U5027 ( .CLK(n5145), .C(n5146) );
  BUFFD0 U5028 ( .I(n5146), .Z(n5147) );
  CKBD0 U5029 ( .CLK(n5147), .C(n5148) );
  CKBD0 U5030 ( .CLK(n5148), .C(n5149) );
  CKBD0 U5031 ( .CLK(n5149), .C(n5150) );
  CKBD0 U5032 ( .CLK(n5150), .C(n5151) );
  CKBD0 U5033 ( .CLK(n5151), .C(n5152) );
  CKBD0 U5034 ( .CLK(n5152), .C(n5153) );
  CKBD0 U5035 ( .CLK(n5153), .C(n5154) );
  CKBD0 U5036 ( .CLK(n5154), .C(n5155) );
  CKBD0 U5037 ( .CLK(n5155), .C(n5156) );
  CKBD0 U5038 ( .CLK(n5156), .C(n5157) );
  BUFFD0 U5039 ( .I(n5157), .Z(n5158) );
  CKBD0 U5040 ( .CLK(n5158), .C(n5159) );
  CKBD0 U5041 ( .CLK(n5159), .C(n5160) );
  CKBD0 U5042 ( .CLK(n5160), .C(n5161) );
  CKBD0 U5043 ( .CLK(n5161), .C(n5162) );
  CKBD0 U5044 ( .CLK(n5162), .C(n5163) );
  CKBD0 U5045 ( .CLK(n5163), .C(n5164) );
  CKBD0 U5046 ( .CLK(n5164), .C(n5165) );
  CKBD0 U5047 ( .CLK(n5165), .C(n5166) );
  CKBD0 U5048 ( .CLK(n5166), .C(n5167) );
  BUFFD0 U5049 ( .I(n5167), .Z(n5168) );
  CKBD0 U5050 ( .CLK(n5168), .C(n5169) );
  CKBD0 U5051 ( .CLK(n5169), .C(n5170) );
  CKBD0 U5052 ( .CLK(n5170), .C(n5171) );
  CKBD0 U5053 ( .CLK(n5171), .C(n5172) );
  CKBD0 U5054 ( .CLK(n5172), .C(n5173) );
  CKBD0 U5055 ( .CLK(n5173), .C(n5174) );
  CKBD0 U5056 ( .CLK(n5174), .C(n5175) );
  CKBD0 U5057 ( .CLK(n5175), .C(n5176) );
  CKBD0 U5058 ( .CLK(n5176), .C(n5177) );
  CKBD0 U5059 ( .CLK(n5177), .C(n5178) );
  BUFFD0 U5060 ( .I(n5178), .Z(n5179) );
  CKBD0 U5061 ( .CLK(n5179), .C(n5180) );
  CKBD0 U5062 ( .CLK(n5180), .C(n5181) );
  CKBD0 U5063 ( .CLK(n5181), .C(n5182) );
  CKBD0 U5064 ( .CLK(n5182), .C(n5183) );
  CKBD0 U5065 ( .CLK(n5183), .C(n5184) );
  CKBD0 U5066 ( .CLK(n5184), .C(n5185) );
  CKBD0 U5067 ( .CLK(n5185), .C(n5186) );
  CKBD0 U5068 ( .CLK(n5186), .C(n5187) );
  CKBD0 U5069 ( .CLK(n5187), .C(n5188) );
  CKBD0 U5070 ( .CLK(n5188), .C(n5189) );
  BUFFD0 U5071 ( .I(n5189), .Z(n5190) );
  CKBD0 U5072 ( .CLK(n5190), .C(n5191) );
  CKBD0 U5073 ( .CLK(n5191), .C(n5192) );
  CKBD0 U5074 ( .CLK(n5192), .C(n5193) );
  CKBD0 U5075 ( .CLK(n5193), .C(n5194) );
  CKBD0 U5076 ( .CLK(n5194), .C(n5195) );
  CKBD0 U5077 ( .CLK(n5195), .C(n5196) );
  CKBD0 U5078 ( .CLK(n5196), .C(n5197) );
  CKBD0 U5079 ( .CLK(n5197), .C(n5198) );
  CKBD0 U5080 ( .CLK(n5198), .C(n5199) );
  CKBD0 U5081 ( .CLK(n5199), .C(n5200) );
  BUFFD0 U5082 ( .I(n5200), .Z(n5201) );
  CKBD0 U5083 ( .CLK(n5201), .C(n5202) );
  CKBD0 U5084 ( .CLK(n5202), .C(n5203) );
  CKBD0 U5085 ( .CLK(n5203), .C(n5204) );
  CKBD0 U5086 ( .CLK(n5204), .C(n5205) );
  CKBD0 U5087 ( .CLK(n5205), .C(n5206) );
  CKBD0 U5088 ( .CLK(n5206), .C(n5207) );
  CKBD0 U5089 ( .CLK(n5207), .C(n5208) );
  CKBD0 U5090 ( .CLK(n5208), .C(n5209) );
  CKBD0 U5091 ( .CLK(n5209), .C(n5210) );
  CKBD0 U5092 ( .CLK(n5210), .C(n5211) );
  BUFFD0 U5093 ( .I(n5211), .Z(n5212) );
  CKBD0 U5094 ( .CLK(n5212), .C(n5213) );
  CKBD0 U5095 ( .CLK(n5213), .C(n5214) );
  CKBD0 U5096 ( .CLK(n5214), .C(n5215) );
  CKBD0 U5097 ( .CLK(n5215), .C(n5216) );
  CKBD0 U5098 ( .CLK(n5216), .C(n5217) );
  CKBD0 U5099 ( .CLK(n5217), .C(n5218) );
  CKBD0 U5100 ( .CLK(n5218), .C(n5219) );
  CKBD0 U5101 ( .CLK(n5219), .C(n5220) );
  CKBD0 U5102 ( .CLK(n5220), .C(n5221) );
  CKBD0 U5103 ( .CLK(n5221), .C(n5222) );
  BUFFD0 U5104 ( .I(n5222), .Z(n5223) );
  CKBD0 U5105 ( .CLK(n5223), .C(n5224) );
  CKBD0 U5106 ( .CLK(n5224), .C(n5225) );
  CKBD0 U5107 ( .CLK(n5225), .C(n5226) );
  CKBD0 U5108 ( .CLK(n5226), .C(n5227) );
  CKBD0 U5109 ( .CLK(n5227), .C(n5228) );
  CKBD0 U5110 ( .CLK(n5228), .C(n5229) );
  CKBD0 U5111 ( .CLK(n5229), .C(n5230) );
  CKBD0 U5112 ( .CLK(n5230), .C(n5231) );
  CKBD0 U5113 ( .CLK(n5231), .C(n5232) );
  CKBD0 U5114 ( .CLK(n5232), .C(n5233) );
  BUFFD0 U5115 ( .I(n5233), .Z(n5234) );
  CKBD0 U5116 ( .CLK(n5234), .C(n5235) );
  CKBD0 U5117 ( .CLK(n5235), .C(n5236) );
  CKBD0 U5118 ( .CLK(n5236), .C(n5237) );
  CKBD0 U5119 ( .CLK(n5237), .C(n5238) );
  CKBD0 U5120 ( .CLK(n5238), .C(n5239) );
  CKBD0 U5121 ( .CLK(n5239), .C(n5240) );
  CKBD0 U5122 ( .CLK(n5240), .C(n5241) );
  CKBD0 U5123 ( .CLK(n5241), .C(n5242) );
  CKBD0 U5124 ( .CLK(n5242), .C(n5243) );
  BUFFD0 U5125 ( .I(n5243), .Z(n5244) );
  CKBD0 U5126 ( .CLK(n5244), .C(n5245) );
  CKBD0 U5127 ( .CLK(n5245), .C(n5246) );
  CKBD0 U5128 ( .CLK(n5246), .C(n5247) );
  CKBD0 U5129 ( .CLK(n5247), .C(n5248) );
  CKBD0 U5130 ( .CLK(n5248), .C(n5249) );
  CKBD0 U5131 ( .CLK(n5249), .C(n5250) );
  CKBD0 U5132 ( .CLK(n5250), .C(n5251) );
  CKBD0 U5133 ( .CLK(n5251), .C(n5252) );
  CKBD0 U5134 ( .CLK(n5252), .C(n5253) );
  CKBD0 U5135 ( .CLK(n5253), .C(n5254) );
  BUFFD0 U5136 ( .I(n5254), .Z(n5255) );
  CKBD0 U5137 ( .CLK(n5255), .C(n5256) );
  CKBD0 U5138 ( .CLK(n5256), .C(n5257) );
  CKBD0 U5139 ( .CLK(n5257), .C(n5258) );
  CKBD0 U5140 ( .CLK(n5258), .C(n5259) );
  CKBD0 U5141 ( .CLK(n5259), .C(n5260) );
  CKBD0 U5142 ( .CLK(n5260), .C(n5261) );
  BUFFD0 U5143 ( .I(n5261), .Z(n5262) );
  CKBD0 U5144 ( .CLK(n5262), .C(n5263) );
  BUFFD0 U5145 ( .I(n5263), .Z(n5264) );
  CKBD0 U5146 ( .CLK(n5264), .C(n5265) );
  BUFFD0 U5147 ( .I(n5265), .Z(n5266) );
  CKBD0 U5148 ( .CLK(n5266), .C(n5267) );
  BUFFD0 U5149 ( .I(n5267), .Z(n5268) );
  CKBD0 U5150 ( .CLK(n5268), .C(n5269) );
  BUFFD0 U5151 ( .I(n5269), .Z(n5270) );
  CKBD0 U5152 ( .CLK(n5270), .C(n5271) );
  BUFFD0 U5153 ( .I(n5271), .Z(n5272) );
  CKBD0 U5154 ( .CLK(n5272), .C(n5273) );
  BUFFD0 U5155 ( .I(n5273), .Z(n5274) );
  CKBD0 U5156 ( .CLK(n5274), .C(n5275) );
  BUFFD0 U5157 ( .I(n5275), .Z(n5276) );
  BUFFD0 U5158 ( .I(n5278), .Z(n5277) );
  BUFFD0 U5159 ( .I(n5279), .Z(n5278) );
  BUFFD0 U5160 ( .I(n9178), .Z(n5279) );
  CKBD0 U5161 ( .CLK(n1136), .C(n5280) );
  CKBD0 U5162 ( .CLK(n5280), .C(n5281) );
  CKBD0 U5163 ( .CLK(n5281), .C(n5282) );
  BUFFD0 U5164 ( .I(n5282), .Z(n5283) );
  CKBD0 U5165 ( .CLK(n5283), .C(n5284) );
  CKBD0 U5166 ( .CLK(n5284), .C(n5285) );
  CKBD0 U5167 ( .CLK(n5285), .C(n5286) );
  CKBD0 U5168 ( .CLK(n5286), .C(n5287) );
  CKBD0 U5169 ( .CLK(n5287), .C(n5288) );
  CKBD0 U5170 ( .CLK(n5288), .C(n5289) );
  CKBD0 U5171 ( .CLK(n5289), .C(n5290) );
  CKBD0 U5172 ( .CLK(n5290), .C(n5291) );
  CKBD0 U5173 ( .CLK(n5291), .C(n5292) );
  CKBD0 U5174 ( .CLK(n5292), .C(n5293) );
  BUFFD0 U5175 ( .I(n5293), .Z(n5294) );
  CKBD0 U5176 ( .CLK(n5294), .C(n5295) );
  CKBD0 U5177 ( .CLK(n5295), .C(n5296) );
  CKBD0 U5178 ( .CLK(n5296), .C(n5297) );
  CKBD0 U5179 ( .CLK(n5297), .C(n5298) );
  CKBD0 U5180 ( .CLK(n5298), .C(n5299) );
  CKBD0 U5181 ( .CLK(n5299), .C(n5300) );
  CKBD0 U5182 ( .CLK(n5300), .C(n5301) );
  CKBD0 U5183 ( .CLK(n5301), .C(n5302) );
  CKBD0 U5184 ( .CLK(n5302), .C(n5303) );
  BUFFD0 U5185 ( .I(n5303), .Z(n5304) );
  CKBD0 U5186 ( .CLK(n5304), .C(n5305) );
  CKBD0 U5187 ( .CLK(n5305), .C(n5306) );
  CKBD0 U5188 ( .CLK(n5306), .C(n5307) );
  CKBD0 U5189 ( .CLK(n5307), .C(n5308) );
  CKBD0 U5190 ( .CLK(n5308), .C(n5309) );
  CKBD0 U5191 ( .CLK(n5309), .C(n5310) );
  CKBD0 U5192 ( .CLK(n5310), .C(n5311) );
  CKBD0 U5193 ( .CLK(n5311), .C(n5312) );
  CKBD0 U5194 ( .CLK(n5312), .C(n5313) );
  CKBD0 U5195 ( .CLK(n5313), .C(n5314) );
  BUFFD0 U5196 ( .I(n5314), .Z(n5315) );
  CKBD0 U5197 ( .CLK(n5315), .C(n5316) );
  CKBD0 U5198 ( .CLK(n5316), .C(n5317) );
  CKBD0 U5199 ( .CLK(n5317), .C(n5318) );
  CKBD0 U5200 ( .CLK(n5318), .C(n5319) );
  CKBD0 U5201 ( .CLK(n5319), .C(n5320) );
  CKBD0 U5202 ( .CLK(n5320), .C(n5321) );
  CKBD0 U5203 ( .CLK(n5321), .C(n5322) );
  CKBD0 U5204 ( .CLK(n5322), .C(n5323) );
  CKBD0 U5205 ( .CLK(n5323), .C(n5324) );
  CKBD0 U5206 ( .CLK(n5324), .C(n5325) );
  BUFFD0 U5207 ( .I(n5325), .Z(n5326) );
  CKBD0 U5208 ( .CLK(n5326), .C(n5327) );
  CKBD0 U5209 ( .CLK(n5327), .C(n5328) );
  CKBD0 U5210 ( .CLK(n5328), .C(n5329) );
  CKBD0 U5211 ( .CLK(n5329), .C(n5330) );
  CKBD0 U5212 ( .CLK(n5330), .C(n5331) );
  CKBD0 U5213 ( .CLK(n5331), .C(n5332) );
  CKBD0 U5214 ( .CLK(n5332), .C(n5333) );
  CKBD0 U5215 ( .CLK(n5333), .C(n5334) );
  CKBD0 U5216 ( .CLK(n5334), .C(n5335) );
  CKBD0 U5217 ( .CLK(n5335), .C(n5336) );
  BUFFD0 U5218 ( .I(n5336), .Z(n5337) );
  CKBD0 U5219 ( .CLK(n5337), .C(n5338) );
  CKBD0 U5220 ( .CLK(n5338), .C(n5339) );
  CKBD0 U5221 ( .CLK(n5339), .C(n5340) );
  CKBD0 U5222 ( .CLK(n5340), .C(n5341) );
  CKBD0 U5223 ( .CLK(n5341), .C(n5342) );
  CKBD0 U5224 ( .CLK(n5342), .C(n5343) );
  CKBD0 U5225 ( .CLK(n5343), .C(n5344) );
  CKBD0 U5226 ( .CLK(n5344), .C(n5345) );
  CKBD0 U5227 ( .CLK(n5345), .C(n5346) );
  CKBD0 U5228 ( .CLK(n5346), .C(n5347) );
  BUFFD0 U5229 ( .I(n5347), .Z(n5348) );
  CKBD0 U5230 ( .CLK(n5348), .C(n5349) );
  CKBD0 U5231 ( .CLK(n5349), .C(n5350) );
  CKBD0 U5232 ( .CLK(n5350), .C(n5351) );
  CKBD0 U5233 ( .CLK(n5351), .C(n5352) );
  CKBD0 U5234 ( .CLK(n5352), .C(n5353) );
  CKBD0 U5235 ( .CLK(n5353), .C(n5354) );
  CKBD0 U5236 ( .CLK(n5354), .C(n5355) );
  CKBD0 U5237 ( .CLK(n5355), .C(n5356) );
  CKBD0 U5238 ( .CLK(n5356), .C(n5357) );
  CKBD0 U5239 ( .CLK(n5357), .C(n5358) );
  BUFFD0 U5240 ( .I(n5358), .Z(n5359) );
  CKBD0 U5241 ( .CLK(n5359), .C(n5360) );
  CKBD0 U5242 ( .CLK(n5360), .C(n5361) );
  CKBD0 U5243 ( .CLK(n5361), .C(n5362) );
  CKBD0 U5244 ( .CLK(n5362), .C(n5363) );
  CKBD0 U5245 ( .CLK(n5363), .C(n5364) );
  CKBD0 U5246 ( .CLK(n5364), .C(n5365) );
  CKBD0 U5247 ( .CLK(n5365), .C(n5366) );
  CKBD0 U5248 ( .CLK(n5366), .C(n5367) );
  CKBD0 U5249 ( .CLK(n5367), .C(n5368) );
  CKBD0 U5250 ( .CLK(n5368), .C(n5369) );
  BUFFD0 U5251 ( .I(n5369), .Z(n5370) );
  CKBD0 U5252 ( .CLK(n5370), .C(n5371) );
  CKBD0 U5253 ( .CLK(n5371), .C(n5372) );
  CKBD0 U5254 ( .CLK(n5372), .C(n5373) );
  CKBD0 U5255 ( .CLK(n5373), .C(n5374) );
  CKBD0 U5256 ( .CLK(n5374), .C(n5375) );
  CKBD0 U5257 ( .CLK(n5375), .C(n5376) );
  CKBD0 U5258 ( .CLK(n5376), .C(n5377) );
  CKBD0 U5259 ( .CLK(n5377), .C(n5378) );
  CKBD0 U5260 ( .CLK(n5378), .C(n5379) );
  BUFFD0 U5261 ( .I(n5379), .Z(n5380) );
  CKBD0 U5262 ( .CLK(n5380), .C(n5381) );
  CKBD0 U5263 ( .CLK(n5381), .C(n5382) );
  CKBD0 U5264 ( .CLK(n5382), .C(n5383) );
  CKBD0 U5265 ( .CLK(n5383), .C(n5384) );
  CKBD0 U5266 ( .CLK(n5384), .C(n5385) );
  CKBD0 U5267 ( .CLK(n5385), .C(n5386) );
  CKBD0 U5268 ( .CLK(n5386), .C(n5387) );
  CKBD0 U5269 ( .CLK(n5387), .C(n5388) );
  CKBD0 U5270 ( .CLK(n5388), .C(n5389) );
  CKBD0 U5271 ( .CLK(n5389), .C(n5390) );
  BUFFD0 U5272 ( .I(n5390), .Z(n5391) );
  CKBD0 U5273 ( .CLK(n5391), .C(n5392) );
  CKBD0 U5274 ( .CLK(n5392), .C(n5393) );
  CKBD0 U5275 ( .CLK(n5393), .C(n5394) );
  CKBD0 U5276 ( .CLK(n5394), .C(n5395) );
  CKBD0 U5277 ( .CLK(n5395), .C(n5396) );
  CKBD0 U5278 ( .CLK(n5396), .C(n5397) );
  BUFFD0 U5279 ( .I(n5397), .Z(n5398) );
  CKBD0 U5280 ( .CLK(n5398), .C(n5399) );
  BUFFD0 U5281 ( .I(n5399), .Z(n5400) );
  CKBD0 U5282 ( .CLK(n5400), .C(n5401) );
  BUFFD0 U5283 ( .I(n5401), .Z(n5402) );
  CKBD0 U5284 ( .CLK(n5402), .C(n5403) );
  BUFFD0 U5285 ( .I(n5403), .Z(n5404) );
  CKBD0 U5286 ( .CLK(n5404), .C(n5405) );
  BUFFD0 U5287 ( .I(n5405), .Z(n5406) );
  CKBD0 U5288 ( .CLK(n5406), .C(n5407) );
  BUFFD0 U5289 ( .I(n5407), .Z(n5408) );
  CKBD0 U5290 ( .CLK(n5408), .C(n5409) );
  BUFFD0 U5291 ( .I(n5409), .Z(n5410) );
  CKBD0 U5292 ( .CLK(n5410), .C(n5411) );
  BUFFD0 U5293 ( .I(n5411), .Z(n5412) );
  BUFFD0 U5294 ( .I(n5414), .Z(n5413) );
  BUFFD0 U5295 ( .I(n5415), .Z(n5414) );
  BUFFD0 U5296 ( .I(n9179), .Z(n5415) );
  CKBD0 U5297 ( .CLK(n1134), .C(n5416) );
  CKBD0 U5298 ( .CLK(n5416), .C(n5417) );
  CKBD0 U5299 ( .CLK(n5417), .C(n5418) );
  BUFFD0 U5300 ( .I(n5418), .Z(n5419) );
  CKBD0 U5301 ( .CLK(n5419), .C(n5420) );
  CKBD0 U5302 ( .CLK(n5420), .C(n5421) );
  CKBD0 U5303 ( .CLK(n5421), .C(n5422) );
  CKBD0 U5304 ( .CLK(n5422), .C(n5423) );
  CKBD0 U5305 ( .CLK(n5423), .C(n5424) );
  CKBD0 U5306 ( .CLK(n5424), .C(n5425) );
  CKBD0 U5307 ( .CLK(n5425), .C(n5426) );
  CKBD0 U5308 ( .CLK(n5426), .C(n5427) );
  CKBD0 U5309 ( .CLK(n5427), .C(n5428) );
  CKBD0 U5310 ( .CLK(n5428), .C(n5429) );
  BUFFD0 U5311 ( .I(n5429), .Z(n5430) );
  CKBD0 U5312 ( .CLK(n5430), .C(n5431) );
  CKBD0 U5313 ( .CLK(n5431), .C(n5432) );
  CKBD0 U5314 ( .CLK(n5432), .C(n5433) );
  CKBD0 U5315 ( .CLK(n5433), .C(n5434) );
  CKBD0 U5316 ( .CLK(n5434), .C(n5435) );
  CKBD0 U5317 ( .CLK(n5435), .C(n5436) );
  CKBD0 U5318 ( .CLK(n5436), .C(n5437) );
  CKBD0 U5319 ( .CLK(n5437), .C(n5438) );
  CKBD0 U5320 ( .CLK(n5438), .C(n5439) );
  BUFFD0 U5321 ( .I(n5439), .Z(n5440) );
  CKBD0 U5322 ( .CLK(n5440), .C(n5441) );
  CKBD0 U5323 ( .CLK(n5441), .C(n5442) );
  CKBD0 U5324 ( .CLK(n5442), .C(n5443) );
  CKBD0 U5325 ( .CLK(n5443), .C(n5444) );
  CKBD0 U5326 ( .CLK(n5444), .C(n5445) );
  CKBD0 U5327 ( .CLK(n5445), .C(n5446) );
  CKBD0 U5328 ( .CLK(n5446), .C(n5447) );
  CKBD0 U5329 ( .CLK(n5447), .C(n5448) );
  CKBD0 U5330 ( .CLK(n5448), .C(n5449) );
  CKBD0 U5331 ( .CLK(n5449), .C(n5450) );
  BUFFD0 U5332 ( .I(n5450), .Z(n5451) );
  CKBD0 U5333 ( .CLK(n5451), .C(n5452) );
  CKBD0 U5334 ( .CLK(n5452), .C(n5453) );
  CKBD0 U5335 ( .CLK(n5453), .C(n5454) );
  CKBD0 U5336 ( .CLK(n5454), .C(n5455) );
  CKBD0 U5337 ( .CLK(n5455), .C(n5456) );
  CKBD0 U5338 ( .CLK(n5456), .C(n5457) );
  CKBD0 U5339 ( .CLK(n5457), .C(n5458) );
  CKBD0 U5340 ( .CLK(n5458), .C(n5459) );
  CKBD0 U5341 ( .CLK(n5459), .C(n5460) );
  CKBD0 U5342 ( .CLK(n5460), .C(n5461) );
  BUFFD0 U5343 ( .I(n5461), .Z(n5462) );
  CKBD0 U5344 ( .CLK(n5462), .C(n5463) );
  CKBD0 U5345 ( .CLK(n5463), .C(n5464) );
  CKBD0 U5346 ( .CLK(n5464), .C(n5465) );
  CKBD0 U5347 ( .CLK(n5465), .C(n5466) );
  CKBD0 U5348 ( .CLK(n5466), .C(n5467) );
  CKBD0 U5349 ( .CLK(n5467), .C(n5468) );
  CKBD0 U5350 ( .CLK(n5468), .C(n5469) );
  CKBD0 U5351 ( .CLK(n5469), .C(n5470) );
  CKBD0 U5352 ( .CLK(n5470), .C(n5471) );
  CKBD0 U5353 ( .CLK(n5471), .C(n5472) );
  BUFFD0 U5354 ( .I(n5472), .Z(n5473) );
  CKBD0 U5355 ( .CLK(n5473), .C(n5474) );
  CKBD0 U5356 ( .CLK(n5474), .C(n5475) );
  CKBD0 U5357 ( .CLK(n5475), .C(n5476) );
  CKBD0 U5358 ( .CLK(n5476), .C(n5477) );
  CKBD0 U5359 ( .CLK(n5477), .C(n5478) );
  CKBD0 U5360 ( .CLK(n5478), .C(n5479) );
  CKBD0 U5361 ( .CLK(n5479), .C(n5480) );
  CKBD0 U5362 ( .CLK(n5480), .C(n5481) );
  CKBD0 U5363 ( .CLK(n5481), .C(n5482) );
  CKBD0 U5364 ( .CLK(n5482), .C(n5483) );
  BUFFD0 U5365 ( .I(n5483), .Z(n5484) );
  CKBD0 U5366 ( .CLK(n5484), .C(n5485) );
  CKBD0 U5367 ( .CLK(n5485), .C(n5486) );
  CKBD0 U5368 ( .CLK(n5486), .C(n5487) );
  CKBD0 U5369 ( .CLK(n5487), .C(n5488) );
  CKBD0 U5370 ( .CLK(n5488), .C(n5489) );
  CKBD0 U5371 ( .CLK(n5489), .C(n5490) );
  CKBD0 U5372 ( .CLK(n5490), .C(n5491) );
  CKBD0 U5373 ( .CLK(n5491), .C(n5492) );
  CKBD0 U5374 ( .CLK(n5492), .C(n5493) );
  CKBD0 U5375 ( .CLK(n5493), .C(n5494) );
  BUFFD0 U5376 ( .I(n5494), .Z(n5495) );
  CKBD0 U5377 ( .CLK(n5495), .C(n5496) );
  CKBD0 U5378 ( .CLK(n5496), .C(n5497) );
  CKBD0 U5379 ( .CLK(n5497), .C(n5498) );
  CKBD0 U5380 ( .CLK(n5498), .C(n5499) );
  CKBD0 U5381 ( .CLK(n5499), .C(n5500) );
  CKBD0 U5382 ( .CLK(n5500), .C(n5501) );
  CKBD0 U5383 ( .CLK(n5501), .C(n5502) );
  CKBD0 U5384 ( .CLK(n5502), .C(n5503) );
  CKBD0 U5385 ( .CLK(n5503), .C(n5504) );
  BUFFD0 U5386 ( .I(n5504), .Z(n5505) );
  CKBD0 U5387 ( .CLK(n5505), .C(n5506) );
  CKBD0 U5388 ( .CLK(n5506), .C(n5507) );
  CKBD0 U5389 ( .CLK(n5507), .C(n5508) );
  CKBD0 U5390 ( .CLK(n5508), .C(n5509) );
  CKBD0 U5391 ( .CLK(n5509), .C(n5510) );
  CKBD0 U5392 ( .CLK(n5510), .C(n5511) );
  CKBD0 U5393 ( .CLK(n5511), .C(n5512) );
  CKBD0 U5394 ( .CLK(n5512), .C(n5513) );
  CKBD0 U5395 ( .CLK(n5513), .C(n5514) );
  CKBD0 U5396 ( .CLK(n5514), .C(n5515) );
  BUFFD0 U5397 ( .I(n5515), .Z(n5516) );
  CKBD0 U5398 ( .CLK(n5516), .C(n5517) );
  CKBD0 U5399 ( .CLK(n5517), .C(n5518) );
  CKBD0 U5400 ( .CLK(n5518), .C(n5519) );
  CKBD0 U5401 ( .CLK(n5519), .C(n5520) );
  CKBD0 U5402 ( .CLK(n5520), .C(n5521) );
  CKBD0 U5403 ( .CLK(n5521), .C(n5522) );
  CKBD0 U5404 ( .CLK(n5522), .C(n5523) );
  CKBD0 U5405 ( .CLK(n5523), .C(n5524) );
  CKBD0 U5406 ( .CLK(n5524), .C(n5525) );
  CKBD0 U5407 ( .CLK(n5525), .C(n5526) );
  BUFFD0 U5408 ( .I(n5526), .Z(n5527) );
  CKBD0 U5409 ( .CLK(n5527), .C(n5528) );
  CKBD0 U5410 ( .CLK(n5528), .C(n5529) );
  CKBD0 U5411 ( .CLK(n5529), .C(n5530) );
  CKBD0 U5412 ( .CLK(n5530), .C(n5531) );
  CKBD0 U5413 ( .CLK(n5531), .C(n5532) );
  CKBD0 U5414 ( .CLK(n5532), .C(n5533) );
  BUFFD0 U5415 ( .I(n5533), .Z(n5534) );
  CKBD0 U5416 ( .CLK(n5534), .C(n5535) );
  BUFFD0 U5417 ( .I(n5535), .Z(n5536) );
  CKBD0 U5418 ( .CLK(n5536), .C(n5537) );
  BUFFD0 U5419 ( .I(n5537), .Z(n5538) );
  CKBD0 U5420 ( .CLK(n5538), .C(n5539) );
  BUFFD0 U5421 ( .I(n5539), .Z(n5540) );
  CKBD0 U5422 ( .CLK(n5540), .C(n5541) );
  BUFFD0 U5423 ( .I(n5541), .Z(n5542) );
  CKBD0 U5424 ( .CLK(n5542), .C(n5543) );
  BUFFD0 U5425 ( .I(n5543), .Z(n5544) );
  CKBD0 U5426 ( .CLK(n5544), .C(n5545) );
  BUFFD0 U5427 ( .I(n5545), .Z(n5546) );
  CKBD0 U5428 ( .CLK(n5546), .C(n5547) );
  BUFFD0 U5429 ( .I(n5547), .Z(n5548) );
  BUFFD0 U5430 ( .I(n5550), .Z(n5549) );
  BUFFD0 U5431 ( .I(n5551), .Z(n5550) );
  BUFFD0 U5432 ( .I(n9180), .Z(n5551) );
  CKBD0 U5433 ( .CLK(n1132), .C(n5552) );
  CKBD0 U5434 ( .CLK(n5552), .C(n5553) );
  CKBD0 U5435 ( .CLK(n5553), .C(n5554) );
  BUFFD0 U5436 ( .I(n5554), .Z(n5555) );
  CKBD0 U5437 ( .CLK(n5555), .C(n5556) );
  CKBD0 U5438 ( .CLK(n5556), .C(n5557) );
  CKBD0 U5439 ( .CLK(n5557), .C(n5558) );
  CKBD0 U5440 ( .CLK(n5558), .C(n5559) );
  CKBD0 U5441 ( .CLK(n5559), .C(n5560) );
  CKBD0 U5442 ( .CLK(n5560), .C(n5561) );
  CKBD0 U5443 ( .CLK(n5561), .C(n5562) );
  CKBD0 U5444 ( .CLK(n5562), .C(n5563) );
  CKBD0 U5445 ( .CLK(n5563), .C(n5564) );
  CKBD0 U5446 ( .CLK(n5564), .C(n5565) );
  BUFFD0 U5447 ( .I(n5565), .Z(n5566) );
  CKBD0 U5448 ( .CLK(n5566), .C(n5567) );
  CKBD0 U5449 ( .CLK(n5567), .C(n5568) );
  CKBD0 U5450 ( .CLK(n5568), .C(n5569) );
  CKBD0 U5451 ( .CLK(n5569), .C(n5570) );
  CKBD0 U5452 ( .CLK(n5570), .C(n5571) );
  CKBD0 U5453 ( .CLK(n5571), .C(n5572) );
  CKBD0 U5454 ( .CLK(n5572), .C(n5573) );
  CKBD0 U5455 ( .CLK(n5573), .C(n5574) );
  CKBD0 U5456 ( .CLK(n5574), .C(n5575) );
  BUFFD0 U5457 ( .I(n5575), .Z(n5576) );
  CKBD0 U5458 ( .CLK(n5576), .C(n5577) );
  CKBD0 U5459 ( .CLK(n5577), .C(n5578) );
  CKBD0 U5460 ( .CLK(n5578), .C(n5579) );
  CKBD0 U5461 ( .CLK(n5579), .C(n5580) );
  CKBD0 U5462 ( .CLK(n5580), .C(n5581) );
  CKBD0 U5463 ( .CLK(n5581), .C(n5582) );
  CKBD0 U5464 ( .CLK(n5582), .C(n5583) );
  CKBD0 U5465 ( .CLK(n5583), .C(n5584) );
  CKBD0 U5466 ( .CLK(n5584), .C(n5585) );
  CKBD0 U5467 ( .CLK(n5585), .C(n5586) );
  BUFFD0 U5468 ( .I(n5586), .Z(n5587) );
  CKBD0 U5469 ( .CLK(n5587), .C(n5588) );
  CKBD0 U5470 ( .CLK(n5588), .C(n5589) );
  CKBD0 U5471 ( .CLK(n5589), .C(n5590) );
  CKBD0 U5472 ( .CLK(n5590), .C(n5591) );
  CKBD0 U5473 ( .CLK(n5591), .C(n5592) );
  CKBD0 U5474 ( .CLK(n5592), .C(n5593) );
  CKBD0 U5475 ( .CLK(n5593), .C(n5594) );
  CKBD0 U5476 ( .CLK(n5594), .C(n5595) );
  CKBD0 U5477 ( .CLK(n5595), .C(n5596) );
  CKBD0 U5478 ( .CLK(n5596), .C(n5597) );
  BUFFD0 U5479 ( .I(n5597), .Z(n5598) );
  CKBD0 U5480 ( .CLK(n5598), .C(n5599) );
  CKBD0 U5481 ( .CLK(n5599), .C(n5600) );
  CKBD0 U5482 ( .CLK(n5600), .C(n5601) );
  CKBD0 U5483 ( .CLK(n5601), .C(n5602) );
  CKBD0 U5484 ( .CLK(n5602), .C(n5603) );
  CKBD0 U5485 ( .CLK(n5603), .C(n5604) );
  CKBD0 U5486 ( .CLK(n5604), .C(n5605) );
  CKBD0 U5487 ( .CLK(n5605), .C(n5606) );
  CKBD0 U5488 ( .CLK(n5606), .C(n5607) );
  CKBD0 U5489 ( .CLK(n5607), .C(n5608) );
  BUFFD0 U5490 ( .I(n5608), .Z(n5609) );
  CKBD0 U5491 ( .CLK(n5609), .C(n5610) );
  CKBD0 U5492 ( .CLK(n5610), .C(n5611) );
  CKBD0 U5493 ( .CLK(n5611), .C(n5612) );
  CKBD0 U5494 ( .CLK(n5612), .C(n5613) );
  CKBD0 U5495 ( .CLK(n5613), .C(n5614) );
  CKBD0 U5496 ( .CLK(n5614), .C(n5615) );
  CKBD0 U5497 ( .CLK(n5615), .C(n5616) );
  CKBD0 U5498 ( .CLK(n5616), .C(n5617) );
  CKBD0 U5499 ( .CLK(n5617), .C(n5618) );
  CKBD0 U5500 ( .CLK(n5618), .C(n5619) );
  BUFFD0 U5501 ( .I(n5619), .Z(n5620) );
  CKBD0 U5502 ( .CLK(n5620), .C(n5621) );
  CKBD0 U5503 ( .CLK(n5621), .C(n5622) );
  CKBD0 U5504 ( .CLK(n5622), .C(n5623) );
  CKBD0 U5505 ( .CLK(n5623), .C(n5624) );
  CKBD0 U5506 ( .CLK(n5624), .C(n5625) );
  CKBD0 U5507 ( .CLK(n5625), .C(n5626) );
  CKBD0 U5508 ( .CLK(n5626), .C(n5627) );
  CKBD0 U5509 ( .CLK(n5627), .C(n5628) );
  CKBD0 U5510 ( .CLK(n5628), .C(n5629) );
  CKBD0 U5511 ( .CLK(n5629), .C(n5630) );
  BUFFD0 U5512 ( .I(n5630), .Z(n5631) );
  CKBD0 U5513 ( .CLK(n5631), .C(n5632) );
  CKBD0 U5514 ( .CLK(n5632), .C(n5633) );
  CKBD0 U5515 ( .CLK(n5633), .C(n5634) );
  CKBD0 U5516 ( .CLK(n5634), .C(n5635) );
  CKBD0 U5517 ( .CLK(n5635), .C(n5636) );
  CKBD0 U5518 ( .CLK(n5636), .C(n5637) );
  CKBD0 U5519 ( .CLK(n5637), .C(n5638) );
  CKBD0 U5520 ( .CLK(n5638), .C(n5639) );
  CKBD0 U5521 ( .CLK(n5639), .C(n5640) );
  BUFFD0 U5522 ( .I(n5640), .Z(n5641) );
  CKBD0 U5523 ( .CLK(n5641), .C(n5642) );
  CKBD0 U5524 ( .CLK(n5642), .C(n5643) );
  CKBD0 U5525 ( .CLK(n5643), .C(n5644) );
  CKBD0 U5526 ( .CLK(n5644), .C(n5645) );
  CKBD0 U5527 ( .CLK(n5645), .C(n5646) );
  CKBD0 U5528 ( .CLK(n5646), .C(n5647) );
  CKBD0 U5529 ( .CLK(n5647), .C(n5648) );
  CKBD0 U5530 ( .CLK(n5648), .C(n5649) );
  CKBD0 U5531 ( .CLK(n5649), .C(n5650) );
  CKBD0 U5532 ( .CLK(n5650), .C(n5651) );
  BUFFD0 U5533 ( .I(n5651), .Z(n5652) );
  CKBD0 U5534 ( .CLK(n5652), .C(n5653) );
  CKBD0 U5535 ( .CLK(n5653), .C(n5654) );
  CKBD0 U5536 ( .CLK(n5654), .C(n5655) );
  CKBD0 U5537 ( .CLK(n5655), .C(n5656) );
  CKBD0 U5538 ( .CLK(n5656), .C(n5657) );
  CKBD0 U5539 ( .CLK(n5657), .C(n5658) );
  CKBD0 U5540 ( .CLK(n5658), .C(n5659) );
  CKBD0 U5541 ( .CLK(n5659), .C(n5660) );
  CKBD0 U5542 ( .CLK(n5660), .C(n5661) );
  CKBD0 U5543 ( .CLK(n5661), .C(n5662) );
  BUFFD0 U5544 ( .I(n5662), .Z(n5663) );
  CKBD0 U5545 ( .CLK(n5663), .C(n5664) );
  CKBD0 U5546 ( .CLK(n5664), .C(n5665) );
  CKBD0 U5547 ( .CLK(n5665), .C(n5666) );
  CKBD0 U5548 ( .CLK(n5666), .C(n5667) );
  CKBD0 U5549 ( .CLK(n5667), .C(n5668) );
  CKBD0 U5550 ( .CLK(n5668), .C(n5669) );
  BUFFD0 U5551 ( .I(n5669), .Z(n5670) );
  CKBD0 U5552 ( .CLK(n5670), .C(n5671) );
  BUFFD0 U5553 ( .I(n5671), .Z(n5672) );
  CKBD0 U5554 ( .CLK(n5672), .C(n5673) );
  BUFFD0 U5555 ( .I(n5673), .Z(n5674) );
  CKBD0 U5556 ( .CLK(n5674), .C(n5675) );
  BUFFD0 U5557 ( .I(n5675), .Z(n5676) );
  CKBD0 U5558 ( .CLK(n5676), .C(n5677) );
  BUFFD0 U5559 ( .I(n5677), .Z(n5678) );
  CKBD0 U5560 ( .CLK(n5678), .C(n5679) );
  BUFFD0 U5561 ( .I(n5679), .Z(n5680) );
  CKBD0 U5562 ( .CLK(n5680), .C(n5681) );
  BUFFD0 U5563 ( .I(n5681), .Z(n5682) );
  CKBD0 U5564 ( .CLK(n5682), .C(n5683) );
  BUFFD0 U5565 ( .I(n5683), .Z(n5684) );
  BUFFD0 U5566 ( .I(n5686), .Z(n5685) );
  BUFFD0 U5567 ( .I(n5687), .Z(n5686) );
  BUFFD0 U5568 ( .I(n9181), .Z(n5687) );
  CKBD0 U5569 ( .CLK(n1130), .C(n5688) );
  CKBD0 U5570 ( .CLK(n5688), .C(n5689) );
  CKBD0 U5571 ( .CLK(n5689), .C(n5690) );
  BUFFD0 U5572 ( .I(n5690), .Z(n5691) );
  CKBD0 U5573 ( .CLK(n5691), .C(n5692) );
  CKBD0 U5574 ( .CLK(n5692), .C(n5693) );
  CKBD0 U5575 ( .CLK(n5693), .C(n5694) );
  CKBD0 U5576 ( .CLK(n5694), .C(n5695) );
  CKBD0 U5577 ( .CLK(n5695), .C(n5696) );
  CKBD0 U5578 ( .CLK(n5696), .C(n5697) );
  CKBD0 U5579 ( .CLK(n5697), .C(n5698) );
  CKBD0 U5580 ( .CLK(n5698), .C(n5699) );
  CKBD0 U5581 ( .CLK(n5699), .C(n5700) );
  CKBD0 U5582 ( .CLK(n5700), .C(n5701) );
  BUFFD0 U5583 ( .I(n5701), .Z(n5702) );
  CKBD0 U5584 ( .CLK(n5702), .C(n5703) );
  CKBD0 U5585 ( .CLK(n5703), .C(n5704) );
  CKBD0 U5586 ( .CLK(n5704), .C(n5705) );
  CKBD0 U5587 ( .CLK(n5705), .C(n5706) );
  CKBD0 U5588 ( .CLK(n5706), .C(n5707) );
  CKBD0 U5589 ( .CLK(n5707), .C(n5708) );
  CKBD0 U5590 ( .CLK(n5708), .C(n5709) );
  CKBD0 U5591 ( .CLK(n5709), .C(n5710) );
  CKBD0 U5592 ( .CLK(n5710), .C(n5711) );
  BUFFD0 U5593 ( .I(n5711), .Z(n5712) );
  CKBD0 U5594 ( .CLK(n5712), .C(n5713) );
  CKBD0 U5595 ( .CLK(n5713), .C(n5714) );
  CKBD0 U5596 ( .CLK(n5714), .C(n5715) );
  CKBD0 U5597 ( .CLK(n5715), .C(n5716) );
  CKBD0 U5598 ( .CLK(n5716), .C(n5717) );
  CKBD0 U5599 ( .CLK(n5717), .C(n5718) );
  CKBD0 U5600 ( .CLK(n5718), .C(n5719) );
  CKBD0 U5601 ( .CLK(n5719), .C(n5720) );
  CKBD0 U5602 ( .CLK(n5720), .C(n5721) );
  CKBD0 U5603 ( .CLK(n5721), .C(n5722) );
  BUFFD0 U5604 ( .I(n5722), .Z(n5723) );
  CKBD0 U5605 ( .CLK(n5723), .C(n5724) );
  CKBD0 U5606 ( .CLK(n5724), .C(n5725) );
  CKBD0 U5607 ( .CLK(n5725), .C(n5726) );
  CKBD0 U5608 ( .CLK(n5726), .C(n5727) );
  CKBD0 U5609 ( .CLK(n5727), .C(n5728) );
  CKBD0 U5610 ( .CLK(n5728), .C(n5729) );
  CKBD0 U5611 ( .CLK(n5729), .C(n5730) );
  CKBD0 U5612 ( .CLK(n5730), .C(n5731) );
  CKBD0 U5613 ( .CLK(n5731), .C(n5732) );
  CKBD0 U5614 ( .CLK(n5732), .C(n5733) );
  BUFFD0 U5615 ( .I(n5733), .Z(n5734) );
  CKBD0 U5616 ( .CLK(n5734), .C(n5735) );
  CKBD0 U5617 ( .CLK(n5735), .C(n5736) );
  CKBD0 U5618 ( .CLK(n5736), .C(n5737) );
  CKBD0 U5619 ( .CLK(n5737), .C(n5738) );
  CKBD0 U5620 ( .CLK(n5738), .C(n5739) );
  CKBD0 U5621 ( .CLK(n5739), .C(n5740) );
  CKBD0 U5622 ( .CLK(n5740), .C(n5741) );
  CKBD0 U5623 ( .CLK(n5741), .C(n5742) );
  CKBD0 U5624 ( .CLK(n5742), .C(n5743) );
  CKBD0 U5625 ( .CLK(n5743), .C(n5744) );
  BUFFD0 U5626 ( .I(n5744), .Z(n5745) );
  CKBD0 U5627 ( .CLK(n5745), .C(n5746) );
  CKBD0 U5628 ( .CLK(n5746), .C(n5747) );
  CKBD0 U5629 ( .CLK(n5747), .C(n5748) );
  CKBD0 U5630 ( .CLK(n5748), .C(n5749) );
  CKBD0 U5631 ( .CLK(n5749), .C(n5750) );
  CKBD0 U5632 ( .CLK(n5750), .C(n5751) );
  CKBD0 U5633 ( .CLK(n5751), .C(n5752) );
  CKBD0 U5634 ( .CLK(n5752), .C(n5753) );
  CKBD0 U5635 ( .CLK(n5753), .C(n5754) );
  CKBD0 U5636 ( .CLK(n5754), .C(n5755) );
  BUFFD0 U5637 ( .I(n5755), .Z(n5756) );
  CKBD0 U5638 ( .CLK(n5756), .C(n5757) );
  CKBD0 U5639 ( .CLK(n5757), .C(n5758) );
  CKBD0 U5640 ( .CLK(n5758), .C(n5759) );
  CKBD0 U5641 ( .CLK(n5759), .C(n5760) );
  CKBD0 U5642 ( .CLK(n5760), .C(n5761) );
  CKBD0 U5643 ( .CLK(n5761), .C(n5762) );
  CKBD0 U5644 ( .CLK(n5762), .C(n5763) );
  CKBD0 U5645 ( .CLK(n5763), .C(n5764) );
  CKBD0 U5646 ( .CLK(n5764), .C(n5765) );
  CKBD0 U5647 ( .CLK(n5765), .C(n5766) );
  BUFFD0 U5648 ( .I(n5766), .Z(n5767) );
  CKBD0 U5649 ( .CLK(n5767), .C(n5768) );
  CKBD0 U5650 ( .CLK(n5768), .C(n5769) );
  CKBD0 U5651 ( .CLK(n5769), .C(n5770) );
  CKBD0 U5652 ( .CLK(n5770), .C(n5771) );
  CKBD0 U5653 ( .CLK(n5771), .C(n5772) );
  CKBD0 U5654 ( .CLK(n5772), .C(n5773) );
  CKBD0 U5655 ( .CLK(n5773), .C(n5774) );
  CKBD0 U5656 ( .CLK(n5774), .C(n5775) );
  CKBD0 U5657 ( .CLK(n5775), .C(n5776) );
  CKBD0 U5658 ( .CLK(n5776), .C(n5777) );
  BUFFD0 U5659 ( .I(n5777), .Z(n5778) );
  CKBD0 U5660 ( .CLK(n5778), .C(n5779) );
  CKBD0 U5661 ( .CLK(n5779), .C(n5780) );
  CKBD0 U5662 ( .CLK(n5780), .C(n5781) );
  CKBD0 U5663 ( .CLK(n5781), .C(n5782) );
  CKBD0 U5664 ( .CLK(n5782), .C(n5783) );
  CKBD0 U5665 ( .CLK(n5783), .C(n5784) );
  CKBD0 U5666 ( .CLK(n5784), .C(n5785) );
  CKBD0 U5667 ( .CLK(n5785), .C(n5786) );
  CKBD0 U5668 ( .CLK(n5786), .C(n5787) );
  BUFFD0 U5669 ( .I(n5787), .Z(n5788) );
  CKBD0 U5670 ( .CLK(n5788), .C(n5789) );
  CKBD0 U5671 ( .CLK(n5789), .C(n5790) );
  CKBD0 U5672 ( .CLK(n5790), .C(n5791) );
  CKBD0 U5673 ( .CLK(n5791), .C(n5792) );
  CKBD0 U5674 ( .CLK(n5792), .C(n5793) );
  CKBD0 U5675 ( .CLK(n5793), .C(n5794) );
  CKBD0 U5676 ( .CLK(n5794), .C(n5795) );
  CKBD0 U5677 ( .CLK(n5795), .C(n5796) );
  CKBD0 U5678 ( .CLK(n5796), .C(n5797) );
  CKBD0 U5679 ( .CLK(n5797), .C(n5798) );
  BUFFD0 U5680 ( .I(n5798), .Z(n5799) );
  CKBD0 U5681 ( .CLK(n5799), .C(n5800) );
  CKBD0 U5682 ( .CLK(n5800), .C(n5801) );
  CKBD0 U5683 ( .CLK(n5801), .C(n5802) );
  CKBD0 U5684 ( .CLK(n5802), .C(n5803) );
  CKBD0 U5685 ( .CLK(n5803), .C(n5804) );
  CKBD0 U5686 ( .CLK(n5804), .C(n5805) );
  BUFFD0 U5687 ( .I(n5805), .Z(n5806) );
  CKBD0 U5688 ( .CLK(n5806), .C(n5807) );
  BUFFD0 U5689 ( .I(n5807), .Z(n5808) );
  CKBD0 U5690 ( .CLK(n5808), .C(n5809) );
  BUFFD0 U5691 ( .I(n5809), .Z(n5810) );
  CKBD0 U5692 ( .CLK(n5810), .C(n5811) );
  BUFFD0 U5693 ( .I(n5811), .Z(n5812) );
  CKBD0 U5694 ( .CLK(n5812), .C(n5813) );
  BUFFD0 U5695 ( .I(n5813), .Z(n5814) );
  CKBD0 U5696 ( .CLK(n5814), .C(n5815) );
  BUFFD0 U5697 ( .I(n5815), .Z(n5816) );
  CKBD0 U5698 ( .CLK(n5816), .C(n5817) );
  BUFFD0 U5699 ( .I(n5817), .Z(n5818) );
  CKBD0 U5700 ( .CLK(n5818), .C(n5819) );
  BUFFD0 U5701 ( .I(n5819), .Z(n5820) );
  BUFFD0 U5702 ( .I(n5822), .Z(n5821) );
  BUFFD0 U5703 ( .I(n5823), .Z(n5822) );
  BUFFD0 U5704 ( .I(n9182), .Z(n5823) );
  CKBD0 U5705 ( .CLK(n2555), .C(n5824) );
  CKBD0 U5706 ( .CLK(n5824), .C(n5825) );
  CKBD0 U5707 ( .CLK(n5825), .C(n5826) );
  BUFFD0 U5708 ( .I(n5826), .Z(n5827) );
  CKBD0 U5709 ( .CLK(n5827), .C(n5828) );
  CKBD0 U5710 ( .CLK(n5828), .C(n5829) );
  CKBD0 U5711 ( .CLK(n5829), .C(n5830) );
  CKBD0 U5712 ( .CLK(n5830), .C(n5831) );
  CKBD0 U5713 ( .CLK(n5831), .C(n5832) );
  CKBD0 U5714 ( .CLK(n5832), .C(n5833) );
  CKBD0 U5715 ( .CLK(n5833), .C(n5834) );
  CKBD0 U5716 ( .CLK(n5834), .C(n5835) );
  CKBD0 U5717 ( .CLK(n5835), .C(n5836) );
  CKBD0 U5718 ( .CLK(n5836), .C(n5837) );
  BUFFD0 U5719 ( .I(n5837), .Z(n5838) );
  CKBD0 U5720 ( .CLK(n5838), .C(n5839) );
  CKBD0 U5721 ( .CLK(n5839), .C(n5840) );
  CKBD0 U5722 ( .CLK(n5840), .C(n5841) );
  CKBD0 U5723 ( .CLK(n5841), .C(n5842) );
  CKBD0 U5724 ( .CLK(n5842), .C(n5843) );
  CKBD0 U5725 ( .CLK(n5843), .C(n5844) );
  CKBD0 U5726 ( .CLK(n5844), .C(n5845) );
  CKBD0 U5727 ( .CLK(n5845), .C(n5846) );
  CKBD0 U5728 ( .CLK(n5846), .C(n5847) );
  BUFFD0 U5729 ( .I(n5847), .Z(n5848) );
  CKBD0 U5730 ( .CLK(n5848), .C(n5849) );
  CKBD0 U5731 ( .CLK(n5849), .C(n5850) );
  CKBD0 U5732 ( .CLK(n5850), .C(n5851) );
  CKBD0 U5733 ( .CLK(n5851), .C(n5852) );
  CKBD0 U5734 ( .CLK(n5852), .C(n5853) );
  CKBD0 U5735 ( .CLK(n5853), .C(n5854) );
  CKBD0 U5736 ( .CLK(n5854), .C(n5855) );
  CKBD0 U5737 ( .CLK(n5855), .C(n5856) );
  CKBD0 U5738 ( .CLK(n5856), .C(n5857) );
  CKBD0 U5739 ( .CLK(n5857), .C(n5858) );
  BUFFD0 U5740 ( .I(n5858), .Z(n5859) );
  CKBD0 U5741 ( .CLK(n5859), .C(n5860) );
  CKBD0 U5742 ( .CLK(n5860), .C(n5861) );
  CKBD0 U5743 ( .CLK(n5861), .C(n5862) );
  CKBD0 U5744 ( .CLK(n5862), .C(n5863) );
  CKBD0 U5745 ( .CLK(n5863), .C(n5864) );
  CKBD0 U5746 ( .CLK(n5864), .C(n5865) );
  CKBD0 U5747 ( .CLK(n5865), .C(n5866) );
  CKBD0 U5748 ( .CLK(n5866), .C(n5867) );
  CKBD0 U5749 ( .CLK(n5867), .C(n5868) );
  CKBD0 U5750 ( .CLK(n5868), .C(n5869) );
  BUFFD0 U5751 ( .I(n5869), .Z(n5870) );
  CKBD0 U5752 ( .CLK(n5870), .C(n5871) );
  CKBD0 U5753 ( .CLK(n5871), .C(n5872) );
  CKBD0 U5754 ( .CLK(n5872), .C(n5873) );
  CKBD0 U5755 ( .CLK(n5873), .C(n5874) );
  CKBD0 U5756 ( .CLK(n5874), .C(n5875) );
  CKBD0 U5757 ( .CLK(n5875), .C(n5876) );
  CKBD0 U5758 ( .CLK(n5876), .C(n5877) );
  CKBD0 U5759 ( .CLK(n5877), .C(n5878) );
  CKBD0 U5760 ( .CLK(n5878), .C(n5879) );
  CKBD0 U5761 ( .CLK(n5879), .C(n5880) );
  BUFFD0 U5762 ( .I(n5880), .Z(n5881) );
  CKBD0 U5763 ( .CLK(n5881), .C(n5882) );
  CKBD0 U5764 ( .CLK(n5882), .C(n5883) );
  CKBD0 U5765 ( .CLK(n5883), .C(n5884) );
  CKBD0 U5766 ( .CLK(n5884), .C(n5885) );
  CKBD0 U5767 ( .CLK(n5885), .C(n5886) );
  CKBD0 U5768 ( .CLK(n5886), .C(n5887) );
  CKBD0 U5769 ( .CLK(n5887), .C(n5888) );
  CKBD0 U5770 ( .CLK(n5888), .C(n5889) );
  CKBD0 U5771 ( .CLK(n5889), .C(n5890) );
  CKBD0 U5772 ( .CLK(n5890), .C(n5891) );
  BUFFD0 U5773 ( .I(n5891), .Z(n5892) );
  CKBD0 U5774 ( .CLK(n5892), .C(n5893) );
  CKBD0 U5775 ( .CLK(n5893), .C(n5894) );
  CKBD0 U5776 ( .CLK(n5894), .C(n5895) );
  CKBD0 U5777 ( .CLK(n5895), .C(n5896) );
  CKBD0 U5778 ( .CLK(n5896), .C(n5897) );
  CKBD0 U5779 ( .CLK(n5897), .C(n5898) );
  CKBD0 U5780 ( .CLK(n5898), .C(n5899) );
  CKBD0 U5781 ( .CLK(n5899), .C(n5900) );
  CKBD0 U5782 ( .CLK(n5900), .C(n5901) );
  CKBD0 U5783 ( .CLK(n5901), .C(n5902) );
  BUFFD0 U5784 ( .I(n5902), .Z(n5903) );
  CKBD0 U5785 ( .CLK(n5903), .C(n5904) );
  CKBD0 U5786 ( .CLK(n5904), .C(n5905) );
  CKBD0 U5787 ( .CLK(n5905), .C(n5906) );
  CKBD0 U5788 ( .CLK(n5906), .C(n5907) );
  CKBD0 U5789 ( .CLK(n5907), .C(n5908) );
  CKBD0 U5790 ( .CLK(n5908), .C(n5909) );
  CKBD0 U5791 ( .CLK(n5909), .C(n5910) );
  CKBD0 U5792 ( .CLK(n5910), .C(n5911) );
  CKBD0 U5793 ( .CLK(n5911), .C(n5912) );
  CKBD0 U5794 ( .CLK(n5912), .C(n5913) );
  BUFFD0 U5795 ( .I(n5913), .Z(n5914) );
  CKBD0 U5796 ( .CLK(n5914), .C(n5915) );
  CKBD0 U5797 ( .CLK(n5915), .C(n5916) );
  CKBD0 U5798 ( .CLK(n5916), .C(n5917) );
  CKBD0 U5799 ( .CLK(n5917), .C(n5918) );
  CKBD0 U5800 ( .CLK(n5918), .C(n5919) );
  CKBD0 U5801 ( .CLK(n5919), .C(n5920) );
  CKBD0 U5802 ( .CLK(n5920), .C(n5921) );
  CKBD0 U5803 ( .CLK(n5921), .C(n5922) );
  CKBD0 U5804 ( .CLK(n5922), .C(n5923) );
  BUFFD0 U5805 ( .I(n5923), .Z(n5924) );
  CKBD0 U5806 ( .CLK(n5924), .C(n5925) );
  CKBD0 U5807 ( .CLK(n5925), .C(n5926) );
  CKBD0 U5808 ( .CLK(n5926), .C(n5927) );
  CKBD0 U5809 ( .CLK(n5927), .C(n5928) );
  CKBD0 U5810 ( .CLK(n5928), .C(n5929) );
  CKBD0 U5811 ( .CLK(n5929), .C(n5930) );
  CKBD0 U5812 ( .CLK(n5930), .C(n5931) );
  CKBD0 U5813 ( .CLK(n5931), .C(n5932) );
  CKBD0 U5814 ( .CLK(n5932), .C(n5933) );
  CKBD0 U5815 ( .CLK(n5933), .C(n5934) );
  BUFFD0 U5816 ( .I(n5934), .Z(n5935) );
  CKBD0 U5817 ( .CLK(n5935), .C(n5936) );
  CKBD0 U5818 ( .CLK(n5936), .C(n5937) );
  CKBD0 U5819 ( .CLK(n5937), .C(n5938) );
  CKBD0 U5820 ( .CLK(n5938), .C(n5939) );
  CKBD0 U5821 ( .CLK(n5939), .C(n5940) );
  CKBD0 U5822 ( .CLK(n5940), .C(n5941) );
  BUFFD0 U5823 ( .I(n5941), .Z(n5942) );
  CKBD0 U5824 ( .CLK(n5942), .C(n5943) );
  BUFFD0 U5825 ( .I(n5943), .Z(n5944) );
  CKBD0 U5826 ( .CLK(n5944), .C(n5945) );
  BUFFD0 U5827 ( .I(n5945), .Z(n5946) );
  CKBD0 U5828 ( .CLK(n5946), .C(n5947) );
  BUFFD0 U5829 ( .I(n5947), .Z(n5948) );
  CKBD0 U5830 ( .CLK(n5948), .C(n5949) );
  BUFFD0 U5831 ( .I(n5949), .Z(n5950) );
  CKBD0 U5832 ( .CLK(n5950), .C(n5951) );
  BUFFD0 U5833 ( .I(n5951), .Z(n5952) );
  CKBD0 U5834 ( .CLK(n5952), .C(n5953) );
  BUFFD0 U5835 ( .I(n5953), .Z(n5954) );
  CKBD0 U5836 ( .CLK(n5954), .C(n5955) );
  BUFFD0 U5837 ( .I(n5955), .Z(n5956) );
  BUFFD0 U5838 ( .I(Decoder[6]), .Z(n5957) );
  BUFFD0 U5839 ( .I(n5959), .Z(n5958) );
  BUFFD0 U5840 ( .I(n5960), .Z(n5959) );
  BUFFD0 U5841 ( .I(n9183), .Z(n5960) );
  CKBD0 U5842 ( .CLK(n933), .C(n5961) );
  CKBD0 U5843 ( .CLK(n5961), .C(n5962) );
  CKBD0 U5844 ( .CLK(n5962), .C(n5963) );
  BUFFD0 U5845 ( .I(n5963), .Z(n5964) );
  CKBD0 U5846 ( .CLK(n5964), .C(n5965) );
  CKBD0 U5847 ( .CLK(n5965), .C(n5966) );
  CKBD0 U5848 ( .CLK(n5966), .C(n5967) );
  CKBD0 U5849 ( .CLK(n5967), .C(n5968) );
  CKBD0 U5850 ( .CLK(n5968), .C(n5969) );
  CKBD0 U5851 ( .CLK(n5969), .C(n5970) );
  CKBD0 U5852 ( .CLK(n5970), .C(n5971) );
  CKBD0 U5853 ( .CLK(n5971), .C(n5972) );
  CKBD0 U5854 ( .CLK(n5972), .C(n5973) );
  CKBD0 U5855 ( .CLK(n5973), .C(n5974) );
  BUFFD0 U5856 ( .I(n5974), .Z(n5975) );
  CKBD0 U5857 ( .CLK(n5975), .C(n5976) );
  CKBD0 U5858 ( .CLK(n5976), .C(n5977) );
  CKBD0 U5859 ( .CLK(n5977), .C(n5978) );
  CKBD0 U5860 ( .CLK(n5978), .C(n5979) );
  CKBD0 U5861 ( .CLK(n5979), .C(n5980) );
  CKBD0 U5862 ( .CLK(n5980), .C(n5981) );
  CKBD0 U5863 ( .CLK(n5981), .C(n5982) );
  CKBD0 U5864 ( .CLK(n5982), .C(n5983) );
  CKBD0 U5865 ( .CLK(n5983), .C(n5984) );
  BUFFD0 U5866 ( .I(n5984), .Z(n5985) );
  CKBD0 U5867 ( .CLK(n5985), .C(n5986) );
  CKBD0 U5868 ( .CLK(n5986), .C(n5987) );
  CKBD0 U5869 ( .CLK(n5987), .C(n5988) );
  CKBD0 U5870 ( .CLK(n5988), .C(n5989) );
  CKBD0 U5871 ( .CLK(n5989), .C(n5990) );
  CKBD0 U5872 ( .CLK(n5990), .C(n5991) );
  CKBD0 U5873 ( .CLK(n5991), .C(n5992) );
  CKBD0 U5874 ( .CLK(n5992), .C(n5993) );
  CKBD0 U5875 ( .CLK(n5993), .C(n5994) );
  CKBD0 U5876 ( .CLK(n5994), .C(n5995) );
  BUFFD0 U5877 ( .I(n5995), .Z(n5996) );
  CKBD0 U5878 ( .CLK(n5996), .C(n5997) );
  CKBD0 U5879 ( .CLK(n5997), .C(n5998) );
  CKBD0 U5880 ( .CLK(n5998), .C(n5999) );
  CKBD0 U5881 ( .CLK(n5999), .C(n6000) );
  CKBD0 U5882 ( .CLK(n6000), .C(n6001) );
  CKBD0 U5883 ( .CLK(n6001), .C(n6002) );
  CKBD0 U5884 ( .CLK(n6002), .C(n6003) );
  CKBD0 U5885 ( .CLK(n6003), .C(n6004) );
  CKBD0 U5886 ( .CLK(n6004), .C(n6005) );
  CKBD0 U5887 ( .CLK(n6005), .C(n6006) );
  BUFFD0 U5888 ( .I(n6006), .Z(n6007) );
  CKBD0 U5889 ( .CLK(n6007), .C(n6008) );
  CKBD0 U5890 ( .CLK(n6008), .C(n6009) );
  CKBD0 U5891 ( .CLK(n6009), .C(n6010) );
  CKBD0 U5892 ( .CLK(n6010), .C(n6011) );
  CKBD0 U5893 ( .CLK(n6011), .C(n6012) );
  CKBD0 U5894 ( .CLK(n6012), .C(n6013) );
  CKBD0 U5895 ( .CLK(n6013), .C(n6014) );
  CKBD0 U5896 ( .CLK(n6014), .C(n6015) );
  CKBD0 U5897 ( .CLK(n6015), .C(n6016) );
  CKBD0 U5898 ( .CLK(n6016), .C(n6017) );
  BUFFD0 U5899 ( .I(n6017), .Z(n6018) );
  CKBD0 U5900 ( .CLK(n6018), .C(n6019) );
  CKBD0 U5901 ( .CLK(n6019), .C(n6020) );
  CKBD0 U5902 ( .CLK(n6020), .C(n6021) );
  CKBD0 U5903 ( .CLK(n6021), .C(n6022) );
  CKBD0 U5904 ( .CLK(n6022), .C(n6023) );
  CKBD0 U5905 ( .CLK(n6023), .C(n6024) );
  CKBD0 U5906 ( .CLK(n6024), .C(n6025) );
  CKBD0 U5907 ( .CLK(n6025), .C(n6026) );
  CKBD0 U5908 ( .CLK(n6026), .C(n6027) );
  CKBD0 U5909 ( .CLK(n6027), .C(n6028) );
  BUFFD0 U5910 ( .I(n6028), .Z(n6029) );
  CKBD0 U5911 ( .CLK(n6029), .C(n6030) );
  CKBD0 U5912 ( .CLK(n6030), .C(n6031) );
  CKBD0 U5913 ( .CLK(n6031), .C(n6032) );
  CKBD0 U5914 ( .CLK(n6032), .C(n6033) );
  CKBD0 U5915 ( .CLK(n6033), .C(n6034) );
  CKBD0 U5916 ( .CLK(n6034), .C(n6035) );
  CKBD0 U5917 ( .CLK(n6035), .C(n6036) );
  CKBD0 U5918 ( .CLK(n6036), .C(n6037) );
  CKBD0 U5919 ( .CLK(n6037), .C(n6038) );
  CKBD0 U5920 ( .CLK(n6038), .C(n6039) );
  BUFFD0 U5921 ( .I(n6039), .Z(n6040) );
  CKBD0 U5922 ( .CLK(n6040), .C(n6041) );
  CKBD0 U5923 ( .CLK(n6041), .C(n6042) );
  CKBD0 U5924 ( .CLK(n6042), .C(n6043) );
  CKBD0 U5925 ( .CLK(n6043), .C(n6044) );
  CKBD0 U5926 ( .CLK(n6044), .C(n6045) );
  CKBD0 U5927 ( .CLK(n6045), .C(n6046) );
  CKBD0 U5928 ( .CLK(n6046), .C(n6047) );
  CKBD0 U5929 ( .CLK(n6047), .C(n6048) );
  CKBD0 U5930 ( .CLK(n6048), .C(n6049) );
  BUFFD0 U5931 ( .I(n6049), .Z(n6050) );
  CKBD0 U5932 ( .CLK(n6050), .C(n6051) );
  CKBD0 U5933 ( .CLK(n6051), .C(n6052) );
  CKBD0 U5934 ( .CLK(n6052), .C(n6053) );
  CKBD0 U5935 ( .CLK(n6053), .C(n6054) );
  CKBD0 U5936 ( .CLK(n6054), .C(n6055) );
  CKBD0 U5937 ( .CLK(n6055), .C(n6056) );
  CKBD0 U5938 ( .CLK(n6056), .C(n6057) );
  CKBD0 U5939 ( .CLK(n6057), .C(n6058) );
  CKBD0 U5940 ( .CLK(n6058), .C(n6059) );
  CKBD0 U5941 ( .CLK(n6059), .C(n6060) );
  BUFFD0 U5942 ( .I(n6060), .Z(n6061) );
  CKBD0 U5943 ( .CLK(n6061), .C(n6062) );
  CKBD0 U5944 ( .CLK(n6062), .C(n6063) );
  CKBD0 U5945 ( .CLK(n6063), .C(n6064) );
  CKBD0 U5946 ( .CLK(n6064), .C(n6065) );
  CKBD0 U5947 ( .CLK(n6065), .C(n6066) );
  CKBD0 U5948 ( .CLK(n6066), .C(n6067) );
  CKBD0 U5949 ( .CLK(n6067), .C(n6068) );
  CKBD0 U5950 ( .CLK(n6068), .C(n6069) );
  CKBD0 U5951 ( .CLK(n6069), .C(n6070) );
  CKBD0 U5952 ( .CLK(n6070), .C(n6071) );
  BUFFD0 U5953 ( .I(n6071), .Z(n6072) );
  CKBD0 U5954 ( .CLK(n6072), .C(n6073) );
  CKBD0 U5955 ( .CLK(n6073), .C(n6074) );
  CKBD0 U5956 ( .CLK(n6074), .C(n6075) );
  CKBD0 U5957 ( .CLK(n6075), .C(n6076) );
  CKBD0 U5958 ( .CLK(n6076), .C(n6077) );
  CKBD0 U5959 ( .CLK(n6077), .C(n6078) );
  BUFFD0 U5960 ( .I(n6078), .Z(n6079) );
  CKBD0 U5961 ( .CLK(n6079), .C(n6080) );
  BUFFD0 U5962 ( .I(n6080), .Z(n6081) );
  CKBD0 U5963 ( .CLK(n6081), .C(n6082) );
  BUFFD0 U5964 ( .I(n6082), .Z(n6083) );
  CKBD0 U5965 ( .CLK(n6083), .C(n6084) );
  BUFFD0 U5966 ( .I(n6084), .Z(n6085) );
  CKBD0 U5967 ( .CLK(n6085), .C(n6086) );
  BUFFD0 U5968 ( .I(n6086), .Z(n6087) );
  CKBD0 U5969 ( .CLK(n6087), .C(n6088) );
  BUFFD0 U5970 ( .I(n6088), .Z(n6089) );
  CKBD0 U5971 ( .CLK(n6089), .C(n6090) );
  BUFFD0 U5972 ( .I(n6090), .Z(n6091) );
  CKBD0 U5973 ( .CLK(n6091), .C(n6092) );
  BUFFD0 U5974 ( .I(n6092), .Z(n6093) );
  BUFFD0 U5975 ( .I(n9184), .Z(n6094) );
  BUFFD0 U5976 ( .I(n6096), .Z(n6095) );
  BUFFD0 U5977 ( .I(n6097), .Z(n6096) );
  BUFFD0 U5978 ( .I(Decoder[5]), .Z(n6097) );
  CKBD0 U5979 ( .CLK(n931), .C(n6098) );
  CKBD0 U5980 ( .CLK(n6098), .C(n6099) );
  CKBD0 U5981 ( .CLK(n6099), .C(n6100) );
  BUFFD0 U5982 ( .I(n6100), .Z(n6101) );
  CKBD0 U5983 ( .CLK(n6101), .C(n6102) );
  CKBD0 U5984 ( .CLK(n6102), .C(n6103) );
  CKBD0 U5985 ( .CLK(n6103), .C(n6104) );
  CKBD0 U5986 ( .CLK(n6104), .C(n6105) );
  CKBD0 U5987 ( .CLK(n6105), .C(n6106) );
  CKBD0 U5988 ( .CLK(n6106), .C(n6107) );
  CKBD0 U5989 ( .CLK(n6107), .C(n6108) );
  CKBD0 U5990 ( .CLK(n6108), .C(n6109) );
  CKBD0 U5991 ( .CLK(n6109), .C(n6110) );
  CKBD0 U5992 ( .CLK(n6110), .C(n6111) );
  BUFFD0 U5993 ( .I(n6111), .Z(n6112) );
  CKBD0 U5994 ( .CLK(n6112), .C(n6113) );
  CKBD0 U5995 ( .CLK(n6113), .C(n6114) );
  CKBD0 U5996 ( .CLK(n6114), .C(n6115) );
  CKBD0 U5997 ( .CLK(n6115), .C(n6116) );
  CKBD0 U5998 ( .CLK(n6116), .C(n6117) );
  CKBD0 U5999 ( .CLK(n6117), .C(n6118) );
  CKBD0 U6000 ( .CLK(n6118), .C(n6119) );
  CKBD0 U6001 ( .CLK(n6119), .C(n6120) );
  CKBD0 U6002 ( .CLK(n6120), .C(n6121) );
  BUFFD0 U6003 ( .I(n6121), .Z(n6122) );
  CKBD0 U6004 ( .CLK(n6122), .C(n6123) );
  CKBD0 U6005 ( .CLK(n6123), .C(n6124) );
  CKBD0 U6006 ( .CLK(n6124), .C(n6125) );
  CKBD0 U6007 ( .CLK(n6125), .C(n6126) );
  CKBD0 U6008 ( .CLK(n6126), .C(n6127) );
  CKBD0 U6009 ( .CLK(n6127), .C(n6128) );
  CKBD0 U6010 ( .CLK(n6128), .C(n6129) );
  CKBD0 U6011 ( .CLK(n6129), .C(n6130) );
  CKBD0 U6012 ( .CLK(n6130), .C(n6131) );
  CKBD0 U6013 ( .CLK(n6131), .C(n6132) );
  BUFFD0 U6014 ( .I(n6132), .Z(n6133) );
  CKBD0 U6015 ( .CLK(n6133), .C(n6134) );
  CKBD0 U6016 ( .CLK(n6134), .C(n6135) );
  CKBD0 U6017 ( .CLK(n6135), .C(n6136) );
  CKBD0 U6018 ( .CLK(n6136), .C(n6137) );
  CKBD0 U6019 ( .CLK(n6137), .C(n6138) );
  CKBD0 U6020 ( .CLK(n6138), .C(n6139) );
  CKBD0 U6021 ( .CLK(n6139), .C(n6140) );
  CKBD0 U6022 ( .CLK(n6140), .C(n6141) );
  CKBD0 U6023 ( .CLK(n6141), .C(n6142) );
  CKBD0 U6024 ( .CLK(n6142), .C(n6143) );
  BUFFD0 U6025 ( .I(n6143), .Z(n6144) );
  CKBD0 U6026 ( .CLK(n6144), .C(n6145) );
  CKBD0 U6027 ( .CLK(n6145), .C(n6146) );
  CKBD0 U6028 ( .CLK(n6146), .C(n6147) );
  CKBD0 U6029 ( .CLK(n6147), .C(n6148) );
  CKBD0 U6030 ( .CLK(n6148), .C(n6149) );
  CKBD0 U6031 ( .CLK(n6149), .C(n6150) );
  CKBD0 U6032 ( .CLK(n6150), .C(n6151) );
  CKBD0 U6033 ( .CLK(n6151), .C(n6152) );
  CKBD0 U6034 ( .CLK(n6152), .C(n6153) );
  CKBD0 U6035 ( .CLK(n6153), .C(n6154) );
  BUFFD0 U6036 ( .I(n6154), .Z(n6155) );
  CKBD0 U6037 ( .CLK(n6155), .C(n6156) );
  CKBD0 U6038 ( .CLK(n6156), .C(n6157) );
  CKBD0 U6039 ( .CLK(n6157), .C(n6158) );
  CKBD0 U6040 ( .CLK(n6158), .C(n6159) );
  CKBD0 U6041 ( .CLK(n6159), .C(n6160) );
  CKBD0 U6042 ( .CLK(n6160), .C(n6161) );
  CKBD0 U6043 ( .CLK(n6161), .C(n6162) );
  CKBD0 U6044 ( .CLK(n6162), .C(n6163) );
  CKBD0 U6045 ( .CLK(n6163), .C(n6164) );
  CKBD0 U6046 ( .CLK(n6164), .C(n6165) );
  BUFFD0 U6047 ( .I(n6165), .Z(n6166) );
  CKBD0 U6048 ( .CLK(n6166), .C(n6167) );
  CKBD0 U6049 ( .CLK(n6167), .C(n6168) );
  CKBD0 U6050 ( .CLK(n6168), .C(n6169) );
  CKBD0 U6051 ( .CLK(n6169), .C(n6170) );
  CKBD0 U6052 ( .CLK(n6170), .C(n6171) );
  CKBD0 U6053 ( .CLK(n6171), .C(n6172) );
  CKBD0 U6054 ( .CLK(n6172), .C(n6173) );
  CKBD0 U6055 ( .CLK(n6173), .C(n6174) );
  CKBD0 U6056 ( .CLK(n6174), .C(n6175) );
  CKBD0 U6057 ( .CLK(n6175), .C(n6176) );
  BUFFD0 U6058 ( .I(n6176), .Z(n6177) );
  CKBD0 U6059 ( .CLK(n6177), .C(n6178) );
  CKBD0 U6060 ( .CLK(n6178), .C(n6179) );
  CKBD0 U6061 ( .CLK(n6179), .C(n6180) );
  CKBD0 U6062 ( .CLK(n6180), .C(n6181) );
  CKBD0 U6063 ( .CLK(n6181), .C(n6182) );
  CKBD0 U6064 ( .CLK(n6182), .C(n6183) );
  CKBD0 U6065 ( .CLK(n6183), .C(n6184) );
  CKBD0 U6066 ( .CLK(n6184), .C(n6185) );
  CKBD0 U6067 ( .CLK(n6185), .C(n6186) );
  CKBD0 U6068 ( .CLK(n6186), .C(n6187) );
  BUFFD0 U6069 ( .I(n6187), .Z(n6188) );
  CKBD0 U6070 ( .CLK(n6188), .C(n6189) );
  CKBD0 U6071 ( .CLK(n6189), .C(n6190) );
  CKBD0 U6072 ( .CLK(n6190), .C(n6191) );
  CKBD0 U6073 ( .CLK(n6191), .C(n6192) );
  CKBD0 U6074 ( .CLK(n6192), .C(n6193) );
  CKBD0 U6075 ( .CLK(n6193), .C(n6194) );
  CKBD0 U6076 ( .CLK(n6194), .C(n6195) );
  CKBD0 U6077 ( .CLK(n6195), .C(n6196) );
  CKBD0 U6078 ( .CLK(n6196), .C(n6197) );
  BUFFD0 U6079 ( .I(n6197), .Z(n6198) );
  CKBD0 U6080 ( .CLK(n6198), .C(n6199) );
  CKBD0 U6081 ( .CLK(n6199), .C(n6200) );
  CKBD0 U6082 ( .CLK(n6200), .C(n6201) );
  CKBD0 U6083 ( .CLK(n6201), .C(n6202) );
  CKBD0 U6084 ( .CLK(n6202), .C(n6203) );
  CKBD0 U6085 ( .CLK(n6203), .C(n6204) );
  CKBD0 U6086 ( .CLK(n6204), .C(n6205) );
  CKBD0 U6087 ( .CLK(n6205), .C(n6206) );
  CKBD0 U6088 ( .CLK(n6206), .C(n6207) );
  CKBD0 U6089 ( .CLK(n6207), .C(n6208) );
  BUFFD0 U6090 ( .I(n6208), .Z(n6209) );
  CKBD0 U6091 ( .CLK(n6209), .C(n6210) );
  CKBD0 U6092 ( .CLK(n6210), .C(n6211) );
  CKBD0 U6093 ( .CLK(n6211), .C(n6212) );
  CKBD0 U6094 ( .CLK(n6212), .C(n6213) );
  CKBD0 U6095 ( .CLK(n6213), .C(n6214) );
  CKBD0 U6096 ( .CLK(n6214), .C(n6215) );
  BUFFD0 U6097 ( .I(n6215), .Z(n6216) );
  CKBD0 U6098 ( .CLK(n6216), .C(n6217) );
  BUFFD0 U6099 ( .I(n6217), .Z(n6218) );
  CKBD0 U6100 ( .CLK(n6218), .C(n6219) );
  BUFFD0 U6101 ( .I(n6219), .Z(n6220) );
  CKBD0 U6102 ( .CLK(n6220), .C(n6221) );
  BUFFD0 U6103 ( .I(n6221), .Z(n6222) );
  CKBD0 U6104 ( .CLK(n6222), .C(n6223) );
  BUFFD0 U6105 ( .I(n6223), .Z(n6224) );
  CKBD0 U6106 ( .CLK(n6224), .C(n6225) );
  BUFFD0 U6107 ( .I(n6225), .Z(n6226) );
  CKBD0 U6108 ( .CLK(n6226), .C(n6227) );
  BUFFD0 U6109 ( .I(n6227), .Z(n6228) );
  CKBD0 U6110 ( .CLK(n6228), .C(n6229) );
  BUFFD0 U6111 ( .I(n6229), .Z(n6230) );
  BUFFD0 U6112 ( .I(n9185), .Z(n6231) );
  BUFFD0 U6113 ( .I(n6233), .Z(n6232) );
  BUFFD0 U6114 ( .I(n6234), .Z(n6233) );
  BUFFD0 U6115 ( .I(Decoder[4]), .Z(n6234) );
  CKBD0 U6116 ( .CLK(n929), .C(n6235) );
  CKBD0 U6117 ( .CLK(n6235), .C(n6236) );
  CKBD0 U6118 ( .CLK(n6236), .C(n6237) );
  BUFFD0 U6119 ( .I(n6237), .Z(n6238) );
  CKBD0 U6120 ( .CLK(n6238), .C(n6239) );
  CKBD0 U6121 ( .CLK(n6239), .C(n6240) );
  CKBD0 U6122 ( .CLK(n6240), .C(n6241) );
  CKBD0 U6123 ( .CLK(n6241), .C(n6242) );
  CKBD0 U6124 ( .CLK(n6242), .C(n6243) );
  CKBD0 U6125 ( .CLK(n6243), .C(n6244) );
  CKBD0 U6126 ( .CLK(n6244), .C(n6245) );
  CKBD0 U6127 ( .CLK(n6245), .C(n6246) );
  CKBD0 U6128 ( .CLK(n6246), .C(n6247) );
  CKBD0 U6129 ( .CLK(n6247), .C(n6248) );
  BUFFD0 U6130 ( .I(n6248), .Z(n6249) );
  CKBD0 U6131 ( .CLK(n6249), .C(n6250) );
  CKBD0 U6132 ( .CLK(n6250), .C(n6251) );
  CKBD0 U6133 ( .CLK(n6251), .C(n6252) );
  CKBD0 U6134 ( .CLK(n6252), .C(n6253) );
  CKBD0 U6135 ( .CLK(n6253), .C(n6254) );
  CKBD0 U6136 ( .CLK(n6254), .C(n6255) );
  CKBD0 U6137 ( .CLK(n6255), .C(n6256) );
  CKBD0 U6138 ( .CLK(n6256), .C(n6257) );
  CKBD0 U6139 ( .CLK(n6257), .C(n6258) );
  CKBD0 U6140 ( .CLK(n6258), .C(n6259) );
  BUFFD0 U6141 ( .I(n6259), .Z(n6260) );
  CKBD0 U6142 ( .CLK(n6260), .C(n6261) );
  CKBD0 U6143 ( .CLK(n6261), .C(n6262) );
  CKBD0 U6144 ( .CLK(n6262), .C(n6263) );
  CKBD0 U6145 ( .CLK(n6263), .C(n6264) );
  CKBD0 U6146 ( .CLK(n6264), .C(n6265) );
  CKBD0 U6147 ( .CLK(n6265), .C(n6266) );
  CKBD0 U6148 ( .CLK(n6266), .C(n6267) );
  CKBD0 U6149 ( .CLK(n6267), .C(n6268) );
  CKBD0 U6150 ( .CLK(n6268), .C(n6269) );
  BUFFD0 U6151 ( .I(n6269), .Z(n6270) );
  CKBD0 U6152 ( .CLK(n6270), .C(n6271) );
  CKBD0 U6153 ( .CLK(n6271), .C(n6272) );
  CKBD0 U6154 ( .CLK(n6272), .C(n6273) );
  CKBD0 U6155 ( .CLK(n6273), .C(n6274) );
  CKBD0 U6156 ( .CLK(n6274), .C(n6275) );
  CKBD0 U6157 ( .CLK(n6275), .C(n6276) );
  CKBD0 U6158 ( .CLK(n6276), .C(n6277) );
  CKBD0 U6159 ( .CLK(n6277), .C(n6278) );
  CKBD0 U6160 ( .CLK(n6278), .C(n6279) );
  CKBD0 U6161 ( .CLK(n6279), .C(n6280) );
  BUFFD0 U6162 ( .I(n6280), .Z(n6281) );
  CKBD0 U6163 ( .CLK(n6281), .C(n6282) );
  CKBD0 U6164 ( .CLK(n6282), .C(n6283) );
  CKBD0 U6165 ( .CLK(n6283), .C(n6284) );
  CKBD0 U6166 ( .CLK(n6284), .C(n6285) );
  CKBD0 U6167 ( .CLK(n6285), .C(n6286) );
  CKBD0 U6168 ( .CLK(n6286), .C(n6287) );
  CKBD0 U6169 ( .CLK(n6287), .C(n6288) );
  CKBD0 U6170 ( .CLK(n6288), .C(n6289) );
  CKBD0 U6171 ( .CLK(n6289), .C(n6290) );
  CKBD0 U6172 ( .CLK(n6290), .C(n6291) );
  BUFFD0 U6173 ( .I(n6291), .Z(n6292) );
  CKBD0 U6174 ( .CLK(n6292), .C(n6293) );
  CKBD0 U6175 ( .CLK(n6293), .C(n6294) );
  CKBD0 U6176 ( .CLK(n6294), .C(n6295) );
  CKBD0 U6177 ( .CLK(n6295), .C(n6296) );
  CKBD0 U6178 ( .CLK(n6296), .C(n6297) );
  CKBD0 U6179 ( .CLK(n6297), .C(n6298) );
  CKBD0 U6180 ( .CLK(n6298), .C(n6299) );
  CKBD0 U6181 ( .CLK(n6299), .C(n6300) );
  CKBD0 U6182 ( .CLK(n6300), .C(n6301) );
  CKBD0 U6183 ( .CLK(n6301), .C(n6302) );
  BUFFD0 U6184 ( .I(n6302), .Z(n6303) );
  CKBD0 U6185 ( .CLK(n6303), .C(n6304) );
  CKBD0 U6186 ( .CLK(n6304), .C(n6305) );
  CKBD0 U6187 ( .CLK(n6305), .C(n6306) );
  CKBD0 U6188 ( .CLK(n6306), .C(n6307) );
  CKBD0 U6189 ( .CLK(n6307), .C(n6308) );
  CKBD0 U6190 ( .CLK(n6308), .C(n6309) );
  CKBD0 U6191 ( .CLK(n6309), .C(n6310) );
  CKBD0 U6192 ( .CLK(n6310), .C(n6311) );
  CKBD0 U6193 ( .CLK(n6311), .C(n6312) );
  CKBD0 U6194 ( .CLK(n6312), .C(n6313) );
  BUFFD0 U6195 ( .I(n6313), .Z(n6314) );
  CKBD0 U6196 ( .CLK(n6314), .C(n6315) );
  CKBD0 U6197 ( .CLK(n6315), .C(n6316) );
  CKBD0 U6198 ( .CLK(n6316), .C(n6317) );
  CKBD0 U6199 ( .CLK(n6317), .C(n6318) );
  CKBD0 U6200 ( .CLK(n6318), .C(n6319) );
  CKBD0 U6201 ( .CLK(n6319), .C(n6320) );
  CKBD0 U6202 ( .CLK(n6320), .C(n6321) );
  CKBD0 U6203 ( .CLK(n6321), .C(n6322) );
  CKBD0 U6204 ( .CLK(n6322), .C(n6323) );
  BUFFD0 U6205 ( .I(n6323), .Z(n6324) );
  CKBD0 U6206 ( .CLK(n6324), .C(n6325) );
  CKBD0 U6207 ( .CLK(n6325), .C(n6326) );
  CKBD0 U6208 ( .CLK(n6326), .C(n6327) );
  CKBD0 U6209 ( .CLK(n6327), .C(n6328) );
  CKBD0 U6210 ( .CLK(n6328), .C(n6329) );
  CKBD0 U6211 ( .CLK(n6329), .C(n6330) );
  CKBD0 U6212 ( .CLK(n6330), .C(n6331) );
  CKBD0 U6213 ( .CLK(n6331), .C(n6332) );
  CKBD0 U6214 ( .CLK(n6332), .C(n6333) );
  CKBD0 U6215 ( .CLK(n6333), .C(n6334) );
  CKBD0 U6216 ( .CLK(n6334), .C(n6335) );
  BUFFD0 U6217 ( .I(n6335), .Z(n6336) );
  CKBD0 U6218 ( .CLK(n6336), .C(n6337) );
  CKBD0 U6219 ( .CLK(n6337), .C(n6338) );
  CKBD0 U6220 ( .CLK(n6338), .C(n6339) );
  CKBD0 U6221 ( .CLK(n6339), .C(n6340) );
  CKBD0 U6222 ( .CLK(n6340), .C(n6341) );
  CKBD0 U6223 ( .CLK(n6341), .C(n6342) );
  CKBD0 U6224 ( .CLK(n6342), .C(n6343) );
  CKBD0 U6225 ( .CLK(n6343), .C(n6344) );
  CKBD0 U6226 ( .CLK(n6344), .C(n6345) );
  BUFFD0 U6227 ( .I(n6345), .Z(n6346) );
  CKBD0 U6228 ( .CLK(n6346), .C(n6347) );
  CKBD0 U6229 ( .CLK(n6347), .C(n6348) );
  CKBD0 U6230 ( .CLK(n6348), .C(n6349) );
  CKBD0 U6231 ( .CLK(n6349), .C(n6350) );
  CKBD0 U6232 ( .CLK(n6350), .C(n6351) );
  CKBD0 U6233 ( .CLK(n6351), .C(n6352) );
  BUFFD0 U6234 ( .I(n6352), .Z(n6353) );
  CKBD0 U6235 ( .CLK(n6353), .C(n6354) );
  BUFFD0 U6236 ( .I(n6354), .Z(n6355) );
  CKBD0 U6237 ( .CLK(n6355), .C(n6356) );
  BUFFD0 U6238 ( .I(n6356), .Z(n6357) );
  CKBD0 U6239 ( .CLK(n6357), .C(n6358) );
  BUFFD0 U6240 ( .I(n6358), .Z(n6359) );
  CKBD0 U6241 ( .CLK(n6359), .C(n6360) );
  BUFFD0 U6242 ( .I(n6360), .Z(n6361) );
  CKBD0 U6243 ( .CLK(n6361), .C(n6362) );
  BUFFD0 U6244 ( .I(n6362), .Z(n6363) );
  CKBD0 U6245 ( .CLK(n6363), .C(n6364) );
  BUFFD0 U6246 ( .I(n6364), .Z(n6365) );
  CKBD0 U6247 ( .CLK(n6365), .C(n6366) );
  BUFFD0 U6248 ( .I(n6366), .Z(n6367) );
  BUFFD0 U6249 ( .I(n9186), .Z(n6368) );
  BUFFD0 U6250 ( .I(n6370), .Z(n6369) );
  BUFFD0 U6251 ( .I(n6371), .Z(n6370) );
  BUFFD0 U6252 ( .I(Decoder[3]), .Z(n6371) );
  CKBD0 U6253 ( .CLK(n927), .C(n6372) );
  CKBD0 U6254 ( .CLK(n6372), .C(n6373) );
  CKBD0 U6255 ( .CLK(n6373), .C(n6374) );
  BUFFD0 U6256 ( .I(n6374), .Z(n6375) );
  CKBD0 U6257 ( .CLK(n6375), .C(n6376) );
  CKBD0 U6258 ( .CLK(n6376), .C(n6377) );
  CKBD0 U6259 ( .CLK(n6377), .C(n6378) );
  CKBD0 U6260 ( .CLK(n6378), .C(n6379) );
  CKBD0 U6261 ( .CLK(n6379), .C(n6380) );
  CKBD0 U6262 ( .CLK(n6380), .C(n6381) );
  CKBD0 U6263 ( .CLK(n6381), .C(n6382) );
  CKBD0 U6264 ( .CLK(n6382), .C(n6383) );
  CKBD0 U6265 ( .CLK(n6383), .C(n6384) );
  CKBD0 U6266 ( .CLK(n6384), .C(n6385) );
  BUFFD0 U6267 ( .I(n6385), .Z(n6386) );
  CKBD0 U6268 ( .CLK(n6386), .C(n6387) );
  CKBD0 U6269 ( .CLK(n6387), .C(n6388) );
  CKBD0 U6270 ( .CLK(n6388), .C(n6389) );
  CKBD0 U6271 ( .CLK(n6389), .C(n6390) );
  CKBD0 U6272 ( .CLK(n6390), .C(n6391) );
  CKBD0 U6273 ( .CLK(n6391), .C(n6392) );
  CKBD0 U6274 ( .CLK(n6392), .C(n6393) );
  CKBD0 U6275 ( .CLK(n6393), .C(n6394) );
  CKBD0 U6276 ( .CLK(n6394), .C(n6395) );
  BUFFD0 U6277 ( .I(n6395), .Z(n6396) );
  CKBD0 U6278 ( .CLK(n6396), .C(n6397) );
  CKBD0 U6279 ( .CLK(n6397), .C(n6398) );
  CKBD0 U6280 ( .CLK(n6398), .C(n6399) );
  CKBD0 U6281 ( .CLK(n6399), .C(n6400) );
  CKBD0 U6282 ( .CLK(n6400), .C(n6401) );
  CKBD0 U6283 ( .CLK(n6401), .C(n6402) );
  CKBD0 U6284 ( .CLK(n6402), .C(n6403) );
  CKBD0 U6285 ( .CLK(n6403), .C(n6404) );
  CKBD0 U6286 ( .CLK(n6404), .C(n6405) );
  CKBD0 U6287 ( .CLK(n6405), .C(n6406) );
  BUFFD0 U6288 ( .I(n6406), .Z(n6407) );
  CKBD0 U6289 ( .CLK(n6407), .C(n6408) );
  CKBD0 U6290 ( .CLK(n6408), .C(n6409) );
  CKBD0 U6291 ( .CLK(n6409), .C(n6410) );
  CKBD0 U6292 ( .CLK(n6410), .C(n6411) );
  CKBD0 U6293 ( .CLK(n6411), .C(n6412) );
  CKBD0 U6294 ( .CLK(n6412), .C(n6413) );
  CKBD0 U6295 ( .CLK(n6413), .C(n6414) );
  CKBD0 U6296 ( .CLK(n6414), .C(n6415) );
  CKBD0 U6297 ( .CLK(n6415), .C(n6416) );
  CKBD0 U6298 ( .CLK(n6416), .C(n6417) );
  BUFFD0 U6299 ( .I(n6417), .Z(n6418) );
  CKBD0 U6300 ( .CLK(n6418), .C(n6419) );
  CKBD0 U6301 ( .CLK(n6419), .C(n6420) );
  CKBD0 U6302 ( .CLK(n6420), .C(n6421) );
  CKBD0 U6303 ( .CLK(n6421), .C(n6422) );
  CKBD0 U6304 ( .CLK(n6422), .C(n6423) );
  CKBD0 U6305 ( .CLK(n6423), .C(n6424) );
  CKBD0 U6306 ( .CLK(n6424), .C(n6425) );
  CKBD0 U6307 ( .CLK(n6425), .C(n6426) );
  CKBD0 U6308 ( .CLK(n6426), .C(n6427) );
  CKBD0 U6309 ( .CLK(n6427), .C(n6428) );
  BUFFD0 U6310 ( .I(n6428), .Z(n6429) );
  CKBD0 U6311 ( .CLK(n6429), .C(n6430) );
  CKBD0 U6312 ( .CLK(n6430), .C(n6431) );
  CKBD0 U6313 ( .CLK(n6431), .C(n6432) );
  CKBD0 U6314 ( .CLK(n6432), .C(n6433) );
  CKBD0 U6315 ( .CLK(n6433), .C(n6434) );
  CKBD0 U6316 ( .CLK(n6434), .C(n6435) );
  CKBD0 U6317 ( .CLK(n6435), .C(n6436) );
  CKBD0 U6318 ( .CLK(n6436), .C(n6437) );
  CKBD0 U6319 ( .CLK(n6437), .C(n6438) );
  CKBD0 U6320 ( .CLK(n6438), .C(n6439) );
  BUFFD0 U6321 ( .I(n6439), .Z(n6440) );
  CKBD0 U6322 ( .CLK(n6440), .C(n6441) );
  CKBD0 U6323 ( .CLK(n6441), .C(n6442) );
  CKBD0 U6324 ( .CLK(n6442), .C(n6443) );
  CKBD0 U6325 ( .CLK(n6443), .C(n6444) );
  CKBD0 U6326 ( .CLK(n6444), .C(n6445) );
  CKBD0 U6327 ( .CLK(n6445), .C(n6446) );
  CKBD0 U6328 ( .CLK(n6446), .C(n6447) );
  CKBD0 U6329 ( .CLK(n6447), .C(n6448) );
  CKBD0 U6330 ( .CLK(n6448), .C(n6449) );
  CKBD0 U6331 ( .CLK(n6449), .C(n6450) );
  BUFFD0 U6332 ( .I(n6450), .Z(n6451) );
  CKBD0 U6333 ( .CLK(n6451), .C(n6452) );
  CKBD0 U6334 ( .CLK(n6452), .C(n6453) );
  CKBD0 U6335 ( .CLK(n6453), .C(n6454) );
  CKBD0 U6336 ( .CLK(n6454), .C(n6455) );
  CKBD0 U6337 ( .CLK(n6455), .C(n6456) );
  CKBD0 U6338 ( .CLK(n6456), .C(n6457) );
  CKBD0 U6339 ( .CLK(n6457), .C(n6458) );
  CKBD0 U6340 ( .CLK(n6458), .C(n6459) );
  CKBD0 U6341 ( .CLK(n6459), .C(n6460) );
  CKBD0 U6342 ( .CLK(n6460), .C(n6461) );
  BUFFD0 U6343 ( .I(n6461), .Z(n6462) );
  CKBD0 U6344 ( .CLK(n6462), .C(n6463) );
  CKBD0 U6345 ( .CLK(n6463), .C(n6464) );
  CKBD0 U6346 ( .CLK(n6464), .C(n6465) );
  CKBD0 U6347 ( .CLK(n6465), .C(n6466) );
  CKBD0 U6348 ( .CLK(n6466), .C(n6467) );
  CKBD0 U6349 ( .CLK(n6467), .C(n6468) );
  CKBD0 U6350 ( .CLK(n6468), .C(n6469) );
  CKBD0 U6351 ( .CLK(n6469), .C(n6470) );
  CKBD0 U6352 ( .CLK(n6470), .C(n6471) );
  BUFFD0 U6353 ( .I(n6471), .Z(n6472) );
  CKBD0 U6354 ( .CLK(n6472), .C(n6473) );
  CKBD0 U6355 ( .CLK(n6473), .C(n6474) );
  CKBD0 U6356 ( .CLK(n6474), .C(n6475) );
  CKBD0 U6357 ( .CLK(n6475), .C(n6476) );
  CKBD0 U6358 ( .CLK(n6476), .C(n6477) );
  CKBD0 U6359 ( .CLK(n6477), .C(n6478) );
  CKBD0 U6360 ( .CLK(n6478), .C(n6479) );
  CKBD0 U6361 ( .CLK(n6479), .C(n6480) );
  CKBD0 U6362 ( .CLK(n6480), .C(n6481) );
  CKBD0 U6363 ( .CLK(n6481), .C(n6482) );
  BUFFD0 U6364 ( .I(n6482), .Z(n6483) );
  CKBD0 U6365 ( .CLK(n6483), .C(n6484) );
  CKBD0 U6366 ( .CLK(n6484), .C(n6485) );
  CKBD0 U6367 ( .CLK(n6485), .C(n6486) );
  CKBD0 U6368 ( .CLK(n6486), .C(n6487) );
  CKBD0 U6369 ( .CLK(n6487), .C(n6488) );
  CKBD0 U6370 ( .CLK(n6488), .C(n6489) );
  BUFFD0 U6371 ( .I(n6489), .Z(n6490) );
  CKBD0 U6372 ( .CLK(n6490), .C(n6491) );
  BUFFD0 U6373 ( .I(n6491), .Z(n6492) );
  CKBD0 U6374 ( .CLK(n6492), .C(n6493) );
  BUFFD0 U6375 ( .I(n6493), .Z(n6494) );
  CKBD0 U6376 ( .CLK(n6494), .C(n6495) );
  BUFFD0 U6377 ( .I(n6495), .Z(n6496) );
  CKBD0 U6378 ( .CLK(n6496), .C(n6497) );
  BUFFD0 U6379 ( .I(n6497), .Z(n6498) );
  CKBD0 U6380 ( .CLK(n6498), .C(n6499) );
  BUFFD0 U6381 ( .I(n6499), .Z(n6500) );
  CKBD0 U6382 ( .CLK(n6500), .C(n6501) );
  BUFFD0 U6383 ( .I(n6501), .Z(n6502) );
  CKBD0 U6384 ( .CLK(n6502), .C(n6503) );
  BUFFD0 U6385 ( .I(n6503), .Z(n6504) );
  BUFFD0 U6386 ( .I(n9187), .Z(n6505) );
  BUFFD0 U6387 ( .I(n6507), .Z(n6506) );
  BUFFD0 U6388 ( .I(n6508), .Z(n6507) );
  BUFFD0 U6389 ( .I(Decoder[2]), .Z(n6508) );
  CKBD0 U6390 ( .CLK(n925), .C(n6509) );
  CKBD0 U6391 ( .CLK(n6509), .C(n6510) );
  CKBD0 U6392 ( .CLK(n6510), .C(n6511) );
  BUFFD0 U6393 ( .I(n6511), .Z(n6512) );
  CKBD0 U6394 ( .CLK(n6512), .C(n6513) );
  CKBD0 U6395 ( .CLK(n6513), .C(n6514) );
  CKBD0 U6396 ( .CLK(n6514), .C(n6515) );
  CKBD0 U6397 ( .CLK(n6515), .C(n6516) );
  CKBD0 U6398 ( .CLK(n6516), .C(n6517) );
  CKBD0 U6399 ( .CLK(n6517), .C(n6518) );
  CKBD0 U6400 ( .CLK(n6518), .C(n6519) );
  CKBD0 U6401 ( .CLK(n6519), .C(n6520) );
  CKBD0 U6402 ( .CLK(n6520), .C(n6521) );
  CKBD0 U6403 ( .CLK(n6521), .C(n6522) );
  BUFFD0 U6404 ( .I(n6522), .Z(n6523) );
  CKBD0 U6405 ( .CLK(n6523), .C(n6524) );
  CKBD0 U6406 ( .CLK(n6524), .C(n6525) );
  CKBD0 U6407 ( .CLK(n6525), .C(n6526) );
  CKBD0 U6408 ( .CLK(n6526), .C(n6527) );
  CKBD0 U6409 ( .CLK(n6527), .C(n6528) );
  CKBD0 U6410 ( .CLK(n6528), .C(n6529) );
  CKBD0 U6411 ( .CLK(n6529), .C(n6530) );
  CKBD0 U6412 ( .CLK(n6530), .C(n6531) );
  CKBD0 U6413 ( .CLK(n6531), .C(n6532) );
  CKBD0 U6414 ( .CLK(n6532), .C(n6533) );
  BUFFD0 U6415 ( .I(n6533), .Z(n6534) );
  CKBD0 U6416 ( .CLK(n6534), .C(n6535) );
  CKBD0 U6417 ( .CLK(n6535), .C(n6536) );
  CKBD0 U6418 ( .CLK(n6536), .C(n6537) );
  CKBD0 U6419 ( .CLK(n6537), .C(n6538) );
  CKBD0 U6420 ( .CLK(n6538), .C(n6539) );
  CKBD0 U6421 ( .CLK(n6539), .C(n6540) );
  CKBD0 U6422 ( .CLK(n6540), .C(n6541) );
  CKBD0 U6423 ( .CLK(n6541), .C(n6542) );
  CKBD0 U6424 ( .CLK(n6542), .C(n6543) );
  BUFFD0 U6425 ( .I(n6543), .Z(n6544) );
  CKBD0 U6426 ( .CLK(n6544), .C(n6545) );
  CKBD0 U6427 ( .CLK(n6545), .C(n6546) );
  CKBD0 U6428 ( .CLK(n6546), .C(n6547) );
  CKBD0 U6429 ( .CLK(n6547), .C(n6548) );
  CKBD0 U6430 ( .CLK(n6548), .C(n6549) );
  CKBD0 U6431 ( .CLK(n6549), .C(n6550) );
  CKBD0 U6432 ( .CLK(n6550), .C(n6551) );
  CKBD0 U6433 ( .CLK(n6551), .C(n6552) );
  CKBD0 U6434 ( .CLK(n6552), .C(n6553) );
  CKBD0 U6435 ( .CLK(n6553), .C(n6554) );
  BUFFD0 U6436 ( .I(n6554), .Z(n6555) );
  CKBD0 U6437 ( .CLK(n6555), .C(n6556) );
  CKBD0 U6438 ( .CLK(n6556), .C(n6557) );
  CKBD0 U6439 ( .CLK(n6557), .C(n6558) );
  CKBD0 U6440 ( .CLK(n6558), .C(n6559) );
  CKBD0 U6441 ( .CLK(n6559), .C(n6560) );
  CKBD0 U6442 ( .CLK(n6560), .C(n6561) );
  CKBD0 U6443 ( .CLK(n6561), .C(n6562) );
  CKBD0 U6444 ( .CLK(n6562), .C(n6563) );
  CKBD0 U6445 ( .CLK(n6563), .C(n6564) );
  CKBD0 U6446 ( .CLK(n6564), .C(n6565) );
  BUFFD0 U6447 ( .I(n6565), .Z(n6566) );
  CKBD0 U6448 ( .CLK(n6566), .C(n6567) );
  CKBD0 U6449 ( .CLK(n6567), .C(n6568) );
  CKBD0 U6450 ( .CLK(n6568), .C(n6569) );
  CKBD0 U6451 ( .CLK(n6569), .C(n6570) );
  CKBD0 U6452 ( .CLK(n6570), .C(n6571) );
  CKBD0 U6453 ( .CLK(n6571), .C(n6572) );
  CKBD0 U6454 ( .CLK(n6572), .C(n6573) );
  CKBD0 U6455 ( .CLK(n6573), .C(n6574) );
  CKBD0 U6456 ( .CLK(n6574), .C(n6575) );
  CKBD0 U6457 ( .CLK(n6575), .C(n6576) );
  BUFFD0 U6458 ( .I(n6576), .Z(n6577) );
  CKBD0 U6459 ( .CLK(n6577), .C(n6578) );
  CKBD0 U6460 ( .CLK(n6578), .C(n6579) );
  CKBD0 U6461 ( .CLK(n6579), .C(n6580) );
  CKBD0 U6462 ( .CLK(n6580), .C(n6581) );
  CKBD0 U6463 ( .CLK(n6581), .C(n6582) );
  CKBD0 U6464 ( .CLK(n6582), .C(n6583) );
  CKBD0 U6465 ( .CLK(n6583), .C(n6584) );
  CKBD0 U6466 ( .CLK(n6584), .C(n6585) );
  CKBD0 U6467 ( .CLK(n6585), .C(n6586) );
  CKBD0 U6468 ( .CLK(n6586), .C(n6587) );
  BUFFD0 U6469 ( .I(n6587), .Z(n6588) );
  CKBD0 U6470 ( .CLK(n6588), .C(n6589) );
  CKBD0 U6471 ( .CLK(n6589), .C(n6590) );
  CKBD0 U6472 ( .CLK(n6590), .C(n6591) );
  CKBD0 U6473 ( .CLK(n6591), .C(n6592) );
  CKBD0 U6474 ( .CLK(n6592), .C(n6593) );
  CKBD0 U6475 ( .CLK(n6593), .C(n6594) );
  CKBD0 U6476 ( .CLK(n6594), .C(n6595) );
  CKBD0 U6477 ( .CLK(n6595), .C(n6596) );
  CKBD0 U6478 ( .CLK(n6596), .C(n6597) );
  CKBD0 U6479 ( .CLK(n6597), .C(n6598) );
  BUFFD0 U6480 ( .I(n6598), .Z(n6599) );
  CKBD0 U6481 ( .CLK(n6599), .C(n6600) );
  CKBD0 U6482 ( .CLK(n6600), .C(n6601) );
  CKBD0 U6483 ( .CLK(n6601), .C(n6602) );
  CKBD0 U6484 ( .CLK(n6602), .C(n6603) );
  CKBD0 U6485 ( .CLK(n6603), .C(n6604) );
  CKBD0 U6486 ( .CLK(n6604), .C(n6605) );
  CKBD0 U6487 ( .CLK(n6605), .C(n6606) );
  CKBD0 U6488 ( .CLK(n6606), .C(n6607) );
  CKBD0 U6489 ( .CLK(n6607), .C(n6608) );
  BUFFD0 U6490 ( .I(n6608), .Z(n6609) );
  CKBD0 U6491 ( .CLK(n6609), .C(n6610) );
  CKBD0 U6492 ( .CLK(n6610), .C(n6611) );
  CKBD0 U6493 ( .CLK(n6611), .C(n6612) );
  CKBD0 U6494 ( .CLK(n6612), .C(n6613) );
  CKBD0 U6495 ( .CLK(n6613), .C(n6614) );
  CKBD0 U6496 ( .CLK(n6614), .C(n6615) );
  CKBD0 U6497 ( .CLK(n6615), .C(n6616) );
  CKBD0 U6498 ( .CLK(n6616), .C(n6617) );
  CKBD0 U6499 ( .CLK(n6617), .C(n6618) );
  CKBD0 U6500 ( .CLK(n6618), .C(n6619) );
  BUFFD0 U6501 ( .I(n6619), .Z(n6620) );
  CKBD0 U6502 ( .CLK(n6620), .C(n6621) );
  CKBD0 U6503 ( .CLK(n6621), .C(n6622) );
  CKBD0 U6504 ( .CLK(n6622), .C(n6623) );
  CKBD0 U6505 ( .CLK(n6623), .C(n6624) );
  CKBD0 U6506 ( .CLK(n6624), .C(n6625) );
  CKBD0 U6507 ( .CLK(n6625), .C(n6626) );
  BUFFD0 U6508 ( .I(n6626), .Z(n6627) );
  CKBD0 U6509 ( .CLK(n6627), .C(n6628) );
  BUFFD0 U6510 ( .I(n6628), .Z(n6629) );
  CKBD0 U6511 ( .CLK(n6629), .C(n6630) );
  BUFFD0 U6512 ( .I(n6630), .Z(n6631) );
  CKBD0 U6513 ( .CLK(n6631), .C(n6632) );
  BUFFD0 U6514 ( .I(n6632), .Z(n6633) );
  CKBD0 U6515 ( .CLK(n6633), .C(n6634) );
  BUFFD0 U6516 ( .I(n6634), .Z(n6635) );
  CKBD0 U6517 ( .CLK(n6635), .C(n6636) );
  BUFFD0 U6518 ( .I(n6636), .Z(n6637) );
  CKBD0 U6519 ( .CLK(n6637), .C(n6638) );
  BUFFD0 U6520 ( .I(n6638), .Z(n6639) );
  CKBD0 U6521 ( .CLK(n6639), .C(n6640) );
  BUFFD0 U6522 ( .I(n6640), .Z(n6641) );
  BUFFD0 U6523 ( .I(n9188), .Z(n6642) );
  BUFFD0 U6524 ( .I(n6644), .Z(n6643) );
  BUFFD0 U6525 ( .I(n6645), .Z(n6644) );
  BUFFD0 U6526 ( .I(Decoder[1]), .Z(n6645) );
  CKBD0 U6527 ( .CLK(n923), .C(n6646) );
  CKBD0 U6528 ( .CLK(n6646), .C(n6647) );
  CKBD0 U6529 ( .CLK(n6647), .C(n6648) );
  BUFFD0 U6530 ( .I(n6648), .Z(n6649) );
  CKBD0 U6531 ( .CLK(n6649), .C(n6650) );
  CKBD0 U6532 ( .CLK(n6650), .C(n6651) );
  CKBD0 U6533 ( .CLK(n6651), .C(n6652) );
  CKBD0 U6534 ( .CLK(n6652), .C(n6653) );
  CKBD0 U6535 ( .CLK(n6653), .C(n6654) );
  CKBD0 U6536 ( .CLK(n6654), .C(n6655) );
  CKBD0 U6537 ( .CLK(n6655), .C(n6656) );
  CKBD0 U6538 ( .CLK(n6656), .C(n6657) );
  CKBD0 U6539 ( .CLK(n6657), .C(n6658) );
  CKBD0 U6540 ( .CLK(n6658), .C(n6659) );
  BUFFD0 U6541 ( .I(n6659), .Z(n6660) );
  CKBD0 U6542 ( .CLK(n6660), .C(n6661) );
  CKBD0 U6543 ( .CLK(n6661), .C(n6662) );
  CKBD0 U6544 ( .CLK(n6662), .C(n6663) );
  CKBD0 U6545 ( .CLK(n6663), .C(n6664) );
  CKBD0 U6546 ( .CLK(n6664), .C(n6665) );
  CKBD0 U6547 ( .CLK(n6665), .C(n6666) );
  CKBD0 U6548 ( .CLK(n6666), .C(n6667) );
  CKBD0 U6549 ( .CLK(n6667), .C(n6668) );
  CKBD0 U6550 ( .CLK(n6668), .C(n6669) );
  BUFFD0 U6551 ( .I(n6669), .Z(n6670) );
  CKBD0 U6552 ( .CLK(n6670), .C(n6671) );
  CKBD0 U6553 ( .CLK(n6671), .C(n6672) );
  CKBD0 U6554 ( .CLK(n6672), .C(n6673) );
  CKBD0 U6555 ( .CLK(n6673), .C(n6674) );
  CKBD0 U6556 ( .CLK(n6674), .C(n6675) );
  CKBD0 U6557 ( .CLK(n6675), .C(n6676) );
  CKBD0 U6558 ( .CLK(n6676), .C(n6677) );
  CKBD0 U6559 ( .CLK(n6677), .C(n6678) );
  CKBD0 U6560 ( .CLK(n6678), .C(n6679) );
  CKBD0 U6561 ( .CLK(n6679), .C(n6680) );
  BUFFD0 U6562 ( .I(n6680), .Z(n6681) );
  CKBD0 U6563 ( .CLK(n6681), .C(n6682) );
  CKBD0 U6564 ( .CLK(n6682), .C(n6683) );
  CKBD0 U6565 ( .CLK(n6683), .C(n6684) );
  CKBD0 U6566 ( .CLK(n6684), .C(n6685) );
  CKBD0 U6567 ( .CLK(n6685), .C(n6686) );
  CKBD0 U6568 ( .CLK(n6686), .C(n6687) );
  CKBD0 U6569 ( .CLK(n6687), .C(n6688) );
  CKBD0 U6570 ( .CLK(n6688), .C(n6689) );
  CKBD0 U6571 ( .CLK(n6689), .C(n6690) );
  CKBD0 U6572 ( .CLK(n6690), .C(n6691) );
  BUFFD0 U6573 ( .I(n6691), .Z(n6692) );
  CKBD0 U6574 ( .CLK(n6692), .C(n6693) );
  CKBD0 U6575 ( .CLK(n6693), .C(n6694) );
  CKBD0 U6576 ( .CLK(n6694), .C(n6695) );
  CKBD0 U6577 ( .CLK(n6695), .C(n6696) );
  CKBD0 U6578 ( .CLK(n6696), .C(n6697) );
  CKBD0 U6579 ( .CLK(n6697), .C(n6698) );
  CKBD0 U6580 ( .CLK(n6698), .C(n6699) );
  CKBD0 U6581 ( .CLK(n6699), .C(n6700) );
  CKBD0 U6582 ( .CLK(n6700), .C(n6701) );
  CKBD0 U6583 ( .CLK(n6701), .C(n6702) );
  BUFFD0 U6584 ( .I(n6702), .Z(n6703) );
  CKBD0 U6585 ( .CLK(n6703), .C(n6704) );
  CKBD0 U6586 ( .CLK(n6704), .C(n6705) );
  CKBD0 U6587 ( .CLK(n6705), .C(n6706) );
  CKBD0 U6588 ( .CLK(n6706), .C(n6707) );
  CKBD0 U6589 ( .CLK(n6707), .C(n6708) );
  CKBD0 U6590 ( .CLK(n6708), .C(n6709) );
  CKBD0 U6591 ( .CLK(n6709), .C(n6710) );
  CKBD0 U6592 ( .CLK(n6710), .C(n6711) );
  CKBD0 U6593 ( .CLK(n6711), .C(n6712) );
  CKBD0 U6594 ( .CLK(n6712), .C(n6713) );
  BUFFD0 U6595 ( .I(n6713), .Z(n6714) );
  CKBD0 U6596 ( .CLK(n6714), .C(n6715) );
  CKBD0 U6597 ( .CLK(n6715), .C(n6716) );
  CKBD0 U6598 ( .CLK(n6716), .C(n6717) );
  CKBD0 U6599 ( .CLK(n6717), .C(n6718) );
  CKBD0 U6600 ( .CLK(n6718), .C(n6719) );
  CKBD0 U6601 ( .CLK(n6719), .C(n6720) );
  CKBD0 U6602 ( .CLK(n6720), .C(n6721) );
  CKBD0 U6603 ( .CLK(n6721), .C(n6722) );
  CKBD0 U6604 ( .CLK(n6722), .C(n6723) );
  CKBD0 U6605 ( .CLK(n6723), .C(n6724) );
  BUFFD0 U6606 ( .I(n6724), .Z(n6725) );
  CKBD0 U6607 ( .CLK(n6725), .C(n6726) );
  CKBD0 U6608 ( .CLK(n6726), .C(n6727) );
  CKBD0 U6609 ( .CLK(n6727), .C(n6728) );
  CKBD0 U6610 ( .CLK(n6728), .C(n6729) );
  CKBD0 U6611 ( .CLK(n6729), .C(n6730) );
  CKBD0 U6612 ( .CLK(n6730), .C(n6731) );
  CKBD0 U6613 ( .CLK(n6731), .C(n6732) );
  CKBD0 U6614 ( .CLK(n6732), .C(n6733) );
  CKBD0 U6615 ( .CLK(n6733), .C(n6734) );
  BUFFD0 U6616 ( .I(n6734), .Z(n6735) );
  CKBD0 U6617 ( .CLK(n6735), .C(n6736) );
  CKBD0 U6618 ( .CLK(n6736), .C(n6737) );
  CKBD0 U6619 ( .CLK(n6737), .C(n6738) );
  CKBD0 U6620 ( .CLK(n6738), .C(n6739) );
  CKBD0 U6621 ( .CLK(n6739), .C(n6740) );
  CKBD0 U6622 ( .CLK(n6740), .C(n6741) );
  CKBD0 U6623 ( .CLK(n6741), .C(n6742) );
  CKBD0 U6624 ( .CLK(n6742), .C(n6743) );
  CKBD0 U6625 ( .CLK(n6743), .C(n6744) );
  CKBD0 U6626 ( .CLK(n6744), .C(n6745) );
  BUFFD0 U6627 ( .I(n6745), .Z(n6746) );
  CKBD0 U6628 ( .CLK(n6746), .C(n6747) );
  CKBD0 U6629 ( .CLK(n6747), .C(n6748) );
  CKBD0 U6630 ( .CLK(n6748), .C(n6749) );
  CKBD0 U6631 ( .CLK(n6749), .C(n6750) );
  CKBD0 U6632 ( .CLK(n6750), .C(n6751) );
  CKBD0 U6633 ( .CLK(n6751), .C(n6752) );
  CKBD0 U6634 ( .CLK(n6752), .C(n6753) );
  CKBD0 U6635 ( .CLK(n6753), .C(n6754) );
  CKBD0 U6636 ( .CLK(n6754), .C(n6755) );
  CKBD0 U6637 ( .CLK(n6755), .C(n6756) );
  BUFFD0 U6638 ( .I(n6756), .Z(n6757) );
  CKBD0 U6639 ( .CLK(n6757), .C(n6758) );
  CKBD0 U6640 ( .CLK(n6758), .C(n6759) );
  CKBD0 U6641 ( .CLK(n6759), .C(n6760) );
  CKBD0 U6642 ( .CLK(n6760), .C(n6761) );
  CKBD0 U6643 ( .CLK(n6761), .C(n6762) );
  CKBD0 U6644 ( .CLK(n6762), .C(n6763) );
  BUFFD0 U6645 ( .I(n6763), .Z(n6764) );
  CKBD0 U6646 ( .CLK(n6764), .C(n6765) );
  BUFFD0 U6647 ( .I(n6765), .Z(n6766) );
  CKBD0 U6648 ( .CLK(n6766), .C(n6767) );
  BUFFD0 U6649 ( .I(n6767), .Z(n6768) );
  CKBD0 U6650 ( .CLK(n6768), .C(n6769) );
  BUFFD0 U6651 ( .I(n6769), .Z(n6770) );
  CKBD0 U6652 ( .CLK(n6770), .C(n6771) );
  BUFFD0 U6653 ( .I(n6771), .Z(n6772) );
  CKBD0 U6654 ( .CLK(n6772), .C(n6773) );
  BUFFD0 U6655 ( .I(n6773), .Z(n6774) );
  CKBD0 U6656 ( .CLK(n6774), .C(n6775) );
  BUFFD0 U6657 ( .I(n6775), .Z(n6776) );
  CKBD0 U6658 ( .CLK(n6776), .C(n6777) );
  BUFFD0 U6659 ( .I(n6777), .Z(n6778) );
  BUFFD0 U6660 ( .I(n9189), .Z(n6779) );
  BUFFD0 U6661 ( .I(n6781), .Z(n6780) );
  BUFFD0 U6662 ( .I(n6782), .Z(n6781) );
  BUFFD0 U6663 ( .I(Decoder[0]), .Z(n6782) );
  CKBD0 U6664 ( .CLK(n921), .C(n6783) );
  CKBD0 U6665 ( .CLK(n6783), .C(n6784) );
  CKBD0 U6666 ( .CLK(n6784), .C(n6785) );
  BUFFD0 U6667 ( .I(n6785), .Z(n6786) );
  CKBD0 U6668 ( .CLK(n6786), .C(n6787) );
  CKBD0 U6669 ( .CLK(n6787), .C(n6788) );
  CKBD0 U6670 ( .CLK(n6788), .C(n6789) );
  CKBD0 U6671 ( .CLK(n6789), .C(n6790) );
  CKBD0 U6672 ( .CLK(n6790), .C(n6791) );
  CKBD0 U6673 ( .CLK(n6791), .C(n6792) );
  CKBD0 U6674 ( .CLK(n6792), .C(n6793) );
  CKBD0 U6675 ( .CLK(n6793), .C(n6794) );
  CKBD0 U6676 ( .CLK(n6794), .C(n6795) );
  CKBD0 U6677 ( .CLK(n6795), .C(n6796) );
  BUFFD0 U6678 ( .I(n6796), .Z(n6797) );
  CKBD0 U6679 ( .CLK(n6797), .C(n6798) );
  CKBD0 U6680 ( .CLK(n6798), .C(n6799) );
  CKBD0 U6681 ( .CLK(n6799), .C(n6800) );
  CKBD0 U6682 ( .CLK(n6800), .C(n6801) );
  CKBD0 U6683 ( .CLK(n6801), .C(n6802) );
  CKBD0 U6684 ( .CLK(n6802), .C(n6803) );
  CKBD0 U6685 ( .CLK(n6803), .C(n6804) );
  CKBD0 U6686 ( .CLK(n6804), .C(n6805) );
  CKBD0 U6687 ( .CLK(n6805), .C(n6806) );
  BUFFD0 U6688 ( .I(n6806), .Z(n6807) );
  CKBD0 U6689 ( .CLK(n6807), .C(n6808) );
  CKBD0 U6690 ( .CLK(n6808), .C(n6809) );
  CKBD0 U6691 ( .CLK(n6809), .C(n6810) );
  CKBD0 U6692 ( .CLK(n6810), .C(n6811) );
  CKBD0 U6693 ( .CLK(n6811), .C(n6812) );
  CKBD0 U6694 ( .CLK(n6812), .C(n6813) );
  CKBD0 U6695 ( .CLK(n6813), .C(n6814) );
  CKBD0 U6696 ( .CLK(n6814), .C(n6815) );
  CKBD0 U6697 ( .CLK(n6815), .C(n6816) );
  CKBD0 U6698 ( .CLK(n6816), .C(n6817) );
  BUFFD0 U6699 ( .I(n6817), .Z(n6818) );
  CKBD0 U6700 ( .CLK(n6818), .C(n6819) );
  CKBD0 U6701 ( .CLK(n6819), .C(n6820) );
  CKBD0 U6702 ( .CLK(n6820), .C(n6821) );
  CKBD0 U6703 ( .CLK(n6821), .C(n6822) );
  CKBD0 U6704 ( .CLK(n6822), .C(n6823) );
  CKBD0 U6705 ( .CLK(n6823), .C(n6824) );
  CKBD0 U6706 ( .CLK(n6824), .C(n6825) );
  CKBD0 U6707 ( .CLK(n6825), .C(n6826) );
  CKBD0 U6708 ( .CLK(n6826), .C(n6827) );
  CKBD0 U6709 ( .CLK(n6827), .C(n6828) );
  BUFFD0 U6710 ( .I(n6828), .Z(n6829) );
  CKBD0 U6711 ( .CLK(n6829), .C(n6830) );
  CKBD0 U6712 ( .CLK(n6830), .C(n6831) );
  CKBD0 U6713 ( .CLK(n6831), .C(n6832) );
  CKBD0 U6714 ( .CLK(n6832), .C(n6833) );
  CKBD0 U6715 ( .CLK(n6833), .C(n6834) );
  CKBD0 U6716 ( .CLK(n6834), .C(n6835) );
  CKBD0 U6717 ( .CLK(n6835), .C(n6836) );
  CKBD0 U6718 ( .CLK(n6836), .C(n6837) );
  CKBD0 U6719 ( .CLK(n6837), .C(n6838) );
  CKBD0 U6720 ( .CLK(n6838), .C(n6839) );
  BUFFD0 U6721 ( .I(n6839), .Z(n6840) );
  CKBD0 U6722 ( .CLK(n6840), .C(n6841) );
  CKBD0 U6723 ( .CLK(n6841), .C(n6842) );
  CKBD0 U6724 ( .CLK(n6842), .C(n6843) );
  CKBD0 U6725 ( .CLK(n6843), .C(n6844) );
  CKBD0 U6726 ( .CLK(n6844), .C(n6845) );
  CKBD0 U6727 ( .CLK(n6845), .C(n6846) );
  CKBD0 U6728 ( .CLK(n6846), .C(n6847) );
  CKBD0 U6729 ( .CLK(n6847), .C(n6848) );
  CKBD0 U6730 ( .CLK(n6848), .C(n6849) );
  CKBD0 U6731 ( .CLK(n6849), .C(n6850) );
  BUFFD0 U6732 ( .I(n6850), .Z(n6851) );
  CKBD0 U6733 ( .CLK(n6851), .C(n6852) );
  CKBD0 U6734 ( .CLK(n6852), .C(n6853) );
  CKBD0 U6735 ( .CLK(n6853), .C(n6854) );
  CKBD0 U6736 ( .CLK(n6854), .C(n6855) );
  CKBD0 U6737 ( .CLK(n6855), .C(n6856) );
  CKBD0 U6738 ( .CLK(n6856), .C(n6857) );
  CKBD0 U6739 ( .CLK(n6857), .C(n6858) );
  CKBD0 U6740 ( .CLK(n6858), .C(n6859) );
  CKBD0 U6741 ( .CLK(n6859), .C(n6860) );
  CKBD0 U6742 ( .CLK(n6860), .C(n6861) );
  BUFFD0 U6743 ( .I(n6861), .Z(n6862) );
  CKBD0 U6744 ( .CLK(n6862), .C(n6863) );
  CKBD0 U6745 ( .CLK(n6863), .C(n6864) );
  CKBD0 U6746 ( .CLK(n6864), .C(n6865) );
  CKBD0 U6747 ( .CLK(n6865), .C(n6866) );
  CKBD0 U6748 ( .CLK(n6866), .C(n6867) );
  CKBD0 U6749 ( .CLK(n6867), .C(n6868) );
  CKBD0 U6750 ( .CLK(n6868), .C(n6869) );
  CKBD0 U6751 ( .CLK(n6869), .C(n6870) );
  CKBD0 U6752 ( .CLK(n6870), .C(n6871) );
  CKBD0 U6753 ( .CLK(n6871), .C(n6872) );
  BUFFD0 U6754 ( .I(n6872), .Z(n6873) );
  CKBD0 U6755 ( .CLK(n6873), .C(n6874) );
  CKBD0 U6756 ( .CLK(n6874), .C(n6875) );
  CKBD0 U6757 ( .CLK(n6875), .C(n6876) );
  CKBD0 U6758 ( .CLK(n6876), .C(n6877) );
  CKBD0 U6759 ( .CLK(n6877), .C(n6878) );
  CKBD0 U6760 ( .CLK(n6878), .C(n6879) );
  CKBD0 U6761 ( .CLK(n6879), .C(n6880) );
  CKBD0 U6762 ( .CLK(n6880), .C(n6881) );
  CKBD0 U6763 ( .CLK(n6881), .C(n6882) );
  BUFFD0 U6764 ( .I(n6882), .Z(n6883) );
  CKBD0 U6765 ( .CLK(n6883), .C(n6884) );
  CKBD0 U6766 ( .CLK(n6884), .C(n6885) );
  CKBD0 U6767 ( .CLK(n6885), .C(n6886) );
  CKBD0 U6768 ( .CLK(n6886), .C(n6887) );
  CKBD0 U6769 ( .CLK(n6887), .C(n6888) );
  CKBD0 U6770 ( .CLK(n6888), .C(n6889) );
  CKBD0 U6771 ( .CLK(n6889), .C(n6890) );
  CKBD0 U6772 ( .CLK(n6890), .C(n6891) );
  CKBD0 U6773 ( .CLK(n6891), .C(n6892) );
  CKBD0 U6774 ( .CLK(n6892), .C(n6893) );
  BUFFD0 U6775 ( .I(n6893), .Z(n6894) );
  CKBD0 U6776 ( .CLK(n6894), .C(n6895) );
  CKBD0 U6777 ( .CLK(n6895), .C(n6896) );
  CKBD0 U6778 ( .CLK(n6896), .C(n6897) );
  CKBD0 U6779 ( .CLK(n6897), .C(n6898) );
  CKBD0 U6780 ( .CLK(n6898), .C(n6899) );
  CKBD0 U6781 ( .CLK(n6899), .C(n6900) );
  BUFFD0 U6782 ( .I(n6900), .Z(n6901) );
  CKBD0 U6783 ( .CLK(n6901), .C(n6902) );
  BUFFD0 U6784 ( .I(n6902), .Z(n6903) );
  CKBD0 U6785 ( .CLK(n6903), .C(n6904) );
  BUFFD0 U6786 ( .I(n6904), .Z(n6905) );
  CKBD0 U6787 ( .CLK(n6905), .C(n6906) );
  BUFFD0 U6788 ( .I(n6906), .Z(n6907) );
  CKBD0 U6789 ( .CLK(n6907), .C(n6908) );
  BUFFD0 U6790 ( .I(n6908), .Z(n6909) );
  CKBD0 U6791 ( .CLK(n6909), .C(n6910) );
  BUFFD0 U6792 ( .I(n6910), .Z(n6911) );
  CKBD0 U6793 ( .CLK(n6911), .C(n6912) );
  BUFFD0 U6794 ( .I(n6912), .Z(n6913) );
  CKBD0 U6795 ( .CLK(n6913), .C(n6914) );
  BUFFD0 U6796 ( .I(n6914), .Z(n6915) );
  BUFFD0 U6797 ( .I(n6917), .Z(n6916) );
  BUFFD0 U6798 ( .I(n9223), .Z(n6917) );
  CKND2D0 U6799 ( .A1(n9155), .A2(ParValidTimer[0]), .ZN(n9278) );
  XOR2D0 U6800 ( .A1(n9021), .A2(n9278), .Z(n9277) );
  BUFFD0 U6801 ( .I(N39), .Z(n6918) );
  CKBD0 U6802 ( .CLK(Count32[0]), .C(n6927) );
  BUFFD0 U6803 ( .I(Count32[1]), .Z(n6919) );
  BUFFD0 U6804 ( .I(n9222), .Z(n6920) );
  BUFFD0 U6805 ( .I(n9276), .Z(n6921) );
  CKXOR2D0 U6806 ( .A1(n9155), .A2(n9282), .Z(n9276) );
  BUFFD0 U6807 ( .I(n6923), .Z(n6922) );
  BUFFD0 U6808 ( .I(N41), .Z(n6923) );
  BUFFD0 U6809 ( .I(n6925), .Z(n6924) );
  BUFFD0 U6810 ( .I(N40), .Z(n6925) );
  BUFFD0 U6811 ( .I(N38), .Z(n6926) );
  BUFFD0 U6812 ( .I(n6929), .Z(n6928) );
  BUFFD0 U6813 ( .I(n6930), .Z(n6929) );
  BUFFD0 U6814 ( .I(n6931), .Z(n6930) );
  BUFFD0 U6815 ( .I(n9192), .Z(n6931) );
  IOA22D0 U6816 ( .B1(n9127), .B2(n9229), .A1(n1), .A2(Decoder[2]), .ZN(n9192)
         );
  BUFFD0 U6817 ( .I(n6933), .Z(n6932) );
  BUFFD0 U6818 ( .I(n6934), .Z(n6933) );
  BUFFD0 U6819 ( .I(n6935), .Z(n6934) );
  BUFFD0 U6820 ( .I(n9191), .Z(n6935) );
  IOA22D0 U6821 ( .B1(n9127), .B2(n9228), .A1(n1), .A2(Decoder[1]), .ZN(n9191)
         );
  BUFFD0 U6822 ( .I(n6937), .Z(n6936) );
  BUFFD0 U6823 ( .I(N37), .Z(n6937) );
  BUFFD0 U6824 ( .I(n6939), .Z(n6938) );
  BUFFD0 U6825 ( .I(N43), .Z(n6939) );
  BUFFD0 U6826 ( .I(n6941), .Z(n6940) );
  BUFFD0 U6827 ( .I(n6942), .Z(n6941) );
  BUFFD0 U6828 ( .I(n6943), .Z(n6942) );
  BUFFD0 U6829 ( .I(n9190), .Z(n6943) );
  IOA22D0 U6830 ( .B1(n9128), .B2(n9227), .A1(n1), .A2(Decoder[0]), .ZN(n9190)
         );
  BUFFD0 U6831 ( .I(n6945), .Z(n6944) );
  BUFFD0 U6832 ( .I(n6946), .Z(n6945) );
  BUFFD0 U6833 ( .I(n6947), .Z(n6946) );
  BUFFD0 U6834 ( .I(n9195), .Z(n6947) );
  IOA22D0 U6835 ( .B1(n9127), .B2(n9232), .A1(n1), .A2(Decoder[5]), .ZN(n9195)
         );
  CKBD0 U6836 ( .CLK(n9202), .C(n6951) );
  BUFFD0 U6837 ( .I(n6949), .Z(n6948) );
  BUFFD0 U6838 ( .I(n6950), .Z(n6949) );
  BUFFD0 U6839 ( .I(n6951), .Z(n6950) );
  CKBD0 U6840 ( .CLK(n9209), .C(n6955) );
  BUFFD0 U6841 ( .I(n6953), .Z(n6952) );
  BUFFD0 U6842 ( .I(n6954), .Z(n6953) );
  BUFFD0 U6843 ( .I(n6955), .Z(n6954) );
  CKBD0 U6844 ( .CLK(n9196), .C(n6959) );
  MOAI22D1 U6845 ( .A1(n9127), .A2(n9233), .B1(n9129), .B2(Decoder[6]), .ZN(
        n9196) );
  BUFFD0 U6846 ( .I(n6957), .Z(n6956) );
  BUFFD0 U6847 ( .I(n6958), .Z(n6957) );
  BUFFD0 U6848 ( .I(n6959), .Z(n6958) );
  IOA22D4 U6849 ( .B1(n9127), .B2(n9236), .A1(n9129), .A2(Decoder[9]), .ZN(
        n9199) );
  BUFFD0 U6850 ( .I(n6961), .Z(n6960) );
  BUFFD0 U6851 ( .I(n6962), .Z(n6961) );
  BUFFD0 U6852 ( .I(n6963), .Z(n6962) );
  BUFFD0 U6853 ( .I(n9199), .Z(n6963) );
  IOA22D4 U6854 ( .B1(n9127), .B2(n9240), .A1(n9129), .A2(Decoder[13]), .ZN(
        n9203) );
  BUFFD0 U6855 ( .I(n6965), .Z(n6964) );
  BUFFD0 U6856 ( .I(n6966), .Z(n6965) );
  BUFFD0 U6857 ( .I(n6967), .Z(n6966) );
  BUFFD0 U6858 ( .I(n9203), .Z(n6967) );
  IOA22D4 U6859 ( .B1(n9128), .B2(n9243), .A1(n9129), .A2(Decoder[16]), .ZN(
        n9206) );
  BUFFD0 U6860 ( .I(n6969), .Z(n6968) );
  BUFFD0 U6861 ( .I(n6970), .Z(n6969) );
  BUFFD0 U6862 ( .I(n6971), .Z(n6970) );
  BUFFD0 U6863 ( .I(n9206), .Z(n6971) );
  IOA22D4 U6864 ( .B1(n9128), .B2(n9247), .A1(n9128), .A2(Decoder[20]), .ZN(
        n9210) );
  BUFFD0 U6865 ( .I(n6973), .Z(n6972) );
  BUFFD0 U6866 ( .I(n6974), .Z(n6973) );
  BUFFD0 U6867 ( .I(n6975), .Z(n6974) );
  BUFFD0 U6868 ( .I(n9210), .Z(n6975) );
  IOA22D4 U6869 ( .B1(n9128), .B2(n9250), .A1(n9129), .A2(Decoder[23]), .ZN(
        n9213) );
  BUFFD0 U6870 ( .I(n6977), .Z(n6976) );
  BUFFD0 U6871 ( .I(n6978), .Z(n6977) );
  BUFFD0 U6872 ( .I(n6979), .Z(n6978) );
  BUFFD0 U6873 ( .I(n9213), .Z(n6979) );
  IOA22D4 U6874 ( .B1(n9128), .B2(n9251), .A1(n9129), .A2(Decoder[24]), .ZN(
        n9214) );
  BUFFD0 U6875 ( .I(n6981), .Z(n6980) );
  BUFFD0 U6876 ( .I(n6982), .Z(n6981) );
  BUFFD0 U6877 ( .I(n6983), .Z(n6982) );
  BUFFD0 U6878 ( .I(n9214), .Z(n6983) );
  IOA22D4 U6879 ( .B1(n9128), .B2(n9254), .A1(n9129), .A2(Decoder[27]), .ZN(
        n9217) );
  BUFFD0 U6880 ( .I(n6985), .Z(n6984) );
  BUFFD0 U6881 ( .I(n6986), .Z(n6985) );
  BUFFD0 U6882 ( .I(n6987), .Z(n6986) );
  BUFFD0 U6883 ( .I(n9217), .Z(n6987) );
  IOA22D4 U6884 ( .B1(n9128), .B2(n9255), .A1(n1), .A2(Decoder[28]), .ZN(n9218) );
  BUFFD0 U6885 ( .I(n6989), .Z(n6988) );
  BUFFD0 U6886 ( .I(n6990), .Z(n6989) );
  BUFFD0 U6887 ( .I(n6991), .Z(n6990) );
  BUFFD0 U6888 ( .I(n9218), .Z(n6991) );
  BUFFD0 U6889 ( .I(n6993), .Z(n6992) );
  BUFFD0 U6890 ( .I(n6994), .Z(n6993) );
  BUFFD0 U6891 ( .I(n6995), .Z(n6994) );
  BUFFD0 U6892 ( .I(n9221), .Z(n6995) );
  BUFFD0 U6893 ( .I(n6997), .Z(n6996) );
  BUFFD0 U6894 ( .I(n6998), .Z(n6997) );
  BUFFD0 U6895 ( .I(n6999), .Z(n6998) );
  BUFFD0 U6896 ( .I(n9193), .Z(n6999) );
  IOA22D0 U6897 ( .B1(n9127), .B2(n9230), .A1(n1), .A2(Decoder[3]), .ZN(n9193)
         );
  BUFFD0 U6898 ( .I(n7001), .Z(n7000) );
  BUFFD0 U6899 ( .I(n7002), .Z(n7001) );
  BUFFD0 U6900 ( .I(n7003), .Z(n7002) );
  BUFFD0 U6901 ( .I(n9194), .Z(n7003) );
  IOA22D0 U6902 ( .B1(n9127), .B2(n9231), .A1(n1), .A2(Decoder[4]), .ZN(n9194)
         );
  IOA22D4 U6903 ( .B1(n9127), .B2(n9237), .A1(n9129), .A2(Decoder[10]), .ZN(
        n9200) );
  BUFFD0 U6904 ( .I(n7005), .Z(n7004) );
  BUFFD0 U6905 ( .I(n7006), .Z(n7005) );
  BUFFD0 U6906 ( .I(n7007), .Z(n7006) );
  BUFFD0 U6907 ( .I(n9200), .Z(n7007) );
  IOA22D4 U6908 ( .B1(n9127), .B2(n9238), .A1(n9129), .A2(Decoder[11]), .ZN(
        n9201) );
  BUFFD0 U6909 ( .I(n7009), .Z(n7008) );
  BUFFD0 U6910 ( .I(n7010), .Z(n7009) );
  BUFFD0 U6911 ( .I(n7011), .Z(n7010) );
  BUFFD0 U6912 ( .I(n9201), .Z(n7011) );
  IOA22D4 U6913 ( .B1(n9128), .B2(n9244), .A1(n9129), .A2(Decoder[17]), .ZN(
        n9207) );
  BUFFD0 U6914 ( .I(n7013), .Z(n7012) );
  BUFFD0 U6915 ( .I(n7014), .Z(n7013) );
  BUFFD0 U6916 ( .I(n7015), .Z(n7014) );
  BUFFD0 U6917 ( .I(n9207), .Z(n7015) );
  IOA22D4 U6918 ( .B1(n9128), .B2(n9245), .A1(n9129), .A2(Decoder[18]), .ZN(
        n9208) );
  BUFFD0 U6919 ( .I(n7017), .Z(n7016) );
  BUFFD0 U6920 ( .I(n7018), .Z(n7017) );
  BUFFD0 U6921 ( .I(n7019), .Z(n7018) );
  BUFFD0 U6922 ( .I(n9208), .Z(n7019) );
  IOA22D4 U6923 ( .B1(n9127), .B2(n9234), .A1(n1), .A2(Decoder[7]), .ZN(n9197)
         );
  BUFFD0 U6924 ( .I(n7021), .Z(n7020) );
  BUFFD0 U6925 ( .I(n7022), .Z(n7021) );
  BUFFD0 U6926 ( .I(n7023), .Z(n7022) );
  BUFFD0 U6927 ( .I(n9197), .Z(n7023) );
  IOA22D4 U6928 ( .B1(n9127), .B2(n9235), .A1(n9129), .A2(Decoder[8]), .ZN(
        n9198) );
  BUFFD0 U6929 ( .I(n7025), .Z(n7024) );
  BUFFD0 U6930 ( .I(n7026), .Z(n7025) );
  BUFFD0 U6931 ( .I(n7027), .Z(n7026) );
  BUFFD0 U6932 ( .I(n9198), .Z(n7027) );
  IOA22D4 U6933 ( .B1(n9128), .B2(n9241), .A1(n9129), .A2(Decoder[14]), .ZN(
        n9204) );
  BUFFD0 U6934 ( .I(n7029), .Z(n7028) );
  BUFFD0 U6935 ( .I(n7030), .Z(n7029) );
  BUFFD0 U6936 ( .I(n7031), .Z(n7030) );
  BUFFD0 U6937 ( .I(n9204), .Z(n7031) );
  IOA22D4 U6938 ( .B1(n9128), .B2(n9242), .A1(n9129), .A2(Decoder[15]), .ZN(
        n9205) );
  BUFFD0 U6939 ( .I(n7033), .Z(n7032) );
  BUFFD0 U6940 ( .I(n7034), .Z(n7033) );
  BUFFD0 U6941 ( .I(n7035), .Z(n7034) );
  BUFFD0 U6942 ( .I(n9205), .Z(n7035) );
  IOA22D4 U6943 ( .B1(n9128), .B2(n9248), .A1(n9129), .A2(Decoder[21]), .ZN(
        n9211) );
  BUFFD0 U6944 ( .I(n7037), .Z(n7036) );
  BUFFD0 U6945 ( .I(n7038), .Z(n7037) );
  BUFFD0 U6946 ( .I(n7039), .Z(n7038) );
  BUFFD0 U6947 ( .I(n9211), .Z(n7039) );
  IOA22D4 U6948 ( .B1(n9128), .B2(n9249), .A1(n9129), .A2(Decoder[22]), .ZN(
        n9212) );
  BUFFD0 U6949 ( .I(n7041), .Z(n7040) );
  BUFFD0 U6950 ( .I(n7042), .Z(n7041) );
  BUFFD0 U6951 ( .I(n7043), .Z(n7042) );
  BUFFD0 U6952 ( .I(n9212), .Z(n7043) );
  IOA22D4 U6953 ( .B1(n9128), .B2(n9252), .A1(n9129), .A2(Decoder[25]), .ZN(
        n9215) );
  BUFFD0 U6954 ( .I(n7045), .Z(n7044) );
  BUFFD0 U6955 ( .I(n7046), .Z(n7045) );
  BUFFD0 U6956 ( .I(n7047), .Z(n7046) );
  BUFFD0 U6957 ( .I(n9215), .Z(n7047) );
  IOA22D4 U6958 ( .B1(n9128), .B2(n9253), .A1(n9129), .A2(Decoder[26]), .ZN(
        n9216) );
  BUFFD0 U6959 ( .I(n7049), .Z(n7048) );
  BUFFD0 U6960 ( .I(n7050), .Z(n7049) );
  BUFFD0 U6961 ( .I(n7051), .Z(n7050) );
  BUFFD0 U6962 ( .I(n9216), .Z(n7051) );
  IOA22D4 U6963 ( .B1(n9128), .B2(n9256), .A1(n1), .A2(Decoder[29]), .ZN(n9219) );
  BUFFD0 U6964 ( .I(n7053), .Z(n7052) );
  BUFFD0 U6965 ( .I(n7054), .Z(n7053) );
  BUFFD0 U6966 ( .I(n7055), .Z(n7054) );
  BUFFD0 U6967 ( .I(n9219), .Z(n7055) );
  IOA22D4 U6968 ( .B1(n9128), .B2(n9257), .A1(n1), .A2(Decoder[30]), .ZN(n9220) );
  BUFFD0 U6969 ( .I(n7057), .Z(n7056) );
  BUFFD0 U6970 ( .I(n7058), .Z(n7057) );
  BUFFD0 U6971 ( .I(n7059), .Z(n7058) );
  BUFFD0 U6972 ( .I(n9220), .Z(n7059) );
  OAI21D0 U6973 ( .A1(n9283), .A2(n9259), .B(n9156), .ZN(n9226) );
  BUFFD0 U6974 ( .I(n7061), .Z(n7060) );
  BUFFD0 U6975 ( .I(n7062), .Z(n7061) );
  BUFFD0 U6976 ( .I(n7063), .Z(n7062) );
  BUFFD0 U6977 ( .I(n9226), .Z(n7063) );
  NR2D0 U6978 ( .A1(n9273), .A2(n9274), .ZN(N47) );
  CKND2D0 U6979 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  CKBD0 U6980 ( .CLK(n2165), .C(n7064) );
  CKBD0 U6981 ( .CLK(n2068), .C(n7065) );
  CKBD0 U6982 ( .CLK(n2262), .C(n7066) );
  CKBD0 U6983 ( .CLK(n1352), .C(n7067) );
  CKBD0 U6984 ( .CLK(n1971), .C(n7068) );
  CKBD0 U6985 ( .CLK(n1366), .C(n7069) );
  CKBD0 U6986 ( .CLK(n2359), .C(n7070) );
  CKBD0 U6987 ( .CLK(n1657), .C(n7071) );
  CKBD0 U6988 ( .CLK(n1240), .C(n7072) );
  CKBD0 U6989 ( .CLK(n916), .C(n7073) );
  CKBD0 U6990 ( .CLK(n227), .C(n7074) );
  CKBD0 U6991 ( .CLK(n1560), .C(n7075) );
  CKBD0 U6992 ( .CLK(n919), .C(n7076) );
  CKBD0 U6993 ( .CLK(n1859), .C(n7077) );
  CKBD0 U6994 ( .CLK(n818), .C(n7078) );
  CKBD0 U6995 ( .CLK(n1030), .C(n7079) );
  CKBD0 U6996 ( .CLK(n718), .C(n7080) );
  CKBD0 U6997 ( .CLK(n1761), .C(n7081) );
  CKBD0 U6998 ( .CLK(n1128), .C(n7082) );
  CKBD0 U6999 ( .CLK(n523), .C(n7083) );
  CKBD0 U7000 ( .CLK(n2553), .C(n7084) );
  BUFFD0 U7001 ( .I(n620), .Z(n7085) );
  CKBD0 U7002 ( .CLK(n328), .C(n7086) );
  BUFFD0 U7003 ( .I(n425), .Z(n7087) );
  CKBD0 U7004 ( .CLK(n2456), .C(n7088) );
  CKBD0 U7005 ( .CLK(n1463), .C(n7089) );
  CKBD0 U7006 ( .CLK(n1864), .C(n7090) );
  CKBD0 U7007 ( .CLK(n1660), .C(n7091) );
  CKBD0 U7008 ( .CLK(n1870), .C(n7092) );
  CKBD0 U7009 ( .CLK(n1664), .C(n7093) );
  CKBD0 U7010 ( .CLK(n1867), .C(n7094) );
  CKBD0 U7011 ( .CLK(n1874), .C(n7095) );
  CKBD0 U7012 ( .CLK(n7064), .C(n7096) );
  CKBD0 U7013 ( .CLK(n7065), .C(n7097) );
  CKBD0 U7014 ( .CLK(n7066), .C(n7098) );
  BUFFD0 U7015 ( .I(n7067), .Z(n7099) );
  CKBD0 U7016 ( .CLK(n7068), .C(n7100) );
  CKBD0 U7017 ( .CLK(n7070), .C(n7101) );
  CKBD0 U7018 ( .CLK(n7069), .C(n7102) );
  CKBD0 U7019 ( .CLK(n7071), .C(n7103) );
  BUFFD0 U7020 ( .I(n7072), .Z(n7104) );
  CKBD0 U7021 ( .CLK(n7073), .C(n7105) );
  CKBD0 U7022 ( .CLK(n7074), .C(n7106) );
  CKBD0 U7023 ( .CLK(n7077), .C(n7107) );
  CKBD0 U7024 ( .CLK(n7075), .C(n7108) );
  CKBD0 U7025 ( .CLK(n7076), .C(n7109) );
  CKBD0 U7026 ( .CLK(n7078), .C(n7110) );
  CKBD0 U7027 ( .CLK(n7080), .C(n7111) );
  CKBD0 U7028 ( .CLK(n7079), .C(n7112) );
  CKBD0 U7029 ( .CLK(n7081), .C(n7113) );
  CKBD0 U7030 ( .CLK(n7082), .C(n7114) );
  CKBD0 U7031 ( .CLK(n7083), .C(n7115) );
  CKBD0 U7032 ( .CLK(n7084), .C(n7116) );
  CKBD0 U7033 ( .CLK(n7086), .C(n7117) );
  CKBD0 U7034 ( .CLK(n7085), .C(n7118) );
  CKBD0 U7035 ( .CLK(n7087), .C(n7119) );
  CKBD0 U7036 ( .CLK(n7088), .C(n7120) );
  CKBD0 U7037 ( .CLK(n7089), .C(n7121) );
  CKBD0 U7038 ( .CLK(n7090), .C(n7122) );
  CKBD0 U7039 ( .CLK(n7091), .C(n7123) );
  CKBD0 U7040 ( .CLK(n7092), .C(n7124) );
  CKBD0 U7041 ( .CLK(n7093), .C(n7125) );
  CKBD0 U7042 ( .CLK(n7094), .C(n7126) );
  CKBD0 U7043 ( .CLK(n7095), .C(n7127) );
  CKBD0 U7044 ( .CLK(n7096), .C(n7128) );
  CKBD0 U7045 ( .CLK(n7097), .C(n7129) );
  CKBD0 U7046 ( .CLK(n7098), .C(n7130) );
  CKBD0 U7047 ( .CLK(n7099), .C(n7131) );
  CKBD0 U7048 ( .CLK(n7100), .C(n7132) );
  CKBD0 U7049 ( .CLK(n7103), .C(n7133) );
  CKBD0 U7050 ( .CLK(n7101), .C(n7134) );
  CKBD0 U7051 ( .CLK(n7102), .C(n7135) );
  CKBD0 U7052 ( .CLK(n7104), .C(n7136) );
  BUFFD0 U7053 ( .I(n7105), .Z(n7137) );
  CKBD0 U7054 ( .CLK(n7106), .C(n7138) );
  CKBD0 U7055 ( .CLK(n7108), .C(n7139) );
  BUFFD0 U7056 ( .I(n7107), .Z(n7140) );
  CKBD0 U7057 ( .CLK(n7109), .C(n7141) );
  BUFFD0 U7058 ( .I(n7110), .Z(n7142) );
  CKBD0 U7059 ( .CLK(n7112), .C(n7143) );
  BUFFD0 U7060 ( .I(n7111), .Z(n7144) );
  CKBD0 U7061 ( .CLK(n7113), .C(n7145) );
  BUFFD0 U7062 ( .I(n7114), .Z(n7146) );
  BUFFD0 U7063 ( .I(n7115), .Z(n7147) );
  CKBD0 U7064 ( .CLK(n7116), .C(n7148) );
  BUFFD0 U7065 ( .I(n7117), .Z(n7149) );
  CKBD0 U7066 ( .CLK(n7118), .C(n7150) );
  CKBD0 U7067 ( .CLK(n7119), .C(n7151) );
  CKBD0 U7068 ( .CLK(n7120), .C(n7152) );
  CKBD0 U7069 ( .CLK(n7121), .C(n7153) );
  CKBD0 U7070 ( .CLK(n7122), .C(n7154) );
  CKBD0 U7071 ( .CLK(n7123), .C(n7155) );
  CKBD0 U7072 ( .CLK(n7124), .C(n7156) );
  CKBD0 U7073 ( .CLK(n7125), .C(n7157) );
  CKBD0 U7074 ( .CLK(n7126), .C(n7158) );
  CKBD0 U7075 ( .CLK(n7127), .C(n7159) );
  BUFFD0 U7076 ( .I(n7128), .Z(n7160) );
  BUFFD0 U7077 ( .I(n7129), .Z(n7161) );
  CKBD0 U7078 ( .CLK(n7130), .C(n7162) );
  CKBD0 U7079 ( .CLK(n7131), .C(n7163) );
  CKBD0 U7080 ( .CLK(n7132), .C(n7164) );
  CKBD0 U7081 ( .CLK(n7134), .C(n7165) );
  BUFFD0 U7082 ( .I(n7133), .Z(n7166) );
  CKBD0 U7083 ( .CLK(n7135), .C(n7167) );
  CKBD0 U7084 ( .CLK(n7136), .C(n7168) );
  CKBD0 U7085 ( .CLK(n7138), .C(n7169) );
  CKBD0 U7086 ( .CLK(n7137), .C(n7170) );
  BUFFD0 U7087 ( .I(n7139), .Z(n7171) );
  CKBD0 U7088 ( .CLK(n7140), .C(n7172) );
  CKBD0 U7089 ( .CLK(n7142), .C(n7173) );
  CKBD0 U7090 ( .CLK(n7141), .C(n7174) );
  CKBD0 U7091 ( .CLK(n7143), .C(n7175) );
  CKBD0 U7092 ( .CLK(n7144), .C(n7176) );
  BUFFD0 U7093 ( .I(n7145), .Z(n7177) );
  CKBD0 U7094 ( .CLK(n7146), .C(n7178) );
  CKBD0 U7095 ( .CLK(n7147), .C(n7179) );
  BUFFD0 U7096 ( .I(n7148), .Z(n7180) );
  CKBD0 U7097 ( .CLK(n7149), .C(n7181) );
  CKBD0 U7098 ( .CLK(n7150), .C(n7182) );
  CKBD0 U7099 ( .CLK(n7151), .C(n7183) );
  CKBD0 U7100 ( .CLK(n7152), .C(n7184) );
  CKBD0 U7101 ( .CLK(n7153), .C(n7185) );
  CKBD0 U7102 ( .CLK(n7154), .C(n7186) );
  CKBD0 U7103 ( .CLK(n7155), .C(n7187) );
  CKBD0 U7104 ( .CLK(n7156), .C(n7188) );
  CKBD0 U7105 ( .CLK(n7157), .C(n7189) );
  CKBD0 U7106 ( .CLK(n7158), .C(n7190) );
  CKBD0 U7107 ( .CLK(n7159), .C(n7191) );
  CKBD0 U7108 ( .CLK(n7160), .C(n7192) );
  CKBD0 U7109 ( .CLK(n7161), .C(n7193) );
  BUFFD0 U7110 ( .I(n7162), .Z(n7194) );
  CKBD0 U7111 ( .CLK(n7163), .C(n7195) );
  BUFFD0 U7112 ( .I(n7164), .Z(n7196) );
  BUFFD0 U7113 ( .I(n7165), .Z(n7197) );
  CKBD0 U7114 ( .CLK(n7166), .C(n7198) );
  CKBD0 U7115 ( .CLK(n7168), .C(n7199) );
  CKBD0 U7116 ( .CLK(n7167), .C(n7200) );
  CKBD0 U7117 ( .CLK(n7170), .C(n7201) );
  BUFFD0 U7118 ( .I(n7169), .Z(n7202) );
  CKBD0 U7119 ( .CLK(n7171), .C(n7203) );
  CKBD0 U7120 ( .CLK(n7172), .C(n7204) );
  CKBD0 U7121 ( .CLK(n7173), .C(n7205) );
  CKBD0 U7122 ( .CLK(n7174), .C(n7206) );
  BUFFD0 U7123 ( .I(n7175), .Z(n7207) );
  CKBD0 U7124 ( .CLK(n7176), .C(n7208) );
  CKBD0 U7125 ( .CLK(n7177), .C(n7209) );
  CKBD0 U7126 ( .CLK(n7178), .C(n7210) );
  CKBD0 U7127 ( .CLK(n7179), .C(n7211) );
  CKBD0 U7128 ( .CLK(n7180), .C(n7212) );
  CKBD0 U7129 ( .CLK(n7181), .C(n7213) );
  CKBD0 U7130 ( .CLK(n7182), .C(n7214) );
  CKBD0 U7131 ( .CLK(n7183), .C(n7215) );
  CKBD0 U7132 ( .CLK(n7184), .C(n7216) );
  BUFFD0 U7133 ( .I(n7185), .Z(n7217) );
  CKBD0 U7134 ( .CLK(n7186), .C(n7218) );
  CKBD0 U7135 ( .CLK(n7187), .C(n7219) );
  CKBD0 U7136 ( .CLK(n7188), .C(n7220) );
  CKBD0 U7137 ( .CLK(n7189), .C(n7221) );
  CKBD0 U7138 ( .CLK(n7190), .C(n7222) );
  CKBD0 U7139 ( .CLK(n7191), .C(n7223) );
  CKBD0 U7140 ( .CLK(n7192), .C(n7224) );
  CKBD0 U7141 ( .CLK(n7193), .C(n7225) );
  CKBD0 U7142 ( .CLK(n7194), .C(n7226) );
  CKBD0 U7143 ( .CLK(n7195), .C(n7227) );
  CKBD0 U7144 ( .CLK(n7196), .C(n7228) );
  CKBD0 U7145 ( .CLK(n7197), .C(n7229) );
  CKBD0 U7146 ( .CLK(n7198), .C(n7230) );
  CKBD0 U7147 ( .CLK(n7199), .C(n7231) );
  CKBD0 U7148 ( .CLK(n7200), .C(n7232) );
  CKBD0 U7149 ( .CLK(n7201), .C(n7233) );
  CKBD0 U7150 ( .CLK(n7202), .C(n7234) );
  CKBD0 U7151 ( .CLK(n7203), .C(n7235) );
  CKBD0 U7152 ( .CLK(n7204), .C(n7236) );
  CKBD0 U7153 ( .CLK(n7205), .C(n7237) );
  CKBD0 U7154 ( .CLK(n7207), .C(n7238) );
  CKBD0 U7155 ( .CLK(n7206), .C(n7239) );
  CKBD0 U7156 ( .CLK(n7208), .C(n7240) );
  CKBD0 U7157 ( .CLK(n7209), .C(n7241) );
  CKBD0 U7158 ( .CLK(n7210), .C(n7242) );
  CKBD0 U7159 ( .CLK(n7211), .C(n7243) );
  CKBD0 U7160 ( .CLK(n7212), .C(n7244) );
  CKBD0 U7161 ( .CLK(n7213), .C(n7245) );
  CKBD0 U7162 ( .CLK(n7214), .C(n7246) );
  CKBD0 U7163 ( .CLK(n7215), .C(n7247) );
  CKBD0 U7164 ( .CLK(n7216), .C(n7248) );
  CKBD0 U7165 ( .CLK(n7217), .C(n7249) );
  CKBD0 U7166 ( .CLK(n7218), .C(n7250) );
  CKBD0 U7167 ( .CLK(n7219), .C(n7251) );
  CKBD0 U7168 ( .CLK(n7220), .C(n7252) );
  CKBD0 U7169 ( .CLK(n7221), .C(n7253) );
  CKBD0 U7170 ( .CLK(n7222), .C(n7254) );
  CKBD0 U7171 ( .CLK(n7223), .C(n7255) );
  CKBD0 U7172 ( .CLK(n7224), .C(n7256) );
  CKBD0 U7173 ( .CLK(n7225), .C(n7257) );
  CKBD0 U7174 ( .CLK(n7226), .C(n7258) );
  CKBD0 U7175 ( .CLK(n7227), .C(n7259) );
  CKBD0 U7176 ( .CLK(n7228), .C(n7260) );
  CKBD0 U7177 ( .CLK(n7229), .C(n7261) );
  CKBD0 U7178 ( .CLK(n7230), .C(n7262) );
  CKBD0 U7179 ( .CLK(n7231), .C(n7263) );
  CKBD0 U7180 ( .CLK(n7233), .C(n7264) );
  CKBD0 U7181 ( .CLK(n7234), .C(n7265) );
  CKBD0 U7182 ( .CLK(n7232), .C(n7266) );
  CKBD0 U7183 ( .CLK(n7235), .C(n7267) );
  CKBD0 U7184 ( .CLK(n7236), .C(n7268) );
  CKBD0 U7185 ( .CLK(n7237), .C(n7269) );
  CKBD0 U7186 ( .CLK(n7238), .C(n7270) );
  CKBD0 U7187 ( .CLK(n7239), .C(n7271) );
  CKBD0 U7188 ( .CLK(n7240), .C(n7272) );
  CKBD0 U7189 ( .CLK(n7241), .C(n7273) );
  CKBD0 U7190 ( .CLK(n7242), .C(n7274) );
  CKBD0 U7191 ( .CLK(n7243), .C(n7275) );
  CKBD0 U7192 ( .CLK(n7244), .C(n7276) );
  CKBD0 U7193 ( .CLK(n7245), .C(n7277) );
  CKBD0 U7194 ( .CLK(n7246), .C(n7278) );
  CKBD0 U7195 ( .CLK(n7247), .C(n7279) );
  CKBD0 U7196 ( .CLK(n7248), .C(n7280) );
  CKBD0 U7197 ( .CLK(n7249), .C(n7281) );
  CKBD0 U7198 ( .CLK(n7250), .C(n7282) );
  CKBD0 U7199 ( .CLK(n7251), .C(n7283) );
  CKBD0 U7200 ( .CLK(n7252), .C(n7284) );
  CKBD0 U7201 ( .CLK(n7253), .C(n7285) );
  CKBD0 U7202 ( .CLK(n7254), .C(n7286) );
  CKBD0 U7203 ( .CLK(n7255), .C(n7287) );
  CKBD0 U7204 ( .CLK(n7256), .C(n7288) );
  CKBD0 U7205 ( .CLK(n7257), .C(n7289) );
  CKBD0 U7206 ( .CLK(n7258), .C(n7290) );
  CKBD0 U7207 ( .CLK(n7259), .C(n7291) );
  CKBD0 U7208 ( .CLK(n7260), .C(n7292) );
  CKBD0 U7209 ( .CLK(n7261), .C(n7293) );
  CKBD0 U7210 ( .CLK(n7262), .C(n7294) );
  CKBD0 U7211 ( .CLK(n7263), .C(n7295) );
  CKBD0 U7212 ( .CLK(n7266), .C(n7296) );
  CKBD0 U7213 ( .CLK(n7264), .C(n7297) );
  CKBD0 U7214 ( .CLK(n7265), .C(n7298) );
  CKBD0 U7215 ( .CLK(n7267), .C(n7299) );
  CKBD0 U7216 ( .CLK(n7268), .C(n7300) );
  CKBD0 U7217 ( .CLK(n7269), .C(n7301) );
  CKBD0 U7218 ( .CLK(n7270), .C(n7302) );
  CKBD0 U7219 ( .CLK(n7272), .C(n7303) );
  CKBD0 U7220 ( .CLK(n7273), .C(n7304) );
  CKBD0 U7221 ( .CLK(n7271), .C(n7305) );
  CKBD0 U7222 ( .CLK(n7274), .C(n7306) );
  CKBD0 U7223 ( .CLK(n7275), .C(n7307) );
  CKBD0 U7224 ( .CLK(n7276), .C(n7308) );
  CKBD0 U7225 ( .CLK(n7277), .C(n7309) );
  CKBD0 U7226 ( .CLK(n7278), .C(n7310) );
  CKBD0 U7227 ( .CLK(n7279), .C(n7311) );
  CKBD0 U7228 ( .CLK(n7280), .C(n7312) );
  CKBD0 U7229 ( .CLK(n7281), .C(n7313) );
  CKBD0 U7230 ( .CLK(n7282), .C(n7314) );
  CKBD0 U7231 ( .CLK(n7283), .C(n7315) );
  CKBD0 U7232 ( .CLK(n7284), .C(n7316) );
  CKBD0 U7233 ( .CLK(n7285), .C(n7317) );
  CKBD0 U7234 ( .CLK(n7286), .C(n7318) );
  CKBD0 U7235 ( .CLK(n7288), .C(n7319) );
  CKBD0 U7236 ( .CLK(n7287), .C(n7320) );
  CKBD0 U7237 ( .CLK(n7289), .C(n7321) );
  CKBD0 U7238 ( .CLK(n7290), .C(n7322) );
  BUFFD0 U7239 ( .I(n7296), .Z(n7323) );
  CKBD0 U7240 ( .CLK(n7291), .C(n7324) );
  CKBD0 U7241 ( .CLK(n7292), .C(n7325) );
  CKBD0 U7242 ( .CLK(n7293), .C(n7326) );
  CKBD0 U7243 ( .CLK(n7294), .C(n7327) );
  CKBD0 U7244 ( .CLK(n7295), .C(n7328) );
  CKBD0 U7245 ( .CLK(n7297), .C(n7329) );
  CKBD0 U7246 ( .CLK(n7298), .C(n7330) );
  CKBD0 U7247 ( .CLK(n7299), .C(n7331) );
  CKBD0 U7248 ( .CLK(n7300), .C(n7332) );
  CKBD0 U7249 ( .CLK(n7301), .C(n7333) );
  CKBD0 U7250 ( .CLK(n7302), .C(n7334) );
  CKBD0 U7251 ( .CLK(n7303), .C(n7335) );
  CKBD0 U7252 ( .CLK(n7304), .C(n7336) );
  CKBD0 U7253 ( .CLK(n7305), .C(n7337) );
  CKBD0 U7254 ( .CLK(n7306), .C(n7338) );
  CKBD0 U7255 ( .CLK(n7307), .C(n7339) );
  CKBD0 U7256 ( .CLK(n7308), .C(n7340) );
  CKBD0 U7257 ( .CLK(n7309), .C(n7341) );
  CKBD0 U7258 ( .CLK(n7310), .C(n7342) );
  CKBD0 U7259 ( .CLK(n7311), .C(n7343) );
  CKBD0 U7260 ( .CLK(n7312), .C(n7344) );
  CKBD0 U7261 ( .CLK(n7313), .C(n7345) );
  BUFFD0 U7262 ( .I(n7314), .Z(n7346) );
  BUFFD0 U7263 ( .I(n7315), .Z(n7347) );
  BUFFD0 U7264 ( .I(n7316), .Z(n7348) );
  CKBD0 U7265 ( .CLK(n7317), .C(n7349) );
  BUFFD0 U7266 ( .I(n7318), .Z(n7350) );
  CKBD0 U7267 ( .CLK(n7319), .C(n7351) );
  CKBD0 U7268 ( .CLK(n7320), .C(n7352) );
  CKBD0 U7269 ( .CLK(n7321), .C(n7353) );
  CKBD0 U7270 ( .CLK(n7322), .C(n7354) );
  CKBD0 U7271 ( .CLK(n7324), .C(n7355) );
  CKBD0 U7272 ( .CLK(n7323), .C(n7356) );
  CKBD0 U7273 ( .CLK(n7325), .C(n7357) );
  CKBD0 U7274 ( .CLK(n7326), .C(n7358) );
  CKBD0 U7275 ( .CLK(n7327), .C(n7359) );
  CKBD0 U7276 ( .CLK(n7328), .C(n7360) );
  CKBD0 U7277 ( .CLK(n7329), .C(n7361) );
  CKBD0 U7278 ( .CLK(n7330), .C(n7362) );
  CKBD0 U7279 ( .CLK(n7331), .C(n7363) );
  CKBD0 U7280 ( .CLK(n7332), .C(n7364) );
  CKBD0 U7281 ( .CLK(n7333), .C(n7365) );
  CKBD0 U7282 ( .CLK(n7334), .C(n7366) );
  CKBD0 U7283 ( .CLK(n7335), .C(n7367) );
  CKBD0 U7284 ( .CLK(n7336), .C(n7368) );
  CKBD0 U7285 ( .CLK(n7337), .C(n7369) );
  CKBD0 U7286 ( .CLK(n7338), .C(n7370) );
  CKBD0 U7287 ( .CLK(n7339), .C(n7371) );
  CKBD0 U7288 ( .CLK(n7340), .C(n7372) );
  CKBD0 U7289 ( .CLK(n7341), .C(n7373) );
  CKBD0 U7290 ( .CLK(n7342), .C(n7374) );
  CKBD0 U7291 ( .CLK(n7343), .C(n7375) );
  CKBD0 U7292 ( .CLK(n7344), .C(n7376) );
  CKBD0 U7293 ( .CLK(n7345), .C(n7377) );
  CKBD0 U7294 ( .CLK(n7346), .C(n7378) );
  CKBD0 U7295 ( .CLK(n7347), .C(n7379) );
  CKBD0 U7296 ( .CLK(n7348), .C(n7380) );
  CKBD0 U7297 ( .CLK(n7349), .C(n7381) );
  CKBD0 U7298 ( .CLK(n7350), .C(n7382) );
  CKBD0 U7299 ( .CLK(n7351), .C(n7383) );
  CKBD0 U7300 ( .CLK(n7352), .C(n7384) );
  CKBD0 U7301 ( .CLK(n7353), .C(n7385) );
  CKBD0 U7302 ( .CLK(n7354), .C(n7386) );
  CKBD0 U7303 ( .CLK(n7355), .C(n7387) );
  CKBD0 U7304 ( .CLK(n7356), .C(n7388) );
  CKBD0 U7305 ( .CLK(n7357), .C(n7389) );
  CKBD0 U7306 ( .CLK(n7358), .C(n7390) );
  CKBD0 U7307 ( .CLK(n7359), .C(n7391) );
  CKBD0 U7308 ( .CLK(n7360), .C(n7392) );
  CKBD0 U7309 ( .CLK(n7361), .C(n7393) );
  CKBD0 U7310 ( .CLK(n7362), .C(n7394) );
  BUFFD0 U7311 ( .I(n7369), .Z(n7395) );
  CKBD0 U7312 ( .CLK(n7363), .C(n7396) );
  CKBD0 U7313 ( .CLK(n7364), .C(n7397) );
  CKBD0 U7314 ( .CLK(n7365), .C(n7398) );
  CKBD0 U7315 ( .CLK(n7366), .C(n7399) );
  CKBD0 U7316 ( .CLK(n7367), .C(n7400) );
  CKBD0 U7317 ( .CLK(n7368), .C(n7401) );
  CKBD0 U7318 ( .CLK(n7370), .C(n7402) );
  CKBD0 U7319 ( .CLK(n7371), .C(n7403) );
  CKBD0 U7320 ( .CLK(n7372), .C(n7404) );
  CKBD0 U7321 ( .CLK(n7373), .C(n7405) );
  CKBD0 U7322 ( .CLK(n7374), .C(n7406) );
  CKBD0 U7323 ( .CLK(n7375), .C(n7407) );
  CKBD0 U7324 ( .CLK(n7376), .C(n7408) );
  CKBD0 U7325 ( .CLK(n7377), .C(n7409) );
  CKBD0 U7326 ( .CLK(n7378), .C(n7410) );
  CKBD0 U7327 ( .CLK(n7379), .C(n7411) );
  CKBD0 U7328 ( .CLK(n7380), .C(n7412) );
  BUFFD0 U7329 ( .I(n7381), .Z(n7413) );
  CKBD0 U7330 ( .CLK(n7382), .C(n7414) );
  BUFFD0 U7331 ( .I(n7384), .Z(n7415) );
  CKBD0 U7332 ( .CLK(n7383), .C(n7416) );
  CKBD0 U7333 ( .CLK(n7385), .C(n7417) );
  CKBD0 U7334 ( .CLK(n7386), .C(n7418) );
  CKBD0 U7335 ( .CLK(n7387), .C(n7419) );
  CKBD0 U7336 ( .CLK(n7389), .C(n7420) );
  CKBD0 U7337 ( .CLK(n7388), .C(n7421) );
  CKBD0 U7338 ( .CLK(n7390), .C(n7422) );
  CKBD0 U7339 ( .CLK(n7391), .C(n7423) );
  CKBD0 U7340 ( .CLK(n7392), .C(n7424) );
  CKBD0 U7341 ( .CLK(n7393), .C(n7425) );
  CKBD0 U7342 ( .CLK(n7394), .C(n7426) );
  CKBD0 U7343 ( .CLK(n7397), .C(n7427) );
  CKBD0 U7344 ( .CLK(n7396), .C(n7428) );
  CKBD0 U7345 ( .CLK(n7395), .C(n7429) );
  CKBD0 U7346 ( .CLK(n7398), .C(n7430) );
  CKBD0 U7347 ( .CLK(n7399), .C(n7431) );
  CKBD0 U7348 ( .CLK(n7400), .C(n7432) );
  CKBD0 U7349 ( .CLK(n7401), .C(n7433) );
  CKBD0 U7350 ( .CLK(n7402), .C(n7434) );
  CKBD0 U7351 ( .CLK(n7403), .C(n7435) );
  CKBD0 U7352 ( .CLK(n7404), .C(n7436) );
  CKBD0 U7353 ( .CLK(n7405), .C(n7437) );
  BUFFD0 U7354 ( .I(n7408), .Z(n7438) );
  CKBD0 U7355 ( .CLK(n7406), .C(n7439) );
  CKBD0 U7356 ( .CLK(n7407), .C(n7440) );
  CKBD0 U7357 ( .CLK(n7409), .C(n7441) );
  CKBD0 U7358 ( .CLK(n7416), .C(n7442) );
  CKBD0 U7359 ( .CLK(n7417), .C(n7443) );
  CKBD0 U7360 ( .CLK(n7418), .C(n7444) );
  BUFFD0 U7361 ( .I(n7419), .Z(n7445) );
  CKBD0 U7362 ( .CLK(n7420), .C(n7446) );
  CKBD0 U7363 ( .CLK(n7422), .C(n7447) );
  CKBD0 U7364 ( .CLK(n7423), .C(n7448) );
  BUFFD0 U7365 ( .I(n7424), .Z(n7449) );
  CKBD0 U7366 ( .CLK(n7425), .C(n7450) );
  CKBD0 U7367 ( .CLK(n7426), .C(n7451) );
  CKBD0 U7368 ( .CLK(n7428), .C(n7452) );
  BUFFD0 U7369 ( .I(n7427), .Z(n7453) );
  CKBD0 U7370 ( .CLK(n7430), .C(n7454) );
  CKBD0 U7371 ( .CLK(n7432), .C(n7455) );
  CKBD0 U7372 ( .CLK(n7431), .C(n7456) );
  CKBD0 U7373 ( .CLK(n7433), .C(n7457) );
  CKBD0 U7374 ( .CLK(n7434), .C(n7458) );
  CKBD0 U7375 ( .CLK(n7435), .C(n7459) );
  CKBD0 U7376 ( .CLK(n7436), .C(n7460) );
  CKBD0 U7377 ( .CLK(n7437), .C(n7461) );
  BUFFD0 U7378 ( .I(n7439), .Z(n7462) );
  BUFFD0 U7379 ( .I(n7440), .Z(n7463) );
  CKBD0 U7380 ( .CLK(n7438), .C(n7464) );
  CKBD0 U7381 ( .CLK(n7441), .C(n7465) );
  CKBD0 U7382 ( .CLK(n7410), .C(n7466) );
  CKBD0 U7383 ( .CLK(n7442), .C(n7467) );
  CKBD0 U7384 ( .CLK(n7443), .C(n7468) );
  CKBD0 U7385 ( .CLK(n7444), .C(n7469) );
  CKBD0 U7386 ( .CLK(n7411), .C(n7470) );
  CKBD0 U7387 ( .CLK(n7412), .C(n7471) );
  CKBD0 U7388 ( .CLK(n7445), .C(n7472) );
  CKBD0 U7389 ( .CLK(n7446), .C(n7473) );
  CKBD0 U7390 ( .CLK(n7447), .C(n7474) );
  CKBD0 U7391 ( .CLK(n7413), .C(n7475) );
  CKBD0 U7392 ( .CLK(n7448), .C(n7476) );
  CKBD0 U7393 ( .CLK(n7449), .C(n7477) );
  CKBD0 U7394 ( .CLK(n7451), .C(n7478) );
  BUFFD0 U7395 ( .I(n7450), .Z(n7479) );
  CKBD0 U7396 ( .CLK(n7414), .C(n7480) );
  CKBD0 U7397 ( .CLK(n7415), .C(n7481) );
  CKBD0 U7398 ( .CLK(n7421), .C(n7482) );
  CKBD0 U7399 ( .CLK(n7429), .C(n7483) );
  CKBD0 U7400 ( .CLK(n7466), .C(n7484) );
  CKBD0 U7401 ( .CLK(n7452), .C(n7485) );
  CKBD0 U7402 ( .CLK(n7453), .C(n7486) );
  BUFFD0 U7403 ( .I(n7454), .Z(n7487) );
  CKBD0 U7404 ( .CLK(n7456), .C(n7488) );
  BUFFD0 U7405 ( .I(n7455), .Z(n7489) );
  CKBD0 U7406 ( .CLK(n7457), .C(n7490) );
  CKBD0 U7407 ( .CLK(n7470), .C(n7491) );
  CKBD0 U7408 ( .CLK(n7471), .C(n7492) );
  BUFFD0 U7409 ( .I(n7458), .Z(n7493) );
  CKBD0 U7410 ( .CLK(n7475), .C(n7494) );
  CKBD0 U7411 ( .CLK(n7480), .C(n7495) );
  CKBD0 U7412 ( .CLK(n7481), .C(n7496) );
  CKBD0 U7413 ( .CLK(n7482), .C(n7497) );
  CKBD0 U7414 ( .CLK(n7483), .C(n7498) );
  CKBD0 U7415 ( .CLK(n7484), .C(n7499) );
  BUFFD0 U7416 ( .I(n7459), .Z(n7500) );
  CKBD0 U7417 ( .CLK(n7460), .C(n7501) );
  CKBD0 U7418 ( .CLK(n7491), .C(n7502) );
  BUFFD0 U7419 ( .I(n7461), .Z(n7503) );
  CKBD0 U7420 ( .CLK(n7492), .C(n7504) );
  CKBD0 U7421 ( .CLK(n7462), .C(n7505) );
  CKBD0 U7422 ( .CLK(n7494), .C(n7506) );
  CKBD0 U7423 ( .CLK(n7495), .C(n7507) );
  CKBD0 U7424 ( .CLK(n7496), .C(n7508) );
  CKBD0 U7425 ( .CLK(n7497), .C(n7509) );
  CKBD0 U7426 ( .CLK(n7498), .C(n7510) );
  CKBD0 U7427 ( .CLK(n7499), .C(n7511) );
  CKBD0 U7428 ( .CLK(n7463), .C(n7512) );
  CKBD0 U7429 ( .CLK(n7464), .C(n7513) );
  CKBD0 U7430 ( .CLK(n7502), .C(n7514) );
  CKBD0 U7431 ( .CLK(n7504), .C(n7515) );
  CKBD0 U7432 ( .CLK(n7506), .C(n7516) );
  CKBD0 U7433 ( .CLK(n7507), .C(n7517) );
  CKBD0 U7434 ( .CLK(n7508), .C(n7518) );
  CKBD0 U7435 ( .CLK(n7509), .C(n7519) );
  CKBD0 U7436 ( .CLK(n7510), .C(n7520) );
  CKBD0 U7437 ( .CLK(n7511), .C(n7521) );
  CKBD0 U7438 ( .CLK(n7514), .C(n7522) );
  CKBD0 U7439 ( .CLK(n7515), .C(n7523) );
  CKBD0 U7440 ( .CLK(n7465), .C(n7524) );
  CKBD0 U7441 ( .CLK(n7516), .C(n7525) );
  CKBD0 U7442 ( .CLK(n7517), .C(n7526) );
  CKBD0 U7443 ( .CLK(n7518), .C(n7527) );
  CKBD0 U7444 ( .CLK(n7467), .C(n7528) );
  CKBD0 U7445 ( .CLK(n7519), .C(n7529) );
  BUFFD0 U7446 ( .I(n7468), .Z(n7530) );
  BUFFD0 U7447 ( .I(n7469), .Z(n7531) );
  CKBD0 U7448 ( .CLK(n7472), .C(n7532) );
  BUFFD0 U7449 ( .I(n7473), .Z(n7533) );
  BUFFD0 U7450 ( .I(n7474), .Z(n7534) );
  CKBD0 U7451 ( .CLK(n7476), .C(n7535) );
  CKBD0 U7452 ( .CLK(n7520), .C(n7536) );
  CKBD0 U7453 ( .CLK(n7521), .C(n7537) );
  CKBD0 U7454 ( .CLK(n7522), .C(n7538) );
  CKBD0 U7455 ( .CLK(n7523), .C(n7539) );
  CKBD0 U7456 ( .CLK(n7525), .C(n7540) );
  CKBD0 U7457 ( .CLK(n7526), .C(n7541) );
  CKBD0 U7458 ( .CLK(n7527), .C(n7542) );
  CKBD0 U7459 ( .CLK(n7529), .C(n7543) );
  CKBD0 U7460 ( .CLK(n7477), .C(n7544) );
  CKBD0 U7461 ( .CLK(n7479), .C(n7545) );
  BUFFD0 U7462 ( .I(n7478), .Z(n7546) );
  CKBD0 U7463 ( .CLK(n7485), .C(n7547) );
  CKBD0 U7464 ( .CLK(n7486), .C(n7548) );
  CKBD0 U7465 ( .CLK(n7536), .C(n7549) );
  CKBD0 U7466 ( .CLK(n7537), .C(n7550) );
  CKBD0 U7467 ( .CLK(n7538), .C(n7551) );
  CKBD0 U7468 ( .CLK(n7539), .C(n7552) );
  CKBD0 U7469 ( .CLK(n7540), .C(n7553) );
  CKBD0 U7470 ( .CLK(n7541), .C(n7554) );
  CKBD0 U7471 ( .CLK(n7542), .C(n7555) );
  CKBD0 U7472 ( .CLK(n7543), .C(n7556) );
  CKBD0 U7473 ( .CLK(n7487), .C(n7557) );
  BUFFD0 U7474 ( .I(n7488), .Z(n7558) );
  CKBD0 U7475 ( .CLK(n7489), .C(n7559) );
  BUFFD0 U7476 ( .I(n7490), .Z(n7560) );
  CKBD0 U7477 ( .CLK(n7493), .C(n7561) );
  CKBD0 U7478 ( .CLK(n7500), .C(n7562) );
  CKBD0 U7479 ( .CLK(n7549), .C(n7563) );
  BUFFD0 U7480 ( .I(n7501), .Z(n7564) );
  CKBD0 U7481 ( .CLK(n7503), .C(n7565) );
  CKBD0 U7482 ( .CLK(n7505), .C(n7566) );
  CKBD0 U7483 ( .CLK(n7512), .C(n7567) );
  CKBD0 U7484 ( .CLK(n7513), .C(n7568) );
  CKBD0 U7485 ( .CLK(n7524), .C(n7569) );
  CKBD0 U7486 ( .CLK(n7550), .C(n7570) );
  BUFFD0 U7487 ( .I(n7551), .Z(n7571) );
  BUFFD0 U7488 ( .I(n7552), .Z(n7572) );
  CKBD0 U7489 ( .CLK(n7553), .C(n7573) );
  CKBD0 U7490 ( .CLK(n7554), .C(n7574) );
  BUFFD0 U7491 ( .I(n7528), .Z(n7575) );
  CKBD0 U7492 ( .CLK(n7555), .C(n7576) );
  CKBD0 U7493 ( .CLK(n7530), .C(n7577) );
  CKBD0 U7494 ( .CLK(n7531), .C(n7578) );
  CKBD0 U7495 ( .CLK(n7532), .C(n7579) );
  CKBD0 U7496 ( .CLK(n7533), .C(n7580) );
  CKBD0 U7497 ( .CLK(n7534), .C(n7581) );
  BUFFD0 U7498 ( .I(n7535), .Z(n7582) );
  BUFFD0 U7499 ( .I(n7556), .Z(n7583) );
  CKBD0 U7500 ( .CLK(n7563), .C(n7584) );
  BUFFD0 U7501 ( .I(n7570), .Z(n7585) );
  CKBD0 U7502 ( .CLK(n7571), .C(n7586) );
  CKBD0 U7503 ( .CLK(n7572), .C(n7587) );
  CKBD0 U7504 ( .CLK(n7573), .C(n7588) );
  BUFFD0 U7505 ( .I(n7574), .Z(n7589) );
  CKBD0 U7506 ( .CLK(n7576), .C(n7590) );
  CKBD0 U7507 ( .CLK(n7544), .C(n7591) );
  CKBD0 U7508 ( .CLK(n7545), .C(n7592) );
  CKBD0 U7509 ( .CLK(n7546), .C(n7593) );
  BUFFD0 U7510 ( .I(n7547), .Z(n7594) );
  CKBD0 U7511 ( .CLK(n7548), .C(n7595) );
  CKBD0 U7512 ( .CLK(n7583), .C(n7596) );
  CKBD0 U7513 ( .CLK(n7584), .C(n7597) );
  CKBD0 U7514 ( .CLK(n7585), .C(n7598) );
  CKBD0 U7515 ( .CLK(n7586), .C(n7599) );
  CKBD0 U7516 ( .CLK(n7587), .C(n7600) );
  CKBD0 U7517 ( .CLK(n7588), .C(n7601) );
  CKBD0 U7518 ( .CLK(n7589), .C(n7602) );
  CKBD0 U7519 ( .CLK(n7590), .C(n7603) );
  CKBD0 U7520 ( .CLK(n7557), .C(n7604) );
  CKBD0 U7521 ( .CLK(n7558), .C(n7605) );
  CKBD0 U7522 ( .CLK(n7559), .C(n7606) );
  CKBD0 U7523 ( .CLK(n7560), .C(n7607) );
  CKBD0 U7524 ( .CLK(n7561), .C(n7608) );
  CKBD0 U7525 ( .CLK(n7562), .C(n7609) );
  CKBD0 U7526 ( .CLK(n7596), .C(n7610) );
  CKBD0 U7527 ( .CLK(n7564), .C(n7611) );
  CKBD0 U7528 ( .CLK(n7565), .C(n7612) );
  CKBD0 U7529 ( .CLK(n7566), .C(n7613) );
  CKBD0 U7530 ( .CLK(n7567), .C(n7614) );
  BUFFD0 U7531 ( .I(n7597), .Z(n7615) );
  CKBD0 U7532 ( .CLK(n7598), .C(n7616) );
  CKBD0 U7533 ( .CLK(n7599), .C(n7617) );
  CKBD0 U7534 ( .CLK(n7600), .C(n7618) );
  BUFFD0 U7535 ( .I(n7601), .Z(n7619) );
  CKBD0 U7536 ( .CLK(n7602), .C(n7620) );
  BUFFD0 U7537 ( .I(n7603), .Z(n7621) );
  CKBD0 U7538 ( .CLK(n7610), .C(n7622) );
  CKBD0 U7539 ( .CLK(n7568), .C(n7623) );
  BUFFD0 U7540 ( .I(n7569), .Z(n7624) );
  CKBD0 U7541 ( .CLK(n7615), .C(n7625) );
  CKBD0 U7542 ( .CLK(n7616), .C(n7626) );
  CKBD0 U7543 ( .CLK(n7617), .C(n7627) );
  CKBD0 U7544 ( .CLK(n7618), .C(n7628) );
  CKBD0 U7545 ( .CLK(n7619), .C(n7629) );
  CKBD0 U7546 ( .CLK(n7620), .C(n7630) );
  CKBD0 U7547 ( .CLK(n7621), .C(n7631) );
  CKBD0 U7548 ( .CLK(n7622), .C(n7632) );
  CKBD0 U7549 ( .CLK(n7625), .C(n7633) );
  CKBD0 U7550 ( .CLK(n7626), .C(n7634) );
  CKBD0 U7551 ( .CLK(n7575), .C(n7635) );
  CKBD0 U7552 ( .CLK(n7577), .C(n7636) );
  CKBD0 U7553 ( .CLK(n7578), .C(n7637) );
  CKBD0 U7554 ( .CLK(n7627), .C(n7638) );
  CKBD0 U7555 ( .CLK(n7628), .C(n7639) );
  CKBD0 U7556 ( .CLK(n7629), .C(n7640) );
  CKBD0 U7557 ( .CLK(n7630), .C(n7641) );
  CKBD0 U7558 ( .CLK(n7631), .C(n7642) );
  CKBD0 U7559 ( .CLK(n7632), .C(n7643) );
  CKBD0 U7560 ( .CLK(n7633), .C(n7644) );
  CKBD0 U7561 ( .CLK(n7634), .C(n7645) );
  CKBD0 U7562 ( .CLK(n7579), .C(n7646) );
  CKBD0 U7563 ( .CLK(n7580), .C(n7647) );
  CKBD0 U7564 ( .CLK(n7581), .C(n7648) );
  CKBD0 U7565 ( .CLK(n7582), .C(n7649) );
  CKBD0 U7566 ( .CLK(n7591), .C(n7650) );
  CKBD0 U7567 ( .CLK(n7638), .C(n7651) );
  CKBD0 U7568 ( .CLK(n7639), .C(n7652) );
  CKBD0 U7569 ( .CLK(n7640), .C(n7653) );
  CKBD0 U7570 ( .CLK(n7641), .C(n7654) );
  CKBD0 U7571 ( .CLK(n7642), .C(n7655) );
  CKBD0 U7572 ( .CLK(n7643), .C(n7656) );
  CKBD0 U7573 ( .CLK(n7644), .C(n7657) );
  CKBD0 U7574 ( .CLK(n7645), .C(n7658) );
  CKBD0 U7575 ( .CLK(n7592), .C(n7659) );
  CKBD0 U7576 ( .CLK(n7593), .C(n7660) );
  CKBD0 U7577 ( .CLK(n7594), .C(n7661) );
  CKBD0 U7578 ( .CLK(n7595), .C(n7662) );
  CKBD0 U7579 ( .CLK(n7604), .C(n7663) );
  CKBD0 U7580 ( .CLK(n7605), .C(n7664) );
  CKBD0 U7581 ( .CLK(n7651), .C(n7665) );
  CKBD0 U7582 ( .CLK(n7652), .C(n7666) );
  CKBD0 U7583 ( .CLK(n7606), .C(n7667) );
  CKBD0 U7584 ( .CLK(n7607), .C(n7668) );
  CKBD0 U7585 ( .CLK(n7653), .C(n7669) );
  CKBD0 U7586 ( .CLK(n7654), .C(n7670) );
  CKBD0 U7587 ( .CLK(n7655), .C(n7671) );
  CKBD0 U7588 ( .CLK(n7656), .C(n7672) );
  CKBD0 U7589 ( .CLK(n7657), .C(n7673) );
  CKBD0 U7590 ( .CLK(n7658), .C(n7674) );
  CKBD0 U7591 ( .CLK(n7608), .C(n7675) );
  CKBD0 U7592 ( .CLK(n7609), .C(n7676) );
  CKBD0 U7593 ( .CLK(n7611), .C(n7677) );
  CKBD0 U7594 ( .CLK(n7665), .C(n7678) );
  CKBD0 U7595 ( .CLK(n7666), .C(n7679) );
  CKBD0 U7596 ( .CLK(n7669), .C(n7680) );
  CKBD0 U7597 ( .CLK(n7670), .C(n7681) );
  CKBD0 U7598 ( .CLK(n7671), .C(n7682) );
  CKBD0 U7599 ( .CLK(n7672), .C(n7683) );
  CKBD0 U7600 ( .CLK(n7673), .C(n7684) );
  CKBD0 U7601 ( .CLK(n7674), .C(n7685) );
  CKBD0 U7602 ( .CLK(n7612), .C(n7686) );
  CKBD0 U7603 ( .CLK(n7613), .C(n7687) );
  CKBD0 U7604 ( .CLK(n7614), .C(n7688) );
  CKBD0 U7605 ( .CLK(n7678), .C(n7689) );
  CKBD0 U7606 ( .CLK(n7679), .C(n7690) );
  CKBD0 U7607 ( .CLK(n7680), .C(n7691) );
  CKBD0 U7608 ( .CLK(n7681), .C(n7692) );
  CKBD0 U7609 ( .CLK(n7682), .C(n7693) );
  CKBD0 U7610 ( .CLK(n7683), .C(n7694) );
  CKBD0 U7611 ( .CLK(n7684), .C(n7695) );
  CKBD0 U7612 ( .CLK(n7685), .C(n7696) );
  CKBD0 U7613 ( .CLK(n7689), .C(n7697) );
  CKBD0 U7614 ( .CLK(n7690), .C(n7698) );
  CKBD0 U7615 ( .CLK(n7691), .C(n7699) );
  CKBD0 U7616 ( .CLK(n7692), .C(n7700) );
  CKBD0 U7617 ( .CLK(n7693), .C(n7701) );
  BUFFD0 U7618 ( .I(n7694), .Z(n7702) );
  CKBD0 U7619 ( .CLK(n7695), .C(n7703) );
  BUFFD0 U7620 ( .I(n7696), .Z(n7704) );
  CKBD0 U7621 ( .CLK(n7623), .C(n7705) );
  CKBD0 U7622 ( .CLK(n7624), .C(n7706) );
  BUFFD0 U7623 ( .I(n7697), .Z(n7707) );
  BUFFD0 U7624 ( .I(n7698), .Z(n7708) );
  CKBD0 U7625 ( .CLK(n7699), .C(n7709) );
  BUFFD0 U7626 ( .I(n7700), .Z(n7710) );
  CKBD0 U7627 ( .CLK(n7701), .C(n7711) );
  CKBD0 U7628 ( .CLK(n7702), .C(n7712) );
  CKBD0 U7629 ( .CLK(n7703), .C(n7713) );
  CKBD0 U7630 ( .CLK(n7704), .C(n7714) );
  CKBD0 U7631 ( .CLK(n7707), .C(n7715) );
  CKBD0 U7632 ( .CLK(n7708), .C(n7716) );
  CKBD0 U7633 ( .CLK(n7709), .C(n7717) );
  CKBD0 U7634 ( .CLK(n7710), .C(n7718) );
  CKBD0 U7635 ( .CLK(n7635), .C(n7719) );
  CKBD0 U7636 ( .CLK(n7711), .C(n7720) );
  CKBD0 U7637 ( .CLK(n7636), .C(n7721) );
  CKBD0 U7638 ( .CLK(n7637), .C(n7722) );
  CKBD0 U7639 ( .CLK(n7646), .C(n7723) );
  CKBD0 U7640 ( .CLK(n7712), .C(n7724) );
  CKBD0 U7641 ( .CLK(n7713), .C(n7725) );
  CKBD0 U7642 ( .CLK(n7714), .C(n7726) );
  CKBD0 U7643 ( .CLK(n7715), .C(n7727) );
  CKBD0 U7644 ( .CLK(n7716), .C(n7728) );
  BUFFD0 U7645 ( .I(n7717), .Z(n7729) );
  CKBD0 U7646 ( .CLK(n7718), .C(n7730) );
  CKBD0 U7647 ( .CLK(n7720), .C(n7731) );
  CKBD0 U7648 ( .CLK(n7647), .C(n7732) );
  CKBD0 U7649 ( .CLK(n7648), .C(n7733) );
  CKBD0 U7650 ( .CLK(n7649), .C(n7734) );
  CKBD0 U7651 ( .CLK(n7650), .C(n7735) );
  CKBD0 U7652 ( .CLK(n7659), .C(n7736) );
  CKBD0 U7653 ( .CLK(n7660), .C(n7737) );
  CKBD0 U7654 ( .CLK(n7661), .C(n7738) );
  CKBD0 U7655 ( .CLK(n7662), .C(n7739) );
  CKBD0 U7656 ( .CLK(n7724), .C(n7740) );
  CKBD0 U7657 ( .CLK(n7663), .C(n7741) );
  CKBD0 U7658 ( .CLK(n7664), .C(n7742) );
  CKBD0 U7659 ( .CLK(n7667), .C(n7743) );
  CKBD0 U7660 ( .CLK(n7668), .C(n7744) );
  CKBD0 U7661 ( .CLK(n7675), .C(n7745) );
  BUFFD0 U7662 ( .I(n7725), .Z(n7746) );
  CKBD0 U7663 ( .CLK(n7726), .C(n7747) );
  CKBD0 U7664 ( .CLK(n7727), .C(n7748) );
  CKBD0 U7665 ( .CLK(n7728), .C(n7749) );
  CKBD0 U7666 ( .CLK(n7729), .C(n7750) );
  CKBD0 U7667 ( .CLK(n7730), .C(n7751) );
  BUFFD0 U7668 ( .I(n7731), .Z(n7752) );
  CKBD0 U7669 ( .CLK(n7740), .C(n7753) );
  CKBD0 U7670 ( .CLK(n7676), .C(n7754) );
  CKBD0 U7671 ( .CLK(n7677), .C(n7755) );
  CKBD0 U7672 ( .CLK(n7686), .C(n7756) );
  CKBD0 U7673 ( .CLK(n7746), .C(n7757) );
  CKBD0 U7674 ( .CLK(n7747), .C(n7758) );
  CKBD0 U7675 ( .CLK(n7748), .C(n7759) );
  CKBD0 U7676 ( .CLK(n7749), .C(n7760) );
  CKBD0 U7677 ( .CLK(n7750), .C(n7761) );
  CKBD0 U7678 ( .CLK(n7751), .C(n7762) );
  CKBD0 U7679 ( .CLK(n7752), .C(n7763) );
  CKBD0 U7680 ( .CLK(n7753), .C(n7764) );
  CKBD0 U7681 ( .CLK(n7687), .C(n7765) );
  CKBD0 U7682 ( .CLK(n7688), .C(n7766) );
  CKBD0 U7683 ( .CLK(n7757), .C(n7767) );
  CKBD0 U7684 ( .CLK(n7758), .C(n7768) );
  CKBD0 U7685 ( .CLK(n7759), .C(n7769) );
  CKBD0 U7686 ( .CLK(n7760), .C(n7770) );
  CKBD0 U7687 ( .CLK(n7761), .C(n7771) );
  CKBD0 U7688 ( .CLK(n7762), .C(n7772) );
  CKBD0 U7689 ( .CLK(n7763), .C(n7773) );
  CKBD0 U7690 ( .CLK(n7705), .C(n7774) );
  CKBD0 U7691 ( .CLK(n7764), .C(n7775) );
  CKBD0 U7692 ( .CLK(n7706), .C(n7776) );
  CKBD0 U7693 ( .CLK(n7767), .C(n7777) );
  CKBD0 U7694 ( .CLK(n7768), .C(n7778) );
  CKBD0 U7695 ( .CLK(n7769), .C(n7779) );
  CKBD0 U7696 ( .CLK(n7770), .C(n7780) );
  CKBD0 U7697 ( .CLK(n7771), .C(n7781) );
  CKBD0 U7698 ( .CLK(n7772), .C(n7782) );
  CKBD0 U7699 ( .CLK(n7773), .C(n7783) );
  CKBD0 U7700 ( .CLK(n7775), .C(n7784) );
  CKBD0 U7701 ( .CLK(n7777), .C(n7785) );
  CKBD0 U7702 ( .CLK(n7719), .C(n7786) );
  CKBD0 U7703 ( .CLK(n7778), .C(n7787) );
  CKBD0 U7704 ( .CLK(n7721), .C(n7788) );
  CKBD0 U7705 ( .CLK(n7722), .C(n7789) );
  CKBD0 U7706 ( .CLK(n7723), .C(n7790) );
  CKBD0 U7707 ( .CLK(n7732), .C(n7791) );
  CKBD0 U7708 ( .CLK(n7733), .C(n7792) );
  CKBD0 U7709 ( .CLK(n7779), .C(n7793) );
  CKBD0 U7710 ( .CLK(n7780), .C(n7794) );
  CKBD0 U7711 ( .CLK(n7734), .C(n7795) );
  CKBD0 U7712 ( .CLK(n7781), .C(n7796) );
  CKBD0 U7713 ( .CLK(n7782), .C(n7797) );
  CKBD0 U7714 ( .CLK(n7783), .C(n7798) );
  CKBD0 U7715 ( .CLK(n7784), .C(n7799) );
  CKBD0 U7716 ( .CLK(n7785), .C(n7800) );
  CKBD0 U7717 ( .CLK(n7787), .C(n7801) );
  CKBD0 U7718 ( .CLK(n7735), .C(n7802) );
  CKBD0 U7719 ( .CLK(n7736), .C(n7803) );
  CKBD0 U7720 ( .CLK(n7737), .C(n7804) );
  CKBD0 U7721 ( .CLK(n7738), .C(n7805) );
  CKBD0 U7722 ( .CLK(n7739), .C(n7806) );
  CKBD0 U7723 ( .CLK(n7793), .C(n7807) );
  CKBD0 U7724 ( .CLK(n7794), .C(n7808) );
  CKBD0 U7725 ( .CLK(n7741), .C(n7809) );
  CKBD0 U7726 ( .CLK(n7796), .C(n7810) );
  CKBD0 U7727 ( .CLK(n7797), .C(n7811) );
  CKBD0 U7728 ( .CLK(n7798), .C(n7812) );
  CKBD0 U7729 ( .CLK(n7799), .C(n7813) );
  CKBD0 U7730 ( .CLK(n7800), .C(n7814) );
  CKBD0 U7731 ( .CLK(n7801), .C(n7815) );
  CKBD0 U7732 ( .CLK(n7742), .C(n7816) );
  CKBD0 U7733 ( .CLK(n7743), .C(n7817) );
  CKBD0 U7734 ( .CLK(n7744), .C(n7818) );
  CKBD0 U7735 ( .CLK(n7745), .C(n7819) );
  CKBD0 U7736 ( .CLK(n7807), .C(n7820) );
  CKBD0 U7737 ( .CLK(n7808), .C(n7821) );
  CKBD0 U7738 ( .CLK(n7810), .C(n7822) );
  CKBD0 U7739 ( .CLK(n7811), .C(n7823) );
  CKBD0 U7740 ( .CLK(n7812), .C(n7824) );
  CKBD0 U7741 ( .CLK(n7813), .C(n7825) );
  CKBD0 U7742 ( .CLK(n7814), .C(n7826) );
  CKBD0 U7743 ( .CLK(n7815), .C(n7827) );
  CKBD0 U7744 ( .CLK(n7754), .C(n7828) );
  CKBD0 U7745 ( .CLK(n7820), .C(n7829) );
  CKBD0 U7746 ( .CLK(n7821), .C(n7830) );
  CKBD0 U7747 ( .CLK(n7822), .C(n7831) );
  CKBD0 U7748 ( .CLK(n7823), .C(n7832) );
  CKBD0 U7749 ( .CLK(n7824), .C(n7833) );
  BUFFD0 U7750 ( .I(n7825), .Z(n7834) );
  CKBD0 U7751 ( .CLK(n7826), .C(n7835) );
  BUFFD0 U7752 ( .I(n7827), .Z(n7836) );
  CKBD0 U7753 ( .CLK(n7755), .C(n7837) );
  CKBD0 U7754 ( .CLK(n7756), .C(n7838) );
  BUFFD0 U7755 ( .I(n7829), .Z(n7839) );
  BUFFD0 U7756 ( .I(n7830), .Z(n7840) );
  CKBD0 U7757 ( .CLK(n7831), .C(n7841) );
  BUFFD0 U7758 ( .I(n7832), .Z(n7842) );
  CKBD0 U7759 ( .CLK(n7833), .C(n7843) );
  CKBD0 U7760 ( .CLK(n7834), .C(n7844) );
  CKBD0 U7761 ( .CLK(n7835), .C(n7845) );
  CKBD0 U7762 ( .CLK(n7836), .C(n7846) );
  CKBD0 U7763 ( .CLK(n7765), .C(n7847) );
  CKBD0 U7764 ( .CLK(n7766), .C(n7848) );
  CKBD0 U7765 ( .CLK(n7774), .C(n7849) );
  CKBD0 U7766 ( .CLK(n7839), .C(n7850) );
  CKBD0 U7767 ( .CLK(n7840), .C(n7851) );
  CKBD0 U7768 ( .CLK(n7776), .C(n7852) );
  CKBD0 U7769 ( .CLK(n7841), .C(n7853) );
  CKBD0 U7770 ( .CLK(n7842), .C(n7854) );
  CKBD0 U7771 ( .CLK(n7843), .C(n7855) );
  CKBD0 U7772 ( .CLK(n7844), .C(n7856) );
  CKBD0 U7773 ( .CLK(n7786), .C(n7857) );
  CKBD0 U7774 ( .CLK(n7788), .C(n7858) );
  CKBD0 U7775 ( .CLK(n7789), .C(n7859) );
  CKBD0 U7776 ( .CLK(n7845), .C(n7860) );
  CKBD0 U7777 ( .CLK(n7846), .C(n7861) );
  CKBD0 U7778 ( .CLK(n7850), .C(n7862) );
  CKBD0 U7779 ( .CLK(n7851), .C(n7863) );
  BUFFD0 U7780 ( .I(n7853), .Z(n7864) );
  CKBD0 U7781 ( .CLK(n7854), .C(n7865) );
  BUFFD0 U7782 ( .I(n7855), .Z(n7866) );
  CKBD0 U7783 ( .CLK(n7856), .C(n7867) );
  CKBD0 U7784 ( .CLK(n7790), .C(n7868) );
  CKBD0 U7785 ( .CLK(n7791), .C(n7869) );
  CKBD0 U7786 ( .CLK(n7792), .C(n7870) );
  CKBD0 U7787 ( .CLK(n7795), .C(n7871) );
  CKBD0 U7788 ( .CLK(n7802), .C(n7872) );
  BUFFD0 U7789 ( .I(n7860), .Z(n7873) );
  CKBD0 U7790 ( .CLK(n7803), .C(n7874) );
  CKBD0 U7791 ( .CLK(n7804), .C(n7875) );
  CKBD0 U7792 ( .CLK(n7861), .C(n7876) );
  CKBD0 U7793 ( .CLK(n7862), .C(n7877) );
  CKBD0 U7794 ( .CLK(n7863), .C(n7878) );
  CKBD0 U7795 ( .CLK(n7864), .C(n7879) );
  CKBD0 U7796 ( .CLK(n7865), .C(n7880) );
  CKBD0 U7797 ( .CLK(n7866), .C(n7881) );
  CKBD0 U7798 ( .CLK(n7867), .C(n7882) );
  CKBD0 U7799 ( .CLK(n7805), .C(n7883) );
  CKBD0 U7800 ( .CLK(n7806), .C(n7884) );
  CKBD0 U7801 ( .CLK(n7809), .C(n7885) );
  CKBD0 U7802 ( .CLK(n7816), .C(n7886) );
  CKBD0 U7803 ( .CLK(n7817), .C(n7887) );
  CKBD0 U7804 ( .CLK(n7873), .C(n7888) );
  CKBD0 U7805 ( .CLK(n7818), .C(n7889) );
  CKBD0 U7806 ( .CLK(n7876), .C(n7890) );
  CKBD0 U7807 ( .CLK(n7877), .C(n7891) );
  CKBD0 U7808 ( .CLK(n7878), .C(n7892) );
  CKBD0 U7809 ( .CLK(n7879), .C(n7893) );
  CKBD0 U7810 ( .CLK(n7880), .C(n7894) );
  CKBD0 U7811 ( .CLK(n7881), .C(n7895) );
  CKBD0 U7812 ( .CLK(n7882), .C(n7896) );
  CKBD0 U7813 ( .CLK(n7819), .C(n7897) );
  CKBD0 U7814 ( .CLK(n7828), .C(n7898) );
  CKBD0 U7815 ( .CLK(n7837), .C(n7899) );
  CKBD0 U7816 ( .CLK(n7888), .C(n7900) );
  CKBD0 U7817 ( .CLK(n7890), .C(n7901) );
  CKBD0 U7818 ( .CLK(n7891), .C(n7902) );
  CKBD0 U7819 ( .CLK(n7892), .C(n7903) );
  CKBD0 U7820 ( .CLK(n7893), .C(n7904) );
  CKBD0 U7821 ( .CLK(n7894), .C(n7905) );
  CKBD0 U7822 ( .CLK(n7895), .C(n7906) );
  CKBD0 U7823 ( .CLK(n7896), .C(n7907) );
  CKBD0 U7824 ( .CLK(n7838), .C(n7908) );
  CKBD0 U7825 ( .CLK(n7847), .C(n7909) );
  CKBD0 U7826 ( .CLK(n7848), .C(n7910) );
  CKBD0 U7827 ( .CLK(n7900), .C(n7911) );
  CKBD0 U7828 ( .CLK(n7901), .C(n7912) );
  CKBD0 U7829 ( .CLK(n7902), .C(n7913) );
  CKBD0 U7830 ( .CLK(n7903), .C(n7914) );
  CKBD0 U7831 ( .CLK(n7904), .C(n7915) );
  CKBD0 U7832 ( .CLK(n7905), .C(n7916) );
  CKBD0 U7833 ( .CLK(n7906), .C(n7917) );
  CKBD0 U7834 ( .CLK(n7907), .C(n7918) );
  CKBD0 U7835 ( .CLK(n7849), .C(n7919) );
  CKBD0 U7836 ( .CLK(n7852), .C(n7920) );
  CKBD0 U7837 ( .CLK(n7911), .C(n7921) );
  CKBD0 U7838 ( .CLK(n7912), .C(n7922) );
  CKBD0 U7839 ( .CLK(n7913), .C(n7923) );
  CKBD0 U7840 ( .CLK(n7914), .C(n7924) );
  CKBD0 U7841 ( .CLK(n7915), .C(n7925) );
  CKBD0 U7842 ( .CLK(n7916), .C(n7926) );
  CKBD0 U7843 ( .CLK(n7917), .C(n7927) );
  CKBD0 U7844 ( .CLK(n7918), .C(n7928) );
  CKBD0 U7845 ( .CLK(n7921), .C(n7929) );
  CKBD0 U7846 ( .CLK(n7857), .C(n7930) );
  CKBD0 U7847 ( .CLK(n7922), .C(n7931) );
  CKBD0 U7848 ( .CLK(n7858), .C(n7932) );
  CKBD0 U7849 ( .CLK(n7859), .C(n7933) );
  CKBD0 U7850 ( .CLK(n7923), .C(n7934) );
  CKBD0 U7851 ( .CLK(n7868), .C(n7935) );
  CKBD0 U7852 ( .CLK(n7924), .C(n7936) );
  CKBD0 U7853 ( .CLK(n7925), .C(n7937) );
  CKBD0 U7854 ( .CLK(n7926), .C(n7938) );
  CKBD0 U7855 ( .CLK(n7927), .C(n7939) );
  CKBD0 U7856 ( .CLK(n7928), .C(n7940) );
  CKBD0 U7857 ( .CLK(n7929), .C(n7941) );
  CKBD0 U7858 ( .CLK(n7931), .C(n7942) );
  CKBD0 U7859 ( .CLK(n7869), .C(n7943) );
  CKBD0 U7860 ( .CLK(n7870), .C(n7944) );
  CKBD0 U7861 ( .CLK(n7871), .C(n7945) );
  CKBD0 U7862 ( .CLK(n7872), .C(n7946) );
  CKBD0 U7863 ( .CLK(n7874), .C(n7947) );
  CKBD0 U7864 ( .CLK(n7875), .C(n7948) );
  CKBD0 U7865 ( .CLK(n7934), .C(n7949) );
  CKBD0 U7866 ( .CLK(n7936), .C(n7950) );
  CKBD0 U7867 ( .CLK(n7937), .C(n7951) );
  CKBD0 U7868 ( .CLK(n7938), .C(n7952) );
  CKBD0 U7869 ( .CLK(n7939), .C(n7953) );
  CKBD0 U7870 ( .CLK(n7940), .C(n7954) );
  CKBD0 U7871 ( .CLK(n7941), .C(n7955) );
  CKBD0 U7872 ( .CLK(n7942), .C(n7956) );
  CKBD0 U7873 ( .CLK(n7883), .C(n7957) );
  CKBD0 U7874 ( .CLK(n7949), .C(n7958) );
  CKBD0 U7875 ( .CLK(n7950), .C(n7959) );
  CKBD0 U7876 ( .CLK(n7951), .C(n7960) );
  CKBD0 U7877 ( .CLK(n7952), .C(n7961) );
  CKBD0 U7878 ( .CLK(n7953), .C(n7962) );
  BUFFD0 U7879 ( .I(n7954), .Z(n7963) );
  CKBD0 U7880 ( .CLK(n7955), .C(n7964) );
  BUFFD0 U7881 ( .I(n7956), .Z(n7965) );
  CKBD0 U7882 ( .CLK(n7884), .C(n7966) );
  CKBD0 U7883 ( .CLK(n7885), .C(n7967) );
  CKBD0 U7884 ( .CLK(n7886), .C(n7968) );
  CKBD0 U7885 ( .CLK(n7887), .C(n7969) );
  CKBD0 U7886 ( .CLK(n7889), .C(n7970) );
  BUFFD0 U7887 ( .I(n7958), .Z(n7971) );
  BUFFD0 U7888 ( .I(n7959), .Z(n7972) );
  CKBD0 U7889 ( .CLK(n7897), .C(n7973) );
  CKBD0 U7890 ( .CLK(n7960), .C(n7974) );
  BUFFD0 U7891 ( .I(n7961), .Z(n7975) );
  CKBD0 U7892 ( .CLK(n7962), .C(n7976) );
  CKBD0 U7893 ( .CLK(n7963), .C(n7977) );
  CKBD0 U7894 ( .CLK(n7964), .C(n7978) );
  CKBD0 U7895 ( .CLK(n7965), .C(n7979) );
  CKBD0 U7896 ( .CLK(n7898), .C(n7980) );
  CKBD0 U7897 ( .CLK(n7899), .C(n7981) );
  CKBD0 U7898 ( .CLK(n7908), .C(n7982) );
  CKBD0 U7899 ( .CLK(n7971), .C(n7983) );
  CKBD0 U7900 ( .CLK(n7972), .C(n7984) );
  CKBD0 U7901 ( .CLK(n7974), .C(n7985) );
  CKBD0 U7902 ( .CLK(n7975), .C(n7986) );
  CKBD0 U7903 ( .CLK(n7976), .C(n7987) );
  CKBD0 U7904 ( .CLK(n7977), .C(n7988) );
  BUFFD0 U7905 ( .I(n7978), .Z(n7989) );
  CKBD0 U7906 ( .CLK(n7979), .C(n7990) );
  CKBD0 U7907 ( .CLK(n7909), .C(n7991) );
  CKBD0 U7908 ( .CLK(n7910), .C(n7992) );
  CKBD0 U7909 ( .CLK(n7983), .C(n7993) );
  CKBD0 U7910 ( .CLK(n7984), .C(n7994) );
  BUFFD0 U7911 ( .I(n7985), .Z(n7995) );
  CKBD0 U7912 ( .CLK(n7986), .C(n7996) );
  BUFFD0 U7913 ( .I(n7987), .Z(n7997) );
  CKBD0 U7914 ( .CLK(n7988), .C(n7998) );
  CKBD0 U7915 ( .CLK(n7989), .C(n7999) );
  CKBD0 U7916 ( .CLK(n7990), .C(n8000) );
  CKBD0 U7917 ( .CLK(n7919), .C(n8001) );
  CKBD0 U7918 ( .CLK(n7920), .C(n8002) );
  CKBD0 U7919 ( .CLK(n7993), .C(n8003) );
  CKBD0 U7920 ( .CLK(n7994), .C(n8004) );
  CKBD0 U7921 ( .CLK(n7995), .C(n8005) );
  CKBD0 U7922 ( .CLK(n7996), .C(n8006) );
  CKBD0 U7923 ( .CLK(n7997), .C(n8007) );
  CKBD0 U7924 ( .CLK(n7930), .C(n8008) );
  CKBD0 U7925 ( .CLK(n7998), .C(n8009) );
  CKBD0 U7926 ( .CLK(n7932), .C(n8010) );
  CKBD0 U7927 ( .CLK(n7933), .C(n8011) );
  CKBD0 U7928 ( .CLK(n7935), .C(n8012) );
  CKBD0 U7929 ( .CLK(n7943), .C(n8013) );
  CKBD0 U7930 ( .CLK(n7944), .C(n8014) );
  CKBD0 U7931 ( .CLK(n7945), .C(n8015) );
  CKBD0 U7932 ( .CLK(n7999), .C(n8016) );
  CKBD0 U7933 ( .CLK(n7946), .C(n8017) );
  CKBD0 U7934 ( .CLK(n8000), .C(n8018) );
  CKBD0 U7935 ( .CLK(n8003), .C(n8019) );
  CKBD0 U7936 ( .CLK(n8004), .C(n8020) );
  CKBD0 U7937 ( .CLK(n8005), .C(n8021) );
  CKBD0 U7938 ( .CLK(n8006), .C(n8022) );
  CKBD0 U7939 ( .CLK(n8007), .C(n8023) );
  CKBD0 U7940 ( .CLK(n8009), .C(n8024) );
  CKBD0 U7941 ( .CLK(n7947), .C(n8025) );
  CKBD0 U7942 ( .CLK(n7948), .C(n8026) );
  CKBD0 U7943 ( .CLK(n7966), .C(n8027) );
  CKBD0 U7944 ( .CLK(n7957), .C(n8028) );
  CKBD0 U7945 ( .CLK(n7967), .C(n8029) );
  CKBD0 U7946 ( .CLK(n8016), .C(n8030) );
  CKBD0 U7947 ( .CLK(n8018), .C(n8031) );
  CKBD0 U7948 ( .CLK(n8019), .C(n8032) );
  CKBD0 U7949 ( .CLK(n8020), .C(n8033) );
  CKBD0 U7950 ( .CLK(n8021), .C(n8034) );
  CKBD0 U7951 ( .CLK(n8022), .C(n8035) );
  CKBD0 U7952 ( .CLK(n8023), .C(n8036) );
  CKBD0 U7953 ( .CLK(n8024), .C(n8037) );
  CKBD0 U7954 ( .CLK(n7969), .C(n8038) );
  CKBD0 U7955 ( .CLK(n7968), .C(n8039) );
  CKBD0 U7956 ( .CLK(n7970), .C(n8040) );
  CKBD0 U7957 ( .CLK(n7973), .C(n8041) );
  CKBD0 U7958 ( .CLK(n7980), .C(n8042) );
  CKBD0 U7959 ( .CLK(n8030), .C(n8043) );
  CKBD0 U7960 ( .CLK(n8031), .C(n8044) );
  CKBD0 U7961 ( .CLK(n8032), .C(n8045) );
  CKBD0 U7962 ( .CLK(n8033), .C(n8046) );
  CKBD0 U7963 ( .CLK(n8034), .C(n8047) );
  CKBD0 U7964 ( .CLK(n8035), .C(n8048) );
  CKBD0 U7965 ( .CLK(n8036), .C(n8049) );
  CKBD0 U7966 ( .CLK(n8037), .C(n8050) );
  CKBD0 U7967 ( .CLK(n7981), .C(n8051) );
  CKBD0 U7968 ( .CLK(n7982), .C(n8052) );
  CKBD0 U7969 ( .CLK(n8043), .C(n8053) );
  CKBD0 U7970 ( .CLK(n8044), .C(n8054) );
  CKBD0 U7971 ( .CLK(n8045), .C(n8055) );
  CKBD0 U7972 ( .CLK(n8046), .C(n8056) );
  CKBD0 U7973 ( .CLK(n8047), .C(n8057) );
  CKBD0 U7974 ( .CLK(n8048), .C(n8058) );
  CKBD0 U7975 ( .CLK(n8049), .C(n8059) );
  CKBD0 U7976 ( .CLK(n8050), .C(n8060) );
  CKBD0 U7977 ( .CLK(n7991), .C(n8061) );
  CKBD0 U7978 ( .CLK(n7992), .C(n8062) );
  CKBD0 U7979 ( .CLK(n8001), .C(n8063) );
  CKBD0 U7980 ( .CLK(n8053), .C(n8064) );
  CKBD0 U7981 ( .CLK(n8054), .C(n8065) );
  CKBD0 U7982 ( .CLK(n8055), .C(n8066) );
  CKBD0 U7983 ( .CLK(n8056), .C(n8067) );
  CKBD0 U7984 ( .CLK(n8057), .C(n8068) );
  CKBD0 U7985 ( .CLK(n8058), .C(n8069) );
  CKBD0 U7986 ( .CLK(n8059), .C(n8070) );
  CKBD0 U7987 ( .CLK(n8060), .C(n8071) );
  CKBD0 U7988 ( .CLK(n8002), .C(n8072) );
  CKBD0 U7989 ( .CLK(n8064), .C(n8073) );
  CKBD0 U7990 ( .CLK(n8008), .C(n8074) );
  CKBD0 U7991 ( .CLK(n8065), .C(n8075) );
  CKBD0 U7992 ( .CLK(n8010), .C(n8076) );
  CKBD0 U7993 ( .CLK(n8011), .C(n8077) );
  CKBD0 U7994 ( .CLK(n8066), .C(n8078) );
  CKBD0 U7995 ( .CLK(n8067), .C(n8079) );
  CKBD0 U7996 ( .CLK(n8068), .C(n8080) );
  CKBD0 U7997 ( .CLK(n8069), .C(n8081) );
  CKBD0 U7998 ( .CLK(n8070), .C(n8082) );
  CKBD0 U7999 ( .CLK(n8071), .C(n8083) );
  CKBD0 U8000 ( .CLK(n8073), .C(n8084) );
  CKBD0 U8001 ( .CLK(n8075), .C(n8085) );
  BUFFD0 U8002 ( .I(n8012), .Z(n8086) );
  CKBD0 U8003 ( .CLK(n8013), .C(n8087) );
  CKBD0 U8004 ( .CLK(n8014), .C(n8088) );
  CKBD0 U8005 ( .CLK(n8015), .C(n8089) );
  CKBD0 U8006 ( .CLK(n8078), .C(n8090) );
  CKBD0 U8007 ( .CLK(n8079), .C(n8091) );
  BUFFD0 U8008 ( .I(n8017), .Z(n8092) );
  CKBD0 U8009 ( .CLK(n8026), .C(n8093) );
  BUFFD0 U8010 ( .I(n8025), .Z(n8094) );
  CKBD0 U8011 ( .CLK(n8028), .C(n8095) );
  BUFFD0 U8012 ( .I(n8027), .Z(n8096) );
  BUFFD0 U8013 ( .I(n8029), .Z(n8097) );
  CKBD0 U8014 ( .CLK(n8039), .C(n8098) );
  CKBD0 U8015 ( .CLK(n8080), .C(n8099) );
  BUFFD0 U8016 ( .I(n8038), .Z(n8100) );
  CKBD0 U8017 ( .CLK(n8040), .C(n8101) );
  CKBD0 U8018 ( .CLK(n8081), .C(n8102) );
  CKBD0 U8019 ( .CLK(n8082), .C(n8103) );
  BUFFD0 U8020 ( .I(n8083), .Z(n8104) );
  CKBD0 U8021 ( .CLK(n8084), .C(n8105) );
  BUFFD0 U8022 ( .I(n8085), .Z(n8106) );
  BUFFD0 U8023 ( .I(n8090), .Z(n8107) );
  BUFFD0 U8024 ( .I(n8091), .Z(n8108) );
  CKBD0 U8025 ( .CLK(n8099), .C(n8109) );
  BUFFD0 U8026 ( .I(n8102), .Z(n8110) );
  CKBD0 U8027 ( .CLK(n8103), .C(n8111) );
  CKBD0 U8028 ( .CLK(n8104), .C(n8112) );
  CKBD0 U8029 ( .CLK(n8105), .C(n8113) );
  CKBD0 U8030 ( .CLK(n8106), .C(n8114) );
  CKBD0 U8031 ( .CLK(n8107), .C(n8115) );
  CKBD0 U8032 ( .CLK(n8108), .C(n8116) );
  CKBD0 U8033 ( .CLK(n8109), .C(n8117) );
  CKBD0 U8034 ( .CLK(n8110), .C(n8118) );
  CKBD0 U8035 ( .CLK(n8111), .C(n8119) );
  CKBD0 U8036 ( .CLK(n8112), .C(n8120) );
  BUFFD0 U8037 ( .I(n8113), .Z(n8121) );
  CKBD0 U8038 ( .CLK(n8114), .C(n8122) );
  BUFFD0 U8039 ( .I(n8041), .Z(n8123) );
  BUFFD0 U8040 ( .I(n8042), .Z(n8124) );
  CKBD0 U8041 ( .CLK(n8051), .C(n8125) );
  CKBD0 U8042 ( .CLK(n8115), .C(n8126) );
  CKBD0 U8043 ( .CLK(n8116), .C(n8127) );
  BUFFD0 U8044 ( .I(n8052), .Z(n8128) );
  BUFFD0 U8045 ( .I(n8117), .Z(n8129) );
  BUFFD0 U8046 ( .I(n8063), .Z(n8130) );
  CKBD0 U8047 ( .CLK(n8061), .C(n8131) );
  CKBD0 U8048 ( .CLK(n8118), .C(n8132) );
  BUFFD0 U8049 ( .I(n8119), .Z(n8133) );
  CKBD0 U8050 ( .CLK(n8120), .C(n8134) );
  CKBD0 U8051 ( .CLK(n8121), .C(n8135) );
  CKBD0 U8052 ( .CLK(n8122), .C(n8136) );
  CKBD0 U8053 ( .CLK(n8126), .C(n8137) );
  CKBD0 U8054 ( .CLK(n8127), .C(n8138) );
  CKBD0 U8055 ( .CLK(n8129), .C(n8139) );
  CKBD0 U8056 ( .CLK(n8132), .C(n8140) );
  CKBD0 U8057 ( .CLK(n8133), .C(n8141) );
  CKBD0 U8058 ( .CLK(n8134), .C(n8142) );
  CKBD0 U8059 ( .CLK(n8135), .C(n8143) );
  CKBD0 U8060 ( .CLK(n8136), .C(n8144) );
  CKBD0 U8061 ( .CLK(n8062), .C(n8145) );
  CKBD0 U8062 ( .CLK(n8072), .C(n8146) );
  CKBD0 U8063 ( .CLK(n8137), .C(n8147) );
  CKBD0 U8064 ( .CLK(n8138), .C(n8148) );
  CKBD0 U8065 ( .CLK(n8139), .C(n8149) );
  CKBD0 U8066 ( .CLK(n8140), .C(n8150) );
  CKBD0 U8067 ( .CLK(n8141), .C(n8151) );
  BUFFD0 U8068 ( .I(n8074), .Z(n8152) );
  CKBD0 U8069 ( .CLK(n8142), .C(n8153) );
  BUFFD0 U8070 ( .I(n8076), .Z(n8154) );
  BUFFD0 U8071 ( .I(n8077), .Z(n8155) );
  CKBD0 U8072 ( .CLK(n8086), .C(n8156) );
  BUFFD0 U8073 ( .I(n8087), .Z(n8157) );
  CKBD0 U8074 ( .CLK(n8143), .C(n8158) );
  BUFFD0 U8075 ( .I(n8088), .Z(n8159) );
  CKBD0 U8076 ( .CLK(n8144), .C(n8160) );
  CKBD0 U8077 ( .CLK(n8147), .C(n8161) );
  CKBD0 U8078 ( .CLK(n8148), .C(n8162) );
  CKBD0 U8079 ( .CLK(n8149), .C(n8163) );
  CKBD0 U8080 ( .CLK(n8150), .C(n8164) );
  CKBD0 U8081 ( .CLK(n8151), .C(n8165) );
  CKBD0 U8082 ( .CLK(n8153), .C(n8166) );
  BUFFD0 U8083 ( .I(n8089), .Z(n8167) );
  CKBD0 U8084 ( .CLK(n8092), .C(n8168) );
  CKBD0 U8085 ( .CLK(n8094), .C(n8169) );
  BUFFD0 U8086 ( .I(n8093), .Z(n8170) );
  CKBD0 U8087 ( .CLK(n8096), .C(n8171) );
  BUFFD0 U8088 ( .I(n8095), .Z(n8172) );
  CKBD0 U8089 ( .CLK(n8158), .C(n8173) );
  CKBD0 U8090 ( .CLK(n8097), .C(n8174) );
  CKBD0 U8091 ( .CLK(n8160), .C(n8175) );
  CKBD0 U8092 ( .CLK(n8161), .C(n8176) );
  CKBD0 U8093 ( .CLK(n8162), .C(n8177) );
  CKBD0 U8094 ( .CLK(n8163), .C(n8178) );
  CKBD0 U8095 ( .CLK(n8164), .C(n8179) );
  CKBD0 U8096 ( .CLK(n8165), .C(n8180) );
  CKBD0 U8097 ( .CLK(n8166), .C(n8181) );
  CKBD0 U8098 ( .CLK(n8100), .C(n8182) );
  BUFFD0 U8099 ( .I(n8098), .Z(n8183) );
  BUFFD0 U8100 ( .I(n8101), .Z(n8184) );
  CKBD0 U8101 ( .CLK(n8123), .C(n8185) );
  CKBD0 U8102 ( .CLK(n8124), .C(n8186) );
  CKBD0 U8103 ( .CLK(n8173), .C(n8187) );
  CKBD0 U8104 ( .CLK(n8175), .C(n8188) );
  CKBD0 U8105 ( .CLK(n8176), .C(n8189) );
  CKBD0 U8106 ( .CLK(n8177), .C(n8190) );
  CKBD0 U8107 ( .CLK(n8178), .C(n8191) );
  CKBD0 U8108 ( .CLK(n8179), .C(n8192) );
  CKBD0 U8109 ( .CLK(n8180), .C(n8193) );
  CKBD0 U8110 ( .CLK(n8181), .C(n8194) );
  BUFFD0 U8111 ( .I(n8125), .Z(n8195) );
  CKBD0 U8112 ( .CLK(n8128), .C(n8196) );
  BUFFD0 U8113 ( .I(n8131), .Z(n8197) );
  BUFFD0 U8114 ( .I(n8145), .Z(n8198) );
  CKBD0 U8115 ( .CLK(n8187), .C(n8199) );
  CKBD0 U8116 ( .CLK(n8188), .C(n8200) );
  CKBD0 U8117 ( .CLK(n8189), .C(n8201) );
  CKBD0 U8118 ( .CLK(n8190), .C(n8202) );
  CKBD0 U8119 ( .CLK(n8191), .C(n8203) );
  CKBD0 U8120 ( .CLK(n8192), .C(n8204) );
  CKBD0 U8121 ( .CLK(n8193), .C(n8205) );
  CKBD0 U8122 ( .CLK(n8194), .C(n8206) );
  CKBD0 U8123 ( .CLK(n8130), .C(n8207) );
  BUFFD0 U8124 ( .I(n8146), .Z(n8208) );
  CKBD0 U8125 ( .CLK(n8199), .C(n8209) );
  CKBD0 U8126 ( .CLK(n8200), .C(n8210) );
  CKBD0 U8127 ( .CLK(n8201), .C(n8211) );
  CKBD0 U8128 ( .CLK(n8202), .C(n8212) );
  CKBD0 U8129 ( .CLK(n8203), .C(n8213) );
  CKBD0 U8130 ( .CLK(n8204), .C(n8214) );
  CKBD0 U8131 ( .CLK(n8205), .C(n8215) );
  CKBD0 U8132 ( .CLK(n8206), .C(n8216) );
  CKBD0 U8133 ( .CLK(n8209), .C(n8217) );
  CKBD0 U8134 ( .CLK(n8210), .C(n8218) );
  CKBD0 U8135 ( .CLK(n8152), .C(n8219) );
  CKBD0 U8136 ( .CLK(n8211), .C(n8220) );
  CKBD0 U8137 ( .CLK(n8212), .C(n8221) );
  CKBD0 U8138 ( .CLK(n8154), .C(n8222) );
  CKBD0 U8139 ( .CLK(n8155), .C(n8223) );
  BUFFD0 U8140 ( .I(n8156), .Z(n8224) );
  CKBD0 U8141 ( .CLK(n8157), .C(n8225) );
  CKBD0 U8142 ( .CLK(n8159), .C(n8226) );
  CKBD0 U8143 ( .CLK(n8167), .C(n8227) );
  CKBD0 U8144 ( .CLK(n8213), .C(n8228) );
  BUFFD0 U8145 ( .I(n8168), .Z(n8229) );
  CKBD0 U8146 ( .CLK(n8170), .C(n8230) );
  BUFFD0 U8147 ( .I(n8169), .Z(n8231) );
  CKBD0 U8148 ( .CLK(n8172), .C(n8232) );
  BUFFD0 U8149 ( .I(n8171), .Z(n8233) );
  BUFFD0 U8150 ( .I(n8174), .Z(n8234) );
  CKBD0 U8151 ( .CLK(n8214), .C(n8235) );
  CKBD0 U8152 ( .CLK(n8183), .C(n8236) );
  BUFFD0 U8153 ( .I(n8182), .Z(n8237) );
  CKBD0 U8154 ( .CLK(n8184), .C(n8238) );
  BUFFD0 U8155 ( .I(n8185), .Z(n8239) );
  BUFFD0 U8156 ( .I(n8186), .Z(n8240) );
  CKBD0 U8157 ( .CLK(n8215), .C(n8241) );
  CKBD0 U8158 ( .CLK(n8195), .C(n8242) );
  BUFFD0 U8159 ( .I(n8196), .Z(n8243) );
  CKBD0 U8160 ( .CLK(n8197), .C(n8244) );
  CKBD0 U8161 ( .CLK(n8198), .C(n8245) );
  BUFFD0 U8162 ( .I(n8216), .Z(n8246) );
  CKBD0 U8163 ( .CLK(n8217), .C(n8247) );
  BUFFD0 U8164 ( .I(n8218), .Z(n8248) );
  BUFFD0 U8165 ( .I(n8220), .Z(n8249) );
  BUFFD0 U8166 ( .I(n8221), .Z(n8250) );
  CKBD0 U8167 ( .CLK(n8228), .C(n8251) );
  BUFFD0 U8168 ( .I(n8235), .Z(n8252) );
  CKBD0 U8169 ( .CLK(n8241), .C(n8253) );
  CKBD0 U8170 ( .CLK(n8207), .C(n8254) );
  CKBD0 U8171 ( .CLK(n8208), .C(n8255) );
  CKBD0 U8172 ( .CLK(n8246), .C(n8256) );
  CKBD0 U8173 ( .CLK(n8247), .C(n8257) );
  CKBD0 U8174 ( .CLK(n8248), .C(n8258) );
  BUFFD0 U8175 ( .I(n8219), .Z(n8259) );
  BUFFD0 U8176 ( .I(n8222), .Z(n8260) );
  BUFFD0 U8177 ( .I(n8223), .Z(n8261) );
  CKBD0 U8178 ( .CLK(n8249), .C(n8262) );
  CKBD0 U8179 ( .CLK(n8250), .C(n8263) );
  CKBD0 U8180 ( .CLK(n8251), .C(n8264) );
  CKBD0 U8181 ( .CLK(n8252), .C(n8265) );
  CKBD0 U8182 ( .CLK(n8253), .C(n8266) );
  CKBD0 U8183 ( .CLK(n8256), .C(n8267) );
  BUFFD0 U8184 ( .I(n8257), .Z(n8268) );
  CKBD0 U8185 ( .CLK(n8258), .C(n8269) );
  CKBD0 U8186 ( .CLK(n8224), .C(n8270) );
  BUFFD0 U8187 ( .I(n8225), .Z(n8271) );
  BUFFD0 U8188 ( .I(n8226), .Z(n8272) );
  BUFFD0 U8189 ( .I(n8227), .Z(n8273) );
  CKBD0 U8190 ( .CLK(n8229), .C(n8274) );
  CKBD0 U8191 ( .CLK(n8231), .C(n8275) );
  CKBD0 U8192 ( .CLK(n8262), .C(n8276) );
  CKBD0 U8193 ( .CLK(n8263), .C(n8277) );
  BUFFD0 U8194 ( .I(n8264), .Z(n8278) );
  CKBD0 U8195 ( .CLK(n8265), .C(n8279) );
  BUFFD0 U8196 ( .I(n8266), .Z(n8280) );
  CKBD0 U8197 ( .CLK(n8267), .C(n8281) );
  CKBD0 U8198 ( .CLK(n8268), .C(n8282) );
  CKBD0 U8199 ( .CLK(n8269), .C(n8283) );
  BUFFD0 U8200 ( .I(n8230), .Z(n8284) );
  CKBD0 U8201 ( .CLK(n8233), .C(n8285) );
  BUFFD0 U8202 ( .I(n8232), .Z(n8286) );
  CKBD0 U8203 ( .CLK(n8234), .C(n8287) );
  CKBD0 U8204 ( .CLK(n8237), .C(n8288) );
  BUFFD0 U8205 ( .I(n8236), .Z(n8289) );
  CKBD0 U8206 ( .CLK(n8276), .C(n8290) );
  CKBD0 U8207 ( .CLK(n8277), .C(n8291) );
  CKBD0 U8208 ( .CLK(n8278), .C(n8292) );
  CKBD0 U8209 ( .CLK(n8279), .C(n8293) );
  CKBD0 U8210 ( .CLK(n8280), .C(n8294) );
  CKBD0 U8211 ( .CLK(n8281), .C(n8295) );
  CKBD0 U8212 ( .CLK(n8282), .C(n8296) );
  CKBD0 U8213 ( .CLK(n8283), .C(n8297) );
  BUFFD0 U8214 ( .I(n8238), .Z(n8298) );
  CKBD0 U8215 ( .CLK(n8239), .C(n8299) );
  CKBD0 U8216 ( .CLK(n8240), .C(n8300) );
  BUFFD0 U8217 ( .I(n8244), .Z(n8301) );
  BUFFD0 U8218 ( .I(n8245), .Z(n8302) );
  BUFFD0 U8219 ( .I(n8242), .Z(n8303) );
  CKBD0 U8220 ( .CLK(n8290), .C(n8304) );
  CKBD0 U8221 ( .CLK(n8291), .C(n8305) );
  CKBD0 U8222 ( .CLK(n8243), .C(n8306) );
  CKBD0 U8223 ( .CLK(n8292), .C(n8307) );
  CKBD0 U8224 ( .CLK(n8293), .C(n8308) );
  CKBD0 U8225 ( .CLK(n8294), .C(n8309) );
  CKBD0 U8226 ( .CLK(n8295), .C(n8310) );
  CKBD0 U8227 ( .CLK(n8296), .C(n8311) );
  CKBD0 U8228 ( .CLK(n8297), .C(n8312) );
  BUFFD0 U8229 ( .I(n8254), .Z(n8313) );
  BUFFD0 U8230 ( .I(n8255), .Z(n8314) );
  CKBD0 U8231 ( .CLK(n8304), .C(n8315) );
  CKBD0 U8232 ( .CLK(n8305), .C(n8316) );
  CKBD0 U8233 ( .CLK(n8307), .C(n8317) );
  CKBD0 U8234 ( .CLK(n8308), .C(n8318) );
  CKBD0 U8235 ( .CLK(n8309), .C(n8319) );
  CKBD0 U8236 ( .CLK(n8310), .C(n8320) );
  CKBD0 U8237 ( .CLK(n8311), .C(n8321) );
  CKBD0 U8238 ( .CLK(n8312), .C(n8322) );
  CKBD0 U8239 ( .CLK(n8315), .C(n8323) );
  CKBD0 U8240 ( .CLK(n8316), .C(n8324) );
  CKBD0 U8241 ( .CLK(n8317), .C(n8325) );
  CKBD0 U8242 ( .CLK(n8318), .C(n8326) );
  CKBD0 U8243 ( .CLK(n8319), .C(n8327) );
  CKBD0 U8244 ( .CLK(n8259), .C(n8328) );
  CKBD0 U8245 ( .CLK(n8320), .C(n8329) );
  CKBD0 U8246 ( .CLK(n8260), .C(n8330) );
  CKBD0 U8247 ( .CLK(n8261), .C(n8331) );
  BUFFD0 U8248 ( .I(n8270), .Z(n8332) );
  CKBD0 U8249 ( .CLK(n8271), .C(n8333) );
  CKBD0 U8250 ( .CLK(n8272), .C(n8334) );
  CKBD0 U8251 ( .CLK(n8321), .C(n8335) );
  CKBD0 U8252 ( .CLK(n8273), .C(n8336) );
  CKBD0 U8253 ( .CLK(n8322), .C(n8337) );
  CKBD0 U8254 ( .CLK(n8323), .C(n8338) );
  CKBD0 U8255 ( .CLK(n8324), .C(n8339) );
  CKBD0 U8256 ( .CLK(n8325), .C(n8340) );
  CKBD0 U8257 ( .CLK(n8326), .C(n8341) );
  CKBD0 U8258 ( .CLK(n8327), .C(n8342) );
  CKBD0 U8259 ( .CLK(n8329), .C(n8343) );
  CKBD0 U8260 ( .CLK(n8335), .C(n8344) );
  CKBD0 U8261 ( .CLK(n8337), .C(n8345) );
  CKBD0 U8262 ( .CLK(n8338), .C(n8346) );
  CKBD0 U8263 ( .CLK(n8339), .C(n8347) );
  CKBD0 U8264 ( .CLK(n8340), .C(n8348) );
  CKBD0 U8265 ( .CLK(n8341), .C(n8349) );
  CKBD0 U8266 ( .CLK(n8342), .C(n8350) );
  CKBD0 U8267 ( .CLK(n8343), .C(n8351) );
  CKBD0 U8268 ( .CLK(n8344), .C(n8352) );
  BUFFD0 U8269 ( .I(n8346), .Z(n8353) );
  CKBD0 U8270 ( .CLK(n8345), .C(n8354) );
  CKBD0 U8271 ( .CLK(n8347), .C(n8355) );
  CKBD0 U8272 ( .CLK(n8348), .C(n8356) );
  CKBD0 U8273 ( .CLK(n8349), .C(n8357) );
  CKBD0 U8274 ( .CLK(n8350), .C(n8358) );
  BUFFD0 U8275 ( .I(n8274), .Z(n8359) );
  CKBD0 U8276 ( .CLK(n8284), .C(n8360) );
  BUFFD0 U8277 ( .I(n8275), .Z(n8361) );
  CKBD0 U8278 ( .CLK(n8286), .C(n8362) );
  BUFFD0 U8279 ( .I(n8285), .Z(n8363) );
  CKBD0 U8280 ( .CLK(n8351), .C(n8364) );
  CKBD0 U8281 ( .CLK(n8352), .C(n8365) );
  CKBD0 U8282 ( .CLK(n8354), .C(n8366) );
  CKBD0 U8283 ( .CLK(n8353), .C(n8367) );
  CKBD0 U8284 ( .CLK(n8355), .C(n8368) );
  CKBD0 U8285 ( .CLK(n8356), .C(n8369) );
  BUFFD0 U8286 ( .I(n8357), .Z(n8370) );
  CKBD0 U8287 ( .CLK(n8358), .C(n8371) );
  BUFFD0 U8288 ( .I(n8287), .Z(n8372) );
  CKBD0 U8289 ( .CLK(n8289), .C(n8373) );
  BUFFD0 U8290 ( .I(n8288), .Z(n8374) );
  CKBD0 U8291 ( .CLK(n8298), .C(n8375) );
  BUFFD0 U8292 ( .I(n8299), .Z(n8376) );
  CKBD0 U8293 ( .CLK(n8301), .C(n8377) );
  BUFFD0 U8294 ( .I(n8364), .Z(n8378) );
  CKBD0 U8295 ( .CLK(n8365), .C(n8379) );
  BUFFD0 U8296 ( .I(n8366), .Z(n8380) );
  CKBD0 U8297 ( .CLK(n8367), .C(n8381) );
  BUFFD0 U8298 ( .I(n8368), .Z(n8382) );
  CKBD0 U8299 ( .CLK(n8369), .C(n8383) );
  CKBD0 U8300 ( .CLK(n8370), .C(n8384) );
  CKBD0 U8301 ( .CLK(n8371), .C(n8385) );
  BUFFD0 U8302 ( .I(n8300), .Z(n8386) );
  CKBD0 U8303 ( .CLK(n8302), .C(n8387) );
  CKBD0 U8304 ( .CLK(n8303), .C(n8388) );
  BUFFD0 U8305 ( .I(n8306), .Z(n8389) );
  CKBD0 U8306 ( .CLK(n8313), .C(n8390) );
  CKBD0 U8307 ( .CLK(n8314), .C(n8391) );
  CKBD0 U8308 ( .CLK(n8378), .C(n8392) );
  CKBD0 U8309 ( .CLK(n8379), .C(n8393) );
  CKBD0 U8310 ( .CLK(n8380), .C(n8394) );
  CKBD0 U8311 ( .CLK(n8381), .C(n8395) );
  CKBD0 U8312 ( .CLK(n8382), .C(n8396) );
  CKBD0 U8313 ( .CLK(n8383), .C(n8397) );
  CKBD0 U8314 ( .CLK(n8384), .C(n8398) );
  CKBD0 U8315 ( .CLK(n8385), .C(n8399) );
  CKBD0 U8316 ( .CLK(n8392), .C(n8400) );
  BUFFD0 U8317 ( .I(n8393), .Z(n8401) );
  CKBD0 U8318 ( .CLK(n8394), .C(n8402) );
  BUFFD0 U8319 ( .I(n8328), .Z(n8403) );
  CKBD0 U8320 ( .CLK(n8395), .C(n8404) );
  CKBD0 U8321 ( .CLK(n8396), .C(n8405) );
  BUFFD0 U8322 ( .I(n8330), .Z(n8406) );
  BUFFD0 U8323 ( .I(n8397), .Z(n8407) );
  CKBD0 U8324 ( .CLK(n8398), .C(n8408) );
  BUFFD0 U8325 ( .I(n8399), .Z(n8409) );
  CKBD0 U8326 ( .CLK(n8400), .C(n8410) );
  CKBD0 U8327 ( .CLK(n8401), .C(n8411) );
  CKBD0 U8328 ( .CLK(n8402), .C(n8412) );
  BUFFD0 U8329 ( .I(n8331), .Z(n8413) );
  CKBD0 U8330 ( .CLK(n8332), .C(n8414) );
  BUFFD0 U8331 ( .I(n8333), .Z(n8415) );
  BUFFD0 U8332 ( .I(n8334), .Z(n8416) );
  BUFFD0 U8333 ( .I(n8336), .Z(n8417) );
  CKBD0 U8334 ( .CLK(n8404), .C(n8418) );
  CKBD0 U8335 ( .CLK(n8359), .C(n8419) );
  CKBD0 U8336 ( .CLK(n8405), .C(n8420) );
  CKBD0 U8337 ( .CLK(n8407), .C(n8421) );
  CKBD0 U8338 ( .CLK(n8408), .C(n8422) );
  CKBD0 U8339 ( .CLK(n8409), .C(n8423) );
  CKBD0 U8340 ( .CLK(n8410), .C(n8424) );
  CKBD0 U8341 ( .CLK(n8411), .C(n8425) );
  CKBD0 U8342 ( .CLK(n8412), .C(n8426) );
  CKBD0 U8343 ( .CLK(n8361), .C(n8427) );
  BUFFD0 U8344 ( .I(n8360), .Z(n8428) );
  CKBD0 U8345 ( .CLK(n8363), .C(n8429) );
  BUFFD0 U8346 ( .I(n8362), .Z(n8430) );
  CKBD0 U8347 ( .CLK(n8372), .C(n8431) );
  CKBD0 U8348 ( .CLK(n8418), .C(n8432) );
  CKBD0 U8349 ( .CLK(n8420), .C(n8433) );
  BUFFD0 U8350 ( .I(n8377), .Z(n8434) );
  CKBD0 U8351 ( .CLK(n8374), .C(n8435) );
  CKBD0 U8352 ( .CLK(n8421), .C(n8436) );
  CKBD0 U8353 ( .CLK(n8422), .C(n8437) );
  CKBD0 U8354 ( .CLK(n8423), .C(n8438) );
  CKBD0 U8355 ( .CLK(n8424), .C(n8439) );
  CKBD0 U8356 ( .CLK(n8425), .C(n8440) );
  CKBD0 U8357 ( .CLK(n8426), .C(n8441) );
  BUFFD0 U8358 ( .I(n8373), .Z(n8442) );
  BUFFD0 U8359 ( .I(n8387), .Z(n8443) );
  BUFFD0 U8360 ( .I(n8375), .Z(n8444) );
  CKBD0 U8361 ( .CLK(n8376), .C(n8445) );
  CKBD0 U8362 ( .CLK(n8386), .C(n8446) );
  BUFFD0 U8363 ( .I(n8390), .Z(n8447) );
  BUFFD0 U8364 ( .I(n8391), .Z(n8448) );
  CKBD0 U8365 ( .CLK(n8432), .C(n8449) );
  CKBD0 U8366 ( .CLK(n8433), .C(n8450) );
  CKBD0 U8367 ( .CLK(n8436), .C(n8451) );
  CKBD0 U8368 ( .CLK(n8437), .C(n8452) );
  CKBD0 U8369 ( .CLK(n8438), .C(n8453) );
  CKBD0 U8370 ( .CLK(n8439), .C(n8454) );
  CKBD0 U8371 ( .CLK(n8440), .C(n8455) );
  CKBD0 U8372 ( .CLK(n8441), .C(n8456) );
  BUFFD0 U8373 ( .I(n8388), .Z(n8457) );
  CKBD0 U8374 ( .CLK(n8389), .C(n8458) );
  CKBD0 U8375 ( .CLK(n8449), .C(n8459) );
  CKBD0 U8376 ( .CLK(n8450), .C(n8460) );
  CKBD0 U8377 ( .CLK(n8451), .C(n8461) );
  CKBD0 U8378 ( .CLK(n8452), .C(n8462) );
  CKBD0 U8379 ( .CLK(n8453), .C(n8463) );
  CKBD0 U8380 ( .CLK(n8454), .C(n8464) );
  CKBD0 U8381 ( .CLK(n8455), .C(n8465) );
  CKBD0 U8382 ( .CLK(n8456), .C(n8466) );
  CKBD0 U8383 ( .CLK(n8459), .C(n8467) );
  CKBD0 U8384 ( .CLK(n8460), .C(n8468) );
  CKBD0 U8385 ( .CLK(n8461), .C(n8469) );
  CKBD0 U8386 ( .CLK(n8462), .C(n8470) );
  CKBD0 U8387 ( .CLK(n8463), .C(n8471) );
  CKBD0 U8388 ( .CLK(n8403), .C(n8472) );
  CKBD0 U8389 ( .CLK(n8464), .C(n8473) );
  CKBD0 U8390 ( .CLK(n8406), .C(n8474) );
  CKBD0 U8391 ( .CLK(n8413), .C(n8475) );
  BUFFD0 U8392 ( .I(n8414), .Z(n8476) );
  CKBD0 U8393 ( .CLK(n8465), .C(n8477) );
  CKBD0 U8394 ( .CLK(n8415), .C(n8478) );
  CKBD0 U8395 ( .CLK(n8466), .C(n8479) );
  CKBD0 U8396 ( .CLK(n8467), .C(n8480) );
  CKBD0 U8397 ( .CLK(n8468), .C(n8481) );
  CKBD0 U8398 ( .CLK(n8469), .C(n8482) );
  CKBD0 U8399 ( .CLK(n8470), .C(n8483) );
  CKBD0 U8400 ( .CLK(n8471), .C(n8484) );
  CKBD0 U8401 ( .CLK(n8473), .C(n8485) );
  CKBD0 U8402 ( .CLK(n8477), .C(n8486) );
  CKBD0 U8403 ( .CLK(n8479), .C(n8487) );
  CKBD0 U8404 ( .CLK(n8480), .C(n8488) );
  CKBD0 U8405 ( .CLK(n8481), .C(n8489) );
  CKBD0 U8406 ( .CLK(n8482), .C(n8490) );
  CKBD0 U8407 ( .CLK(n8483), .C(n8491) );
  CKBD0 U8408 ( .CLK(n8484), .C(n8492) );
  CKBD0 U8409 ( .CLK(n8485), .C(n8493) );
  CKBD0 U8410 ( .CLK(n8486), .C(n8494) );
  BUFFD0 U8411 ( .I(n8487), .Z(n8495) );
  BUFFD0 U8412 ( .I(n8488), .Z(n8496) );
  BUFFD0 U8413 ( .I(n8489), .Z(n8497) );
  CKBD0 U8414 ( .CLK(n8490), .C(n8498) );
  BUFFD0 U8415 ( .I(n8491), .Z(n8499) );
  CKBD0 U8416 ( .CLK(n8492), .C(n8500) );
  CKBD0 U8417 ( .CLK(n8416), .C(n8501) );
  CKBD0 U8418 ( .CLK(n8417), .C(n8502) );
  BUFFD0 U8419 ( .I(n8419), .Z(n8503) );
  CKBD0 U8420 ( .CLK(n8428), .C(n8504) );
  BUFFD0 U8421 ( .I(n8427), .Z(n8505) );
  CKBD0 U8422 ( .CLK(n8430), .C(n8506) );
  BUFFD0 U8423 ( .I(n8493), .Z(n8507) );
  CKBD0 U8424 ( .CLK(n8494), .C(n8508) );
  CKBD0 U8425 ( .CLK(n8495), .C(n8509) );
  CKBD0 U8426 ( .CLK(n8496), .C(n8510) );
  CKBD0 U8427 ( .CLK(n8497), .C(n8511) );
  CKBD0 U8428 ( .CLK(n8498), .C(n8512) );
  CKBD0 U8429 ( .CLK(n8499), .C(n8513) );
  CKBD0 U8430 ( .CLK(n8500), .C(n8514) );
  BUFFD0 U8431 ( .I(n8429), .Z(n8515) );
  BUFFD0 U8432 ( .I(n8431), .Z(n8516) );
  CKBD0 U8433 ( .CLK(n8434), .C(n8517) );
  CKBD0 U8434 ( .CLK(n8442), .C(n8518) );
  BUFFD0 U8435 ( .I(n8435), .Z(n8519) );
  CKBD0 U8436 ( .CLK(n8443), .C(n8520) );
  CKBD0 U8437 ( .CLK(n8444), .C(n8521) );
  CKBD0 U8438 ( .CLK(n8507), .C(n8522) );
  CKBD0 U8439 ( .CLK(n8508), .C(n8523) );
  CKBD0 U8440 ( .CLK(n8509), .C(n8524) );
  CKBD0 U8441 ( .CLK(n8510), .C(n8525) );
  CKBD0 U8442 ( .CLK(n8511), .C(n8526) );
  CKBD0 U8443 ( .CLK(n8512), .C(n8527) );
  CKBD0 U8444 ( .CLK(n8513), .C(n8528) );
  CKBD0 U8445 ( .CLK(n8514), .C(n8529) );
  BUFFD0 U8446 ( .I(n8445), .Z(n8530) );
  CKBD0 U8447 ( .CLK(n8447), .C(n8531) );
  BUFFD0 U8448 ( .I(n8446), .Z(n8532) );
  CKBD0 U8449 ( .CLK(n8448), .C(n8533) );
  CKBD0 U8450 ( .CLK(n8457), .C(n8534) );
  BUFFD0 U8451 ( .I(n8458), .Z(n8535) );
  CKBD0 U8452 ( .CLK(n8522), .C(n8536) );
  BUFFD0 U8453 ( .I(n8523), .Z(n8537) );
  CKBD0 U8454 ( .CLK(n8524), .C(n8538) );
  CKBD0 U8455 ( .CLK(n8525), .C(n8539) );
  CKBD0 U8456 ( .CLK(n8526), .C(n8540) );
  BUFFD0 U8457 ( .I(n8472), .Z(n8541) );
  BUFFD0 U8458 ( .I(n8527), .Z(n8542) );
  BUFFD0 U8459 ( .I(n8474), .Z(n8543) );
  BUFFD0 U8460 ( .I(n8475), .Z(n8544) );
  CKBD0 U8461 ( .CLK(n8476), .C(n8545) );
  BUFFD0 U8462 ( .I(n8478), .Z(n8546) );
  BUFFD0 U8463 ( .I(n8501), .Z(n8547) );
  CKBD0 U8464 ( .CLK(n8528), .C(n8548) );
  BUFFD0 U8465 ( .I(n8502), .Z(n8549) );
  CKBD0 U8466 ( .CLK(n8503), .C(n8550) );
  CKBD0 U8467 ( .CLK(n8505), .C(n8551) );
  BUFFD0 U8468 ( .I(n8517), .Z(n8552) );
  BUFFD0 U8469 ( .I(n8504), .Z(n8553) );
  BUFFD0 U8470 ( .I(n8520), .Z(n8554) );
  CKBD0 U8471 ( .CLK(n8515), .C(n8555) );
  BUFFD0 U8472 ( .I(n8529), .Z(n8556) );
  CKBD0 U8473 ( .CLK(n8536), .C(n8557) );
  CKBD0 U8474 ( .CLK(n8537), .C(n8558) );
  CKBD0 U8475 ( .CLK(n8538), .C(n8559) );
  CKBD0 U8476 ( .CLK(n8539), .C(n8560) );
  CKBD0 U8477 ( .CLK(n8540), .C(n8561) );
  CKBD0 U8478 ( .CLK(n8542), .C(n8562) );
  BUFFD0 U8479 ( .I(n8506), .Z(n8563) );
  CKBD0 U8480 ( .CLK(n8516), .C(n8564) );
  CKBD0 U8481 ( .CLK(n8548), .C(n8565) );
  CKBD0 U8482 ( .CLK(n8519), .C(n8566) );
  BUFFD0 U8483 ( .I(n8531), .Z(n8567) );
  BUFFD0 U8484 ( .I(n8518), .Z(n8568) );
  BUFFD0 U8485 ( .I(n8533), .Z(n8569) );
  BUFFD0 U8486 ( .I(n8521), .Z(n8570) );
  CKBD0 U8487 ( .CLK(n8530), .C(n8571) );
  CKBD0 U8488 ( .CLK(n8532), .C(n8572) );
  CKBD0 U8489 ( .CLK(n8556), .C(n8573) );
  BUFFD0 U8490 ( .I(n8534), .Z(n8574) );
  CKBD0 U8491 ( .CLK(n8535), .C(n8575) );
  CKBD0 U8492 ( .CLK(n8557), .C(n8576) );
  CKBD0 U8493 ( .CLK(n8558), .C(n8577) );
  CKBD0 U8494 ( .CLK(n8559), .C(n8578) );
  CKBD0 U8495 ( .CLK(n8541), .C(n8579) );
  CKBD0 U8496 ( .CLK(n8560), .C(n8580) );
  CKBD0 U8497 ( .CLK(n8561), .C(n8581) );
  CKBD0 U8498 ( .CLK(n8543), .C(n8582) );
  CKBD0 U8499 ( .CLK(n8544), .C(n8583) );
  CKBD0 U8500 ( .CLK(n8562), .C(n8584) );
  CKBD0 U8501 ( .CLK(n8565), .C(n8585) );
  CKBD0 U8502 ( .CLK(n8573), .C(n8586) );
  CKBD0 U8503 ( .CLK(n8576), .C(n8587) );
  CKBD0 U8504 ( .CLK(n8577), .C(n8588) );
  CKBD0 U8505 ( .CLK(n8578), .C(n8589) );
  BUFFD0 U8506 ( .I(n8545), .Z(n8590) );
  CKBD0 U8507 ( .CLK(n8546), .C(n8591) );
  CKBD0 U8508 ( .CLK(n8547), .C(n8592) );
  CKBD0 U8509 ( .CLK(n8549), .C(n8593) );
  CKBD0 U8510 ( .CLK(n8580), .C(n8594) );
  CKBD0 U8511 ( .CLK(n8581), .C(n8595) );
  CKBD0 U8512 ( .CLK(n8584), .C(n8596) );
  CKBD0 U8513 ( .CLK(n8585), .C(n8597) );
  CKBD0 U8514 ( .CLK(n8586), .C(n8598) );
  CKBD0 U8515 ( .CLK(n8587), .C(n8599) );
  CKBD0 U8516 ( .CLK(n8588), .C(n8600) );
  CKBD0 U8517 ( .CLK(n8589), .C(n8601) );
  BUFFD0 U8518 ( .I(n8550), .Z(n8602) );
  CKBD0 U8519 ( .CLK(n8552), .C(n8603) );
  CKBD0 U8520 ( .CLK(n8553), .C(n8604) );
  BUFFD0 U8521 ( .I(n8551), .Z(n8605) );
  CKBD0 U8522 ( .CLK(n8563), .C(n8606) );
  CKBD0 U8523 ( .CLK(n8554), .C(n8607) );
  BUFFD0 U8524 ( .I(n8555), .Z(n8608) );
  BUFFD0 U8525 ( .I(n8564), .Z(n8609) );
  CKBD0 U8526 ( .CLK(n8594), .C(n8610) );
  CKBD0 U8527 ( .CLK(n8595), .C(n8611) );
  CKBD0 U8528 ( .CLK(n8568), .C(n8612) );
  CKBD0 U8529 ( .CLK(n8596), .C(n8613) );
  CKBD0 U8530 ( .CLK(n8597), .C(n8614) );
  CKBD0 U8531 ( .CLK(n8598), .C(n8615) );
  CKBD0 U8532 ( .CLK(n8599), .C(n8616) );
  CKBD0 U8533 ( .CLK(n8600), .C(n8617) );
  CKBD0 U8534 ( .CLK(n8601), .C(n8618) );
  CKBD0 U8535 ( .CLK(n8567), .C(n8619) );
  CKBD0 U8536 ( .CLK(n8569), .C(n8620) );
  BUFFD0 U8537 ( .I(n8566), .Z(n8621) );
  CKBD0 U8538 ( .CLK(n8570), .C(n8622) );
  BUFFD0 U8539 ( .I(n8571), .Z(n8623) );
  BUFFD0 U8540 ( .I(n8572), .Z(n8624) );
  CKBD0 U8541 ( .CLK(n8610), .C(n8625) );
  CKBD0 U8542 ( .CLK(n8611), .C(n8626) );
  CKBD0 U8543 ( .CLK(n8574), .C(n8627) );
  CKBD0 U8544 ( .CLK(n8613), .C(n8628) );
  CKBD0 U8545 ( .CLK(n8614), .C(n8629) );
  CKBD0 U8546 ( .CLK(n8615), .C(n8630) );
  CKBD0 U8547 ( .CLK(n8616), .C(n8631) );
  CKBD0 U8548 ( .CLK(n8617), .C(n8632) );
  CKBD0 U8549 ( .CLK(n8618), .C(n8633) );
  BUFFD0 U8550 ( .I(n8575), .Z(n8634) );
  CKBD0 U8551 ( .CLK(n8625), .C(n8635) );
  CKBD0 U8552 ( .CLK(n8626), .C(n8636) );
  CKBD0 U8553 ( .CLK(n8628), .C(n8637) );
  CKBD0 U8554 ( .CLK(n8629), .C(n8638) );
  CKBD0 U8555 ( .CLK(n8630), .C(n8639) );
  CKBD0 U8556 ( .CLK(n8631), .C(n8640) );
  BUFFD0 U8557 ( .I(n8579), .Z(n8641) );
  CKBD0 U8558 ( .CLK(n8632), .C(n8642) );
  BUFFD0 U8559 ( .I(n8582), .Z(n8643) );
  BUFFD0 U8560 ( .I(n8583), .Z(n8644) );
  CKBD0 U8561 ( .CLK(n8590), .C(n8645) );
  CKBD0 U8562 ( .CLK(n8633), .C(n8646) );
  CKBD0 U8563 ( .CLK(n8635), .C(n8647) );
  CKBD0 U8564 ( .CLK(n8636), .C(n8648) );
  CKBD0 U8565 ( .CLK(n8637), .C(n8649) );
  CKBD0 U8566 ( .CLK(n8638), .C(n8650) );
  CKBD0 U8567 ( .CLK(n8639), .C(n8651) );
  BUFFD0 U8568 ( .I(n8640), .Z(n8652) );
  CKBD0 U8569 ( .CLK(n8642), .C(n8653) );
  BUFFD0 U8570 ( .I(n8603), .Z(n8654) );
  BUFFD0 U8571 ( .I(n8591), .Z(n8655) );
  BUFFD0 U8572 ( .I(n8607), .Z(n8656) );
  BUFFD0 U8573 ( .I(n8592), .Z(n8657) );
  BUFFD0 U8574 ( .I(n8593), .Z(n8658) );
  CKBD0 U8575 ( .CLK(n8602), .C(n8659) );
  CKBD0 U8576 ( .CLK(n8605), .C(n8660) );
  BUFFD0 U8577 ( .I(n8604), .Z(n8661) );
  BUFFD0 U8578 ( .I(n8619), .Z(n8662) );
  BUFFD0 U8579 ( .I(n8620), .Z(n8663) );
  BUFFD0 U8580 ( .I(n8646), .Z(n8664) );
  BUFFD0 U8581 ( .I(n8647), .Z(n8665) );
  BUFFD0 U8582 ( .I(n8648), .Z(n8666) );
  CKBD0 U8583 ( .CLK(n8649), .C(n8667) );
  BUFFD0 U8584 ( .I(n8650), .Z(n8668) );
  CKBD0 U8585 ( .CLK(n8651), .C(n8669) );
  CKBD0 U8586 ( .CLK(n8652), .C(n8670) );
  CKBD0 U8587 ( .CLK(n8653), .C(n8671) );
  CKBD0 U8588 ( .CLK(n8608), .C(n8672) );
  CKBD0 U8589 ( .CLK(n8664), .C(n8673) );
  CKBD0 U8590 ( .CLK(n8665), .C(n8674) );
  CKBD0 U8591 ( .CLK(n8666), .C(n8675) );
  CKBD0 U8592 ( .CLK(n8667), .C(n8676) );
  CKBD0 U8593 ( .CLK(n8668), .C(n8677) );
  CKBD0 U8594 ( .CLK(n8669), .C(n8678) );
  CKBD0 U8595 ( .CLK(n8670), .C(n8679) );
  CKBD0 U8596 ( .CLK(n8671), .C(n8680) );
  CKBD0 U8597 ( .CLK(n8673), .C(n8681) );
  CKBD0 U8598 ( .CLK(n8674), .C(n8682) );
  CKBD0 U8599 ( .CLK(n8675), .C(n8683) );
  CKBD0 U8600 ( .CLK(n8676), .C(n8684) );
  CKBD0 U8601 ( .CLK(n8677), .C(n8685) );
  BUFFD0 U8602 ( .I(n8678), .Z(n8686) );
  CKBD0 U8603 ( .CLK(n8679), .C(n8687) );
  BUFFD0 U8604 ( .I(n8606), .Z(n8688) );
  CKBD0 U8605 ( .CLK(n8609), .C(n8689) );
  CKBD0 U8606 ( .CLK(n8621), .C(n8690) );
  BUFFD0 U8607 ( .I(n8612), .Z(n8691) );
  BUFFD0 U8608 ( .I(n8622), .Z(n8692) );
  CKBD0 U8609 ( .CLK(n8623), .C(n8693) );
  BUFFD0 U8610 ( .I(n8680), .Z(n8694) );
  CKBD0 U8611 ( .CLK(n8681), .C(n8695) );
  CKBD0 U8612 ( .CLK(n8682), .C(n8696) );
  CKBD0 U8613 ( .CLK(n8683), .C(n8697) );
  BUFFD0 U8614 ( .I(n8684), .Z(n8698) );
  CKBD0 U8615 ( .CLK(n8685), .C(n8699) );
  CKBD0 U8616 ( .CLK(n8686), .C(n8700) );
  CKBD0 U8617 ( .CLK(n8687), .C(n8701) );
  CKBD0 U8618 ( .CLK(n8624), .C(n8702) );
  CKBD0 U8619 ( .CLK(n8634), .C(n8703) );
  CKBD0 U8620 ( .CLK(n8694), .C(n8704) );
  BUFFD0 U8621 ( .I(n8627), .Z(n8705) );
  CKBD0 U8622 ( .CLK(n8695), .C(n8706) );
  CKBD0 U8623 ( .CLK(n8696), .C(n8707) );
  CKBD0 U8624 ( .CLK(n8697), .C(n8708) );
  CKBD0 U8625 ( .CLK(n8698), .C(n8709) );
  CKBD0 U8626 ( .CLK(n8641), .C(n8710) );
  CKBD0 U8627 ( .CLK(n8699), .C(n8711) );
  CKBD0 U8628 ( .CLK(n8643), .C(n8712) );
  CKBD0 U8629 ( .CLK(n8644), .C(n8713) );
  BUFFD0 U8630 ( .I(n8645), .Z(n8714) );
  CKBD0 U8631 ( .CLK(n8654), .C(n8715) );
  CKBD0 U8632 ( .CLK(n8655), .C(n8716) );
  CKBD0 U8633 ( .CLK(n8700), .C(n8717) );
  CKBD0 U8634 ( .CLK(n8657), .C(n8718) );
  CKBD0 U8635 ( .CLK(n8656), .C(n8719) );
  CKBD0 U8636 ( .CLK(n8701), .C(n8720) );
  CKBD0 U8637 ( .CLK(n8704), .C(n8721) );
  CKBD0 U8638 ( .CLK(n8706), .C(n8722) );
  CKBD0 U8639 ( .CLK(n8707), .C(n8723) );
  CKBD0 U8640 ( .CLK(n8708), .C(n8724) );
  CKBD0 U8641 ( .CLK(n8709), .C(n8725) );
  CKBD0 U8642 ( .CLK(n8711), .C(n8726) );
  BUFFD0 U8643 ( .I(n8659), .Z(n8727) );
  CKBD0 U8644 ( .CLK(n8661), .C(n8728) );
  BUFFD0 U8645 ( .I(n8660), .Z(n8729) );
  CKBD0 U8646 ( .CLK(n8662), .C(n8730) );
  CKBD0 U8647 ( .CLK(n8663), .C(n8731) );
  BUFFD0 U8648 ( .I(n8672), .Z(n8732) );
  CKBD0 U8649 ( .CLK(n8717), .C(n8733) );
  CKBD0 U8650 ( .CLK(n8658), .C(n8734) );
  BUFFD0 U8651 ( .I(n8689), .Z(n8735) );
  CKBD0 U8652 ( .CLK(n8691), .C(n8736) );
  BUFFD0 U8653 ( .I(n8690), .Z(n8737) );
  CKBD0 U8654 ( .CLK(n8692), .C(n8738) );
  CKBD0 U8655 ( .CLK(n8688), .C(n8739) );
  BUFFD0 U8656 ( .I(n8693), .Z(n8740) );
  BUFFD0 U8657 ( .I(n8702), .Z(n8741) );
  BUFFD0 U8658 ( .I(n8703), .Z(n8742) );
  CKBD0 U8659 ( .CLK(n8720), .C(n8743) );
  CKBD0 U8660 ( .CLK(n8721), .C(n8744) );
  CKBD0 U8661 ( .CLK(n8705), .C(n8745) );
  CKBD0 U8662 ( .CLK(n8722), .C(n8746) );
  CKBD0 U8663 ( .CLK(n8723), .C(n8747) );
  CKBD0 U8664 ( .CLK(n8724), .C(n8748) );
  BUFFD0 U8665 ( .I(n8710), .Z(n8749) );
  CKBD0 U8666 ( .CLK(n8725), .C(n8750) );
  BUFFD0 U8667 ( .I(n8715), .Z(n8751) );
  BUFFD0 U8668 ( .I(n8719), .Z(n8752) );
  BUFFD0 U8669 ( .I(n8712), .Z(n8753) );
  BUFFD0 U8670 ( .I(n8713), .Z(n8754) );
  CKBD0 U8671 ( .CLK(n8714), .C(n8755) );
  BUFFD0 U8672 ( .I(n8730), .Z(n8756) );
  BUFFD0 U8673 ( .I(n8716), .Z(n8757) );
  BUFFD0 U8674 ( .I(n8731), .Z(n8758) );
  BUFFD0 U8675 ( .I(n8718), .Z(n8759) );
  CKBD0 U8676 ( .CLK(n8726), .C(n8760) );
  CKBD0 U8677 ( .CLK(n8727), .C(n8761) );
  BUFFD0 U8678 ( .I(n8734), .Z(n8762) );
  CKBD0 U8679 ( .CLK(n8729), .C(n8763) );
  BUFFD0 U8680 ( .I(n8728), .Z(n8764) );
  CKBD0 U8681 ( .CLK(n8732), .C(n8765) );
  BUFFD0 U8682 ( .I(n8739), .Z(n8766) );
  CKBD0 U8683 ( .CLK(n8735), .C(n8767) );
  CKBD0 U8684 ( .CLK(n8733), .C(n8768) );
  CKBD0 U8685 ( .CLK(n8737), .C(n8769) );
  BUFFD0 U8686 ( .I(n8736), .Z(n8770) );
  BUFFD0 U8687 ( .I(n8738), .Z(n8771) );
  CKBD0 U8688 ( .CLK(n8740), .C(n8772) );
  CKBD0 U8689 ( .CLK(n8741), .C(n8773) );
  CKBD0 U8690 ( .CLK(n8742), .C(n8774) );
  CKBD0 U8691 ( .CLK(n8743), .C(n8775) );
  BUFFD0 U8692 ( .I(n8745), .Z(n8776) );
  CKBD0 U8693 ( .CLK(n8744), .C(n8777) );
  CKBD0 U8694 ( .CLK(n8746), .C(n8778) );
  CKBD0 U8695 ( .CLK(n8747), .C(n8779) );
  CKBD0 U8696 ( .CLK(n8748), .C(n8780) );
  CKBD0 U8697 ( .CLK(n8749), .C(n8781) );
  CKBD0 U8698 ( .CLK(n8751), .C(n8782) );
  CKBD0 U8699 ( .CLK(n8750), .C(n8783) );
  CKBD0 U8700 ( .CLK(n8753), .C(n8784) );
  CKBD0 U8701 ( .CLK(n8752), .C(n8785) );
  CKBD0 U8702 ( .CLK(n8754), .C(n8786) );
  BUFFD0 U8703 ( .I(n8755), .Z(n8787) );
  CKBD0 U8704 ( .CLK(n8757), .C(n8788) );
  CKBD0 U8705 ( .CLK(n8756), .C(n8789) );
  CKBD0 U8706 ( .CLK(n8758), .C(n8790) );
  CKBD0 U8707 ( .CLK(n8759), .C(n8791) );
  CKBD0 U8708 ( .CLK(n8762), .C(n8792) );
  BUFFD0 U8709 ( .I(n8761), .Z(n8793) );
  CKBD0 U8710 ( .CLK(n8760), .C(n8794) );
  CKBD0 U8711 ( .CLK(n8764), .C(n8795) );
  BUFFD0 U8712 ( .I(n8763), .Z(n8796) );
  CKBD0 U8713 ( .CLK(n8766), .C(n8797) );
  BUFFD0 U8714 ( .I(n8765), .Z(n8798) );
  BUFFD0 U8715 ( .I(n8767), .Z(n8799) );
  CKBD0 U8716 ( .CLK(n8768), .C(n8800) );
  CKBD0 U8717 ( .CLK(n8770), .C(n8801) );
  BUFFD0 U8718 ( .I(n8769), .Z(n8802) );
  CKBD0 U8719 ( .CLK(n8771), .C(n8803) );
  BUFFD0 U8720 ( .I(n8772), .Z(n8804) );
  BUFFD0 U8721 ( .I(n8773), .Z(n8805) );
  BUFFD0 U8722 ( .I(n8774), .Z(n8806) );
  CKBD0 U8723 ( .CLK(n8775), .C(n8807) );
  CKBD0 U8724 ( .CLK(n8776), .C(n8808) );
  CKBD0 U8725 ( .CLK(n8777), .C(n8809) );
  CKBD0 U8726 ( .CLK(n8778), .C(n8810) );
  BUFFD0 U8727 ( .I(n8782), .Z(n8811) );
  CKBD0 U8728 ( .CLK(n8779), .C(n8812) );
  CKBD0 U8729 ( .CLK(n8780), .C(n8813) );
  BUFFD0 U8730 ( .I(n8785), .Z(n8814) );
  CKBD0 U8731 ( .CLK(n8783), .C(n8815) );
  CKBD0 U8732 ( .CLK(n8794), .C(n8816) );
  CKBD0 U8733 ( .CLK(n8800), .C(n8817) );
  CKBD0 U8734 ( .CLK(n8807), .C(n8818) );
  CKBD0 U8735 ( .CLK(n8809), .C(n8819) );
  CKBD0 U8736 ( .CLK(n8810), .C(n8820) );
  BUFFD0 U8737 ( .I(n8781), .Z(n8821) );
  BUFFD0 U8738 ( .I(n8789), .Z(n8822) );
  BUFFD0 U8739 ( .I(n8790), .Z(n8823) );
  CKBD0 U8740 ( .CLK(n8812), .C(n8824) );
  CKBD0 U8741 ( .CLK(n8813), .C(n8825) );
  CKBD0 U8742 ( .CLK(n8815), .C(n8826) );
  CKBD0 U8743 ( .CLK(n8816), .C(n8827) );
  CKBD0 U8744 ( .CLK(n8817), .C(n8828) );
  CKBD0 U8745 ( .CLK(n8818), .C(n8829) );
  CKBD0 U8746 ( .CLK(n8819), .C(n8830) );
  CKBD0 U8747 ( .CLK(n8820), .C(n8831) );
  CKBD0 U8748 ( .CLK(n8824), .C(n8832) );
  CKBD0 U8749 ( .CLK(n8825), .C(n8833) );
  CKBD0 U8750 ( .CLK(n8826), .C(n8834) );
  CKBD0 U8751 ( .CLK(n8827), .C(n8835) );
  CKBD0 U8752 ( .CLK(n8828), .C(n8836) );
  BUFFD0 U8753 ( .I(n8829), .Z(n8837) );
  CKBD0 U8754 ( .CLK(n8830), .C(n8838) );
  BUFFD0 U8755 ( .I(n8831), .Z(n8839) );
  CKBD0 U8756 ( .CLK(n8787), .C(n8840) );
  CKBD0 U8757 ( .CLK(n8793), .C(n8841) );
  BUFFD0 U8758 ( .I(n8832), .Z(n8842) );
  BUFFD0 U8759 ( .I(n8833), .Z(n8843) );
  BUFFD0 U8760 ( .I(n8834), .Z(n8844) );
  BUFFD0 U8761 ( .I(n8835), .Z(n8845) );
  BUFFD0 U8762 ( .I(n8836), .Z(n8846) );
  CKBD0 U8763 ( .CLK(n8837), .C(n8847) );
  BUFFD0 U8764 ( .I(n8838), .Z(n8848) );
  CKBD0 U8765 ( .CLK(n8839), .C(n8849) );
  CKBD0 U8766 ( .CLK(n8796), .C(n8850) );
  CKBD0 U8767 ( .CLK(n8842), .C(n8851) );
  CKBD0 U8768 ( .CLK(n8843), .C(n8852) );
  CKBD0 U8769 ( .CLK(n8844), .C(n8853) );
  CKBD0 U8770 ( .CLK(n8845), .C(n8854) );
  CKBD0 U8771 ( .CLK(n8846), .C(n8855) );
  CKBD0 U8772 ( .CLK(n8847), .C(n8856) );
  CKBD0 U8773 ( .CLK(n8848), .C(n8857) );
  BUFFD0 U8774 ( .I(n8849), .Z(n8858) );
  CKBD0 U8775 ( .CLK(n8798), .C(n8859) );
  BUFFD0 U8776 ( .I(n8851), .Z(n8860) );
  BUFFD0 U8777 ( .I(n8852), .Z(n8861) );
  BUFFD0 U8778 ( .I(n8853), .Z(n8862) );
  BUFFD0 U8779 ( .I(n8854), .Z(n8863) );
  BUFFD0 U8780 ( .I(n8855), .Z(n8864) );
  BUFFD0 U8781 ( .I(n8856), .Z(n8865) );
  BUFFD0 U8782 ( .I(n8857), .Z(n8866) );
  CKBD0 U8783 ( .CLK(n8858), .C(n8867) );
  CKBD0 U8784 ( .CLK(n8860), .C(n8868) );
  CKBD0 U8785 ( .CLK(n8861), .C(n8869) );
  CKBD0 U8786 ( .CLK(n8862), .C(n8870) );
  CKBD0 U8787 ( .CLK(n8863), .C(n8871) );
  CKBD0 U8788 ( .CLK(n8864), .C(n8872) );
  CKBD0 U8789 ( .CLK(n8865), .C(n8873) );
  CKBD0 U8790 ( .CLK(n8866), .C(n8874) );
  BUFFD0 U8791 ( .I(n8867), .Z(n8875) );
  CKBD0 U8792 ( .CLK(n8804), .C(n8876) );
  BUFFD0 U8793 ( .I(n8868), .Z(n8877) );
  BUFFD0 U8794 ( .I(n8869), .Z(n8878) );
  BUFFD0 U8795 ( .I(n8870), .Z(n8879) );
  BUFFD0 U8796 ( .I(n8871), .Z(n8880) );
  BUFFD0 U8797 ( .I(n8872), .Z(n8881) );
  BUFFD0 U8798 ( .I(n8873), .Z(n8882) );
  BUFFD0 U8799 ( .I(n8874), .Z(n8883) );
  CKBD0 U8800 ( .CLK(n8875), .C(n8884) );
  CKBD0 U8801 ( .CLK(n8877), .C(n8885) );
  CKBD0 U8802 ( .CLK(n8878), .C(n8886) );
  CKBD0 U8803 ( .CLK(n8879), .C(n8887) );
  CKBD0 U8804 ( .CLK(n8880), .C(n8888) );
  CKBD0 U8805 ( .CLK(n8881), .C(n8889) );
  CKBD0 U8806 ( .CLK(n8882), .C(n8890) );
  CKBD0 U8807 ( .CLK(n8883), .C(n8891) );
  BUFFD0 U8808 ( .I(n8884), .Z(n8892) );
  CKBD0 U8809 ( .CLK(n8799), .C(n8893) );
  BUFFD0 U8810 ( .I(n8788), .Z(n8894) );
  BUFFD0 U8811 ( .I(n8784), .Z(n8895) );
  BUFFD0 U8812 ( .I(n8786), .Z(n8896) );
  BUFFD0 U8813 ( .I(n8885), .Z(n8897) );
  BUFFD0 U8814 ( .I(n8886), .Z(n8898) );
  BUFFD0 U8815 ( .I(n8795), .Z(n8899) );
  BUFFD0 U8816 ( .I(n8791), .Z(n8900) );
  CKBD0 U8817 ( .CLK(n8802), .C(n8901) );
  BUFFD0 U8818 ( .I(n8887), .Z(n8902) );
  CKBD0 U8819 ( .CLK(n8806), .C(n8903) );
  CKBD0 U8820 ( .CLK(n8805), .C(n8904) );
  BUFFD0 U8821 ( .I(n8792), .Z(n8905) );
  BUFFD0 U8822 ( .I(n8888), .Z(n8906) );
  BUFFD0 U8823 ( .I(n8803), .Z(n8907) );
  BUFFD0 U8824 ( .I(n8801), .Z(n8908) );
  BUFFD0 U8825 ( .I(n8797), .Z(n8909) );
  BUFFD0 U8826 ( .I(n8889), .Z(n8910) );
  BUFFD0 U8827 ( .I(n8890), .Z(n8911) );
  CKBD0 U8828 ( .CLK(n8811), .C(n8912) );
  CKBD0 U8829 ( .CLK(n8814), .C(n8913) );
  BUFFD0 U8830 ( .I(n8891), .Z(n8914) );
  CKBD0 U8831 ( .CLK(n8892), .C(n8915) );
  CKBD0 U8832 ( .CLK(n8897), .C(n8916) );
  CKBD0 U8833 ( .CLK(n8898), .C(n8917) );
  CKBD0 U8834 ( .CLK(n8902), .C(n8918) );
  CKBD0 U8835 ( .CLK(n8906), .C(n8919) );
  CKBD0 U8836 ( .CLK(n8910), .C(n8920) );
  CKBD0 U8837 ( .CLK(n8911), .C(n8921) );
  CKBD0 U8838 ( .CLK(n8914), .C(n8922) );
  BUFFD0 U8839 ( .I(n8915), .Z(n8923) );
  BUFFD0 U8840 ( .I(n8916), .Z(n8924) );
  BUFFD0 U8841 ( .I(n8917), .Z(n8925) );
  BUFFD0 U8842 ( .I(n8918), .Z(n8926) );
  BUFFD0 U8843 ( .I(n8919), .Z(n8927) );
  BUFFD0 U8844 ( .I(n8920), .Z(n8928) );
  BUFFD0 U8845 ( .I(n8921), .Z(n8929) );
  CKBD0 U8846 ( .CLK(n8822), .C(n8930) );
  CKBD0 U8847 ( .CLK(n8823), .C(n8931) );
  BUFFD0 U8848 ( .I(n8922), .Z(n8932) );
  CKBD0 U8849 ( .CLK(n8923), .C(n8933) );
  CKBD0 U8850 ( .CLK(n8924), .C(n8934) );
  CKBD0 U8851 ( .CLK(n8925), .C(n8935) );
  CKBD0 U8852 ( .CLK(n8926), .C(n8936) );
  CKBD0 U8853 ( .CLK(n8927), .C(n8937) );
  CKBD0 U8854 ( .CLK(n8928), .C(n8938) );
  CKBD0 U8855 ( .CLK(n8929), .C(n8939) );
  CKBD0 U8856 ( .CLK(n8932), .C(n8940) );
  BUFFD0 U8857 ( .I(n8933), .Z(n8941) );
  BUFFD0 U8858 ( .I(n8934), .Z(n8942) );
  BUFFD0 U8859 ( .I(n8935), .Z(n8943) );
  BUFFD0 U8860 ( .I(n8936), .Z(n8944) );
  BUFFD0 U8861 ( .I(n8937), .Z(n8945) );
  BUFFD0 U8862 ( .I(n8938), .Z(n8946) );
  BUFFD0 U8863 ( .I(n8939), .Z(n8947) );
  BUFFD0 U8864 ( .I(n8940), .Z(n8948) );
  BUFFD0 U8865 ( .I(n8808), .Z(n8949) );
  CKBD0 U8866 ( .CLK(n8941), .C(n8950) );
  CKBD0 U8867 ( .CLK(n8821), .C(n8951) );
  CKBD0 U8868 ( .CLK(n8942), .C(n8952) );
  CKBD0 U8869 ( .CLK(n8943), .C(n8953) );
  CKBD0 U8870 ( .CLK(n8894), .C(n8954) );
  CKBD0 U8871 ( .CLK(n8895), .C(n8955) );
  CKBD0 U8872 ( .CLK(n8896), .C(n8956) );
  CKBD0 U8873 ( .CLK(n8944), .C(n8957) );
  CKBD0 U8874 ( .CLK(n8899), .C(n8958) );
  CKBD0 U8875 ( .CLK(n8900), .C(n8959) );
  BUFFD0 U8876 ( .I(n8840), .Z(n8960) );
  CKBD0 U8877 ( .CLK(n8945), .C(n8961) );
  BUFFD0 U8878 ( .I(n8841), .Z(n8962) );
  BUFFD0 U8879 ( .I(n8850), .Z(n8963) );
  BUFFD0 U8880 ( .I(n8859), .Z(n8964) );
  CKBD0 U8881 ( .CLK(n8905), .C(n8965) );
  BUFFD0 U8882 ( .I(n8893), .Z(n8966) );
  CKBD0 U8883 ( .CLK(n8907), .C(n8967) );
  CKBD0 U8884 ( .CLK(n8946), .C(n8968) );
  CKBD0 U8885 ( .CLK(n8908), .C(n8969) );
  BUFFD0 U8886 ( .I(n8876), .Z(n8970) );
  CKBD0 U8887 ( .CLK(n8909), .C(n8971) );
  BUFFD0 U8888 ( .I(n8901), .Z(n8972) );
  BUFFD0 U8889 ( .I(n8903), .Z(n8973) );
  BUFFD0 U8890 ( .I(n8904), .Z(n8974) );
  CKBD0 U8891 ( .CLK(n8947), .C(n8975) );
  CKBD0 U8892 ( .CLK(n8948), .C(n8976) );
  CKBD0 U8893 ( .CLK(n8949), .C(n8977) );
  BUFFD0 U8894 ( .I(n8912), .Z(n8978) );
  BUFFD0 U8895 ( .I(n8913), .Z(n8979) );
  BUFFD0 U8896 ( .I(n8930), .Z(n8980) );
  BUFFD0 U8897 ( .I(n8950), .Z(n8981) );
  BUFFD0 U8898 ( .I(n8931), .Z(n8982) );
  BUFFD0 U8899 ( .I(n8952), .Z(n8983) );
  BUFFD0 U8900 ( .I(n8953), .Z(n8984) );
  BUFFD0 U8901 ( .I(n8957), .Z(n8985) );
  BUFFD0 U8902 ( .I(n8961), .Z(n8986) );
  BUFFD0 U8903 ( .I(n8968), .Z(n8987) );
  BUFFD0 U8904 ( .I(n8951), .Z(n8988) );
  BUFFD0 U8905 ( .I(n8954), .Z(n8989) );
  BUFFD0 U8906 ( .I(n8955), .Z(n8990) );
  BUFFD0 U8907 ( .I(n8956), .Z(n8991) );
  BUFFD0 U8908 ( .I(n8958), .Z(n8992) );
  BUFFD0 U8909 ( .I(n8959), .Z(n8993) );
  BUFFD0 U8910 ( .I(n8975), .Z(n8994) );
  BUFFD0 U8911 ( .I(n8976), .Z(n8995) );
  BUFFD0 U8912 ( .I(n8965), .Z(n8996) );
  BUFFD0 U8913 ( .I(n8971), .Z(n8997) );
  CKBD0 U8914 ( .CLK(n8981), .C(n8998) );
  CKBD0 U8915 ( .CLK(n8983), .C(n8999) );
  CKBD0 U8916 ( .CLK(n8984), .C(n9000) );
  CKBD0 U8917 ( .CLK(n8985), .C(n9001) );
  CKBD0 U8918 ( .CLK(n8986), .C(n9002) );
  CKBD0 U8919 ( .CLK(n8987), .C(n9003) );
  CKBD0 U8920 ( .CLK(n8994), .C(n9004) );
  CKBD0 U8921 ( .CLK(n8995), .C(n9005) );
  BUFFD0 U8922 ( .I(n9275), .Z(n9006) );
  BUFFD0 U8923 ( .I(n8998), .Z(n9007) );
  BUFFD0 U8924 ( .I(n8969), .Z(n9008) );
  BUFFD0 U8925 ( .I(n8967), .Z(n9009) );
  BUFFD0 U8926 ( .I(n8999), .Z(n9010) );
  BUFFD0 U8927 ( .I(n9000), .Z(n9011) );
  BUFFD0 U8928 ( .I(n9001), .Z(n9012) );
  BUFFD0 U8929 ( .I(n8977), .Z(n9013) );
  BUFFD0 U8930 ( .I(n9002), .Z(n9014) );
  BUFFD0 U8931 ( .I(n9003), .Z(n9015) );
  BUFFD0 U8932 ( .I(n9004), .Z(n9016) );
  BUFFD0 U8933 ( .I(n9005), .Z(n9017) );
  BUFFD0 U8934 ( .I(n9126), .Z(n9018) );
  INR2XD0 U8935 ( .A1(n9027), .B1(n9127), .ZN(n9225) );
  BUFFD0 U8936 ( .I(n9020), .Z(n9019) );
  BUFFD0 U8937 ( .I(n9225), .Z(n9020) );
  CKBD0 U8938 ( .CLK(ParValidTimer[1]), .C(n9021) );
  BUFFD0 U8939 ( .I(n9224), .Z(n9022) );
  BUFFD0 U8940 ( .I(n9024), .Z(n9023) );
  BUFFD0 U8941 ( .I(n9280), .Z(n9024) );
  BUFFD1 U8942 ( .I(n9149), .Z(n9150) );
  BUFFD1 U8943 ( .I(n9151), .Z(n9149) );
  BUFFD1 U8944 ( .I(n9152), .Z(n9148) );
  BUFFD1 U8945 ( .I(n9152), .Z(n9147) );
  BUFFD1 U8946 ( .I(n9153), .Z(n9151) );
  BUFFD1 U8947 ( .I(n9153), .Z(n9152) );
  BUFFD1 U8948 ( .I(n9154), .Z(n9153) );
  INVD1 U8949 ( .I(Reset), .ZN(n9154) );
  INVD1 U8950 ( .I(n9275), .ZN(n9126) );
  BUFFD1 U8951 ( .I(n9130), .Z(n9137) );
  BUFFD1 U8952 ( .I(n9130), .Z(n9138) );
  BUFFD1 U8953 ( .I(n9131), .Z(n9139) );
  BUFFD1 U8954 ( .I(n9131), .Z(n9140) );
  BUFFD1 U8955 ( .I(n9132), .Z(n9141) );
  BUFFD1 U8956 ( .I(n9132), .Z(n9142) );
  BUFFD1 U8957 ( .I(n9133), .Z(n9143) );
  BUFFD1 U8958 ( .I(n9133), .Z(n9144) );
  BUFFD1 U8959 ( .I(n9134), .Z(n9145) );
  BUFFD1 U8960 ( .I(n9134), .Z(n9146) );
  INVD1 U8961 ( .I(n9156), .ZN(n9127) );
  INVD1 U8962 ( .I(n9156), .ZN(n9128) );
  INVD1 U8963 ( .I(n9156), .ZN(n9129) );
  BUFFD1 U8964 ( .I(n9135), .Z(n9132) );
  BUFFD1 U8965 ( .I(n9135), .Z(n9133) );
  BUFFD1 U8966 ( .I(n9131), .Z(n9134) );
  BUFFD1 U8967 ( .I(n9136), .Z(n9130) );
  BUFFD1 U8968 ( .I(n9136), .Z(n9131) );
  IND2D1 U8969 ( .A1(n9274), .B1(n9273), .ZN(n9275) );
  BUFFD1 U8970 ( .I(SerClock), .Z(n9135) );
  BUFFD1 U8971 ( .I(SerClock), .Z(n9136) );
  NR2D1 U8972 ( .A1(ParClk), .A2(n9155), .ZN(n9283) );
  NR2D1 U8973 ( .A1(ParClk), .A2(n9261), .ZN(N37) );
  NR4D0 U8974 ( .A1(n9260), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n9262) );
  AN2D1 U8975 ( .A1(N34), .A2(n9284), .Z(N42) );
  AN2D1 U8976 ( .A1(N33), .A2(n9284), .Z(N41) );
  AN2D1 U8977 ( .A1(N32), .A2(n9284), .Z(N40) );
  AN2D1 U8978 ( .A1(N31), .A2(n9284), .Z(N39) );
  INVD1 U8979 ( .I(n9021), .ZN(n9281) );
  AO22D0 U8980 ( .A1(n6915), .A2(n9018), .B1(n6780), .B2(n9275), .Z(n9189) );
  AO22D0 U8981 ( .A1(n6778), .A2(n9018), .B1(n6643), .B2(n9275), .Z(n9188) );
  AO22D0 U8982 ( .A1(n6641), .A2(n9018), .B1(n6506), .B2(n9275), .Z(n9187) );
  AO22D0 U8983 ( .A1(n6504), .A2(n9018), .B1(n6369), .B2(n9006), .Z(n9186) );
  AO22D0 U8984 ( .A1(n6367), .A2(n9018), .B1(n6232), .B2(n9275), .Z(n9185) );
  AO22D0 U8985 ( .A1(n6230), .A2(n9018), .B1(n6095), .B2(n9275), .Z(n9184) );
  AO22D0 U8986 ( .A1(n6093), .A2(n9018), .B1(n5957), .B2(n9006), .Z(n9183) );
  AO22D0 U8987 ( .A1(n5956), .A2(n9018), .B1(Decoder[7]), .B2(n9275), .Z(n9182) );
  AO22D0 U8988 ( .A1(n5820), .A2(n9126), .B1(Decoder[8]), .B2(n9275), .Z(n9181) );
  AO22D0 U8989 ( .A1(n5684), .A2(n9126), .B1(Decoder[9]), .B2(n9275), .Z(n9180) );
  AO22D0 U8990 ( .A1(n5548), .A2(n9126), .B1(Decoder[10]), .B2(n9275), .Z(
        n9179) );
  AO22D0 U8991 ( .A1(n5412), .A2(n9018), .B1(Decoder[11]), .B2(n9275), .Z(
        n9178) );
  AO22D0 U8992 ( .A1(n5276), .A2(n9018), .B1(n5140), .B2(n9275), .Z(n9177) );
  AO22D0 U8993 ( .A1(n5139), .A2(n9126), .B1(Decoder[13]), .B2(n9275), .Z(
        n9176) );
  AO22D0 U8994 ( .A1(n5003), .A2(n9126), .B1(Decoder[14]), .B2(n9275), .Z(
        n9175) );
  AO22D0 U8995 ( .A1(n4867), .A2(n9126), .B1(Decoder[15]), .B2(n9275), .Z(
        n9174) );
  AO22D0 U8996 ( .A1(n4731), .A2(n9126), .B1(Decoder[16]), .B2(n9006), .Z(
        n9173) );
  AO22D0 U8997 ( .A1(n4595), .A2(n9126), .B1(Decoder[17]), .B2(n9006), .Z(
        n9172) );
  AO22D0 U8998 ( .A1(n4459), .A2(n9126), .B1(Decoder[18]), .B2(n9006), .Z(
        n9171) );
  AO22D0 U8999 ( .A1(n4323), .A2(n9126), .B1(n4187), .B2(n9006), .Z(n9170) );
  AO22D0 U9000 ( .A1(n4186), .A2(n9126), .B1(Decoder[20]), .B2(n9006), .Z(
        n9169) );
  AO22D0 U9001 ( .A1(n4050), .A2(n9018), .B1(Decoder[21]), .B2(n9006), .Z(
        n9168) );
  AO22D0 U9002 ( .A1(n3914), .A2(n9126), .B1(Decoder[22]), .B2(n9006), .Z(
        n9167) );
  AO22D0 U9003 ( .A1(n3778), .A2(n9018), .B1(Decoder[23]), .B2(n9006), .Z(
        n9166) );
  AO22D0 U9004 ( .A1(n3642), .A2(n9126), .B1(Decoder[24]), .B2(n9006), .Z(
        n9165) );
  AO22D0 U9005 ( .A1(n3506), .A2(n9126), .B1(Decoder[25]), .B2(n9006), .Z(
        n9164) );
  AO22D0 U9006 ( .A1(n3370), .A2(n9126), .B1(Decoder[26]), .B2(n9006), .Z(
        n9163) );
  AO22D0 U9007 ( .A1(n3234), .A2(n9126), .B1(Decoder[27]), .B2(n9006), .Z(
        n9162) );
  AO22D0 U9008 ( .A1(n3098), .A2(n9018), .B1(Decoder[28]), .B2(n9275), .Z(
        n9161) );
  AO22D0 U9009 ( .A1(n2962), .A2(n9126), .B1(Decoder[29]), .B2(n9006), .Z(
        n9160) );
  AO22D0 U9010 ( .A1(n2826), .A2(n9126), .B1(Decoder[30]), .B2(n9006), .Z(
        n9159) );
  AO22D0 U9011 ( .A1(n2687), .A2(n9126), .B1(Decoder[31]), .B2(n9006), .Z(
        n9158) );
  OAI31D0 U9012 ( .A1(n9282), .A2(n9157), .A3(n9281), .B(n9155), .ZN(n9027) );
  NR2D1 U9013 ( .A1(n9277), .A2(n9127), .ZN(n9223) );
  NR2D1 U9014 ( .A1(n6921), .A2(n9127), .ZN(n9222) );
  NR2D1 U9015 ( .A1(n9127), .A2(n9023), .ZN(n9224) );
  XOR2D1 U9016 ( .A1(n9157), .A2(n9279), .Z(n9280) );
  NR2D1 U9017 ( .A1(n9281), .A2(n9278), .ZN(n9279) );
  NR4D0 U9018 ( .A1(n9266), .A2(n8996), .A3(n8991), .A4(n8988), .ZN(n9267) );
  NR4D0 U9019 ( .A1(n9016), .A2(n9014), .A3(n9010), .A4(n9007), .ZN(n9272) );
  NR4D0 U9020 ( .A1(n9017), .A2(n9015), .A3(n9012), .A4(n9011), .ZN(n9271) );
  AN4D1 U9021 ( .A1(n9270), .A2(n9269), .A3(n9268), .A4(n9267), .Z(n9273) );
  INR4D0 U9022 ( .A1(n8982), .B1(n9263), .B2(n9009), .B3(n9013), .ZN(n9270) );
  NR4D0 U9023 ( .A1(n9264), .A2(n9008), .A3(n8992), .A4(n8989), .ZN(n9269) );
  NR4D0 U9024 ( .A1(n9265), .A2(n8997), .A3(n8993), .A4(n8990), .ZN(n9268) );
  ND3D1 U9025 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n9263) );
  AN2D1 U9026 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_1 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_1 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N46, N47, N48, N49, N63, N64, N65, N66, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n53, n70, n71,
         n91, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n25), .CPN(StateClock), .Q(FullFIFO), .QN(n30) );
  DFND1 EmptyFIFOr_reg ( .D(n26), .CPN(StateClock), .Q(EmptyFIFO) );
  IAO21D1 U6 ( .A1(n168), .A2(n167), .B(Reset), .ZN(n169) );
  MOAI22D1 U7 ( .A1(n12), .A2(n166), .B1(n166), .B2(OldReadAr[1]), .ZN(n24) );
  MOAI22D1 U8 ( .A1(n13), .A2(n166), .B1(n166), .B2(OldReadAr[2]), .ZN(n23) );
  MOAI22D1 U9 ( .A1(n165), .A2(n164), .B1(n165), .B2(OldWriteAr[1]), .ZN(n22)
         );
  MOAI22D1 U10 ( .A1(n165), .A2(n163), .B1(n165), .B2(OldWriteAr[2]), .ZN(n21)
         );
  MOAI22D1 U11 ( .A1(n10), .A2(n165), .B1(n165), .B2(OldWriteAr[0]), .ZN(n20)
         );
  MOAI22D1 U70 ( .A1(n11), .A2(n166), .B1(n166), .B2(OldReadAr[0]), .ZN(n14)
         );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n14), .CPN(StateClock), .CDN(n9), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n20), .CPN(StateClock), .CDN(n9), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n21), .CPN(StateClock), .CDN(n9), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n22), .CPN(StateClock), .CDN(n9), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n23), .CPN(StateClock), .CDN(n9), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n24), .CPN(StateClock), .CDN(n9), .Q(
        OldReadAr[1]) );
  DFNCND1 ReadCmdr_reg ( .D(n15), .CPN(StateClock), .CDN(n9), .Q(ReadCmd) );
  DFNCND1 WriteCmdr_reg ( .D(n17), .CPN(StateClock), .CDN(n9), .Q(WriteCmd) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n9), .Q(
        CurState[2]), .QN(n140) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n9), .Q(
        CurState[1]), .QN(n156) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n9), .Q(
        CurState[0]), .QN(n131) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N65), .E(N66), .CP(StateClock), .CDN(n9), .Q(
        WriteAddr[2]), .QN(n163) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N64), .E(N66), .CP(StateClock), .CDN(n9), .Q(
        WriteAddr[1]), .QN(n164) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N48), .CP(StateClock), .CDN(n9), .Q(
        ReadAddr[2]), .QN(n13) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N47), .E(N48), .CP(StateClock), .CDN(n9), .Q(
        ReadAddr[1]), .QN(n12) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N46), .E(N48), .CP(StateClock), .CDN(n9), .Q(
        ReadAddr[0]), .QN(n11) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N63), .E(N66), .CP(StateClock), .CDN(n9), .Q(
        WriteAddr[0]), .QN(n10) );
  DFNCND1 \NextState_reg[1]  ( .D(n18), .CPN(StateClock), .CDN(n9), .Q(
        NextState[1]), .QN(n28) );
  DFNCND1 \NextState_reg[0]  ( .D(n16), .CPN(StateClock), .CDN(n9), .Q(
        NextState[0]), .QN(n27) );
  DFNCND1 \NextState_reg[2]  ( .D(n19), .CPN(StateClock), .CDN(n9), .Q(
        NextState[2]), .QN(n29) );
  INVD1 U3 ( .I(Reset), .ZN(n9) );
  INVD1 U4 ( .I(n133), .ZN(n126) );
  INVD1 U5 ( .I(n161), .ZN(n155) );
  MAOI22D0 U12 ( .A1(ReadAddr[0]), .A2(n135), .B1(n164), .B2(n113), .ZN(n110)
         );
  XNR2D1 U13 ( .A1(n163), .A2(n135), .ZN(n133) );
  INVD1 U14 ( .I(n135), .ZN(n129) );
  XNR2D1 U15 ( .A1(n126), .A2(ReadAddr[2]), .ZN(n152) );
  INVD1 U16 ( .I(n167), .ZN(n172) );
  ND2D1 U17 ( .A1(n127), .A2(n170), .ZN(n124) );
  ND3D1 U18 ( .A1(n170), .A2(n172), .A3(n32), .ZN(N66) );
  NR2D1 U19 ( .A1(n140), .A2(n131), .ZN(n168) );
  ND2D1 U20 ( .A1(n127), .A2(n172), .ZN(n162) );
  NR2D1 U21 ( .A1(ReadAddr[0]), .A2(n53), .ZN(N46) );
  NR2D1 U22 ( .A1(n112), .A2(n53), .ZN(N49) );
  NR2D1 U23 ( .A1(n31), .A2(n53), .ZN(N47) );
  XNR2D1 U24 ( .A1(ReadAddr[0]), .A2(ReadAddr[1]), .ZN(n31) );
  OAI211D1 U25 ( .A1(CurState[1]), .A2(n131), .B(n127), .C(n107), .ZN(n161) );
  AOI21D1 U26 ( .A1(WriteReq), .A2(n167), .B(n106), .ZN(n107) );
  AOI21D1 U27 ( .A1(CurState[0]), .A2(n91), .B(n140), .ZN(n106) );
  OAI33D1 U28 ( .A1(n125), .A2(n167), .A3(n124), .B1(n123), .B2(n122), .B3(
        n121), .ZN(n17) );
  INVD1 U29 ( .I(WriteCmd), .ZN(n125) );
  XNR2D1 U30 ( .A1(n163), .A2(OldWriteAr[2]), .ZN(n121) );
  XNR2D1 U31 ( .A1(n164), .A2(OldWriteAr[1]), .ZN(n122) );
  ND2D1 U32 ( .A1(WriteReq), .A2(n162), .ZN(n165) );
  OAI22D0 U33 ( .A1(n161), .A2(n28), .B1(n155), .B2(n149), .ZN(n18) );
  AOI31D0 U34 ( .A1(n148), .A2(n147), .A3(n146), .B(n167), .ZN(n149) );
  IIND4D1 U35 ( .A1(n139), .A2(n137), .B1(n132), .B2(n131), .ZN(n147) );
  AOI31D0 U36 ( .A1(n11), .A2(CurState[0]), .A3(n145), .B(n144), .ZN(n146) );
  OAI22D0 U37 ( .A1(n161), .A2(n27), .B1(n155), .B2(n119), .ZN(n16) );
  AOI21D1 U38 ( .A1(CurState[1]), .A2(n118), .B(n168), .ZN(n119) );
  OAI21D1 U39 ( .A1(CurState[2]), .A2(n117), .B(n116), .ZN(n118) );
  AOI22D0 U40 ( .A1(n153), .A2(ReadAddr[2]), .B1(n13), .B2(n154), .ZN(n117) );
  OAI31D0 U41 ( .A1(n172), .A2(WriteReq), .A3(Reset), .B(n171), .ZN(n26) );
  OAI31D0 U42 ( .A1(CurState[0]), .A2(Reset), .A3(CurState[2]), .B(EmptyFIFO), 
        .ZN(n171) );
  OAI21D1 U43 ( .A1(n161), .A2(n29), .B(n160), .ZN(n19) );
  OAI211D1 U44 ( .A1(CurState[2]), .A2(n159), .B(CurState[0]), .C(n158), .ZN(
        n160) );
  NR4D0 U45 ( .A1(n152), .A2(n151), .A3(n156), .A4(n150), .ZN(n159) );
  AOI21D1 U46 ( .A1(n157), .A2(n156), .B(n155), .ZN(n158) );
  ND3D1 U47 ( .A1(n120), .A2(n162), .A3(WriteReq), .ZN(n123) );
  XNR2D1 U48 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n120) );
  MAOI22D0 U49 ( .A1(WriteAddr[0]), .A2(n108), .B1(n12), .B2(n113), .ZN(n109)
         );
  OAI33D1 U50 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n110), .B1(n163), 
        .B2(WriteAddr[1]), .B3(n109), .ZN(n154) );
  OAI33D1 U51 ( .A1(ReadAddr[1]), .A2(n110), .A3(n163), .B1(n109), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n153) );
  NR2D1 U52 ( .A1(n164), .A2(n10), .ZN(n135) );
  OAI21D1 U53 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n129), .ZN(n111) );
  XOR2D1 U54 ( .A1(n111), .A2(n12), .Z(n151) );
  AOI31D0 U55 ( .A1(n10), .A2(CurState[0]), .A3(n128), .B(n127), .ZN(n148) );
  NR3D0 U56 ( .A1(n151), .A2(n11), .A3(n152), .ZN(n128) );
  OAI31D0 U57 ( .A1(n115), .A2(n114), .A3(n150), .B(CurState[0]), .ZN(n116) );
  XNR2D1 U58 ( .A1(WriteAddr[2]), .A2(n112), .ZN(n114) );
  INVD1 U59 ( .I(n151), .ZN(n115) );
  NR3D0 U60 ( .A1(n151), .A2(n10), .A3(n136), .ZN(n145) );
  AOI21D1 U61 ( .A1(n139), .A2(n135), .B(n134), .ZN(n136) );
  OAI32D1 U62 ( .A1(n163), .A2(n13), .A3(n135), .B1(ReadAddr[2]), .B2(n133), 
        .ZN(n134) );
  AO22D0 U63 ( .A1(ReadAddr[2]), .A2(n154), .B1(n153), .B2(n13), .Z(n157) );
  OAI222D0 U64 ( .A1(n163), .A2(ReadAddr[2]), .B1(n164), .B2(ReadAddr[1]), 
        .C1(n10), .C2(ReadAddr[0]), .ZN(n137) );
  AOI22D0 U65 ( .A1(n140), .A2(CurState[1]), .B1(n156), .B2(n168), .ZN(n127)
         );
  NR3D0 U66 ( .A1(CurState[1]), .A2(CurState[2]), .A3(CurState[0]), .ZN(n167)
         );
  ND2D1 U67 ( .A1(CurState[1]), .A2(n168), .ZN(n170) );
  ND2D1 U68 ( .A1(ReadCmd), .A2(n172), .ZN(n53) );
  OAI21D1 U69 ( .A1(n10), .A2(n11), .B(n113), .ZN(n150) );
  OAI32D0 U71 ( .A1(n170), .A2(Reset), .A3(ReadReq), .B1(n169), .B2(n30), .ZN(
        n25) );
  ND2D1 U72 ( .A1(WriteCmd), .A2(n170), .ZN(n32) );
  OAI211D1 U73 ( .A1(n10), .A2(ReadAddr[1]), .B(n130), .C(n129), .ZN(n132) );
  OAI21D1 U74 ( .A1(WriteAddr[1]), .A2(n12), .B(n11), .ZN(n130) );
  CKND2D0 U75 ( .A1(ReadReq), .A2(n124), .ZN(n166) );
  NR2D1 U76 ( .A1(WriteAddr[2]), .A2(n13), .ZN(n139) );
  ND2D1 U77 ( .A1(n10), .A2(n11), .ZN(n113) );
  OAI22D0 U78 ( .A1(n11), .A2(n170), .B1(WriteAddr[0]), .B2(n32), .ZN(N63) );
  OAI22D0 U79 ( .A1(n13), .A2(n170), .B1(n126), .B2(n32), .ZN(N65) );
  OAI22D0 U80 ( .A1(n12), .A2(n170), .B1(n111), .B2(n32), .ZN(N64) );
  AOI31D0 U81 ( .A1(n143), .A2(n142), .A3(n141), .B(n140), .ZN(n144) );
  AOI22D0 U82 ( .A1(n139), .A2(ReadAddr[1]), .B1(n10), .B2(ReadAddr[0]), .ZN(
        n141) );
  OAI21D1 U83 ( .A1(n139), .A2(n137), .B(n164), .ZN(n143) );
  OAI21D1 U84 ( .A1(ReadAddr[1]), .A2(n138), .B(n137), .ZN(n142) );
  OAI32D1 U85 ( .A1(n71), .A2(n70), .A3(n91), .B1(n124), .B2(n53), .ZN(n15) );
  XNR2D1 U86 ( .A1(n12), .A2(OldReadAr[1]), .ZN(n70) );
  ND3D1 U87 ( .A1(n34), .A2(n124), .A3(n33), .ZN(n71) );
  XNR2D1 U88 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .ZN(n34) );
  IND2D1 U89 ( .A1(ReadCmd), .B1(n172), .ZN(N48) );
  NR2D1 U90 ( .A1(n11), .A2(n12), .ZN(n108) );
  XOR2D1 U91 ( .A1(n108), .A2(n13), .Z(n112) );
  XNR2D1 U92 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n138) );
  XNR2D1 U93 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n33) );
  ND2D1 U94 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U95 ( .I(ReadReq), .ZN(n91) );
endmodule


module DPMem1kx32_AWid3_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockW, Dreadyr, \Storage[7][32] , \Storage[7][31] ,
         \Storage[7][30] , \Storage[7][29] , \Storage[7][28] ,
         \Storage[7][27] , \Storage[7][26] , \Storage[7][25] ,
         \Storage[7][24] , \Storage[7][23] , \Storage[7][22] ,
         \Storage[7][21] , \Storage[7][20] , \Storage[7][19] ,
         \Storage[7][18] , \Storage[7][17] , \Storage[7][16] ,
         \Storage[7][15] , \Storage[7][14] , \Storage[7][13] ,
         \Storage[7][12] , \Storage[7][11] , \Storage[7][10] , \Storage[7][9] ,
         \Storage[7][8] , \Storage[7][7] , \Storage[7][6] , \Storage[7][5] ,
         \Storage[7][4] , \Storage[7][3] , \Storage[7][2] , \Storage[7][1] ,
         \Storage[7][0] , \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N87, N99, N161, N194, N227, N260, N293,
         N326, N359, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n223) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n224) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n227) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n230) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n233) );
  XOR4D1 U21 ( .A1(n218), .A2(N74), .A3(n217), .A4(N77), .Z(n219) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n217) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n211) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n212) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n215) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n221) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(N194), .CP(n174), .CDN(
        n194), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n163), .CP(n185), .CDN(
        n194), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n163), .CP(n174), .CDN(
        n193), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n163), .CP(n179), .CDN(
        n193), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n163), .CP(n183), .CDN(
        n193), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n163), .CP(n185), .CDN(
        n193), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n163), .CP(n177), .CDN(
        n193), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n163), .CP(n180), .CDN(
        n193), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n163), .CP(n181), .CDN(
        n193), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n163), .CP(n176), .CDN(
        n193), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n163), .CP(n178), .CDN(n192), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n163), .CP(n173), .CDN(n192), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n163), .CP(ClockW), .CDN(
        n192), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n163), .CP(n184), .CDN(n192), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n163), .CP(n183), .CDN(n192), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n163), .CP(n182), .CDN(n192), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n163), .CP(n185), .CDN(n192), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n161), .CP(n173), .CDN(n192), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(N194), .CP(n173), .CDN(n192), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(N194), .CP(n173), .CDN(n192), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n169), .CP(n179), .CDN(
        n207), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(N99), .CP(n179), .CDN(n206), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n169), .CP(n180), .CDN(
        n202), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n169), .CP(n180), .CDN(
        n202), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n169), .CP(n180), .CDN(
        n207), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n169), .CP(n180), .CDN(
        n201), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n169), .CP(n180), .CDN(
        n200), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n171), .CP(n180), .CDN(
        n200), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n171), .CP(n181), .CDN(
        n202), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n171), .CP(n181), .CDN(
        n200), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n171), .CP(n181), .CDN(n201), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n171), .CP(n181), .CDN(n201), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n171), .CP(n181), .CDN(n202), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n171), .CP(n181), .CDN(n204), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n171), .CP(n181), .CDN(n201), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n171), .CP(n181), .CDN(n200), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n171), .CP(n181), .CDN(n205), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n169), .CP(n176), .CDN(n202), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n169), .CP(n182), .CDN(n204), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n169), .CP(n179), .CDN(n201), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n145), .CP(n182), .CDN(
        n192), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n147), .CP(n173), .CDN(
        n203), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n147), .CP(n173), .CDN(
        n205), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n147), .CP(n178), .CDN(
        n207), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n147), .CP(n175), .CDN(
        n207), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n147), .CP(ClockW), .CDN(
        n207), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n147), .CP(n176), .CDN(
        n207), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n147), .CP(n178), .CDN(
        n207), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n145), .CP(n175), .CDN(
        n207), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n145), .CP(n185), .CDN(
        n207), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n145), .CP(n175), .CDN(n198), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n145), .CP(n177), .CDN(n198), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n145), .CP(n176), .CDN(n198), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n147), .CP(n174), .CDN(n198), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n147), .CP(n185), .CDN(n198), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n147), .CP(n183), .CDN(n198), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n147), .CP(n184), .CDN(n198), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(N326), .CP(n185), .CDN(n198), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n145), .CP(n182), .CDN(n198), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n145), .CP(n173), .CDN(n198), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(N293), .CP(n182), .CDN(
        n205), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n151), .CP(n174), .CDN(
        n204), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n151), .CP(n183), .CDN(
        n199), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n151), .CP(n185), .CDN(
        n206), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n151), .CP(n183), .CDN(
        n204), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n151), .CP(n178), .CDN(
        n203), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n151), .CP(ClockW), .CDN(
        n205), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n151), .CP(n173), .CDN(
        n206), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n151), .CP(n183), .CDN(
        n203), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n151), .CP(n181), .CDN(
        n195), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n151), .CP(n184), .CDN(n205), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n151), .CP(n181), .CDN(n199), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n151), .CP(n174), .CDN(n204), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n151), .CP(n177), .CDN(n203), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n151), .CP(n178), .CDN(n206), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n151), .CP(n179), .CDN(n206), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n151), .CP(n180), .CDN(n199), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n149), .CP(n185), .CDN(n206), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(N293), .CP(n181), .CDN(n193), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(N293), .CP(n174), .CDN(n199), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(N260), .CP(n183), .CDN(
        n193), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n155), .CP(ClockW), .CDN(
        n195), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n155), .CP(n184), .CDN(
        n197), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n155), .CP(n173), .CDN(
        n199), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n155), .CP(ClockW), .CDN(
        n199), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n155), .CP(n185), .CDN(
        n197), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n155), .CP(n177), .CDN(
        n203), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n155), .CP(n182), .CDN(
        n205), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n155), .CP(ClockW), .CDN(
        n199), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n155), .CP(n177), .CDN(
        n193), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n155), .CP(n174), .CDN(n207), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n155), .CP(n183), .CDN(n207), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n155), .CP(n176), .CDN(n196), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n155), .CP(n174), .CDN(n196), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n155), .CP(n173), .CDN(n204), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n155), .CP(n185), .CDN(n203), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n155), .CP(n184), .CDN(n205), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n153), .CP(n182), .CDN(n205), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(N260), .CP(n184), .CDN(n193), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(N260), .CP(n180), .CDN(n204), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(N227), .CP(n182), .CDN(
        n197), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n159), .CP(n184), .CDN(
        n197), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n159), .CP(n182), .CDN(
        n196), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n159), .CP(n181), .CDN(
        n196), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n159), .CP(n183), .CDN(
        n196), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n159), .CP(n182), .CDN(
        n196), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n159), .CP(n176), .CDN(
        n196), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n159), .CP(n180), .CDN(
        n196), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n159), .CP(n185), .CDN(
        n196), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n159), .CP(n177), .CDN(
        n196), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n159), .CP(n174), .CDN(n195), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n159), .CP(ClockW), .CDN(
        n195), .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n159), .CP(n174), .CDN(n195), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n159), .CP(n183), .CDN(n195), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n159), .CP(n184), .CDN(n195), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n159), .CP(n182), .CDN(n195), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n159), .CP(n181), .CDN(n195), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n157), .CP(n176), .CDN(n195), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n157), .CP(n179), .CDN(n195), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n157), .CP(n181), .CDN(n195), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n165), .CP(n184), .CDN(
        n205), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n167), .CP(n174), .CDN(
        n202), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n167), .CP(n174), .CDN(
        n202), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n167), .CP(n174), .CDN(
        n204), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n167), .CP(n179), .CDN(
        n202), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n167), .CP(n177), .CDN(
        n202), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n167), .CP(n177), .CDN(
        n205), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n167), .CP(n177), .CDN(
        n202), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n167), .CP(n177), .CDN(
        n203), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n167), .CP(n177), .CDN(
        n206), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n167), .CP(n177), .CDN(n201), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n167), .CP(n177), .CDN(n200), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n167), .CP(n177), .CDN(n197), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n167), .CP(n177), .CDN(n203), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n167), .CP(n178), .CDN(n200), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n167), .CP(n178), .CDN(n202), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n167), .CP(n178), .CDN(n201), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n165), .CP(n178), .CDN(n202), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n165), .CP(n178), .CDN(n200), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n165), .CP(n178), .CDN(n206), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(N359), .CP(n176), .CDN(
        n196), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n143), .CP(n176), .CDN(
        n195), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n143), .CP(n176), .CDN(
        n198), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n143), .CP(n176), .CDN(
        n205), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n143), .CP(n176), .CDN(
        n203), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n143), .CP(n184), .CDN(
        n192), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n143), .CP(ClockW), .CDN(
        n198), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n143), .CP(ClockW), .CDN(
        n204), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n143), .CP(n175), .CDN(
        n197), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n143), .CP(n179), .CDN(
        n197), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n143), .CP(n180), .CDN(n192), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n143), .CP(n178), .CDN(n192), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n143), .CP(n176), .CDN(n193), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n143), .CP(n184), .CDN(n204), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n143), .CP(ClockW), .CDN(
        n203), .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n143), .CP(n175), .CDN(n198), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n143), .CP(n178), .CDN(n207), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n141), .CP(n173), .CDN(n195), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(N359), .CP(n184), .CDN(n203), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(N359), .CP(n182), .CDN(n192), 
        .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n2), .CP(n186), .CDN(n202), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N87), .E(N194), .CP(n183), .CDN(n195), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(N194), .CP(ClockW), .CDN(
        n194), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(N194), .CP(n174), .CDN(
        n194), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(N194), .CP(n184), .CDN(
        n194), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n161), .CP(n183), .CDN(
        n194), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n161), .CP(n182), .CDN(
        n194), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n161), .CP(n185), .CDN(
        n194), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n161), .CP(n177), .CDN(
        n194), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n161), .CP(n183), .CDN(
        n194), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n163), .CP(n184), .CDN(
        n194), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n163), .CP(n182), .CDN(
        n193), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n163), .CP(n174), .CDN(
        n193), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n163), .CP(n178), .CDN(
        n193), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N87), .E(n169), .CP(n178), .CDN(n200), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n169), .CP(n178), .CDN(
        n193), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n169), .CP(n178), .CDN(
        n197), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(N99), .CP(n179), .CDN(n194), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(N99), .CP(n179), .CDN(n203), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n169), .CP(n179), .CDN(
        n203), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N99), .CP(n179), .CDN(n205), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n169), .CP(n179), .CDN(
        n196), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n169), .CP(n179), .CDN(
        n205), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n169), .CP(n179), .CDN(
        n207), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(N99), .CP(n180), .CDN(n207), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(N99), .CP(n180), .CDN(n201), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(N99), .CP(n180), .CDN(n200), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N87), .E(n145), .CP(n183), .CDN(n195), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(N326), .CP(n179), .CDN(
        n193), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(N326), .CP(n185), .CDN(
        n198), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(N326), .CP(n184), .CDN(
        n204), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(N326), .CP(n183), .CDN(
        n197), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(N326), .CP(n182), .CDN(
        n193), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(N326), .CP(n185), .CDN(
        n204), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n145), .CP(n180), .CDN(
        n197), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n145), .CP(n177), .CDN(
        n198), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n147), .CP(n177), .CDN(
        n194), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n147), .CP(n179), .CDN(
        n207), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n147), .CP(n180), .CDN(
        n207), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n147), .CP(n178), .CDN(
        n207), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N87), .E(N293), .CP(n180), .CDN(n198), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(N293), .CP(n176), .CDN(
        n204), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(N293), .CP(n181), .CDN(
        n196), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(N293), .CP(n181), .CDN(
        n206), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n149), .CP(n179), .CDN(
        n206), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n149), .CP(n180), .CDN(
        n204), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n149), .CP(n182), .CDN(
        n195), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n149), .CP(n177), .CDN(
        n205), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n149), .CP(n178), .CDN(
        n206), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n151), .CP(n185), .CDN(
        n206), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n151), .CP(n183), .CDN(
        n205), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n151), .CP(n182), .CDN(
        n196), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n151), .CP(n174), .CDN(
        n204), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N87), .E(N260), .CP(n173), .CDN(n206), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(N260), .CP(n185), .CDN(
        n204), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(N260), .CP(n176), .CDN(
        n203), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(N260), .CP(n179), .CDN(
        n205), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n153), .CP(n175), .CDN(
        n204), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n153), .CP(n176), .CDN(
        n206), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n153), .CP(n175), .CDN(
        n199), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n153), .CP(n178), .CDN(
        n203), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n153), .CP(ClockW), .CDN(
        n206), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n155), .CP(n173), .CDN(
        n199), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n155), .CP(n179), .CDN(
        n192), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n155), .CP(n173), .CDN(
        n205), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n155), .CP(n184), .CDN(
        n203), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N87), .E(N227), .CP(n175), .CDN(n203), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(N227), .CP(n177), .CDN(
        n197), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(N227), .CP(n180), .CDN(
        n197), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(N227), .CP(n181), .CDN(
        n197), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(N227), .CP(n173), .CDN(
        n197), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(N227), .CP(n184), .CDN(
        n197), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n157), .CP(ClockW), .CDN(
        n197), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n157), .CP(n174), .CDN(
        n197), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n157), .CP(n184), .CDN(
        n197), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n159), .CP(n183), .CDN(
        n197), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n159), .CP(n173), .CDN(
        n196), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n159), .CP(n174), .CDN(
        n196), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n159), .CP(n175), .CDN(
        n196), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N87), .E(n165), .CP(n185), .CDN(n192), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(N161), .CP(n181), .CDN(
        n196), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(N161), .CP(ClockW), .CDN(
        n202), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(N161), .CP(ClockW), .CDN(
        n206), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(N161), .CP(n180), .CDN(
        n192), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(N161), .CP(n173), .CDN(
        n202), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(N161), .CP(ClockW), .CDN(
        n202), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(N161), .CP(n174), .CDN(
        n195), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n165), .CP(n175), .CDN(
        n202), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n167), .CP(n175), .CDN(
        n205), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n167), .CP(n185), .CDN(
        n202), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n167), .CP(n182), .CDN(
        n201), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n167), .CP(n183), .CDN(
        n207), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N87), .E(N359), .CP(n175), .CDN(n199), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(N359), .CP(n175), .CDN(
        n198), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(N359), .CP(n175), .CDN(
        n196), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(N359), .CP(n175), .CDN(
        n195), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n141), .CP(n175), .CDN(
        n197), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n141), .CP(n175), .CDN(
        n203), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n141), .CP(n175), .CDN(
        n198), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n141), .CP(n175), .CDN(
        n198), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n141), .CP(n175), .CDN(
        n192), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n143), .CP(n176), .CDN(
        n195), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n143), .CP(n176), .CDN(
        n198), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n143), .CP(n176), .CDN(
        n196), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n143), .CP(n176), .CDN(
        n194), .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N53), .E(n188), .CP(n187), .CDN(n202), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N54), .E(n188), .CP(n187), .CDN(n201), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N55), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N56), .E(n188), .CP(n187), .CDN(n201), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N57), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N58), .E(n188), .CP(n187), .CDN(n201), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N59), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N60), .E(n188), .CP(n187), .CDN(n201), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N61), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N62), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N63), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N64), .E(n188), .CP(n186), .CDN(n201), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N65), .E(n188), .CP(n186), .CDN(n200), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N66), .E(n188), .CP(n186), .CDN(n200), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N67), .E(n188), .CP(n186), .CDN(n200), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N68), .E(n188), .CP(n186), .CDN(n200), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N69), .E(n188), .CP(n186), .CDN(n200), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N70), .E(Read), .CP(n186), .CDN(n200), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N71), .E(Read), .CP(n187), .CDN(n200), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N72), .E(Read), .CP(n187), .CDN(n200), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N73), .E(Read), .CP(n187), .CDN(n200), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N74), .E(Read), .CP(n187), .CDN(n200), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N75), .E(Read), .CP(n187), .CDN(n200), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N76), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N77), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N78), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N79), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N80), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N81), .E(Read), .CP(n186), .CDN(n199), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N82), .E(Read), .CP(n186), .CDN(n199), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N83), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N84), .E(Read), .CP(n187), .CDN(n199), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N85), .E(Read), .CP(n186), .CDN(n199), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKBD0 U3 ( .CLK(N49), .C(n191) );
  BUFFD0 U4 ( .I(n190), .Z(n136) );
  CKBD0 U5 ( .CLK(N48), .C(n190) );
  INVD0 U6 ( .I(N99), .ZN(n170) );
  CKND2D0 U7 ( .A1(ClkR), .A2(ChipEna), .ZN(n1) );
  CKNXD0 U8 ( .I(n142), .ZN(n141) );
  INVD0 U9 ( .I(N161), .ZN(n166) );
  CKNXD0 U10 ( .I(n166), .ZN(n165) );
  CKNXD0 U11 ( .I(n154), .ZN(n153) );
  CKNXD0 U12 ( .I(n150), .ZN(n149) );
  CKNXD0 U18 ( .I(n158), .ZN(n157) );
  INVD0 U19 ( .I(N326), .ZN(n146) );
  CKNXD0 U20 ( .I(n146), .ZN(n145) );
  CKNXD0 U23 ( .I(n162), .ZN(n161) );
  CKAN2D0 U24 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U25 ( .I(N50), .ZN(n130) );
  BUFFD1 U26 ( .I(n205), .Z(n192) );
  BUFFD1 U31 ( .I(n205), .Z(n193) );
  BUFFD1 U32 ( .I(n204), .Z(n194) );
  BUFFD1 U33 ( .I(n204), .Z(n195) );
  BUFFD1 U34 ( .I(n203), .Z(n196) );
  BUFFD1 U35 ( .I(n203), .Z(n197) );
  BUFFD1 U36 ( .I(n193), .Z(n198) );
  BUFFD1 U37 ( .I(n194), .Z(n199) );
  BUFFD1 U38 ( .I(n204), .Z(n200) );
  BUFFD1 U39 ( .I(n202), .Z(n201) );
  BUFFD1 U40 ( .I(n206), .Z(n205) );
  BUFFD1 U41 ( .I(n206), .Z(n204) );
  BUFFD1 U42 ( .I(n206), .Z(n203) );
  BUFFD1 U43 ( .I(n207), .Z(n202) );
  BUFFD1 U44 ( .I(n207), .Z(n206) );
  INVD1 U45 ( .I(Reset), .ZN(n207) );
  BUFFD1 U46 ( .I(n185), .Z(n176) );
  BUFFD1 U47 ( .I(n185), .Z(n175) );
  INVD1 U48 ( .I(n164), .ZN(n163) );
  INVD1 U49 ( .I(n160), .ZN(n159) );
  INVD1 U50 ( .I(n148), .ZN(n147) );
  INVD1 U51 ( .I(n144), .ZN(n143) );
  BUFFD1 U52 ( .I(n182), .Z(n181) );
  BUFFD1 U53 ( .I(n183), .Z(n180) );
  BUFFD1 U54 ( .I(n183), .Z(n179) );
  BUFFD1 U55 ( .I(n184), .Z(n178) );
  BUFFD1 U56 ( .I(n184), .Z(n177) );
  BUFFD1 U57 ( .I(n182), .Z(n185) );
  BUFFD1 U58 ( .I(n136), .Z(n140) );
  BUFFD1 U59 ( .I(n136), .Z(n138) );
  BUFFD1 U60 ( .I(n136), .Z(n139) );
  BUFFD1 U61 ( .I(n135), .Z(n133) );
  INVD1 U62 ( .I(n157), .ZN(n160) );
  INVD1 U63 ( .I(n145), .ZN(n148) );
  INVD1 U64 ( .I(n141), .ZN(n144) );
  INVD1 U65 ( .I(n161), .ZN(n164) );
  INVD1 U66 ( .I(n172), .ZN(n171) );
  INVD1 U67 ( .I(n168), .ZN(n167) );
  INVD1 U68 ( .I(n156), .ZN(n155) );
  INVD1 U69 ( .I(n152), .ZN(n151) );
  BUFFD1 U70 ( .I(n173), .Z(n182) );
  BUFFD1 U71 ( .I(n173), .Z(n183) );
  BUFFD1 U72 ( .I(n173), .Z(n184) );
  INVD1 U73 ( .I(n1), .ZN(n187) );
  INVD1 U74 ( .I(n1), .ZN(n186) );
  XOR3D1 U75 ( .A1(N69), .A2(N68), .A3(n216), .Z(n218) );
  XOR3D1 U76 ( .A1(N67), .A2(n215), .A3(n214), .Z(n216) );
  XOR3D1 U77 ( .A1(N62), .A2(N61), .A3(n213), .Z(n214) );
  XOR3D1 U78 ( .A1(n212), .A2(N60), .A3(n211), .Z(n213) );
  XOR3D1 U79 ( .A1(N81), .A2(N76), .A3(n222), .Z(N85) );
  XOR3D1 U80 ( .A1(N75), .A2(n221), .A3(n220), .Z(n222) );
  XOR3D1 U81 ( .A1(N79), .A2(N78), .A3(n219), .Z(n220) );
  BUFFD1 U82 ( .I(n190), .Z(n137) );
  BUFFD1 U83 ( .I(n191), .Z(n135) );
  BUFFD1 U84 ( .I(n191), .Z(n134) );
  INVD1 U85 ( .I(n130), .ZN(n131) );
  INVD1 U86 ( .I(n130), .ZN(n132) );
  INVD1 U87 ( .I(AddrW[0]), .ZN(n208) );
  INVD1 U88 ( .I(n169), .ZN(n172) );
  INVD1 U89 ( .I(n165), .ZN(n168) );
  INVD1 U90 ( .I(n153), .ZN(n156) );
  INVD1 U91 ( .I(n149), .ZN(n152) );
  INVD1 U92 ( .I(N194), .ZN(n162) );
  NR3D0 U93 ( .A1(n210), .A2(AddrW[0]), .A3(n235), .ZN(N194) );
  INVD1 U94 ( .I(N227), .ZN(n158) );
  NR3D0 U95 ( .A1(n210), .A2(n235), .A3(n208), .ZN(N227) );
  NR3D0 U96 ( .A1(n210), .A2(AddrW[0]), .A3(n209), .ZN(N326) );
  INVD1 U97 ( .I(N359), .ZN(n142) );
  NR3D0 U98 ( .A1(n210), .A2(n209), .A3(n208), .ZN(N359) );
  INVD1 U99 ( .I(n189), .ZN(n188) );
  BUFFD1 U100 ( .I(n174), .Z(n173) );
  BUFFD1 U101 ( .I(ClockW), .Z(n174) );
  XOR3D1 U102 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n234), .Z(N87) );
  XOR3D1 U103 ( .A1(DataI[0]), .A2(n233), .A3(n232), .Z(n234) );
  XOR3D1 U104 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n231), .Z(n232) );
  XOR3D1 U105 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n225), .Z(n226) );
  XOR3D1 U106 ( .A1(n224), .A2(DataI[17]), .A3(n223), .Z(n225) );
  XOR3D1 U107 ( .A1(n230), .A2(DataI[3]), .A3(n229), .Z(n231) );
  XOR3D1 U108 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n228), .Z(n229) );
  XOR3D1 U109 ( .A1(n227), .A2(DataI[10]), .A3(n226), .Z(n228) );
  MUX4ND0 U110 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n140), .S1(n134), .ZN(
        n111) );
  MUX4ND0 U111 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n136), .S1(n134), .ZN(
        n114) );
  MUX4ND0 U112 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n140), .S1(n134), .ZN(
        n108) );
  MUX4ND0 U113 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n136), .S1(n134), .ZN(
        n117) );
  MUX4ND0 U114 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(N48), .S1(n191), .ZN(n8)
         );
  MUX4ND0 U115 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(N48), .S1(n191), .ZN(n11)
         );
  MUX4ND0 U116 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(N48), .S1(N49), .ZN(n26)
         );
  MUX4ND0 U117 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n139), .S1(n134), .ZN(
        n41) );
  MUX4ND0 U118 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n140), .S1(n135), .ZN(
        n44) );
  MUX4ND0 U119 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n140), .S1(n134), .ZN(
        n62) );
  MUX4ND0 U120 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n139), .S1(n133), .ZN(
        n65) );
  MUX4ND0 U121 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n139), .S1(n134), .ZN(
        n123) );
  MUX4ND0 U122 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n139), .S1(n134), .ZN(
        n126) );
  MUX4ND0 U123 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n139), .S1(N49), .ZN(n23)
         );
  MUX4ND0 U124 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n140), .S1(N49), .ZN(n29)
         );
  MUX4ND0 U125 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n139), .S1(N49), .ZN(n53) );
  MUX4ND0 U126 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n140), .S1(n133), .ZN(
        n102) );
  MUX4ND0 U127 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n190), .S1(n134), .ZN(
        n105) );
  MUX4ND0 U128 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(N48), .S1(n191), .ZN(n5)
         );
  MUX4ND0 U129 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n140), .S1(n191), .ZN(n17)
         );
  MUX4ND0 U130 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n139), .S1(N49), .ZN(n35) );
  MUX4ND0 U131 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n140), .S1(N49), .ZN(n38) );
  MUX4ND0 U132 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n139), .S1(n191), .ZN(
        n47) );
  MUX4ND0 U133 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n140), .S1(n191), .ZN(
        n59) );
  MUX4ND0 U134 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n140), .S1(n191), .ZN(
        n96) );
  MUX4ND0 U135 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n136), .S1(n133), .ZN(
        n120) );
  MUX4ND0 U136 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(N48), .S1(n191), .ZN(n14)
         );
  MUX4ND0 U137 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n140), .S1(n191), .ZN(n20)
         );
  MUX4ND0 U138 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n139), .S1(N49), .ZN(n32)
         );
  MUX4ND0 U139 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n139), .S1(N49), .ZN(n50) );
  MUX4ND0 U140 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n140), .S1(n134), .ZN(
        n56) );
  MUX4ND0 U141 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n139), .S1(n191), .ZN(
        n99) );
  MUX4ND0 U142 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n136), .S1(n134), .ZN(
        n129) );
  INVD1 U143 ( .I(N260), .ZN(n154) );
  NR3D0 U144 ( .A1(n209), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N260) );
  INVD1 U145 ( .I(n170), .ZN(n169) );
  NR3D0 U146 ( .A1(n235), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N99) );
  INVD1 U147 ( .I(N293), .ZN(n150) );
  NR3D0 U148 ( .A1(n208), .A2(AddrW[1]), .A3(n209), .ZN(N293) );
  INVD1 U149 ( .I(AddrW[1]), .ZN(n210) );
  ND2D1 U150 ( .A1(AddrW[2]), .A2(Write), .ZN(n209) );
  IND2D1 U151 ( .A1(AddrW[2]), .B1(Write), .ZN(n235) );
  NR3D0 U152 ( .A1(n208), .A2(AddrW[1]), .A3(n235), .ZN(N161) );
  INVD1 U153 ( .I(Read), .ZN(n189) );
  OR2D1 U154 ( .A1(Read), .A2(Dreadyr), .Z(n2) );
  CKAN2D0 U155 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX3ND0 U156 ( .I0(n3), .I1(n4), .I2(n5), .S0(n133), .S1(n131), .ZN(N84) );
  MUX3ND0 U157 ( .I0(n6), .I1(n7), .I2(n8), .S0(n133), .S1(n131), .ZN(N83) );
  MUX3ND0 U158 ( .I0(n9), .I1(n10), .I2(n11), .S0(n133), .S1(n131), .ZN(N82)
         );
  MUX3ND0 U159 ( .I0(n12), .I1(n13), .I2(n14), .S0(n133), .S1(n131), .ZN(N81)
         );
  MUX3ND0 U160 ( .I0(n15), .I1(n16), .I2(n17), .S0(n133), .S1(n131), .ZN(N80)
         );
  MUX3ND0 U161 ( .I0(n18), .I1(n19), .I2(n20), .S0(n133), .S1(n131), .ZN(N79)
         );
  MUX3ND0 U162 ( .I0(n21), .I1(n22), .I2(n23), .S0(n133), .S1(n131), .ZN(N78)
         );
  MUX3ND0 U163 ( .I0(n24), .I1(n25), .I2(n26), .S0(n133), .S1(n131), .ZN(N77)
         );
  MUX3ND0 U164 ( .I0(n27), .I1(n28), .I2(n29), .S0(n133), .S1(n131), .ZN(N76)
         );
  MUX3ND0 U165 ( .I0(n30), .I1(n31), .I2(n32), .S0(n133), .S1(n131), .ZN(N75)
         );
  MUX3ND0 U166 ( .I0(n33), .I1(n34), .I2(n35), .S0(n133), .S1(n131), .ZN(N74)
         );
  MUX3ND0 U167 ( .I0(n36), .I1(n37), .I2(n38), .S0(n133), .S1(n131), .ZN(N73)
         );
  MUX3ND0 U168 ( .I0(n39), .I1(n40), .I2(n41), .S0(n133), .S1(n131), .ZN(N72)
         );
  MUX3ND0 U169 ( .I0(n42), .I1(n43), .I2(n44), .S0(n135), .S1(n131), .ZN(N71)
         );
  MUX3ND0 U170 ( .I0(n45), .I1(n46), .I2(n47), .S0(n135), .S1(n131), .ZN(N70)
         );
  MUX3ND0 U171 ( .I0(n48), .I1(n49), .I2(n50), .S0(n135), .S1(n131), .ZN(N69)
         );
  MUX3ND0 U172 ( .I0(n51), .I1(n52), .I2(n53), .S0(n135), .S1(n131), .ZN(N68)
         );
  MUX3ND0 U173 ( .I0(n54), .I1(n55), .I2(n56), .S0(n135), .S1(n131), .ZN(N67)
         );
  MUX3ND0 U174 ( .I0(n57), .I1(n58), .I2(n59), .S0(n135), .S1(n131), .ZN(N66)
         );
  MUX3ND0 U175 ( .I0(n60), .I1(n61), .I2(n62), .S0(n135), .S1(n131), .ZN(N65)
         );
  MUX3ND0 U176 ( .I0(n63), .I1(n64), .I2(n65), .S0(n134), .S1(n132), .ZN(N64)
         );
  MUX3ND0 U177 ( .I0(n94), .I1(n95), .I2(n96), .S0(n135), .S1(n132), .ZN(N63)
         );
  MUX3ND0 U178 ( .I0(n97), .I1(n98), .I2(n99), .S0(n135), .S1(n132), .ZN(N62)
         );
  MUX3ND0 U179 ( .I0(n100), .I1(n101), .I2(n102), .S0(n134), .S1(n132), .ZN(
        N61) );
  MUX3ND0 U180 ( .I0(n103), .I1(n104), .I2(n105), .S0(n135), .S1(n132), .ZN(
        N60) );
  MUX3ND0 U181 ( .I0(n106), .I1(n107), .I2(n108), .S0(n135), .S1(n132), .ZN(
        N59) );
  MUX3ND0 U182 ( .I0(n109), .I1(n110), .I2(n111), .S0(n135), .S1(n132), .ZN(
        N58) );
  MUX3ND0 U183 ( .I0(n112), .I1(n113), .I2(n114), .S0(N49), .S1(n132), .ZN(N57) );
  MUX3ND0 U184 ( .I0(n115), .I1(n116), .I2(n117), .S0(N49), .S1(n132), .ZN(N56) );
  MUX3ND0 U185 ( .I0(n118), .I1(n119), .I2(n120), .S0(n191), .S1(n132), .ZN(
        N55) );
  MUX3ND0 U186 ( .I0(n121), .I1(n122), .I2(n123), .S0(N49), .S1(n132), .ZN(N54) );
  MUX3ND0 U187 ( .I0(n124), .I1(n125), .I2(n126), .S0(N49), .S1(n132), .ZN(N53) );
  MUX3ND0 U188 ( .I0(n127), .I1(n128), .I2(n129), .S0(n191), .S1(n132), .ZN(
        N52) );
  MUX2ND0 U189 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n138), .ZN(n4)
         );
  MUX2ND0 U190 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n138), .ZN(n3)
         );
  MUX2ND0 U191 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(N48), .ZN(n7)
         );
  MUX2ND0 U192 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n138), .ZN(n6)
         );
  MUX2ND0 U193 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n139), .ZN(n10) );
  MUX2ND0 U194 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n138), .ZN(n9)
         );
  MUX2ND0 U195 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n139), .ZN(n13) );
  MUX2ND0 U196 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n139), .ZN(n12) );
  MUX2ND0 U197 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n138), .ZN(n16) );
  MUX2ND0 U198 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n139), .ZN(n15) );
  MUX2ND0 U199 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n138), .ZN(n19) );
  MUX2ND0 U200 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n138), .ZN(n18) );
  MUX2ND0 U201 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n139), .ZN(n22) );
  MUX2ND0 U202 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n138), .ZN(n21) );
  MUX2ND0 U203 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n138), .ZN(n25) );
  MUX2ND0 U204 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n138), .ZN(n24) );
  MUX2ND0 U205 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n138), .ZN(n28) );
  MUX2ND0 U206 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n138), .ZN(n27) );
  MUX2ND0 U207 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n138), .ZN(n31) );
  MUX2ND0 U208 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n138), .ZN(n30) );
  MUX2ND0 U209 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n138), .ZN(
        n34) );
  MUX2ND0 U210 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n138), .ZN(
        n33) );
  MUX2ND0 U211 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n138), .ZN(
        n37) );
  MUX2ND0 U212 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n138), .ZN(
        n36) );
  MUX2ND0 U213 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n138), .ZN(
        n40) );
  MUX2ND0 U214 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n137), .ZN(
        n39) );
  MUX2ND0 U215 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(n137), .ZN(
        n43) );
  MUX2ND0 U216 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n140), .ZN(
        n42) );
  MUX2ND0 U217 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(N48), .ZN(
        n46) );
  MUX2ND0 U218 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n140), .ZN(
        n45) );
  MUX2ND0 U219 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(N48), .ZN(
        n49) );
  MUX2ND0 U220 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(N48), .ZN(
        n48) );
  MUX2ND0 U221 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(N48), .ZN(
        n52) );
  MUX2ND0 U222 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(N48), .ZN(
        n51) );
  MUX2ND0 U223 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n137), .ZN(
        n55) );
  MUX2ND0 U224 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n137), .ZN(
        n54) );
  MUX2ND0 U225 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n137), .ZN(
        n58) );
  MUX2ND0 U226 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n137), .ZN(
        n57) );
  MUX2ND0 U227 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(n137), .ZN(
        n61) );
  MUX2ND0 U228 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n137), .ZN(
        n60) );
  MUX2ND0 U229 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n137), .ZN(
        n64) );
  MUX2ND0 U230 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(n137), .ZN(
        n63) );
  MUX2ND0 U231 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(n137), .ZN(
        n95) );
  MUX2ND0 U232 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(n190), .ZN(
        n94) );
  MUX2ND0 U233 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(n190), .ZN(
        n98) );
  MUX2ND0 U234 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(n190), .ZN(
        n97) );
  MUX2ND0 U235 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(n190), .ZN(
        n101) );
  MUX2ND0 U236 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(n190), .ZN(
        n100) );
  MUX2ND0 U237 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n190), .ZN(
        n104) );
  MUX2ND0 U238 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n190), .ZN(
        n103) );
  MUX2ND0 U239 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n137), .ZN(
        n107) );
  MUX2ND0 U240 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n137), .ZN(
        n106) );
  MUX2ND0 U241 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n137), .ZN(
        n110) );
  MUX2ND0 U242 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n137), .ZN(
        n109) );
  MUX2ND0 U243 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n137), .ZN(
        n113) );
  MUX2ND0 U244 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n137), .ZN(
        n112) );
  MUX2ND0 U245 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n137), .ZN(
        n116) );
  MUX2ND0 U246 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n137), .ZN(
        n115) );
  MUX2ND0 U247 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n139), .ZN(
        n119) );
  MUX2ND0 U248 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n140), .ZN(
        n118) );
  MUX2ND0 U249 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(N48), .ZN(
        n122) );
  MUX2ND0 U250 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n139), .ZN(
        n121) );
  MUX2ND0 U251 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(N48), .ZN(
        n125) );
  MUX2ND0 U252 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n139), .ZN(
        n124) );
  MUX2ND0 U253 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n138), .ZN(
        n128) );
  MUX2ND0 U254 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n137), .ZN(
        n127) );
endmodule


module PLLTop_1 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_1 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_1 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_1 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_2 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_2 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_2 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_2 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_3 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_3 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_3 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_3 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N47, N48, N49, N50, N51, N67, N68, N69,
         N70, N71, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n88, n89,
         n93, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n177,
         n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n33), .CPN(StateClock), .Q(FullFIFO) );
  DFND1 EmptyFIFOr_reg ( .D(n93), .CPN(StateClock), .Q(EmptyFIFO), .QN(n136)
         );
  MOAI22D1 U6 ( .A1(n20), .A2(n225), .B1(n225), .B2(OldReadAr[1]), .ZN(n88) );
  OA21D1 U11 ( .A1(n13), .A2(n15), .B(n230), .Z(n221) );
  MOAI22D1 U12 ( .A1(n17), .A2(n220), .B1(n220), .B2(OldWriteAr[2]), .ZN(n32)
         );
  MOAI22D1 U13 ( .A1(n16), .A2(n220), .B1(n220), .B2(OldWriteAr[0]), .ZN(n31)
         );
  MOAI22D1 U14 ( .A1(n220), .A2(n219), .B1(n220), .B2(OldWriteAr[1]), .ZN(n30)
         );
  MOAI22D1 U15 ( .A1(n18), .A2(n220), .B1(n220), .B2(OldWriteAr[3]), .ZN(n29)
         );
  IAO21D1 U31 ( .A1(n192), .A2(n191), .B(n210), .ZN(n193) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n189), .B(n190), .Z(n184) );
  MOAI22D1 U88 ( .A1(n19), .A2(n225), .B1(n225), .B2(OldReadAr[0]), .ZN(n23)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n34), .CPN(StateClock), .CDN(n12), .QN(n224)
         );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n89), .CPN(StateClock), .CDN(n12), .QN(n226)
         );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n23), .CPN(StateClock), .CDN(n11), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n29), .CPN(StateClock), .CDN(n11), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n30), .CPN(StateClock), .CDN(n12), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n31), .CPN(StateClock), .CDN(n12), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n32), .CPN(StateClock), .CDN(n12), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n88), .CPN(StateClock), .CDN(n12), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n25), .CPN(StateClock), .CDN(n11), .Q(
        NextState[0]), .QN(n133) );
  DFNCND1 \NextState_reg[1]  ( .D(n26), .CPN(StateClock), .CDN(n11), .Q(
        NextState[1]), .QN(n134) );
  DFNCND1 \NextState_reg[2]  ( .D(n28), .CPN(StateClock), .CDN(n11), .Q(
        NextState[2]), .QN(n135) );
  DFNCND1 WriteCmdr_reg ( .D(n27), .CPN(StateClock), .CDN(n11), .Q(WriteCmd)
         );
  DFNCND1 ReadCmdr_reg ( .D(n24), .CPN(StateClock), .CDN(n11), .Q(ReadCmd) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n11), 
        .QN(n15) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n11), .Q(
        n213), .QN(n13) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n11), 
        .QN(n14) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(N68), .E(N71), .CP(StateClock), .CDN(n12), 
        .Q(WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[3]  ( .D(N51), .E(N50), .CP(StateClock), .CDN(n11), .Q(
        ReadAddr[3]), .QN(n22) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N50), .CP(StateClock), .CDN(n12), .Q(
        ReadAddr[2]), .QN(n21) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N48), .E(N50), .CP(StateClock), .CDN(n12), .Q(
        ReadAddr[1]), .QN(n20) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N47), .E(N50), .CP(StateClock), .CDN(n12), .Q(
        ReadAddr[0]), .QN(n19) );
  EDFCND1 \WriteAr_reg[3]  ( .D(N70), .E(N71), .CP(StateClock), .CDN(n12), .Q(
        WriteAddr[3]), .QN(n18) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N69), .E(N71), .CP(StateClock), .CDN(n11), .Q(
        WriteAddr[2]), .QN(n17) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N67), .E(N71), .CP(StateClock), .CDN(n12), .Q(
        WriteAddr[0]), .QN(n16) );
  CKNXD0 U3 ( .I(Reset), .ZN(n12) );
  CKNXD0 U4 ( .I(Reset), .ZN(n11) );
  ND2D1 U5 ( .A1(n199), .A2(n223), .ZN(n149) );
  INVD1 U7 ( .I(n217), .ZN(n216) );
  INVD1 U8 ( .I(n225), .ZN(n227) );
  MAOI22D0 U9 ( .A1(n196), .A2(n15), .B1(n15), .B2(n194), .ZN(n199) );
  OAI211D1 U10 ( .A1(n230), .A2(n202), .B(n199), .C(n153), .ZN(n217) );
  INR2D1 U16 ( .A1(n194), .B1(n152), .ZN(n153) );
  AOI21D1 U17 ( .A1(n213), .A2(n151), .B(n15), .ZN(n152) );
  INVD1 U18 ( .I(n212), .ZN(n223) );
  ND2D1 U19 ( .A1(WriteReq), .A2(n218), .ZN(n220) );
  ND2D1 U20 ( .A1(ReadReq), .A2(n149), .ZN(n225) );
  ND2D1 U21 ( .A1(n199), .A2(n230), .ZN(n218) );
  OAI21D1 U22 ( .A1(n138), .A2(ReadAddr[2]), .B(n139), .ZN(n154) );
  AOI21D1 U23 ( .A1(n189), .A2(n182), .B(ReadAddr[1]), .ZN(n163) );
  INVD1 U24 ( .I(n162), .ZN(n189) );
  OA211D0 U25 ( .A1(n190), .A2(n189), .B(n188), .C(n187), .Z(n210) );
  INVD1 U26 ( .I(n180), .ZN(n188) );
  NR3D0 U27 ( .A1(n186), .A2(n185), .A3(n184), .ZN(n187) );
  NR3D0 U28 ( .A1(WriteAddr[2]), .A2(n219), .A3(ReadAddr[2]), .ZN(n185) );
  ND2D1 U29 ( .A1(n138), .A2(ReadAddr[2]), .ZN(n139) );
  ND2D1 U30 ( .A1(n161), .A2(n160), .ZN(n180) );
  XNR2D1 U32 ( .A1(ReadAddr[1]), .A2(n219), .ZN(n161) );
  INVD1 U33 ( .I(n177), .ZN(n181) );
  XNR2D1 U35 ( .A1(n142), .A2(WriteAddr[3]), .ZN(n169) );
  INVD1 U36 ( .I(n171), .ZN(n160) );
  ND3D1 U37 ( .A1(n223), .A2(n230), .A3(n209), .ZN(N71) );
  ND2D1 U38 ( .A1(n230), .A2(n150), .ZN(N50) );
  NR3D0 U39 ( .A1(n151), .A2(n144), .A3(n143), .ZN(n145) );
  XNR2D1 U40 ( .A1(ReadAddr[3]), .A2(n224), .ZN(n143) );
  XNR2D1 U41 ( .A1(ReadAddr[2]), .A2(n226), .ZN(n144) );
  XNR2D1 U42 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n164) );
  NR2D1 U43 ( .A1(n154), .A2(n150), .ZN(N49) );
  NR2D1 U44 ( .A1(n137), .A2(n150), .ZN(N48) );
  XNR2D1 U45 ( .A1(ReadAddr[1]), .A2(ReadAddr[0]), .ZN(n137) );
  NR2D1 U46 ( .A1(n156), .A2(n150), .ZN(N51) );
  NR2D1 U47 ( .A1(ReadAddr[0]), .A2(n150), .ZN(N47) );
  INVD1 U48 ( .I(ReadReq), .ZN(n151) );
  INVD1 U49 ( .I(WriteReq), .ZN(n202) );
  INVD1 U50 ( .I(WriteAddr[1]), .ZN(n219) );
  OAI211D1 U51 ( .A1(n219), .A2(ReadAddr[1]), .B(n182), .C(n175), .ZN(n191) );
  AOI22D0 U52 ( .A1(n22), .A2(WriteAddr[3]), .B1(n19), .B2(WriteAddr[0]), .ZN(
        n175) );
  ND2D1 U53 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n140) );
  OAI21D1 U54 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n140), .ZN(n155) );
  AOI21D1 U55 ( .A1(n140), .A2(n17), .B(n142), .ZN(n170) );
  OAI211D1 U56 ( .A1(n20), .A2(WriteAddr[1]), .B(n181), .C(n178), .ZN(n192) );
  AOI22D0 U57 ( .A1(n18), .A2(ReadAddr[3]), .B1(n16), .B2(ReadAddr[0]), .ZN(
        n178) );
  ND2D1 U58 ( .A1(n14), .A2(n213), .ZN(n194) );
  OAI22D0 U59 ( .A1(n227), .A2(n226), .B1(n21), .B2(n225), .ZN(n89) );
  OAI22D0 U60 ( .A1(n227), .A2(n224), .B1(n22), .B2(n225), .ZN(n34) );
  NR3D0 U61 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n212) );
  ND2D1 U62 ( .A1(n21), .A2(WriteAddr[2]), .ZN(n182) );
  OAI22D0 U63 ( .A1(n217), .A2(n135), .B1(n216), .B2(n215), .ZN(n28) );
  AOI21D1 U64 ( .A1(n214), .A2(n213), .B(n212), .ZN(n215) );
  OAI22D0 U65 ( .A1(n14), .A2(n211), .B1(n15), .B2(n210), .ZN(n214) );
  OAI22D0 U66 ( .A1(n217), .A2(n134), .B1(n216), .B2(n198), .ZN(n26) );
  AOI31D0 U67 ( .A1(n197), .A2(n196), .A3(n15), .B(n195), .ZN(n198) );
  IOA21D1 U68 ( .A1(n213), .A2(n211), .B(n179), .ZN(n197) );
  OAI31D0 U69 ( .A1(n194), .A2(n15), .A3(n193), .B(n230), .ZN(n195) );
  OAI22D0 U70 ( .A1(n217), .A2(n133), .B1(n216), .B2(n168), .ZN(n25) );
  AOI22D0 U71 ( .A1(n167), .A2(n213), .B1(n166), .B2(n165), .ZN(n168) );
  AOI211D1 U72 ( .A1(n21), .A2(n162), .B(n228), .C(n180), .ZN(n166) );
  AOI221D0 U73 ( .A1(n177), .A2(n189), .B1(n164), .B2(ReadAddr[1]), .C(n163), 
        .ZN(n165) );
  AOI21D1 U74 ( .A1(n182), .A2(n181), .B(WriteAddr[1]), .ZN(n186) );
  INVD1 U75 ( .I(n14), .ZN(n196) );
  NR2D1 U76 ( .A1(WriteAddr[2]), .A2(n21), .ZN(n177) );
  OAI21D1 U77 ( .A1(n150), .A2(n149), .B(n148), .ZN(n24) );
  ND4D1 U78 ( .A1(n147), .A2(n149), .A3(n146), .A4(n145), .ZN(n148) );
  XNR2D1 U79 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n147) );
  XNR2D1 U80 ( .A1(ReadAddr[1]), .A2(OldReadAr[1]), .ZN(n146) );
  OAI21D1 U81 ( .A1(n14), .A2(n159), .B(n15), .ZN(n167) );
  NR4D0 U82 ( .A1(n160), .A2(n158), .A3(n173), .A4(n157), .ZN(n159) );
  XNR2D1 U83 ( .A1(WriteAddr[2]), .A2(n154), .ZN(n158) );
  XNR2D1 U84 ( .A1(WriteAddr[3]), .A2(n156), .ZN(n157) );
  OAI21D1 U85 ( .A1(n209), .A2(n218), .B(n208), .ZN(n27) );
  ND4D1 U86 ( .A1(n207), .A2(n218), .A3(n206), .A4(n205), .ZN(n208) );
  XNR2D1 U87 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n207) );
  XNR2D1 U89 ( .A1(WriteAddr[2]), .A2(OldWriteAr[2]), .ZN(n206) );
  ND4D1 U90 ( .A1(n174), .A2(n173), .A3(n172), .A4(n171), .ZN(n211) );
  XNR2D1 U91 ( .A1(n169), .A2(n22), .ZN(n174) );
  XNR2D1 U92 ( .A1(ReadAddr[2]), .A2(n170), .ZN(n172) );
  NR2D1 U93 ( .A1(n140), .A2(n17), .ZN(n142) );
  NR2D1 U94 ( .A1(n219), .A2(n17), .ZN(n190) );
  XNR2D1 U95 ( .A1(ReadAddr[3]), .A2(n18), .ZN(n162) );
  XNR2D1 U96 ( .A1(WriteAddr[0]), .A2(n19), .ZN(n171) );
  NR2D1 U97 ( .A1(n19), .A2(n20), .ZN(n138) );
  XNR2D1 U98 ( .A1(n155), .A2(n20), .ZN(n173) );
  XNR2D1 U99 ( .A1(n22), .A2(n139), .ZN(n156) );
  ND2D1 U100 ( .A1(ReadCmd), .A2(n230), .ZN(n150) );
  ND2D1 U101 ( .A1(WriteCmd), .A2(n223), .ZN(n209) );
  OAI32D1 U102 ( .A1(n230), .A2(WriteReq), .A3(Reset), .B1(n229), .B2(n136), 
        .ZN(n93) );
  AOI21D1 U103 ( .A1(n228), .A2(n230), .B(Reset), .ZN(n229) );
  ND3D1 U104 ( .A1(n14), .A2(n15), .A3(n13), .ZN(n230) );
  OAI22D0 U105 ( .A1(n20), .A2(n223), .B1(n155), .B2(n209), .ZN(N68) );
  OAI22D0 U106 ( .A1(n22), .A2(n223), .B1(n169), .B2(n209), .ZN(N70) );
  OAI22D0 U107 ( .A1(n21), .A2(n223), .B1(n141), .B2(n209), .ZN(N69) );
  INVD1 U108 ( .I(n170), .ZN(n141) );
  OAI22D0 U109 ( .A1(n19), .A2(n223), .B1(WriteAddr[0]), .B2(n209), .ZN(N67)
         );
  ND3D1 U110 ( .A1(n15), .A2(n196), .A3(n13), .ZN(n228) );
  NR3D0 U111 ( .A1(n204), .A2(n203), .A3(n202), .ZN(n205) );
  XNR2D1 U112 ( .A1(n18), .A2(OldWriteAr[3]), .ZN(n203) );
  XNR2D1 U113 ( .A1(n219), .A2(OldWriteAr[1]), .ZN(n204) );
  OAI21D1 U114 ( .A1(n191), .A2(n192), .B(n13), .ZN(n179) );
  OAI31D0 U115 ( .A1(n223), .A2(Reset), .A3(ReadReq), .B(n222), .ZN(n33) );
  OAI21D1 U116 ( .A1(n221), .A2(Reset), .B(FullFIFO), .ZN(n222) );
  ND2D1 U117 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid4_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, N133, N166, N199, N232, N265, N298, N331, N364, N397,
         N430, N463, N496, N529, N562, N595, N628, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  OR2D1 U3 ( .A1(Read), .A2(Dreadyr), .Z(n374) );
  XNR4D1 U13 ( .A1(n214), .A2(n213), .A3(n216), .A4(n215), .ZN(n400) );
  XOR4D1 U14 ( .A1(n218), .A2(n217), .A3(n220), .A4(n219), .Z(n401) );
  XOR4D1 U15 ( .A1(n210), .A2(n209), .A3(n212), .A4(n211), .Z(n404) );
  XOR4D1 U16 ( .A1(n203), .A2(n202), .A3(n205), .A4(n204), .Z(n407) );
  XNR4D1 U17 ( .A1(n196), .A2(n195), .A3(n198), .A4(n197), .ZN(n410) );
  XOR4D1 U21 ( .A1(n395), .A2(N71), .A3(n394), .A4(N74), .Z(n396) );
  XNR4D1 U22 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n394) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n388) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n389) );
  XNR4D1 U29 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .ZN(n392) );
  XNR4D1 U30 ( .A1(N79), .A2(N77), .A3(N81), .A4(N80), .ZN(n398) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N84), .E(N595), .CP(n290), .CDN(n350), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n220), .E(N595), .CP(n290), .CDN(n349), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n219), .E(N595), .CP(n290), .CDN(n349), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n218), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n213), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n212), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n211), .E(N595), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n210), .E(n227), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n209), .E(n227), .CP(n292), .CDN(n354), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n208), .E(n225), .CP(n292), .CDN(n319), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n207), .E(N595), .CP(n292), .CDN(n320), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n206), .E(N595), .CP(n292), .CDN(n349), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n205), .E(N595), .CP(n292), .CDN(n320), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n204), .E(N595), .CP(n292), .CDN(n346), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n203), .E(N595), .CP(n292), .CDN(n340), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n202), .E(N595), .CP(n292), .CDN(n350), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n201), .E(n227), .CP(n292), .CDN(n349), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n200), .E(n227), .CP(n293), .CDN(n355), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n199), .E(n227), .CP(n293), .CDN(n353), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n198), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n197), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n196), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n195), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n194), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n193), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n192), .E(n227), .CP(n293), .CDN(n348), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n191), .E(n225), .CP(n294), .CDN(n348), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n190), .E(n225), .CP(n294), .CDN(n348), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n189), .E(n225), .CP(n294), .CDN(n348), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N84), .E(N562), .CP(n294), .CDN(n348), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n220), .E(n231), .CP(n294), .CDN(n324), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n219), .E(n231), .CP(n294), .CDN(n347), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n218), .E(n231), .CP(n294), .CDN(n356), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n213), .E(n231), .CP(n295), .CDN(n358), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n212), .E(n231), .CP(n295), .CDN(n356), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n211), .E(N562), .CP(n295), .CDN(n358), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n210), .E(N562), .CP(n295), .CDN(n356), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n209), .E(n229), .CP(n295), .CDN(n347), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n208), .E(n229), .CP(n295), .CDN(n347), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n207), .E(n229), .CP(n295), .CDN(n347), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n206), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n205), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n204), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n203), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n202), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n201), .E(n231), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n200), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n199), .E(n229), .CP(n296), .CDN(n347), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n198), .E(N562), .CP(n296), .CDN(n346), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n197), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n196), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n195), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n194), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n193), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n192), .E(N562), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n191), .E(n231), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n190), .E(n231), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n189), .E(n231), .CP(n297), .CDN(n346), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N84), .E(N463), .CP(n287), .CDN(n329), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n220), .E(n243), .CP(n287), .CDN(n340), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n219), .E(n243), .CP(n290), .CDN(n340), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n218), .E(n243), .CP(n291), .CDN(n340), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n213), .E(n243), .CP(n301), .CDN(n340), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n212), .E(n243), .CP(n300), .CDN(n340), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n211), .E(N463), .CP(n298), .CDN(n340), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n210), .E(n241), .CP(n299), .CDN(n340), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n209), .E(n241), .CP(n306), .CDN(n352), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n208), .E(n241), .CP(n303), .CDN(n353), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n207), .E(n241), .CP(n302), .CDN(n329), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n206), .E(n241), .CP(n294), .CDN(n341), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n205), .E(N463), .CP(n295), .CDN(n342), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n204), .E(N463), .CP(n293), .CDN(n340), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n203), .E(N463), .CP(n292), .CDN(n327), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n202), .E(N463), .CP(n297), .CDN(n359), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n201), .E(n241), .CP(n296), .CDN(n341), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n200), .E(n243), .CP(n298), .CDN(n342), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n199), .E(n241), .CP(n299), .CDN(n340), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n198), .E(n241), .CP(n303), .CDN(n339), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n197), .E(n241), .CP(n295), .CDN(n339), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n196), .E(N463), .CP(n298), .CDN(n339), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n195), .E(N463), .CP(n301), .CDN(n339), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n194), .E(N463), .CP(n310), .CDN(n339), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n193), .E(N463), .CP(n311), .CDN(n339), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n192), .E(n241), .CP(n288), .CDN(n339), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n191), .E(n243), .CP(n292), .CDN(n339), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n190), .E(n243), .CP(n286), .CDN(n339), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n189), .E(n243), .CP(n285), .CDN(n339), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N84), .E(n245), .CP(n301), .CDN(n339), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n220), .E(n247), .CP(n306), .CDN(n348), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n219), .E(N430), .CP(n303), .CDN(n345), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n218), .E(N430), .CP(n302), .CDN(n351), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n213), .E(N430), .CP(n297), .CDN(n353), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n212), .E(N430), .CP(n308), .CDN(n347), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n211), .E(n247), .CP(n292), .CDN(n352), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n210), .E(n247), .CP(n285), .CDN(n359), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n209), .E(n247), .CP(n308), .CDN(n368), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n208), .E(n247), .CP(n307), .CDN(n360), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n207), .E(n247), .CP(n306), .CDN(n358), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n206), .E(n247), .CP(n305), .CDN(n360), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n205), .E(n247), .CP(n304), .CDN(n360), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n204), .E(n247), .CP(n289), .CDN(n360), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n203), .E(n247), .CP(n293), .CDN(n341), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n202), .E(n247), .CP(n285), .CDN(n341), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n201), .E(n245), .CP(n309), .CDN(n368), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n200), .E(n245), .CP(n287), .CDN(n334), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n199), .E(N430), .CP(n289), .CDN(n344), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n198), .E(N430), .CP(n288), .CDN(n338), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n197), .E(N430), .CP(n291), .CDN(n338), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n196), .E(n245), .CP(n290), .CDN(n338), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n195), .E(n245), .CP(n296), .CDN(n338), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n194), .E(n245), .CP(n290), .CDN(n338), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n193), .E(n245), .CP(n293), .CDN(n338), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n192), .E(n245), .CP(n295), .CDN(n338), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n191), .E(n245), .CP(n294), .CDN(n338), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n190), .E(n245), .CP(n297), .CDN(n338), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n189), .E(n247), .CP(n296), .CDN(n338), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N84), .E(N331), .CP(n303), .CDN(n343), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n220), .E(n259), .CP(n304), .CDN(n333), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n219), .E(n259), .CP(n308), .CDN(n333), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n218), .E(n259), .CP(n286), .CDN(n333), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n213), .E(n259), .CP(ClockW), .CDN(n333), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n212), .E(n259), .CP(n307), .CDN(n333), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n211), .E(N331), .CP(n310), .CDN(n333), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n210), .E(N331), .CP(n299), .CDN(n333), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n209), .E(n257), .CP(n290), .CDN(n332), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n208), .E(n257), .CP(n285), .CDN(n332), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n207), .E(n257), .CP(n304), .CDN(n332), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n206), .E(n257), .CP(n305), .CDN(n332), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n205), .E(n257), .CP(n306), .CDN(n332), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n204), .E(n257), .CP(n308), .CDN(n332), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n203), .E(n257), .CP(ClockW), .CDN(n332), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n202), .E(n257), .CP(n295), .CDN(n332), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n201), .E(n259), .CP(n291), .CDN(n332), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n200), .E(n257), .CP(n288), .CDN(n332), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n199), .E(n257), .CP(n297), .CDN(n332), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n198), .E(N331), .CP(n307), .CDN(n331), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n197), .E(N331), .CP(n297), .CDN(n331), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n196), .E(N331), .CP(n296), .CDN(n331), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n195), .E(N331), .CP(n296), .CDN(n331), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n194), .E(N331), .CP(n286), .CDN(n331), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n193), .E(N331), .CP(n289), .CDN(n331), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n192), .E(N331), .CP(n288), .CDN(n331), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n191), .E(n259), .CP(n291), .CDN(n331), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n190), .E(n259), .CP(n290), .CDN(n331), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n189), .E(n259), .CP(n294), .CDN(n331), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N84), .E(N298), .CP(n310), .CDN(n331), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n220), .E(n263), .CP(n285), .CDN(n355), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n219), .E(n263), .CP(n311), .CDN(n330), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n218), .E(n263), .CP(n307), .CDN(n362), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n213), .E(n263), .CP(n289), .CDN(n362), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n212), .E(n263), .CP(n303), .CDN(n321), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n211), .E(N298), .CP(n302), .CDN(n354), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n210), .E(N298), .CP(n300), .CDN(n321), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n209), .E(n261), .CP(n306), .CDN(n330), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n208), .E(n261), .CP(n311), .CDN(n330), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n207), .E(n261), .CP(n294), .CDN(n330), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n206), .E(n261), .CP(n304), .CDN(n330), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n205), .E(n261), .CP(n299), .CDN(n330), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n204), .E(n261), .CP(n290), .CDN(n330), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n203), .E(n261), .CP(n300), .CDN(n330), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n202), .E(n261), .CP(n292), .CDN(n330), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n201), .E(n263), .CP(n302), .CDN(n330), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n200), .E(n261), .CP(n298), .CDN(n330), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n199), .E(n261), .CP(n307), .CDN(n330), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n198), .E(N298), .CP(n310), .CDN(n329), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n197), .E(N298), .CP(n296), .CDN(n329), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n196), .E(N298), .CP(n311), .CDN(n329), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n195), .E(N298), .CP(n303), .CDN(n329), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n194), .E(N298), .CP(n286), .CDN(n329), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n193), .E(N298), .CP(n299), .CDN(n329), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n192), .E(N298), .CP(n286), .CDN(n329), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n191), .E(n263), .CP(n303), .CDN(n329), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n190), .E(n263), .CP(n311), .CDN(n329), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n189), .E(n263), .CP(n285), .CDN(n329), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N84), .E(N199), .CP(n309), .CDN(n324), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n220), .E(n275), .CP(n286), .CDN(n338), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n219), .E(n275), .CP(n306), .CDN(n338), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n218), .E(n275), .CP(n291), .CDN(n352), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n213), .E(n275), .CP(ClockW), .CDN(n365), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n212), .E(n275), .CP(n304), .CDN(n350), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n211), .E(N199), .CP(n300), .CDN(n365), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n210), .E(N199), .CP(n293), .CDN(n351), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n209), .E(n273), .CP(n308), .CDN(n323), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n208), .E(n273), .CP(n310), .CDN(n323), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n207), .E(n273), .CP(n304), .CDN(n323), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n206), .E(n273), .CP(n304), .CDN(n323), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n205), .E(n273), .CP(n310), .CDN(n323), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n204), .E(n273), .CP(n301), .CDN(n323), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n203), .E(n273), .CP(n299), .CDN(n323), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n202), .E(n273), .CP(n304), .CDN(n323), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n201), .E(n275), .CP(n304), .CDN(n323), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n200), .E(n273), .CP(n307), .CDN(n323), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n199), .E(n273), .CP(n305), .CDN(n323), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n198), .E(N199), .CP(n307), .CDN(n322), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n197), .E(N199), .CP(n309), .CDN(n322), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n196), .E(N199), .CP(n292), .CDN(n322), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n195), .E(N199), .CP(n299), .CDN(n322), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n194), .E(N199), .CP(ClockW), .CDN(n322), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n193), .E(N199), .CP(n294), .CDN(n322), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n192), .E(N199), .CP(n304), .CDN(n322), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n191), .E(n275), .CP(n286), .CDN(n322), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n190), .E(n275), .CP(n311), .CDN(n322), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n189), .E(n275), .CP(n304), .CDN(n322), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N84), .E(N166), .CP(n300), .CDN(n322), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n220), .E(n279), .CP(n302), .CDN(n341), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n219), .E(n279), .CP(n303), .CDN(n353), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n218), .E(n279), .CP(n309), .CDN(n354), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n213), .E(n279), .CP(n310), .CDN(n321), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n212), .E(n279), .CP(n287), .CDN(n320), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n211), .E(N166), .CP(n303), .CDN(n321), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n210), .E(N166), .CP(n308), .CDN(n321), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n209), .E(n277), .CP(n310), .CDN(n342), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n208), .E(n277), .CP(ClockW), .CDN(n359), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n207), .E(n277), .CP(n298), .CDN(n353), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n206), .E(n277), .CP(n286), .CDN(n353), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n205), .E(n277), .CP(n305), .CDN(n353), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n204), .E(n277), .CP(n307), .CDN(n326), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n203), .E(n277), .CP(n306), .CDN(n328), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n202), .E(n277), .CP(n290), .CDN(n341), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n201), .E(n279), .CP(n305), .CDN(n323), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n200), .E(n277), .CP(n302), .CDN(n342), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n199), .E(n277), .CP(n311), .CDN(n363), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n198), .E(N166), .CP(n285), .CDN(n321), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n197), .E(N166), .CP(n302), .CDN(n321), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n196), .E(N166), .CP(n309), .CDN(n321), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n195), .E(N166), .CP(n285), .CDN(n321), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n194), .E(N166), .CP(n305), .CDN(n321), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n193), .E(N166), .CP(n311), .CDN(n321), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n192), .E(N166), .CP(n293), .CDN(n321), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n191), .E(n279), .CP(n311), .CDN(n321), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n190), .E(n279), .CP(n304), .CDN(n321), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n189), .E(n279), .CP(n301), .CDN(n321), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N84), .E(n221), .CP(n287), .CDN(n353), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n220), .E(n223), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n219), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n218), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n213), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n212), .E(N628), .CP(n288), .CDN(n352), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n211), .E(n223), .CP(n288), .CDN(n352), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n210), .E(n223), .CP(n288), .CDN(n352), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n209), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n208), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n207), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n206), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n205), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n204), .E(n223), .CP(n288), .CDN(n351), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n203), .E(n223), .CP(n289), .CDN(n351), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n202), .E(n223), .CP(n289), .CDN(n351), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n201), .E(n221), .CP(n289), .CDN(n351), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n200), .E(n221), .CP(n289), .CDN(n351), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n199), .E(N628), .CP(n289), .CDN(n351), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n198), .E(N628), .CP(n289), .CDN(n350), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n197), .E(N628), .CP(n289), .CDN(n350), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n196), .E(n221), .CP(n289), .CDN(n350), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n195), .E(n221), .CP(n289), .CDN(n350), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n194), .E(n221), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n193), .E(n221), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n192), .E(n221), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n191), .E(n221), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n190), .E(n221), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n189), .E(n223), .CP(n290), .CDN(n350), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N84), .E(N529), .CP(n298), .CDN(n346), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n220), .E(N529), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n219), .E(N529), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n218), .E(n233), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n213), .E(n233), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n212), .E(n233), .CP(n299), .CDN(n345), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n211), .E(N529), .CP(n299), .CDN(n345), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n210), .E(n235), .CP(n299), .CDN(n345), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n209), .E(n235), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n208), .E(n233), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n207), .E(N529), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n206), .E(N529), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n205), .E(N529), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n204), .E(N529), .CP(n299), .CDN(n344), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n203), .E(N529), .CP(n300), .CDN(n344), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n202), .E(N529), .CP(n300), .CDN(n344), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n201), .E(n235), .CP(n300), .CDN(n344), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n200), .E(n235), .CP(n300), .CDN(n344), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n199), .E(n235), .CP(n300), .CDN(n344), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n198), .E(n235), .CP(n300), .CDN(n343), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n197), .E(n235), .CP(n300), .CDN(n343), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n196), .E(n235), .CP(n300), .CDN(n343), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n195), .E(n235), .CP(n300), .CDN(n343), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n194), .E(n235), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n193), .E(n235), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n192), .E(n235), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n191), .E(n233), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n190), .E(n233), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n189), .E(n233), .CP(n301), .CDN(n343), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N84), .E(N496), .CP(n301), .CDN(n343), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n220), .E(n239), .CP(n301), .CDN(n342), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n219), .E(n239), .CP(n301), .CDN(n342), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n218), .E(n239), .CP(n305), .CDN(n342), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n213), .E(n239), .CP(n297), .CDN(n342), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n212), .E(n239), .CP(n298), .CDN(n342), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n211), .E(N496), .CP(n300), .CDN(n342), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n210), .E(N496), .CP(n301), .CDN(n342), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n209), .E(n237), .CP(n287), .CDN(n341), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n208), .E(n237), .CP(n291), .CDN(n341), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n207), .E(n237), .CP(n290), .CDN(n341), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n206), .E(n237), .CP(n289), .CDN(n341), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n205), .E(n237), .CP(n288), .CDN(n341), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n204), .E(n237), .CP(n292), .CDN(n341), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n203), .E(n237), .CP(n309), .CDN(n341), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n202), .E(n237), .CP(ClockW), .CDN(n341), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n201), .E(n239), .CP(n286), .CDN(n341), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n200), .E(n237), .CP(n310), .CDN(n341), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n199), .E(n237), .CP(n303), .CDN(n341), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n198), .E(N496), .CP(n310), .CDN(n353), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n197), .E(N496), .CP(n285), .CDN(n342), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n196), .E(N496), .CP(n308), .CDN(n359), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n195), .E(N496), .CP(n307), .CDN(n354), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n194), .E(N496), .CP(n305), .CDN(n348), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n193), .E(N496), .CP(n304), .CDN(n320), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n192), .E(N496), .CP(n285), .CDN(n359), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n191), .E(n239), .CP(n289), .CDN(n354), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n190), .E(n239), .CP(n297), .CDN(n345), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n189), .E(n239), .CP(n296), .CDN(n320), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N84), .E(N397), .CP(n302), .CDN(n338), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n220), .E(n251), .CP(n292), .CDN(n337), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n219), .E(n251), .CP(n295), .CDN(n337), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n218), .E(n251), .CP(n297), .CDN(n337), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n213), .E(n251), .CP(n303), .CDN(n337), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n212), .E(n251), .CP(n302), .CDN(n337), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n211), .E(N397), .CP(n298), .CDN(n337), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n210), .E(N397), .CP(n306), .CDN(n337), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n209), .E(n249), .CP(n285), .CDN(n336), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n208), .E(n249), .CP(n286), .CDN(n336), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n207), .E(n249), .CP(n307), .CDN(n336), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n206), .E(n249), .CP(n301), .CDN(n336), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n205), .E(n249), .CP(n302), .CDN(n336), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n204), .E(n249), .CP(n307), .CDN(n336), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n203), .E(n249), .CP(n291), .CDN(n336), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n202), .E(n249), .CP(n311), .CDN(n336), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n201), .E(n251), .CP(n288), .CDN(n336), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n200), .E(n249), .CP(n296), .CDN(n336), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n199), .E(n249), .CP(n290), .CDN(n336), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n198), .E(N397), .CP(n291), .CDN(n335), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n197), .E(N397), .CP(n288), .CDN(n335), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n196), .E(N397), .CP(n289), .CDN(n335), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n195), .E(N397), .CP(n287), .CDN(n335), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n194), .E(N397), .CP(n292), .CDN(n335), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n193), .E(N397), .CP(n293), .CDN(n335), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n192), .E(N397), .CP(n294), .CDN(n335), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n191), .E(n251), .CP(n307), .CDN(n335), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n190), .E(n251), .CP(n308), .CDN(n335), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n189), .E(n251), .CP(n289), .CDN(n335), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N84), .E(N364), .CP(ClockW), .CDN(n335), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n220), .E(n255), .CP(n309), .CDN(n334), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n219), .E(n255), .CP(n288), .CDN(n334), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n218), .E(n255), .CP(n289), .CDN(n334), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n213), .E(n255), .CP(n294), .CDN(n334), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n212), .E(n255), .CP(n295), .CDN(n334), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n211), .E(N364), .CP(n292), .CDN(n334), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n210), .E(N364), .CP(n293), .CDN(n334), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n209), .E(n253), .CP(n296), .CDN(n321), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n208), .E(n253), .CP(n302), .CDN(n361), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n207), .E(n253), .CP(n287), .CDN(n341), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n206), .E(n253), .CP(n297), .CDN(n361), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n205), .E(n253), .CP(n311), .CDN(n360), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n204), .E(n253), .CP(n311), .CDN(n361), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n203), .E(n253), .CP(n291), .CDN(n362), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n202), .E(n253), .CP(n289), .CDN(n334), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n201), .E(n255), .CP(n310), .CDN(n367), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n200), .E(n253), .CP(n286), .CDN(n367), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n199), .E(n253), .CP(n286), .CDN(n320), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n198), .E(N364), .CP(n303), .CDN(n362), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n197), .E(N364), .CP(n309), .CDN(n354), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n196), .E(N364), .CP(n301), .CDN(n334), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n195), .E(N364), .CP(n308), .CDN(n321), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n194), .E(N364), .CP(n307), .CDN(n354), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n193), .E(N364), .CP(n287), .CDN(n342), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n192), .E(N364), .CP(n301), .CDN(n362), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n191), .E(n255), .CP(n310), .CDN(n361), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n190), .E(n255), .CP(n309), .CDN(n321), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n189), .E(n255), .CP(n308), .CDN(n354), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N84), .E(N265), .CP(n287), .CDN(n329), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n220), .E(n267), .CP(n302), .CDN(n328), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n219), .E(n267), .CP(n300), .CDN(n328), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n218), .E(n267), .CP(n293), .CDN(n328), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n213), .E(n267), .CP(n293), .CDN(n328), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n212), .E(n267), .CP(n298), .CDN(n328), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n211), .E(N265), .CP(n309), .CDN(n328), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n210), .E(N265), .CP(n302), .CDN(n328), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n209), .E(n265), .CP(n310), .CDN(n327), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n208), .E(n265), .CP(n308), .CDN(n327), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n207), .E(n265), .CP(n311), .CDN(n327), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n206), .E(n265), .CP(n298), .CDN(n327), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n205), .E(n265), .CP(n305), .CDN(n327), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n204), .E(n265), .CP(n295), .CDN(n327), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n203), .E(n265), .CP(n285), .CDN(n327), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n202), .E(n265), .CP(n286), .CDN(n327), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n201), .E(n267), .CP(ClockW), .CDN(n327), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n200), .E(n265), .CP(n299), .CDN(n327), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n199), .E(n265), .CP(n291), .CDN(n327), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n198), .E(N265), .CP(ClockW), .CDN(n326), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n197), .E(N265), .CP(n309), .CDN(n326), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n196), .E(N265), .CP(n308), .CDN(n326), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n195), .E(N265), .CP(n307), .CDN(n326), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n194), .E(N265), .CP(n286), .CDN(n326), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n193), .E(N265), .CP(n300), .CDN(n326), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n192), .E(N265), .CP(n303), .CDN(n326), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n191), .E(n267), .CP(n311), .CDN(n326), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n190), .E(n267), .CP(n290), .CDN(n326), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n189), .E(n267), .CP(n305), .CDN(n326), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N84), .E(N232), .CP(n309), .CDN(n326), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n220), .E(n271), .CP(ClockW), .CDN(n348), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n219), .E(n271), .CP(n306), .CDN(n325), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n218), .E(n271), .CP(n305), .CDN(n324), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n213), .E(n271), .CP(n304), .CDN(n324), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n212), .E(n271), .CP(n286), .CDN(n322), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n211), .E(N232), .CP(n306), .CDN(n324), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n210), .E(N232), .CP(n307), .CDN(n365), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n209), .E(n269), .CP(n304), .CDN(n325), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n208), .E(n269), .CP(n305), .CDN(n325), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n207), .E(n269), .CP(n311), .CDN(n325), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n206), .E(n269), .CP(n311), .CDN(n325), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n205), .E(n269), .CP(n287), .CDN(n325), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n204), .E(n269), .CP(ClockW), .CDN(n325), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n203), .E(n269), .CP(n285), .CDN(n325), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n202), .E(n269), .CP(n285), .CDN(n325), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n201), .E(n271), .CP(n288), .CDN(n325), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n200), .E(n269), .CP(n303), .CDN(n325), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n199), .E(n269), .CP(n302), .CDN(n325), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n198), .E(N232), .CP(n285), .CDN(n324), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n197), .E(N232), .CP(n294), .CDN(n324), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n196), .E(N232), .CP(n295), .CDN(n324), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n195), .E(N232), .CP(n302), .CDN(n324), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n194), .E(N232), .CP(n309), .CDN(n324), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n193), .E(N232), .CP(n301), .CDN(n324), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n192), .E(N232), .CP(n295), .CDN(n324), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n191), .E(n271), .CP(ClockW), .CDN(n324), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n190), .E(n271), .CP(n306), .CDN(n324), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n189), .E(n271), .CP(n310), .CDN(n324), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N84), .E(N133), .CP(n305), .CDN(n321), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n220), .E(N133), .CP(n300), .CDN(n320), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n219), .E(n281), .CP(ClockW), .CDN(n320), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n218), .E(n281), .CP(n286), .CDN(n320), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n213), .E(n281), .CP(n285), .CDN(n320), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n212), .E(n281), .CP(n304), .CDN(n320), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n211), .E(n283), .CP(n285), .CDN(n320), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n210), .E(n283), .CP(n306), .CDN(n320), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n209), .E(n283), .CP(n303), .CDN(n342), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n208), .E(n283), .CP(n302), .CDN(n339), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n207), .E(n283), .CP(n306), .CDN(n365), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n206), .E(n283), .CP(n292), .CDN(n356), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n205), .E(n283), .CP(n296), .CDN(n358), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n204), .E(n283), .CP(n287), .CDN(n343), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n203), .E(n283), .CP(n300), .CDN(n359), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n202), .E(n283), .CP(n291), .CDN(n356), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n201), .E(N133), .CP(n304), .CDN(n341), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n200), .E(N133), .CP(n310), .CDN(n342), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n199), .E(N133), .CP(n305), .CDN(n353), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n198), .E(N133), .CP(n309), .CDN(n319), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n197), .E(N133), .CP(n305), .CDN(n319), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n196), .E(N133), .CP(n308), .CDN(n319), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n195), .E(N133), .CP(n310), .CDN(n319), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n194), .E(n281), .CP(n301), .CDN(n319), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n193), .E(n281), .CP(n306), .CDN(n319), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n192), .E(N133), .CP(n293), .CDN(n319), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n191), .E(n281), .CP(n298), .CDN(n319), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n190), .E(n281), .CP(n306), .CDN(n319), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n189), .E(n281), .CP(ClockW), .CDN(n319), 
        .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n374), .CP(ClockR), .CDN(n319), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n217), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n216), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n215), .E(n225), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n214), .E(N595), .CP(n291), .CDN(n349), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n217), .E(n231), .CP(n294), .CDN(n345), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n216), .E(n231), .CP(n294), .CDN(n346), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n215), .E(n229), .CP(n295), .CDN(n358), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n214), .E(N562), .CP(n295), .CDN(n323), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n217), .E(n243), .CP(n294), .CDN(n340), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n216), .E(n243), .CP(n295), .CDN(n340), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n215), .E(n241), .CP(n286), .CDN(n340), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n214), .E(N463), .CP(n309), .CDN(n340), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n217), .E(N430), .CP(n288), .CDN(n344), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n216), .E(N430), .CP(n307), .CDN(n319), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n215), .E(N430), .CP(ClockW), .CDN(n354), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n214), .E(N430), .CP(n309), .CDN(n320), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n217), .E(n259), .CP(n310), .CDN(n333), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n216), .E(n259), .CP(n309), .CDN(n333), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n215), .E(n257), .CP(n288), .CDN(n333), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n214), .E(N331), .CP(n302), .CDN(n333), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n217), .E(n263), .CP(n305), .CDN(n342), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n216), .E(n263), .CP(n294), .CDN(n349), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n215), .E(n261), .CP(n295), .CDN(n350), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n214), .E(N298), .CP(n308), .CDN(n351), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n217), .E(n275), .CP(n286), .CDN(n338), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n216), .E(n275), .CP(n285), .CDN(n328), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n215), .E(n273), .CP(n303), .CDN(n326), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n214), .E(N199), .CP(n309), .CDN(n327), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n217), .E(n279), .CP(n297), .CDN(n320), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n216), .E(n279), .CP(n296), .CDN(n341), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n215), .E(n277), .CP(n308), .CDN(n322), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n214), .E(N166), .CP(n306), .CDN(n321), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n217), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n216), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n215), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n214), .E(N628), .CP(n287), .CDN(n352), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n217), .E(n233), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n216), .E(n233), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n215), .E(n233), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n214), .E(N529), .CP(n298), .CDN(n345), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n217), .E(n239), .CP(n294), .CDN(n342), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n216), .E(n239), .CP(n308), .CDN(n342), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n215), .E(n237), .CP(n306), .CDN(n342), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n214), .E(N496), .CP(n311), .CDN(n342), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n217), .E(n251), .CP(n300), .CDN(n337), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n216), .E(n251), .CP(n308), .CDN(n337), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n215), .E(n249), .CP(n307), .CDN(n337), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n214), .E(N397), .CP(n305), .CDN(n337), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n217), .E(n255), .CP(n303), .CDN(n334), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n216), .E(n255), .CP(n290), .CDN(n334), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n215), .E(n253), .CP(n289), .CDN(n334), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n214), .E(N364), .CP(n298), .CDN(n334), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n217), .E(n267), .CP(n299), .CDN(n328), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n216), .E(n267), .CP(n302), .CDN(n328), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n215), .E(n265), .CP(n292), .CDN(n328), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n214), .E(N265), .CP(n299), .CDN(n328), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n217), .E(n271), .CP(n303), .CDN(n364), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n216), .E(n271), .CP(n286), .CDN(n366), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n215), .E(n269), .CP(n293), .CDN(n366), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n214), .E(N232), .CP(n297), .CDN(n366), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n217), .E(n281), .CP(n307), .CDN(n320), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n216), .E(n283), .CP(n308), .CDN(n320), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n215), .E(N133), .CP(n309), .CDN(n320), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n214), .E(n283), .CP(n306), .CDN(n320), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N50), .E(Read), .CP(n312), .CDN(n320), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N51), .E(Read), .CP(n312), .CDN(n354), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N52), .E(Read), .CP(n312), .CDN(n354), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N53), .E(Read), .CP(ClockR), .CDN(n354), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N54), .E(Read), .CP(ClockR), .CDN(n354), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N55), .E(Read), .CP(n312), .CDN(n354), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N56), .E(Read), .CP(n312), .CDN(n354), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N57), .E(Read), .CP(ClockR), .CDN(n354), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N58), .E(n316), .CP(ClockR), .CDN(n354), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N59), .E(Read), .CP(n312), .CDN(n354), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N60), .E(n314), .CP(ClockR), .CDN(n354), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N61), .E(n314), .CP(ClockR), .CDN(n354), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N62), .E(n314), .CP(n312), .CDN(n360), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N63), .E(n314), .CP(n312), .CDN(n364), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N64), .E(n314), .CP(ClockR), .CDN(n338), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N65), .E(n314), .CP(n312), .CDN(n365), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N66), .E(n314), .CP(n312), .CDN(n319), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N67), .E(n314), .CP(ClockR), .CDN(n338), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N68), .E(n314), .CP(n312), .CDN(n324), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N69), .E(n314), .CP(n312), .CDN(n357), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N70), .E(Read), .CP(n312), .CDN(n346), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N71), .E(Read), .CP(n312), .CDN(n325), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N72), .E(Read), .CP(n312), .CDN(n324), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N73), .E(n316), .CP(n312), .CDN(n353), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N74), .E(n316), .CP(n312), .CDN(n353), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N75), .E(Read), .CP(n312), .CDN(n353), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N76), .E(Read), .CP(n312), .CDN(n353), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N77), .E(Read), .CP(ClockR), .CDN(n353), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N78), .E(n316), .CP(ClockR), .CDN(n353), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N79), .E(Read), .CP(ClockR), .CDN(n353), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N80), .E(Read), .CP(ClockR), .CDN(n353), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N81), .E(n316), .CP(ClockR), .CDN(n353), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N82), .E(Read), .CP(ClockR), .CDN(n353), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKBD0 U4 ( .CLK(N45), .C(n176) );
  CKBD0 U5 ( .CLK(N45), .C(n175) );
  CKBD0 U6 ( .CLK(N44), .C(n182) );
  CKNXD0 U7 ( .I(n233), .ZN(n236) );
  CKNXD0 U8 ( .I(n225), .ZN(n228) );
  CKNXD0 U9 ( .I(n281), .ZN(n284) );
  NR2XD0 U10 ( .A1(n382), .A2(n378), .ZN(N133) );
  INVD0 U11 ( .I(n269), .ZN(n272) );
  INVD0 U12 ( .I(n270), .ZN(n269) );
  CKNXD0 U18 ( .I(n272), .ZN(n271) );
  INVD0 U19 ( .I(n265), .ZN(n268) );
  INVD0 U20 ( .I(n266), .ZN(n265) );
  CKNXD0 U23 ( .I(n268), .ZN(n267) );
  INVD0 U24 ( .I(n253), .ZN(n256) );
  INVD0 U25 ( .I(n254), .ZN(n253) );
  CKNXD0 U26 ( .I(n256), .ZN(n255) );
  INVD0 U31 ( .I(n249), .ZN(n252) );
  INVD0 U32 ( .I(n250), .ZN(n249) );
  CKNXD0 U33 ( .I(n252), .ZN(n251) );
  INVD0 U34 ( .I(n237), .ZN(n240) );
  INVD0 U35 ( .I(n238), .ZN(n237) );
  CKNXD0 U36 ( .I(n240), .ZN(n239) );
  INVD0 U37 ( .I(n277), .ZN(n280) );
  INVD0 U38 ( .I(n278), .ZN(n277) );
  CKNXD0 U39 ( .I(n280), .ZN(n279) );
  INVD0 U40 ( .I(n273), .ZN(n276) );
  INVD0 U41 ( .I(n274), .ZN(n273) );
  CKNXD0 U42 ( .I(n276), .ZN(n275) );
  INVD0 U43 ( .I(n261), .ZN(n264) );
  INVD0 U44 ( .I(n262), .ZN(n261) );
  CKNXD0 U45 ( .I(n264), .ZN(n263) );
  INVD0 U46 ( .I(n257), .ZN(n260) );
  INVD0 U47 ( .I(n258), .ZN(n257) );
  CKNXD0 U48 ( .I(n260), .ZN(n259) );
  INVD0 U49 ( .I(n229), .ZN(n232) );
  INVD0 U50 ( .I(n230), .ZN(n229) );
  CKNXD0 U51 ( .I(n232), .ZN(n231) );
  INVD0 U52 ( .I(n236), .ZN(n235) );
  CKNXD0 U53 ( .I(n234), .ZN(n233) );
  INVD0 U54 ( .I(n241), .ZN(n244) );
  INVD0 U55 ( .I(n228), .ZN(n227) );
  CKNXD0 U56 ( .I(n226), .ZN(n225) );
  INVD0 U57 ( .I(n282), .ZN(n281) );
  INVD0 U58 ( .I(n221), .ZN(n224) );
  INVD0 U59 ( .I(n224), .ZN(n223) );
  INVD0 U60 ( .I(n222), .ZN(n221) );
  NR2XD0 U61 ( .A1(n386), .A2(n379), .ZN(N364) );
  NR2XD0 U62 ( .A1(n386), .A2(n378), .ZN(N331) );
  NR2XD0 U63 ( .A1(n383), .A2(n379), .ZN(N232) );
  NR2XD0 U64 ( .A1(n384), .A2(n378), .ZN(N265) );
  NR2XD0 U65 ( .A1(n387), .A2(n383), .ZN(N496) );
  NR2XD0 U66 ( .A1(n384), .A2(n379), .ZN(N298) );
  NR2XD0 U67 ( .A1(n387), .A2(n384), .ZN(N562) );
  INVD0 U68 ( .I(N595), .ZN(n226) );
  NR2XD0 U69 ( .A1(n386), .A2(n385), .ZN(N595) );
  INVD0 U70 ( .I(N529), .ZN(n234) );
  NR2XD0 U71 ( .A1(n385), .A2(n384), .ZN(N529) );
  NR2XD0 U72 ( .A1(n383), .A2(n378), .ZN(N199) );
  NR2XD0 U73 ( .A1(n382), .A2(n379), .ZN(N166) );
  INVD0 U74 ( .I(N463), .ZN(n242) );
  CKNXD0 U75 ( .I(n244), .ZN(n243) );
  INVD0 U76 ( .I(n242), .ZN(n241) );
  NR2XD0 U77 ( .A1(n385), .A2(n383), .ZN(N463) );
  INVD0 U78 ( .I(N133), .ZN(n282) );
  CKNXD0 U79 ( .I(n284), .ZN(n283) );
  NR2XD0 U80 ( .A1(n385), .A2(n382), .ZN(N397) );
  INVD0 U81 ( .I(n245), .ZN(n248) );
  INVD0 U82 ( .I(n248), .ZN(n247) );
  INVD0 U83 ( .I(n246), .ZN(n245) );
  NR2XD0 U84 ( .A1(n387), .A2(n382), .ZN(N430) );
  INVD0 U85 ( .I(Read), .ZN(n317) );
  CKNXD0 U86 ( .I(n317), .ZN(n316) );
  INVD0 U87 ( .I(n318), .ZN(n173) );
  CKBD0 U88 ( .CLK(N46), .C(n318) );
  CKAN2D0 U89 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  INVD1 U90 ( .I(N47), .ZN(n171) );
  BUFFD1 U91 ( .I(n365), .Z(n322) );
  BUFFD1 U92 ( .I(n365), .Z(n323) );
  BUFFD1 U93 ( .I(n364), .Z(n324) );
  BUFFD1 U94 ( .I(n357), .Z(n325) );
  BUFFD1 U95 ( .I(n363), .Z(n326) );
  BUFFD1 U96 ( .I(n363), .Z(n327) );
  BUFFD1 U97 ( .I(n363), .Z(n328) );
  BUFFD1 U98 ( .I(n363), .Z(n329) );
  BUFFD1 U99 ( .I(n362), .Z(n330) );
  BUFFD1 U100 ( .I(n361), .Z(n331) );
  BUFFD1 U101 ( .I(n361), .Z(n332) );
  BUFFD1 U102 ( .I(n361), .Z(n333) );
  BUFFD1 U103 ( .I(n363), .Z(n334) );
  BUFFD1 U104 ( .I(n360), .Z(n335) );
  BUFFD1 U105 ( .I(n360), .Z(n336) );
  BUFFD1 U106 ( .I(n360), .Z(n337) );
  BUFFD1 U107 ( .I(n364), .Z(n338) );
  BUFFD1 U108 ( .I(n359), .Z(n339) );
  BUFFD1 U109 ( .I(n357), .Z(n340) );
  BUFFD1 U110 ( .I(n368), .Z(n341) );
  BUFFD1 U111 ( .I(n367), .Z(n342) );
  BUFFD1 U112 ( .I(n358), .Z(n343) );
  BUFFD1 U113 ( .I(n358), .Z(n344) );
  BUFFD1 U114 ( .I(n357), .Z(n345) );
  BUFFD1 U115 ( .I(n357), .Z(n346) );
  BUFFD1 U116 ( .I(n356), .Z(n347) );
  BUFFD1 U117 ( .I(n357), .Z(n348) );
  BUFFD1 U118 ( .I(n355), .Z(n349) );
  BUFFD1 U119 ( .I(n355), .Z(n350) );
  BUFFD1 U120 ( .I(n355), .Z(n351) );
  BUFFD1 U121 ( .I(n355), .Z(n352) );
  BUFFD1 U122 ( .I(n371), .Z(n353) );
  BUFFD1 U123 ( .I(n366), .Z(n354) );
  BUFFD1 U124 ( .I(n357), .Z(n319) );
  BUFFD1 U125 ( .I(n370), .Z(n320) );
  BUFFD1 U126 ( .I(n366), .Z(n321) );
  BUFFD1 U127 ( .I(n366), .Z(n365) );
  BUFFD1 U128 ( .I(n366), .Z(n364) );
  BUFFD1 U129 ( .I(n368), .Z(n363) );
  BUFFD1 U130 ( .I(n367), .Z(n362) );
  BUFFD1 U131 ( .I(n367), .Z(n361) );
  BUFFD1 U132 ( .I(n368), .Z(n360) );
  BUFFD1 U133 ( .I(n369), .Z(n359) );
  BUFFD1 U134 ( .I(n369), .Z(n358) );
  BUFFD1 U135 ( .I(n369), .Z(n357) );
  BUFFD1 U136 ( .I(n369), .Z(n356) );
  BUFFD1 U137 ( .I(n369), .Z(n355) );
  BUFFD1 U138 ( .I(n372), .Z(n366) );
  BUFFD1 U139 ( .I(n371), .Z(n367) );
  BUFFD1 U140 ( .I(n371), .Z(n368) );
  BUFFD1 U141 ( .I(n370), .Z(n369) );
  BUFFD1 U142 ( .I(n373), .Z(n371) );
  BUFFD1 U143 ( .I(n373), .Z(n370) );
  BUFFD1 U144 ( .I(n373), .Z(n372) );
  INVD1 U145 ( .I(Reset), .ZN(n373) );
  BUFFD1 U146 ( .I(n302), .Z(n301) );
  BUFFD1 U147 ( .I(n302), .Z(n300) );
  BUFFD1 U148 ( .I(n303), .Z(n299) );
  BUFFD1 U149 ( .I(n303), .Z(n298) );
  BUFFD1 U150 ( .I(n304), .Z(n297) );
  BUFFD1 U151 ( .I(n304), .Z(n296) );
  BUFFD1 U152 ( .I(n305), .Z(n295) );
  BUFFD1 U153 ( .I(n305), .Z(n294) );
  BUFFD1 U154 ( .I(n306), .Z(n293) );
  BUFFD1 U155 ( .I(n306), .Z(n292) );
  BUFFD1 U156 ( .I(n307), .Z(n291) );
  BUFFD1 U157 ( .I(n307), .Z(n290) );
  BUFFD1 U158 ( .I(n308), .Z(n289) );
  BUFFD1 U159 ( .I(n308), .Z(n288) );
  BUFFD1 U160 ( .I(n309), .Z(n287) );
  BUFFD1 U161 ( .I(n310), .Z(n309) );
  BUFFD1 U162 ( .I(n305), .Z(n302) );
  BUFFD1 U163 ( .I(n304), .Z(n303) );
  BUFFD1 U164 ( .I(n311), .Z(n304) );
  BUFFD1 U165 ( .I(n311), .Z(n305) );
  BUFFD1 U166 ( .I(n311), .Z(n306) );
  BUFFD1 U167 ( .I(n310), .Z(n307) );
  BUFFD1 U168 ( .I(n310), .Z(n308) );
  BUFFD1 U169 ( .I(n285), .Z(n311) );
  BUFFD1 U170 ( .I(n285), .Z(n310) );
  BUFFD1 U171 ( .I(n186), .Z(n184) );
  BUFFD1 U172 ( .I(n182), .Z(n185) );
  BUFFD1 U173 ( .I(n183), .Z(n186) );
  BUFFD1 U174 ( .I(n182), .Z(n187) );
  BUFFD1 U175 ( .I(n182), .Z(n188) );
  BUFFD1 U176 ( .I(n176), .Z(n177) );
  BUFFD1 U177 ( .I(n175), .Z(n178) );
  BUFFD1 U178 ( .I(N45), .Z(n179) );
  BUFFD1 U179 ( .I(n175), .Z(n180) );
  BUFFD1 U180 ( .I(n175), .Z(n181) );
  INVD1 U181 ( .I(N397), .ZN(n250) );
  INVD1 U182 ( .I(n315), .ZN(n314) );
  BUFFD1 U183 ( .I(n286), .Z(n285) );
  INVD1 U184 ( .I(n313), .ZN(n312) );
  XOR3D1 U185 ( .A1(n191), .A2(n190), .A3(n411), .Z(N84) );
  XOR3D1 U186 ( .A1(n189), .A2(n410), .A3(n409), .Z(n411) );
  XOR3D1 U187 ( .A1(n194), .A2(n193), .A3(n408), .Z(n409) );
  XOR3D1 U188 ( .A1(n208), .A2(n207), .A3(n402), .Z(n403) );
  XOR3D1 U189 ( .A1(n401), .A2(n206), .A3(n400), .Z(n402) );
  XOR3D1 U190 ( .A1(n407), .A2(n192), .A3(n406), .Z(n408) );
  XOR3D1 U191 ( .A1(n201), .A2(n200), .A3(n405), .Z(n406) );
  XOR3D1 U192 ( .A1(n404), .A2(n199), .A3(n403), .Z(n405) );
  XOR3D1 U193 ( .A1(N66), .A2(N65), .A3(n393), .Z(n395) );
  XOR3D1 U194 ( .A1(N64), .A2(n392), .A3(n391), .Z(n393) );
  XOR3D1 U195 ( .A1(N59), .A2(N58), .A3(n390), .Z(n391) );
  XOR3D1 U196 ( .A1(n389), .A2(N57), .A3(n388), .Z(n390) );
  XOR3D1 U197 ( .A1(N78), .A2(N73), .A3(n399), .Z(N82) );
  XOR3D1 U198 ( .A1(N72), .A2(n398), .A3(n397), .Z(n399) );
  XOR3D1 U199 ( .A1(N76), .A2(N75), .A3(n396), .Z(n397) );
  BUFFD1 U200 ( .I(N44), .Z(n183) );
  INVD1 U201 ( .I(n171), .ZN(n172) );
  INVD1 U202 ( .I(n173), .ZN(n174) );
  ND2D1 U203 ( .A1(n375), .A2(n380), .ZN(n378) );
  ND2D1 U204 ( .A1(n377), .A2(n376), .ZN(n382) );
  ND2D1 U205 ( .A1(n381), .A2(n380), .ZN(n385) );
  INVD1 U206 ( .I(N199), .ZN(n274) );
  INVD1 U207 ( .I(N232), .ZN(n270) );
  INVD1 U208 ( .I(N265), .ZN(n266) );
  INVD1 U209 ( .I(N298), .ZN(n262) );
  INVD1 U210 ( .I(N331), .ZN(n258) );
  INVD1 U211 ( .I(N364), .ZN(n254) );
  INVD1 U212 ( .I(N166), .ZN(n278) );
  INVD1 U213 ( .I(N430), .ZN(n246) );
  INVD1 U214 ( .I(N496), .ZN(n238) );
  INVD1 U215 ( .I(N562), .ZN(n230) );
  INVD1 U216 ( .I(N628), .ZN(n222) );
  NR2D1 U217 ( .A1(n387), .A2(n386), .ZN(N628) );
  INVD1 U218 ( .I(n316), .ZN(n315) );
  INVD1 U219 ( .I(ClockR), .ZN(n313) );
  BUFFD1 U220 ( .I(ClockW), .Z(n286) );
  BUFFD1 U221 ( .I(DataI[14]), .Z(n203) );
  BUFFD1 U222 ( .I(DataI[15]), .Z(n204) );
  BUFFD1 U223 ( .I(DataI[21]), .Z(n210) );
  BUFFD1 U224 ( .I(DataI[22]), .Z(n211) );
  BUFFD1 U225 ( .I(DataI[25]), .Z(n214) );
  BUFFD1 U226 ( .I(DataI[26]), .Z(n215) );
  BUFFD1 U227 ( .I(DataI[29]), .Z(n218) );
  BUFFD1 U228 ( .I(DataI[30]), .Z(n219) );
  BUFFD1 U229 ( .I(DataI[10]), .Z(n199) );
  BUFFD1 U230 ( .I(DataI[17]), .Z(n206) );
  BUFFD1 U231 ( .I(DataI[18]), .Z(n207) );
  BUFFD1 U232 ( .I(DataI[13]), .Z(n202) );
  BUFFD1 U233 ( .I(DataI[16]), .Z(n205) );
  BUFFD1 U234 ( .I(DataI[20]), .Z(n209) );
  BUFFD1 U235 ( .I(DataI[23]), .Z(n212) );
  BUFFD1 U236 ( .I(DataI[24]), .Z(n213) );
  BUFFD1 U237 ( .I(DataI[27]), .Z(n216) );
  BUFFD1 U238 ( .I(DataI[28]), .Z(n217) );
  BUFFD1 U239 ( .I(DataI[31]), .Z(n220) );
  BUFFD1 U240 ( .I(DataI[19]), .Z(n208) );
  BUFFD1 U241 ( .I(DataI[2]), .Z(n191) );
  BUFFD1 U242 ( .I(DataI[1]), .Z(n190) );
  BUFFD1 U243 ( .I(DataI[7]), .Z(n196) );
  BUFFD1 U244 ( .I(DataI[8]), .Z(n197) );
  BUFFD1 U245 ( .I(DataI[3]), .Z(n192) );
  BUFFD1 U246 ( .I(DataI[4]), .Z(n193) );
  BUFFD1 U247 ( .I(DataI[11]), .Z(n200) );
  BUFFD1 U248 ( .I(DataI[6]), .Z(n195) );
  BUFFD1 U249 ( .I(DataI[9]), .Z(n198) );
  BUFFD1 U250 ( .I(DataI[0]), .Z(n189) );
  BUFFD1 U251 ( .I(DataI[5]), .Z(n194) );
  BUFFD1 U252 ( .I(DataI[12]), .Z(n201) );
  MUX4D0 U253 ( .I0(n8), .I1(n6), .I2(n7), .I3(n5), .S0(n172), .S1(n174), .Z(
        N80) );
  MUX4D0 U254 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n182), .S1(n177), .Z(n7)
         );
  MUX4D0 U255 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n186), .S1(n177), .Z(n6)
         );
  MUX4D0 U256 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n185), .S1(n177), .Z(n8)
         );
  MUX4D0 U257 ( .I0(n12), .I1(n10), .I2(n11), .I3(n9), .S0(n172), .S1(n174), 
        .Z(N79) );
  MUX4D0 U258 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n183), .S1(n177), .Z(n11)
         );
  MUX4D0 U259 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n185), .S1(n177), .Z(n10) );
  MUX4D0 U260 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n183), .S1(n177), .Z(n12)
         );
  MUX4D0 U261 ( .I0(n32), .I1(n30), .I2(n31), .I3(n29), .S0(n172), .S1(n174), 
        .Z(N74) );
  MUX4D0 U262 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n185), .S1(n176), .Z(n31)
         );
  MUX4D0 U263 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n185), .S1(n178), .Z(n30) );
  MUX4D0 U264 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n185), .S1(n177), .Z(n32)
         );
  MUX4D0 U265 ( .I0(n52), .I1(n50), .I2(n51), .I3(n49), .S0(n172), .S1(n174), 
        .Z(N69) );
  MUX4D0 U266 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n186), .S1(n178), .Z(n51) );
  MUX4D0 U267 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n186), .S1(N45), .Z(
        n50) );
  MUX4D0 U268 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n183), .S1(n179), .Z(n52) );
  MUX4D0 U269 ( .I0(n56), .I1(n54), .I2(n55), .I3(n53), .S0(n172), .S1(n174), 
        .Z(N68) );
  MUX4D0 U270 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n188), .S1(n181), .Z(n55) );
  MUX4D0 U271 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n183), .S1(n176), .Z(
        n54) );
  MUX4D0 U272 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n182), .S1(n177), .Z(n56) );
  MUX4D0 U273 ( .I0(n118), .I1(n116), .I2(n117), .I3(n115), .S0(n172), .S1(
        n174), .Z(N62) );
  MUX4D0 U274 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n186), .S1(N45), .Z(n117) );
  MUX4D0 U275 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n186), .S1(n176), .Z(
        n116) );
  MUX4D0 U276 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n186), .S1(n176), .Z(
        n118) );
  MUX4D0 U277 ( .I0(n122), .I1(n120), .I2(n121), .I3(n119), .S0(n172), .S1(
        n174), .Z(N61) );
  MUX4D0 U278 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n186), .S1(n176), .Z(
        n121) );
  MUX4D0 U279 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n186), .S1(N45), .Z(
        n120) );
  MUX4D0 U280 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n186), .S1(N45), .Z(n122) );
  MUX4D0 U281 ( .I0(n146), .I1(n144), .I2(n145), .I3(n143), .S0(N47), .S1(n318), .Z(N55) );
  MUX4D0 U282 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(N44), .S1(n179), .Z(n145) );
  MUX4D0 U283 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n188), .S1(n179), .Z(
        n144) );
  MUX4D0 U284 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(N44), .S1(n179), .Z(n146) );
  MUX4D0 U285 ( .I0(n150), .I1(n148), .I2(n149), .I3(n147), .S0(N47), .S1(n318), .Z(N54) );
  MUX4D0 U286 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n187), .S1(n180), .Z(
        n149) );
  MUX4D0 U287 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n187), .S1(n180), .Z(
        n148) );
  MUX4D0 U288 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n187), .S1(n180), .Z(
        n150) );
  MUX4D0 U289 ( .I0(n162), .I1(n160), .I2(n161), .I3(n159), .S0(N47), .S1(N46), 
        .Z(N51) );
  MUX4D0 U290 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n188), .S1(n181), .Z(
        n161) );
  MUX4D0 U291 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n188), .S1(n181), .Z(
        n160) );
  MUX4D0 U292 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n188), .S1(n181), .Z(
        n162) );
  MUX4D0 U293 ( .I0(n166), .I1(n164), .I2(n165), .I3(n163), .S0(N47), .S1(N46), 
        .Z(N50) );
  MUX4D0 U294 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n188), .S1(n181), .Z(
        n165) );
  MUX4D0 U295 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n188), .S1(n181), .Z(
        n164) );
  MUX4D0 U296 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n188), .S1(n181), .Z(
        n166) );
  MUX4D0 U297 ( .I0(n28), .I1(n26), .I2(n27), .I3(n25), .S0(n172), .S1(n174), 
        .Z(N75) );
  MUX4D0 U298 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(N44), .S1(n181), .Z(n27)
         );
  MUX4D0 U299 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n186), .S1(n179), .Z(n26) );
  MUX4D0 U300 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n183), .S1(n179), .Z(n28)
         );
  MUX4D0 U301 ( .I0(n106), .I1(n104), .I2(n105), .I3(n102), .S0(n172), .S1(
        n174), .Z(N65) );
  MUX4D0 U302 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n185), .S1(n178), .Z(
        n105) );
  MUX4D0 U303 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n185), .S1(n178), .Z(
        n104) );
  MUX4D0 U304 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n185), .S1(n180), .Z(
        n106) );
  MUX4D0 U305 ( .I0(n134), .I1(n132), .I2(n133), .I3(n131), .S0(N47), .S1(N46), 
        .Z(N58) );
  MUX4D0 U306 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n182), .S1(n178), .Z(
        n133) );
  MUX4D0 U307 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n182), .S1(n178), .Z(
        n132) );
  MUX4D0 U308 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n183), .S1(n178), .Z(
        n134) );
  MUX4D0 U309 ( .I0(n138), .I1(n136), .I2(n137), .I3(n135), .S0(N47), .S1(N46), 
        .Z(N57) );
  MUX4D0 U310 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n183), .S1(n179), .Z(
        n137) );
  MUX4D0 U311 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n188), .S1(n179), .Z(
        n136) );
  MUX4D0 U312 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(N44), .S1(n179), .Z(n138) );
  MUX4D0 U313 ( .I0(n4), .I1(n2), .I2(n3), .I3(n1), .S0(n172), .S1(n174), .Z(
        N81) );
  MUX4D0 U314 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n186), .S1(n177), .Z(n3)
         );
  MUX4D0 U315 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n185), .S1(n177), .Z(n2)
         );
  MUX4D0 U316 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n185), .S1(n177), .Z(n4)
         );
  MUX4D0 U317 ( .I0(n20), .I1(n18), .I2(n19), .I3(n17), .S0(n172), .S1(n174), 
        .Z(N77) );
  MUX4D0 U318 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n187), .S1(n175), .Z(n19)
         );
  MUX4D0 U319 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n187), .S1(n175), .Z(n18) );
  MUX4D0 U320 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n184), .S1(n175), .Z(n20)
         );
  MUX4D0 U321 ( .I0(n44), .I1(n42), .I2(n43), .I3(n41), .S0(n172), .S1(n174), 
        .Z(N71) );
  MUX4D0 U322 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n184), .S1(n181), .Z(n43) );
  MUX4D0 U323 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n184), .S1(n175), .Z(
        n42) );
  MUX4D0 U324 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n184), .S1(n179), .Z(n44) );
  MUX4D0 U325 ( .I0(n48), .I1(n46), .I2(n47), .I3(n45), .S0(n172), .S1(n174), 
        .Z(N70) );
  MUX4D0 U326 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n184), .S1(n181), .Z(n47) );
  MUX4D0 U327 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n184), .S1(n181), .Z(
        n46) );
  MUX4D0 U328 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n184), .S1(n176), .Z(n48) );
  MUX4D0 U329 ( .I0(n60), .I1(n58), .I2(n59), .I3(n57), .S0(n172), .S1(n174), 
        .Z(N67) );
  MUX4D0 U330 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n183), .S1(n177), .Z(n59) );
  MUX4D0 U331 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n188), .S1(n179), .Z(
        n58) );
  MUX4D0 U332 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n187), .S1(n177), .Z(n60) );
  MUX4D0 U333 ( .I0(n114), .I1(n112), .I2(n113), .I3(n111), .S0(n172), .S1(
        n174), .Z(N63) );
  MUX4D0 U334 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n186), .S1(n179), .Z(
        n113) );
  MUX4D0 U335 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n186), .S1(n176), .Z(
        n112) );
  MUX4D0 U336 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n186), .S1(n176), .Z(
        n114) );
  MUX4D0 U337 ( .I0(n126), .I1(n124), .I2(n125), .I3(n123), .S0(N47), .S1(N46), 
        .Z(N60) );
  MUX4D0 U338 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n183), .S1(n178), .Z(
        n125) );
  MUX4D0 U339 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n183), .S1(n178), .Z(
        n124) );
  MUX4D0 U340 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n187), .S1(n178), .Z(
        n126) );
  MUX4D0 U341 ( .I0(n142), .I1(n140), .I2(n141), .I3(n139), .S0(N47), .S1(n318), .Z(N56) );
  MUX4D0 U342 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n187), .S1(n179), .Z(
        n141) );
  MUX4D0 U343 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n183), .S1(n179), .Z(
        n140) );
  MUX4D0 U344 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(N44), .S1(n179), .Z(n142) );
  MUX4D0 U345 ( .I0(n154), .I1(n152), .I2(n153), .I3(n151), .S0(N47), .S1(n318), .Z(N53) );
  MUX4D0 U346 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n187), .S1(n180), .Z(
        n153) );
  MUX4D0 U347 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n187), .S1(n180), .Z(
        n152) );
  MUX4D0 U348 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n187), .S1(n180), .Z(
        n154) );
  MUX4D0 U349 ( .I0(n158), .I1(n156), .I2(n157), .I3(n155), .S0(N47), .S1(n318), .Z(N52) );
  MUX4D0 U350 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n187), .S1(n180), .Z(
        n157) );
  MUX4D0 U351 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n187), .S1(n180), .Z(
        n156) );
  MUX4D0 U352 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n187), .S1(n180), .Z(
        n158) );
  MUX4D0 U353 ( .I0(n24), .I1(n22), .I2(n23), .I3(n21), .S0(n172), .S1(n174), 
        .Z(N76) );
  MUX4D0 U354 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(N44), .S1(n175), .Z(n23)
         );
  MUX4D0 U355 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n183), .S1(n175), .Z(n22) );
  MUX4D0 U356 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n184), .S1(n175), .Z(n24)
         );
  MUX4D0 U357 ( .I0(n40), .I1(n38), .I2(n39), .I3(n37), .S0(n172), .S1(n174), 
        .Z(N72) );
  MUX4D0 U358 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n184), .S1(n180), .Z(n39)
         );
  MUX4D0 U359 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n184), .S1(n177), .Z(n38) );
  MUX4D0 U360 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n184), .S1(N45), .Z(n40)
         );
  MUX4D0 U361 ( .I0(n64), .I1(n62), .I2(n63), .I3(n61), .S0(n172), .S1(n174), 
        .Z(N66) );
  MUX4D0 U362 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n185), .S1(n177), .Z(n63) );
  MUX4D0 U363 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n185), .S1(n177), .Z(
        n62) );
  MUX4D0 U364 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n185), .S1(n177), .Z(n64) );
  MUX4D0 U365 ( .I0(n110), .I1(n108), .I2(n109), .I3(n107), .S0(n172), .S1(
        n174), .Z(N64) );
  MUX4D0 U366 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n185), .S1(N45), .Z(n109) );
  MUX4D0 U367 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n185), .S1(n178), .Z(
        n108) );
  MUX4D0 U368 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n185), .S1(N45), .Z(n110) );
  MUX4D0 U369 ( .I0(n130), .I1(n128), .I2(n129), .I3(n127), .S0(N47), .S1(N46), 
        .Z(N59) );
  MUX4D0 U370 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n183), .S1(n178), .Z(
        n129) );
  MUX4D0 U371 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n183), .S1(n178), .Z(
        n128) );
  MUX4D0 U372 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n183), .S1(n178), .Z(
        n130) );
  MUX4D0 U373 ( .I0(n170), .I1(n168), .I2(n169), .I3(n167), .S0(N47), .S1(N46), 
        .Z(N49) );
  MUX4D0 U374 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n188), .S1(n181), .Z(
        n169) );
  MUX4D0 U375 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n188), .S1(n181), .Z(
        n168) );
  MUX4D0 U376 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n188), .S1(n181), .Z(
        n170) );
  MUX4D0 U377 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n188), .S1(n181), .Z(
        n167) );
  MUX4D0 U378 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n183), .S1(n177), .Z(n1)
         );
  MUX4D0 U379 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n182), .S1(n177), .Z(n5)
         );
  MUX4D0 U380 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n183), .S1(n177), .Z(n9)
         );
  MUX4D0 U381 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n184), .S1(n175), .Z(n17) );
  MUX4D0 U382 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n188), .S1(n175), .Z(n21) );
  MUX4D0 U383 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n187), .S1(n179), .Z(n25) );
  MUX4D0 U384 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n185), .S1(n175), .Z(n29) );
  MUX4D0 U385 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n184), .S1(n181), .Z(n37) );
  MUX4D0 U386 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n184), .S1(n179), .Z(
        n41) );
  MUX4D0 U387 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n184), .S1(n178), .Z(
        n45) );
  MUX4D0 U388 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n182), .S1(n178), .Z(
        n49) );
  MUX4D0 U389 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n183), .S1(n176), .Z(
        n53) );
  MUX4D0 U390 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n182), .S1(n176), .Z(
        n57) );
  MUX4D0 U391 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n185), .S1(n175), .Z(
        n61) );
  MUX4D0 U392 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n185), .S1(n178), .Z(
        n102) );
  MUX4D0 U393 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n185), .S1(n181), .Z(
        n107) );
  MUX4D0 U394 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n186), .S1(n176), .Z(
        n111) );
  MUX4D0 U395 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n186), .S1(n176), .Z(
        n115) );
  MUX4D0 U396 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n186), .S1(n176), .Z(
        n119) );
  MUX4D0 U397 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n188), .S1(n178), .Z(
        n123) );
  MUX4D0 U398 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n183), .S1(n178), .Z(
        n127) );
  MUX4D0 U399 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n182), .S1(n178), .Z(
        n131) );
  MUX4D0 U400 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(N44), .S1(n179), .Z(
        n135) );
  MUX4D0 U401 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(N44), .S1(n179), .Z(
        n139) );
  MUX4D0 U402 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(N44), .S1(n179), .Z(
        n143) );
  MUX4D0 U403 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n187), .S1(n180), .Z(
        n147) );
  MUX4D0 U404 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n187), .S1(n180), .Z(
        n151) );
  MUX4D0 U405 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n187), .S1(n180), .Z(
        n155) );
  MUX4D0 U406 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n188), .S1(n181), .Z(
        n159) );
  MUX4D0 U407 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n188), .S1(n181), .Z(
        n163) );
  MUX4D0 U408 ( .I0(n36), .I1(n34), .I2(n35), .I3(n33), .S0(n172), .S1(n174), 
        .Z(N73) );
  MUX4D0 U409 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(N44), .S1(N45), .Z(n35) );
  MUX4D0 U410 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(N44), .S1(N45), .Z(n34)
         );
  MUX4D0 U411 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(N44), .S1(N45), .Z(n36) );
  MUX4D0 U412 ( .I0(n16), .I1(n14), .I2(n15), .I3(n13), .S0(N47), .S1(n318), 
        .Z(N78) );
  MUX4D0 U413 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n184), .S1(n180), .Z(n15)
         );
  MUX4D0 U414 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n184), .S1(n180), .Z(n14) );
  MUX4D0 U415 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n186), .S1(n181), .Z(n16)
         );
  MUX4D0 U416 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(N44), .S1(n180), .Z(n13)
         );
  MUX4D0 U417 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(N44), .S1(N45), .Z(n33)
         );
  ND2D1 U418 ( .A1(AddrW[1]), .A2(n376), .ZN(n383) );
  ND2D1 U419 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n386) );
  ND2D1 U420 ( .A1(n375), .A2(AddrW[0]), .ZN(n379) );
  ND2D1 U421 ( .A1(AddrW[2]), .A2(n377), .ZN(n384) );
  ND2D1 U422 ( .A1(AddrW[0]), .A2(n381), .ZN(n387) );
  INR2D1 U423 ( .A1(Write), .B1(AddrW[3]), .ZN(n375) );
  INVD1 U424 ( .I(AddrW[1]), .ZN(n377) );
  INVD1 U425 ( .I(AddrW[0]), .ZN(n380) );
  INVD1 U426 ( .I(AddrW[2]), .ZN(n376) );
  AN2D1 U427 ( .A1(Write), .A2(AddrW[3]), .Z(n381) );
  INR2D1 U428 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INR2D1 U429 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U430 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_1 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n4,
         n6, n9, n10, n11;

  AO211D1 U8 ( .A1(n10), .A2(n9), .B(N8), .C(N5), .Z(n6) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n11), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n11), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n4), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n4), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n11), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n11), .QN(n10) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n4), .QN(n11) );
  INVD1 U3 ( .I(Reset), .ZN(n4) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n10), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n9), .A2(n10), .B(n6), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n9) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_2 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n4,
         n6, n9, n10, n11;

  AO211D1 U8 ( .A1(n10), .A2(n9), .B(N8), .C(N5), .Z(n6) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n11), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n11), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n4), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n4), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n11), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n11), .QN(n10) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n4), .QN(n11) );
  INVD1 U3 ( .I(Reset), .ZN(n4) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n10), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n9), .A2(n10), .B(n6), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n9) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_3 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n4,
         n6, n9, n10, n11;

  AO211D1 U8 ( .A1(n10), .A2(n9), .B(N8), .C(N5), .Z(n6) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n11), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n11), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n4), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n4), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n11), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n11), .QN(n10) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n4), .QN(n11) );
  INVD1 U3 ( .I(Reset), .ZN(n4) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n10), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n9), .A2(n10), .B(n6), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n9) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_1 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_1_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_1_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_1_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n34), .CP(FastClock), .CDN(n2), .Q(ClockOut) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n32), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[4]), .QN(n14) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n33), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[1]), .QN(n30) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n31), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[0]), .QN(n28) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[3]), .QN(n23) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[5]), .QN(n9) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  AO222D0 U4 ( .A1(N27), .A2(n3), .B1(N35), .B2(n4), .C1(DivideFactor[0]), 
        .C2(n5), .Z(n31) );
  AO222D0 U5 ( .A1(N31), .A2(n3), .B1(N39), .B2(n4), .C1(DivideFactor[4]), 
        .C2(n5), .Z(n32) );
  AO222D0 U6 ( .A1(N28), .A2(n3), .B1(N36), .B2(n4), .C1(DivideFactor[1]), 
        .C2(n5), .Z(n33) );
  CKND0 U7 ( .CLK(N54), .CN(n5) );
  AN2D0 U8 ( .A1(n6), .A2(n7), .Z(n4) );
  AN3D0 U9 ( .A1(n8), .A2(n9), .A3(n10), .Z(n3) );
  CKXOR2D0 U10 ( .A1(ClockOut), .A2(n11), .Z(n34) );
  AO22D0 U11 ( .A1(N32), .A2(n10), .B1(N40), .B2(n6), .Z(N55) );
  MUX2ND0 U12 ( .I0(n12), .I1(n13), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U13 ( .A1(AdjustFreq[1]), .A2(n7), .ZN(n13) );
  ND3D0 U14 ( .A1(n14), .A2(n9), .A3(n15), .ZN(n7) );
  ND4D0 U15 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n15) );
  IND3D0 U16 ( .A1(AdjustFreq[1]), .B1(n9), .B2(n8), .ZN(n12) );
  CKND2D0 U17 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n8) );
  AO22D0 U18 ( .A1(N30), .A2(n10), .B1(N38), .B2(n6), .Z(N51) );
  AO22D0 U19 ( .A1(N29), .A2(n10), .B1(N37), .B2(n6), .Z(N49) );
  AN2D0 U20 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n6) );
  NR2D0 U21 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n10) );
  INR2D0 U22 ( .A1(N14), .B1(n11), .ZN(N21) );
  INR2D0 U23 ( .A1(N13), .B1(n11), .ZN(N20) );
  INR2D0 U24 ( .A1(N12), .B1(n11), .ZN(N19) );
  INR2D0 U25 ( .A1(N11), .B1(n11), .ZN(N18) );
  INR2D0 U26 ( .A1(N10), .B1(n11), .ZN(N17) );
  INR2D0 U27 ( .A1(N9), .B1(n11), .ZN(N16) );
  OA21D0 U28 ( .A1(FastDivvy[5]), .A2(n9), .B(n16), .Z(n11) );
  IOA22D0 U29 ( .B1(n20), .B2(n22), .A1(n9), .A2(FastDivvy[5]), .ZN(n16) );
  AOI221D0 U30 ( .A1(FastDivvy[4]), .A2(n14), .B1(FastDivvy[3]), .B2(n23), .C(
        n24), .ZN(n22) );
  AOI221D0 U31 ( .A1(DivideFactor[3]), .A2(n25), .B1(DivideFactor[2]), .B2(n26), .C(n27), .ZN(n24) );
  IAO21D0 U32 ( .A1(n26), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n27) );
  OAI32D0 U33 ( .A1(n28), .A2(FastDivvy[0]), .A3(n29), .B1(FastDivvy[1]), .B2(
        n30), .ZN(n26) );
  AN2D0 U34 ( .A1(FastDivvy[1]), .A2(n30), .Z(n29) );
  CKND0 U35 ( .CLK(FastDivvy[3]), .CN(n25) );
  NR2D0 U36 ( .A1(FastDivvy[4]), .A2(n14), .ZN(n20) );
  CKND0 U37 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U38 ( .A1(WireD[5]), .A2(n2), .ZN(WireD[0]) );
endmodule


module VFO_2 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_2_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_2_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_2_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n1), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n33), .CP(FastClock), .CDN(n1), .Q(ClockOut) );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n1), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n1), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n31), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[4]), .QN(n13) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n32), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[1]), .QN(n29) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n30), .CP(Sample), .SDN(n1), .Q(
        DivideFactor[0]), .QN(n27) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n1), .Q(
        DivideFactor[3]), .QN(n22) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
  AO222D0 U4 ( .A1(N27), .A2(n2), .B1(N35), .B2(n3), .C1(DivideFactor[0]), 
        .C2(n4), .Z(n30) );
  AO222D0 U5 ( .A1(N31), .A2(n2), .B1(N39), .B2(n3), .C1(DivideFactor[4]), 
        .C2(n4), .Z(n31) );
  AO222D0 U6 ( .A1(N28), .A2(n2), .B1(N36), .B2(n3), .C1(DivideFactor[1]), 
        .C2(n4), .Z(n32) );
  CKND0 U7 ( .CLK(N54), .CN(n4) );
  AN2D0 U8 ( .A1(n5), .A2(n6), .Z(n3) );
  AN3D0 U9 ( .A1(n7), .A2(n8), .A3(n9), .Z(n2) );
  CKXOR2D0 U10 ( .A1(ClockOut), .A2(n10), .Z(n33) );
  AO22D0 U11 ( .A1(N32), .A2(n9), .B1(N40), .B2(n5), .Z(N55) );
  MUX2ND0 U12 ( .I0(n11), .I1(n12), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U13 ( .A1(AdjustFreq[1]), .A2(n6), .ZN(n12) );
  ND3D0 U14 ( .A1(n13), .A2(n8), .A3(n14), .ZN(n6) );
  ND4D0 U15 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n14) );
  IND3D0 U16 ( .A1(AdjustFreq[1]), .B1(n8), .B2(n7), .ZN(n11) );
  CKND2D0 U17 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n7) );
  AO22D0 U18 ( .A1(N30), .A2(n9), .B1(N38), .B2(n5), .Z(N51) );
  AO22D0 U19 ( .A1(N29), .A2(n9), .B1(N37), .B2(n5), .Z(N49) );
  AN2D0 U20 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n5) );
  NR2D0 U21 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n9) );
  INR2D0 U22 ( .A1(N14), .B1(n10), .ZN(N21) );
  INR2D0 U23 ( .A1(N13), .B1(n10), .ZN(N20) );
  INR2D0 U24 ( .A1(N12), .B1(n10), .ZN(N19) );
  INR2D0 U25 ( .A1(N11), .B1(n10), .ZN(N18) );
  INR2D0 U26 ( .A1(N10), .B1(n10), .ZN(N17) );
  INR2D0 U27 ( .A1(N9), .B1(n10), .ZN(N16) );
  OA21D0 U28 ( .A1(FastDivvy[5]), .A2(n8), .B(n15), .Z(n10) );
  IOA22D0 U29 ( .B1(n16), .B2(n20), .A1(n8), .A2(FastDivvy[5]), .ZN(n15) );
  AOI221D0 U30 ( .A1(FastDivvy[4]), .A2(n13), .B1(FastDivvy[3]), .B2(n22), .C(
        n23), .ZN(n20) );
  AOI221D0 U31 ( .A1(DivideFactor[3]), .A2(n24), .B1(DivideFactor[2]), .B2(n25), .C(n26), .ZN(n23) );
  IAO21D0 U32 ( .A1(n25), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n26) );
  OAI32D0 U33 ( .A1(n27), .A2(FastDivvy[0]), .A3(n28), .B1(FastDivvy[1]), .B2(
        n29), .ZN(n25) );
  AN2D0 U34 ( .A1(FastDivvy[1]), .A2(n29), .Z(n28) );
  CKND0 U35 ( .CLK(FastDivvy[3]), .CN(n24) );
  NR2D0 U36 ( .A1(FastDivvy[4]), .A2(n13), .ZN(n16) );
  CKND0 U37 ( .CLK(DivideFactor[5]), .CN(n8) );
  CKND0 U38 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U39 ( .A1(WireD[5]), .A2(n1), .ZN(WireD[0]) );
endmodule


module VFO_3 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_3_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_3_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_3_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n34), .CP(FastClock), .CDN(n2), .Q(ClockOut) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[3]), .QN(n23) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n2), .Q(
        DivideFactor[5]), .QN(n9) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n32), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[4]), .QN(n14) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n33), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[1]), .QN(n30) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n31), .CP(Sample), .SDN(n2), .Q(
        DivideFactor[0]), .QN(n28) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  AO222D0 U4 ( .A1(N27), .A2(n3), .B1(N35), .B2(n4), .C1(DivideFactor[0]), 
        .C2(n5), .Z(n31) );
  AO222D0 U5 ( .A1(N31), .A2(n3), .B1(N39), .B2(n4), .C1(DivideFactor[4]), 
        .C2(n5), .Z(n32) );
  AO222D0 U6 ( .A1(N28), .A2(n3), .B1(N36), .B2(n4), .C1(DivideFactor[1]), 
        .C2(n5), .Z(n33) );
  CKND0 U7 ( .CLK(N54), .CN(n5) );
  AN2D0 U8 ( .A1(n6), .A2(n7), .Z(n4) );
  AN3D0 U9 ( .A1(n8), .A2(n9), .A3(n10), .Z(n3) );
  CKXOR2D0 U10 ( .A1(ClockOut), .A2(n11), .Z(n34) );
  AO22D0 U11 ( .A1(N32), .A2(n10), .B1(N40), .B2(n6), .Z(N55) );
  MUX2ND0 U12 ( .I0(n12), .I1(n13), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U13 ( .A1(AdjustFreq[1]), .A2(n7), .ZN(n13) );
  ND3D0 U14 ( .A1(n14), .A2(n9), .A3(n15), .ZN(n7) );
  ND4D0 U15 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n15) );
  IND3D0 U16 ( .A1(AdjustFreq[1]), .B1(n9), .B2(n8), .ZN(n12) );
  CKND2D0 U17 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n8) );
  AO22D0 U18 ( .A1(N30), .A2(n10), .B1(N38), .B2(n6), .Z(N51) );
  AO22D0 U19 ( .A1(N29), .A2(n10), .B1(N37), .B2(n6), .Z(N49) );
  AN2D0 U20 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n6) );
  NR2D0 U21 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n10) );
  INR2D0 U22 ( .A1(N14), .B1(n11), .ZN(N21) );
  INR2D0 U23 ( .A1(N13), .B1(n11), .ZN(N20) );
  INR2D0 U24 ( .A1(N12), .B1(n11), .ZN(N19) );
  INR2D0 U25 ( .A1(N11), .B1(n11), .ZN(N18) );
  INR2D0 U26 ( .A1(N10), .B1(n11), .ZN(N17) );
  INR2D0 U27 ( .A1(N9), .B1(n11), .ZN(N16) );
  OA21D0 U28 ( .A1(FastDivvy[5]), .A2(n9), .B(n16), .Z(n11) );
  IOA22D0 U29 ( .B1(n20), .B2(n22), .A1(n9), .A2(FastDivvy[5]), .ZN(n16) );
  AOI221D0 U30 ( .A1(FastDivvy[4]), .A2(n14), .B1(FastDivvy[3]), .B2(n23), .C(
        n24), .ZN(n22) );
  AOI221D0 U31 ( .A1(DivideFactor[3]), .A2(n25), .B1(DivideFactor[2]), .B2(n26), .C(n27), .ZN(n24) );
  IAO21D0 U32 ( .A1(n26), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n27) );
  OAI32D0 U33 ( .A1(n28), .A2(FastDivvy[0]), .A3(n29), .B1(FastDivvy[1]), .B2(
        n30), .ZN(n26) );
  AN2D0 U34 ( .A1(FastDivvy[1]), .A2(n30), .Z(n29) );
  CKND0 U35 ( .CLK(FastDivvy[3]), .CN(n25) );
  NR2D0 U36 ( .A1(FastDivvy[4]), .A2(n14), .ZN(n20) );
  CKND0 U37 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U38 ( .A1(WireD[5]), .A2(n2), .ZN(WireD[0]) );
endmodule


module MultiCounter_1 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_1_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_2 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_2_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_3 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_3_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n2, \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D1 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(n2) );
  BUFFD0 U2 ( .I(n2), .Z(SUM[4]) );
  CKND0 U3 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_2_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_3_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n2, \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D1 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(n2) );
  BUFFD0 U2 ( .I(n2), .Z(SUM[4]) );
  CKND0 U3 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

