

`ifndef RKV_I2C_CGM_SV
`define RKV_I2C_CGM_SV

// Coverage Model
class rkv_i2c_cgm extends uvm_component;
   
  // TODO
  // Covergroup definition below

  // Analysis import declarion below

  `uvm_component_utils(rkv_i2c_cgm)

  function new(string name = "rkv_i2c_cgm", uvm_component parent = null);
    super.new(name, parent);
  endfunction

endclass


`endif // RKV_I2C_CGM_SV
