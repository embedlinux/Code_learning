`ifndef __MY_TEST__SV__
`define __MY_TEST__SV__

class my_test extends uvm_test;

	`uvm_component_utils(my_test)

	my_env m_env;

	function new(string name = "", uvm_component parent);
		super.new(name, parent);
	endfunction : new


	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		m_env = my_env::type_id::create("m_env", this);
		uvm_config_db#(uvm_object_wrapper)::set(this, "*.m_seqr.run_phase",
								"default_sequence", my_sequence::get_type());
	endfunction : build_phase


	virtual function void start_of_simulation_phase(uvm_phase phase);
		super.start_of_simulation_phase(phase);
		uvm_top.print_topology(uvm_default_table_printer);
	endfunction : start_of_simulation_phase


endclass : my_test

`endif // __MY_TEST__SV__
