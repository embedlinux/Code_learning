
module FIFO_Top ( Dout, Din, ReadIn, WriteIn, Clocker, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, Clocker, Reseter;
  wire   E_FIFO, F_FIFO, ReadWire, WriteWire, _0_net_, n4, n5, Mem_Enable, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38;
  wire   [4:0] SM_MemAddr;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(E_FIFO), .FullFIFO(F_FIFO), .ReadCmd(ReadWire), .WriteCmd(
        WriteWire), .ReadReq(ReadIn), .WriteReq(WriteIn), .Clk(Clocker), 
        .Reset(n6) );
  Mem1kx32 RegFile1 ( .DataO(Dout), .DataI({n38, n37, n36, n35, n34, n33, n32, 
        n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, n18, 
        n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, n7}), .Addr(SM_MemAddr), .ClockIn(_0_net_), .ChipEna(Mem_Enable), .Read(ReadWire), .Write(WriteWire)
         );
  AOI211D1 U10 ( .A1(WriteWire), .A2(ReadWire), .B(F_FIFO), .C(E_FIFO), .ZN(
        Mem_Enable) );
  INR2D1 U11 ( .A1(ReadWire), .B1(WriteWire), .ZN(n5) );
  INVD1 U12 ( .I(n5), .ZN(n4) );
  BUFFD1 U13 ( .I(Din[10]), .Z(n17) );
  BUFFD1 U14 ( .I(Din[11]), .Z(n18) );
  BUFFD1 U15 ( .I(Din[12]), .Z(n19) );
  BUFFD1 U16 ( .I(Din[13]), .Z(n20) );
  BUFFD1 U17 ( .I(Din[14]), .Z(n21) );
  BUFFD1 U18 ( .I(Din[15]), .Z(n22) );
  BUFFD1 U19 ( .I(Din[16]), .Z(n23) );
  BUFFD1 U20 ( .I(Din[17]), .Z(n24) );
  BUFFD1 U21 ( .I(Din[18]), .Z(n25) );
  BUFFD1 U22 ( .I(Din[19]), .Z(n26) );
  BUFFD1 U23 ( .I(Din[20]), .Z(n27) );
  BUFFD1 U24 ( .I(Din[21]), .Z(n28) );
  BUFFD1 U25 ( .I(Din[22]), .Z(n29) );
  BUFFD1 U26 ( .I(Din[23]), .Z(n30) );
  BUFFD1 U27 ( .I(Din[24]), .Z(n31) );
  BUFFD1 U28 ( .I(Din[25]), .Z(n32) );
  BUFFD1 U29 ( .I(Din[26]), .Z(n33) );
  BUFFD1 U30 ( .I(Din[27]), .Z(n34) );
  BUFFD1 U31 ( .I(Din[28]), .Z(n35) );
  BUFFD1 U32 ( .I(Din[29]), .Z(n36) );
  BUFFD1 U33 ( .I(Din[30]), .Z(n37) );
  BUFFD1 U34 ( .I(Din[31]), .Z(n38) );
  BUFFD1 U35 ( .I(Din[0]), .Z(n7) );
  BUFFD1 U36 ( .I(Din[1]), .Z(n8) );
  BUFFD1 U37 ( .I(Din[2]), .Z(n9) );
  BUFFD1 U38 ( .I(Din[3]), .Z(n10) );
  BUFFD1 U39 ( .I(Din[4]), .Z(n11) );
  BUFFD1 U40 ( .I(Din[5]), .Z(n12) );
  BUFFD1 U41 ( .I(Din[6]), .Z(n13) );
  BUFFD1 U42 ( .I(Din[7]), .Z(n14) );
  BUFFD1 U43 ( .I(Din[8]), .Z(n15) );
  BUFFD1 U44 ( .I(Din[9]), .Z(n16) );
  AO22D0 U45 ( .A1(SM_WriteAddr[0]), .A2(n4), .B1(SM_ReadAddr[0]), .B2(n5), 
        .Z(SM_MemAddr[0]) );
  AO22D0 U46 ( .A1(SM_WriteAddr[2]), .A2(n4), .B1(SM_ReadAddr[2]), .B2(n5), 
        .Z(SM_MemAddr[2]) );
  AO22D0 U47 ( .A1(SM_WriteAddr[1]), .A2(n4), .B1(SM_ReadAddr[1]), .B2(n5), 
        .Z(SM_MemAddr[1]) );
  AO22D0 U48 ( .A1(SM_WriteAddr[3]), .A2(n4), .B1(SM_ReadAddr[3]), .B2(n5), 
        .Z(SM_MemAddr[3]) );
  AO22D0 U49 ( .A1(SM_WriteAddr[4]), .A2(n4), .B1(SM_ReadAddr[4]), .B2(n5), 
        .Z(SM_MemAddr[4]) );
  BUFFD1 U50 ( .I(Reseter), .Z(n6) );
  INVD1 U51 ( .I(Clocker), .ZN(_0_net_) );
endmodule


module FIFOStateM ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, Clk, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, Clk, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N72, N73, N74, N75, N76, N88, N89, N90, N91, N92,
         N93, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N144, N146, N148, N150, N152, N155,
         N158, N161, N164, N167, N169, N172, N175, N178, N181, N184, N186,
         N187, N190, N191, N200, N201, N202, N211, N212, N213, N214, N217,
         N220, N223, N226, N229, N232, N235, N238, N241, n2, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n73, n74, n75, n76;
  wire   [2:0] CurState;
  wire   [2:0] NextState;

  LHQD1 \WriteCount_tri_enable_reg[0]  ( .E(N200), .D(N201), .Q(N9) );
  LHQD1 \NextState_reg[0]  ( .E(N190), .D(N144), .Q(NextState[0]) );
  LHQD1 \WriteCount_reg[1]  ( .E(N200), .D(N155), .Q(N238) );
  LHQD1 \ReadCount_reg[1]  ( .E(N211), .D(N172), .Q(N223) );
  LHQD1 \NextState_reg[1]  ( .E(N190), .D(N146), .Q(NextState[1]) );
  LHQD1 \NextState_reg[2]  ( .E(N190), .D(N148), .Q(NextState[2]) );
  LHQD1 WriteCmdReg_reg ( .E(N202), .D(N167), .Q(WriteCmd) );
  LHQD1 FullFIFOReg_reg ( .E(N191), .D(N150), .Q(FullFIFO) );
  LHQD1 \WriteCount_tri_enable_reg[4]  ( .E(N200), .D(N201), .Q(N5) );
  LHQD1 \WriteCount_tri_enable_reg[2]  ( .E(N200), .D(N201), .Q(N7) );
  LHQD1 \WriteCount_tri_enable_reg[1]  ( .E(N200), .D(N201), .Q(N8) );
  LHQD1 \WriteCount_tri_enable_reg[3]  ( .E(N200), .D(N201), .Q(N6) );
  LHQD1 \ReadCount_tri_enable_reg[4]  ( .E(N211), .D(N212), .Q(N0) );
  LHQD1 \ReadCount_tri_enable_reg[2]  ( .E(N211), .D(N212), .Q(N2) );
  LHQD1 \ReadCount_tri_enable_reg[0]  ( .E(N211), .D(N212), .Q(N4) );
  LHQD1 \ReadCount_tri_enable_reg[1]  ( .E(N211), .D(N212), .Q(N3) );
  LHQD1 \ReadCount_tri_enable_reg[3]  ( .E(N211), .D(N212), .Q(N1) );
  LHQD1 \ReadCount_reg[0]  ( .E(N211), .D(N169), .Q(N226) );
  LHQD1 \ReadCount_reg[4]  ( .E(N211), .D(N181), .Q(N214) );
  LHQD1 \WriteCount_reg[4]  ( .E(N200), .D(N164), .Q(N229) );
  LHQD1 \WriteCount_reg[3]  ( .E(N200), .D(N161), .Q(N232) );
  LHQD1 \WriteCount_reg[2]  ( .E(N200), .D(N158), .Q(N235) );
  LHQD1 \ReadCount_reg[2]  ( .E(N211), .D(N175), .Q(N220) );
  LHQD1 \ReadCount_reg[3]  ( .E(N211), .D(N178), .Q(N217) );
  LHQD1 \WriteCount_reg[0]  ( .E(N200), .D(N152), .Q(N241) );
  BUFTD1 \WriteCount_tri[0]  ( .I(N241), .OE(n70), .Z(WriteAddr[0]) );
  BUFTD1 \WriteCount_tri[1]  ( .I(N238), .OE(n69), .Z(WriteAddr[1]) );
  BUFTD1 \WriteCount_tri[2]  ( .I(N235), .OE(n68), .Z(WriteAddr[2]) );
  BUFTD1 \WriteCount_tri[3]  ( .I(N232), .OE(n67), .Z(WriteAddr[3]) );
  BUFTD1 \WriteCount_tri[4]  ( .I(N229), .OE(n66), .Z(WriteAddr[4]) );
  BUFTD1 \ReadCount_tri[0]  ( .I(N226), .OE(n65), .Z(ReadAddr[0]) );
  BUFTD1 \ReadCount_tri[1]  ( .I(N223), .OE(n64), .Z(ReadAddr[1]) );
  BUFTD1 \ReadCount_tri[2]  ( .I(N220), .OE(n63), .Z(ReadAddr[2]) );
  BUFTD1 \ReadCount_tri[3]  ( .I(N217), .OE(n62), .Z(ReadAddr[3]) );
  BUFTD1 \ReadCount_tri[4]  ( .I(N214), .OE(n61), .Z(ReadAddr[4]) );
  MOAI22D1 U25 ( .A1(Clk), .A2(n26), .B1(n20), .B2(N213), .ZN(N200) );
  OA21D1 U27 ( .A1(n29), .A2(n21), .B(n30), .Z(n26) );
  AO222D1 U60 ( .A1(ReadAddr[4]), .A2(n33), .B1(N54), .B2(n43), .C1(N76), .C2(
        n52), .Z(N164) );
  AO222D1 U61 ( .A1(ReadAddr[3]), .A2(n33), .B1(N53), .B2(n43), .C1(N75), .C2(
        n52), .Z(N161) );
  AO222D1 U62 ( .A1(ReadAddr[2]), .A2(n33), .B1(N52), .B2(n43), .C1(N74), .C2(
        n52), .Z(N158) );
  AO222D1 U63 ( .A1(ReadAddr[1]), .A2(n33), .B1(N51), .B2(n43), .C1(N73), .C2(
        n52), .Z(N155) );
  AO222D1 U64 ( .A1(ReadAddr[0]), .A2(n33), .B1(N50), .B2(n43), .C1(N72), .C2(
        n52), .Z(N152) );
  FIFOStateM_DW01_inc_0 add_211 ( .A({n2, N105, N104, N103, N102, N101}), 
        .SUM({N111, N110, N109, N108, N107, N106}) );
  FIFOStateM_DW01_inc_1 add_199 ( .A({n2, N76, N75, N74, N73, N72}), .SUM({N93, 
        N92, N91, N90, N89, N88}) );
  FIFOStateM_DW01_inc_2 add_111_C148 ( .A({N45, N46, N47, N48, N49}), .SUM({
        N54, N53, N52, N51, N50}) );
  FIFOStateM_DW01_inc_3 r109 ( .A(ReadAddr), .SUM({N105, N104, N103, N102, 
        N101}) );
  FIFOStateM_DW01_inc_4 r106 ( .A(WriteAddr), .SUM({N76, N75, N74, N73, N72})
         );
  LHQD2 ReadCmdReg_reg ( .E(N187), .D(N186), .Q(ReadCmd) );
  LHD1 EmptyFIFOReg_reg ( .E(N213), .D(N184), .Q(EmptyFIFO) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(Clk), .CDN(n71), .Q(n58), 
        .QN(n72) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(Clk), .CDN(n71), .Q(
        CurState[2]), .QN(n36) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(Clk), .CDN(n71), .Q(
        CurState[0]), .QN(n41) );
  AOI21D1 U3 ( .A1(ReadAddr[1]), .A2(n7), .B(n8), .ZN(n9) );
  IAO21D1 U4 ( .A1(N107), .A2(n15), .B(n17), .ZN(n18) );
  NR3D0 U5 ( .A1(n41), .A2(n72), .A3(n36), .ZN(n33) );
  NR3D0 U6 ( .A1(CurState[0]), .A2(CurState[2]), .A3(n58), .ZN(n32) );
  INVD1 U7 ( .I(n43), .ZN(n51) );
  INVD1 U8 ( .I(n47), .ZN(n42) );
  NR2D1 U9 ( .A1(n27), .A2(n21), .ZN(n43) );
  OAI21D1 U10 ( .A1(n47), .A2(n46), .B(n51), .ZN(N167) );
  NR2D1 U11 ( .A1(n54), .A2(n46), .ZN(N150) );
  INVD1 U12 ( .I(n25), .ZN(N186) );
  INVD1 U13 ( .I(n53), .ZN(n52) );
  INVD1 U14 ( .I(n50), .ZN(n31) );
  NR2D1 U15 ( .A1(n52), .A2(n50), .ZN(n47) );
  INVD1 U16 ( .I(n38), .ZN(n48) );
  INVD1 U17 ( .I(n23), .ZN(N211) );
  INVD1 U18 ( .I(n39), .ZN(n46) );
  AOI21D1 U19 ( .A1(n42), .A2(n46), .B(n33), .ZN(n25) );
  INVD1 U20 ( .I(n20), .ZN(n21) );
  OAI221D0 U21 ( .A1(n46), .A2(n53), .B1(N112), .B2(n29), .C(n59), .ZN(N144)
         );
  NR2D1 U22 ( .A1(n33), .A2(n50), .ZN(n59) );
  OAI21D1 U23 ( .A1(n46), .A2(n55), .B(n54), .ZN(N148) );
  AOI21D1 U24 ( .A1(N95), .A2(n49), .B(n50), .ZN(n55) );
  NR2D1 U26 ( .A1(n27), .A2(n20), .ZN(N184) );
  ND3D1 U28 ( .A1(n51), .A2(n31), .A3(n56), .ZN(N146) );
  AOI22D0 U29 ( .A1(n49), .A2(n57), .B1(n40), .B2(n39), .ZN(n56) );
  ND2D1 U30 ( .A1(N95), .A2(n39), .ZN(n57) );
  NR3D0 U31 ( .A1(n41), .A2(n58), .A3(n36), .ZN(n50) );
  INVD1 U32 ( .I(n32), .ZN(n27) );
  INVD1 U33 ( .I(n49), .ZN(n29) );
  NR2D1 U34 ( .A1(n40), .A2(n49), .ZN(n53) );
  INVD1 U35 ( .I(n33), .ZN(n54) );
  AN2D1 U36 ( .A1(N150), .A2(n22), .Z(N201) );
  AN2D1 U37 ( .A1(N184), .A2(n22), .Z(N212) );
  AO22D0 U38 ( .A1(n32), .A2(N45), .B1(N105), .B2(n48), .Z(N181) );
  AO22D0 U39 ( .A1(n32), .A2(N49), .B1(N101), .B2(n48), .Z(N169) );
  AO22D0 U40 ( .A1(n32), .A2(N48), .B1(N102), .B2(n48), .Z(N172) );
  AO22D0 U41 ( .A1(n32), .A2(N46), .B1(N104), .B2(n48), .Z(N178) );
  AO22D0 U42 ( .A1(n32), .A2(N47), .B1(N103), .B2(n48), .Z(N175) );
  INVD1 U43 ( .I(Reset), .ZN(n71) );
  NR3D0 U44 ( .A1(n33), .A2(n49), .A3(n50), .ZN(n38) );
  AOI221D0 U45 ( .A1(n42), .A2(n20), .B1(Reset), .B2(n32), .C(n43), .ZN(n24)
         );
  OAI21D1 U46 ( .A1(n45), .A2(n32), .B(n22), .ZN(n23) );
  NR2D1 U47 ( .A1(n38), .A2(n39), .ZN(n45) );
  AOI21D1 U48 ( .A1(Reset), .A2(n32), .B(n33), .ZN(n30) );
  INVD1 U49 ( .I(n40), .ZN(n28) );
  ND2D1 U50 ( .A1(ReadReq), .A2(n60), .ZN(n39) );
  AO22D0 U51 ( .A1(n20), .A2(N73), .B1(n21), .B2(WriteAddr[1]), .Z(N99) );
  INVD1 U52 ( .I(WriteReq), .ZN(n60) );
  AO22D0 U53 ( .A1(n21), .A2(WriteAddr[0]), .B1(n20), .B2(N72), .Z(N100) );
  XNR2D1 U54 ( .A1(n3), .A2(N109), .ZN(n73) );
  AOI22D0 U55 ( .A1(n20), .A2(N75), .B1(n21), .B2(WriteAddr[3]), .ZN(n3) );
  XNR2D1 U56 ( .A1(n4), .A2(N108), .ZN(n74) );
  AOI22D0 U57 ( .A1(n20), .A2(N74), .B1(n21), .B2(WriteAddr[2]), .ZN(n4) );
  AO22D0 U58 ( .A1(n20), .A2(N76), .B1(n21), .B2(WriteAddr[4]), .Z(N96) );
  NR2D1 U59 ( .A1(n60), .A2(ReadReq), .ZN(n20) );
  NR3D0 U65 ( .A1(CurState[2]), .A2(n72), .A3(n41), .ZN(n49) );
  NR3D0 U66 ( .A1(CurState[2]), .A2(n72), .A3(CurState[0]), .ZN(n40) );
  INVD1 U67 ( .I(Clk), .ZN(n22) );
  INVD1 U68 ( .I(N7), .ZN(n68) );
  INVD1 U69 ( .I(N8), .ZN(n69) );
  INVD1 U70 ( .I(N9), .ZN(n70) );
  INR2D1 U71 ( .A1(WriteAddr[1]), .B1(Reset), .ZN(N48) );
  INR2D1 U72 ( .A1(WriteAddr[2]), .B1(Reset), .ZN(N47) );
  INR2D1 U73 ( .A1(WriteAddr[3]), .B1(Reset), .ZN(N46) );
  INR2D1 U74 ( .A1(WriteAddr[4]), .B1(Reset), .ZN(N45) );
  AN2D1 U75 ( .A1(WriteAddr[0]), .A2(n71), .Z(N49) );
  INVD1 U76 ( .I(N0), .ZN(n61) );
  INVD1 U77 ( .I(N1), .ZN(n62) );
  INVD1 U78 ( .I(N2), .ZN(n63) );
  INVD1 U79 ( .I(N3), .ZN(n64) );
  INVD1 U80 ( .I(N4), .ZN(n65) );
  INVD1 U81 ( .I(N5), .ZN(n66) );
  INVD1 U82 ( .I(N6), .ZN(n67) );
  AOI31D0 U83 ( .A1(n24), .A2(n34), .A3(n35), .B(Clk), .ZN(N190) );
  ND2D1 U84 ( .A1(CurState[2]), .A2(n41), .ZN(n34) );
  AOI31D0 U85 ( .A1(n72), .A2(n36), .A3(CurState[0]), .B(n37), .ZN(n35) );
  AOI21D1 U86 ( .A1(n38), .A2(n28), .B(n39), .ZN(n37) );
  AOI21D1 U87 ( .A1(n27), .A2(n28), .B(Clk), .ZN(N213) );
  OAI21D1 U88 ( .A1(Clk), .A2(n44), .B(n23), .ZN(N187) );
  AOI22D0 U89 ( .A1(n20), .A2(n42), .B1(n40), .B2(n46), .ZN(n44) );
  AOI21D1 U90 ( .A1(n30), .A2(n31), .B(Clk), .ZN(N191) );
  AOI21D1 U91 ( .A1(n24), .A2(n25), .B(Clk), .ZN(N202) );
  TIEL U92 ( .ZN(n2) );
  INR2D0 U93 ( .A1(N88), .B1(ReadAddr[0]), .ZN(n6) );
  CKND0 U94 ( .CLK(ReadAddr[1]), .CN(n5) );
  OAI22D0 U95 ( .A1(n6), .A2(n5), .B1(N89), .B2(n6), .ZN(n10) );
  INR2D0 U96 ( .A1(ReadAddr[0]), .B1(N88), .ZN(n8) );
  CKND0 U97 ( .CLK(N89), .CN(n7) );
  IND3D0 U98 ( .A1(N93), .B1(n10), .B2(n9), .ZN(n14) );
  CKXOR2D0 U99 ( .A1(N92), .A2(ReadAddr[4]), .Z(n13) );
  CKXOR2D0 U100 ( .A1(N90), .A2(ReadAddr[2]), .Z(n12) );
  CKXOR2D0 U101 ( .A1(N91), .A2(ReadAddr[3]), .Z(n11) );
  NR4D0 U102 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(N95) );
  INR2D0 U103 ( .A1(N106), .B1(N100), .ZN(n16) );
  CKND0 U104 ( .CLK(N99), .CN(n15) );
  OAI22D0 U105 ( .A1(N107), .A2(n16), .B1(n16), .B2(n15), .ZN(n19) );
  INR2D0 U106 ( .A1(N100), .B1(N106), .ZN(n17) );
  IND3D0 U107 ( .A1(N111), .B1(n19), .B2(n18), .ZN(n76) );
  CKXOR2D0 U108 ( .A1(N96), .A2(N110), .Z(n75) );
  NR4D0 U109 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(N112) );
endmodule


module Mem1kx32 ( Dready, ParityErr, DataO, DataI, Addr, ClockIn, ChipEna, 
        Read, Write );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] Addr;
  input ClockIn, ChipEna, Read, Write;
  output Dready, ParityErr;
  wire   N43, N44, N45, N46, N47, ChipClock, DreadyReg, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N84, N2262, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103, n105,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n102, n104, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762;
  wire   [31:0] DataOreg;
  assign N43 = Addr[0];
  assign N44 = Addr[1];
  assign N45 = Addr[2];
  assign N46 = Addr[3];
  assign N47 = Addr[4];

  XNR4D1 U10 ( .A1(n742), .A2(n739), .A3(n748), .A4(n745), .ZN(n77) );
  XOR4D1 U11 ( .A1(n754), .A2(n751), .A3(n760), .A4(n757), .Z(n76) );
  XOR4D1 U12 ( .A1(n730), .A2(n727), .A3(n736), .A4(n733), .Z(n73) );
  XOR4D1 U13 ( .A1(n709), .A2(n706), .A3(n715), .A4(n712), .Z(n70) );
  XNR4D1 U14 ( .A1(n688), .A2(n685), .A3(n694), .A4(n691), .ZN(n67) );
  XOR4D1 U18 ( .A1(n82), .A2(N71), .A3(n83), .A4(N74), .Z(n81) );
  XNR4D1 U19 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n83) );
  XNR4D1 U24 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n89) );
  XOR4D1 U25 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n88) );
  XNR4D1 U26 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .ZN(n85) );
  XNR4D1 U27 ( .A1(N79), .A2(N77), .A3(N81), .A4(N80), .ZN(n79) );
  AN2D2 U81 ( .A1(ClockIn), .A2(ChipEna), .Z(ChipClock) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOreg[1]), .OE(n659), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOreg[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOreg[21]), .OE(n659), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOreg[20]), .OE(n659), .Z(DataO[20]) );
  EDFQD1 DreadyReg_reg ( .D(Read), .E(ChipEna), .CP(ChipClock), .Q(DreadyReg)
         );
  EDFQD1 \DataOreg_reg[9]  ( .D(N72), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[9]) );
  EDFQD1 \Storage_reg[26][10]  ( .D(n698), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][10] ) );
  EDFQD1 \Storage_reg[26][9]  ( .D(DataI[9]), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][9] ) );
  EDFQD1 \Storage_reg[26][8]  ( .D(n692), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][8] ) );
  EDFQD1 \Storage_reg[26][7]  ( .D(n689), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][7] ) );
  EDFQD1 \Storage_reg[26][6]  ( .D(DataI[6]), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][6] ) );
  EDFQD1 \Storage_reg[26][5]  ( .D(DataI[5]), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][5] ) );
  EDFQD1 \Storage_reg[26][4]  ( .D(n680), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][4] ) );
  EDFQD1 \Storage_reg[26][3]  ( .D(n677), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][3] ) );
  EDFQD1 \Storage_reg[26][2]  ( .D(DataI[2]), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][2] ) );
  EDFQD1 \Storage_reg[26][1]  ( .D(n671), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][1] ) );
  EDFQD1 \Storage_reg[26][0]  ( .D(DataI[0]), .E(n577), .CP(ChipClock), .Q(
        \Storage[26][0] ) );
  EDFQD1 \Storage_reg[24][10]  ( .D(n698), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][10] ) );
  EDFQD1 \Storage_reg[24][9]  ( .D(n695), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][9] ) );
  EDFQD1 \Storage_reg[24][8]  ( .D(n692), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][8] ) );
  EDFQD1 \Storage_reg[24][7]  ( .D(n689), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][7] ) );
  EDFQD1 \Storage_reg[24][6]  ( .D(n686), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][6] ) );
  EDFQD1 \Storage_reg[24][5]  ( .D(n683), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][5] ) );
  EDFQD1 \Storage_reg[24][4]  ( .D(n680), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][4] ) );
  EDFQD1 \Storage_reg[24][3]  ( .D(n677), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][3] ) );
  EDFQD1 \Storage_reg[24][2]  ( .D(n674), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][2] ) );
  EDFQD1 \Storage_reg[24][1]  ( .D(n671), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][1] ) );
  EDFQD1 \Storage_reg[24][0]  ( .D(n668), .E(n583), .CP(ChipClock), .Q(
        \Storage[24][0] ) );
  EDFQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][10] ) );
  EDFQD1 \Storage_reg[30][9]  ( .D(n695), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][9] ) );
  EDFQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][8] ) );
  EDFQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][7] ) );
  EDFQD1 \Storage_reg[30][6]  ( .D(n686), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][6] ) );
  EDFQD1 \Storage_reg[30][5]  ( .D(n683), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][5] ) );
  EDFQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][4] ) );
  EDFQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][3] ) );
  EDFQD1 \Storage_reg[30][2]  ( .D(n674), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][2] ) );
  EDFQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][1] ) );
  EDFQD1 \Storage_reg[30][0]  ( .D(n668), .E(n565), .CP(ChipClock), .Q(
        \Storage[30][0] ) );
  EDFQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][10] ) );
  EDFQD1 \Storage_reg[29][9]  ( .D(n695), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][9] ) );
  EDFQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][8] ) );
  EDFQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][7] ) );
  EDFQD1 \Storage_reg[29][6]  ( .D(n686), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][6] ) );
  EDFQD1 \Storage_reg[29][5]  ( .D(n683), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][5] ) );
  EDFQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][4] ) );
  EDFQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][3] ) );
  EDFQD1 \Storage_reg[29][2]  ( .D(n674), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][2] ) );
  EDFQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][1] ) );
  EDFQD1 \Storage_reg[29][0]  ( .D(n668), .E(n568), .CP(ChipClock), .Q(
        \Storage[29][0] ) );
  EDFQD1 \Storage_reg[28][10]  ( .D(n698), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][10] ) );
  EDFQD1 \Storage_reg[28][9]  ( .D(DataI[9]), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][9] ) );
  EDFQD1 \Storage_reg[28][8]  ( .D(n692), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][8] ) );
  EDFQD1 \Storage_reg[28][7]  ( .D(n689), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][7] ) );
  EDFQD1 \Storage_reg[28][6]  ( .D(DataI[6]), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][6] ) );
  EDFQD1 \Storage_reg[28][5]  ( .D(DataI[5]), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][5] ) );
  EDFQD1 \Storage_reg[28][4]  ( .D(n680), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][4] ) );
  EDFQD1 \Storage_reg[28][3]  ( .D(n677), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][3] ) );
  EDFQD1 \Storage_reg[28][2]  ( .D(DataI[2]), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][2] ) );
  EDFQD1 \Storage_reg[28][1]  ( .D(n671), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][1] ) );
  EDFQD1 \Storage_reg[28][0]  ( .D(DataI[0]), .E(n571), .CP(ChipClock), .Q(
        \Storage[28][0] ) );
  EDFQD1 \Storage_reg[27][10]  ( .D(n698), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][10] ) );
  EDFQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][9] ) );
  EDFQD1 \Storage_reg[27][8]  ( .D(n692), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][8] ) );
  EDFQD1 \Storage_reg[27][7]  ( .D(n689), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][7] ) );
  EDFQD1 \Storage_reg[27][6]  ( .D(DataI[6]), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][6] ) );
  EDFQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][5] ) );
  EDFQD1 \Storage_reg[27][4]  ( .D(n680), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][4] ) );
  EDFQD1 \Storage_reg[27][3]  ( .D(n677), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][3] ) );
  EDFQD1 \Storage_reg[27][2]  ( .D(DataI[2]), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][2] ) );
  EDFQD1 \Storage_reg[27][1]  ( .D(n671), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][1] ) );
  EDFQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(n574), .CP(ChipClock), .Q(
        \Storage[27][0] ) );
  EDFQD1 \Storage_reg[25][10]  ( .D(n698), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][10] ) );
  EDFQD1 \Storage_reg[25][9]  ( .D(DataI[9]), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][9] ) );
  EDFQD1 \Storage_reg[25][8]  ( .D(n692), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][8] ) );
  EDFQD1 \Storage_reg[25][7]  ( .D(n689), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][7] ) );
  EDFQD1 \Storage_reg[25][6]  ( .D(DataI[6]), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][6] ) );
  EDFQD1 \Storage_reg[25][5]  ( .D(DataI[5]), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][5] ) );
  EDFQD1 \Storage_reg[25][4]  ( .D(n680), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][4] ) );
  EDFQD1 \Storage_reg[25][3]  ( .D(n677), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][3] ) );
  EDFQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][2] ) );
  EDFQD1 \Storage_reg[25][1]  ( .D(n671), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][1] ) );
  EDFQD1 \Storage_reg[25][0]  ( .D(DataI[0]), .E(n580), .CP(ChipClock), .Q(
        \Storage[25][0] ) );
  EDFQD1 \Storage_reg[22][10]  ( .D(n698), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][10] ) );
  EDFQD1 \Storage_reg[22][9]  ( .D(n695), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][9] ) );
  EDFQD1 \Storage_reg[22][8]  ( .D(n692), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][8] ) );
  EDFQD1 \Storage_reg[22][7]  ( .D(n689), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][7] ) );
  EDFQD1 \Storage_reg[22][6]  ( .D(n686), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][6] ) );
  EDFQD1 \Storage_reg[22][5]  ( .D(n683), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][5] ) );
  EDFQD1 \Storage_reg[22][4]  ( .D(n680), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][4] ) );
  EDFQD1 \Storage_reg[22][3]  ( .D(n677), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][3] ) );
  EDFQD1 \Storage_reg[22][2]  ( .D(n674), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][2] ) );
  EDFQD1 \Storage_reg[22][1]  ( .D(n671), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][1] ) );
  EDFQD1 \Storage_reg[22][0]  ( .D(n668), .E(n589), .CP(ChipClock), .Q(
        \Storage[22][0] ) );
  EDFQD1 \Storage_reg[21][10]  ( .D(n698), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][10] ) );
  EDFQD1 \Storage_reg[21][9]  ( .D(n695), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][9] ) );
  EDFQD1 \Storage_reg[21][8]  ( .D(n692), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][8] ) );
  EDFQD1 \Storage_reg[21][7]  ( .D(n689), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][7] ) );
  EDFQD1 \Storage_reg[21][6]  ( .D(n686), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][6] ) );
  EDFQD1 \Storage_reg[21][5]  ( .D(n683), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][5] ) );
  EDFQD1 \Storage_reg[21][4]  ( .D(n680), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][4] ) );
  EDFQD1 \Storage_reg[21][3]  ( .D(n677), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][3] ) );
  EDFQD1 \Storage_reg[21][2]  ( .D(n674), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][2] ) );
  EDFQD1 \Storage_reg[21][1]  ( .D(n671), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][1] ) );
  EDFQD1 \Storage_reg[21][0]  ( .D(n668), .E(n592), .CP(ChipClock), .Q(
        \Storage[21][0] ) );
  EDFQD1 \Storage_reg[18][10]  ( .D(n698), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][10] ) );
  EDFQD1 \Storage_reg[18][9]  ( .D(n695), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][9] ) );
  EDFQD1 \Storage_reg[18][8]  ( .D(n692), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][8] ) );
  EDFQD1 \Storage_reg[18][7]  ( .D(n689), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][7] ) );
  EDFQD1 \Storage_reg[18][6]  ( .D(n686), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][6] ) );
  EDFQD1 \Storage_reg[18][5]  ( .D(n683), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][5] ) );
  EDFQD1 \Storage_reg[18][4]  ( .D(n680), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][4] ) );
  EDFQD1 \Storage_reg[18][3]  ( .D(n677), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][3] ) );
  EDFQD1 \Storage_reg[18][2]  ( .D(n674), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][2] ) );
  EDFQD1 \Storage_reg[18][1]  ( .D(n671), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][1] ) );
  EDFQD1 \Storage_reg[18][0]  ( .D(n668), .E(n601), .CP(ChipClock), .Q(
        \Storage[18][0] ) );
  EDFQD1 \Storage_reg[17][10]  ( .D(n698), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][10] ) );
  EDFQD1 \Storage_reg[17][9]  ( .D(n695), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][9] ) );
  EDFQD1 \Storage_reg[17][8]  ( .D(n692), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][8] ) );
  EDFQD1 \Storage_reg[17][7]  ( .D(n689), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][7] ) );
  EDFQD1 \Storage_reg[17][6]  ( .D(n686), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][6] ) );
  EDFQD1 \Storage_reg[17][5]  ( .D(n683), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][5] ) );
  EDFQD1 \Storage_reg[17][4]  ( .D(n680), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][4] ) );
  EDFQD1 \Storage_reg[17][3]  ( .D(n677), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][3] ) );
  EDFQD1 \Storage_reg[17][2]  ( .D(n674), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][2] ) );
  EDFQD1 \Storage_reg[17][1]  ( .D(n671), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][1] ) );
  EDFQD1 \Storage_reg[17][0]  ( .D(n668), .E(n604), .CP(ChipClock), .Q(
        \Storage[17][0] ) );
  EDFQD1 \Storage_reg[14][10]  ( .D(n698), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][10] ) );
  EDFQD1 \Storage_reg[14][9]  ( .D(n695), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][9] ) );
  EDFQD1 \Storage_reg[14][8]  ( .D(n692), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][8] ) );
  EDFQD1 \Storage_reg[14][7]  ( .D(n689), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][7] ) );
  EDFQD1 \Storage_reg[14][6]  ( .D(n686), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][6] ) );
  EDFQD1 \Storage_reg[14][5]  ( .D(n683), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][5] ) );
  EDFQD1 \Storage_reg[14][4]  ( .D(n680), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][4] ) );
  EDFQD1 \Storage_reg[14][3]  ( .D(n677), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][3] ) );
  EDFQD1 \Storage_reg[14][2]  ( .D(n674), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][2] ) );
  EDFQD1 \Storage_reg[14][1]  ( .D(n671), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][1] ) );
  EDFQD1 \Storage_reg[14][0]  ( .D(n668), .E(n613), .CP(ChipClock), .Q(
        \Storage[14][0] ) );
  EDFQD1 \Storage_reg[13][10]  ( .D(n697), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][10] ) );
  EDFQD1 \Storage_reg[13][9]  ( .D(n695), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][9] ) );
  EDFQD1 \Storage_reg[13][8]  ( .D(n691), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][8] ) );
  EDFQD1 \Storage_reg[13][7]  ( .D(n688), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][7] ) );
  EDFQD1 \Storage_reg[13][6]  ( .D(n686), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][6] ) );
  EDFQD1 \Storage_reg[13][5]  ( .D(n683), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][5] ) );
  EDFQD1 \Storage_reg[13][4]  ( .D(n679), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][4] ) );
  EDFQD1 \Storage_reg[13][3]  ( .D(n676), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][3] ) );
  EDFQD1 \Storage_reg[13][2]  ( .D(n674), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][2] ) );
  EDFQD1 \Storage_reg[13][1]  ( .D(n670), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][1] ) );
  EDFQD1 \Storage_reg[13][0]  ( .D(n668), .E(n616), .CP(ChipClock), .Q(
        \Storage[13][0] ) );
  EDFQD1 \Storage_reg[10][10]  ( .D(n697), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][10] ) );
  EDFQD1 \Storage_reg[10][9]  ( .D(n694), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][9] ) );
  EDFQD1 \Storage_reg[10][8]  ( .D(n691), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][8] ) );
  EDFQD1 \Storage_reg[10][7]  ( .D(n688), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][7] ) );
  EDFQD1 \Storage_reg[10][6]  ( .D(n685), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][6] ) );
  EDFQD1 \Storage_reg[10][5]  ( .D(n682), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][5] ) );
  EDFQD1 \Storage_reg[10][4]  ( .D(n679), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][4] ) );
  EDFQD1 \Storage_reg[10][3]  ( .D(n676), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][3] ) );
  EDFQD1 \Storage_reg[10][2]  ( .D(n673), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][2] ) );
  EDFQD1 \Storage_reg[10][1]  ( .D(n670), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][1] ) );
  EDFQD1 \Storage_reg[10][0]  ( .D(n667), .E(n625), .CP(ChipClock), .Q(
        \Storage[10][0] ) );
  EDFQD1 \Storage_reg[9][10]  ( .D(n697), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][10] ) );
  EDFQD1 \Storage_reg[9][9]  ( .D(n694), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][9] ) );
  EDFQD1 \Storage_reg[9][8]  ( .D(n691), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][8] ) );
  EDFQD1 \Storage_reg[9][7]  ( .D(n688), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][7] ) );
  EDFQD1 \Storage_reg[9][6]  ( .D(n685), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][6] ) );
  EDFQD1 \Storage_reg[9][5]  ( .D(n682), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][5] ) );
  EDFQD1 \Storage_reg[9][4]  ( .D(n679), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][4] ) );
  EDFQD1 \Storage_reg[9][3]  ( .D(n676), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][3] ) );
  EDFQD1 \Storage_reg[9][2]  ( .D(n673), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][2] ) );
  EDFQD1 \Storage_reg[9][1]  ( .D(n670), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][1] ) );
  EDFQD1 \Storage_reg[9][0]  ( .D(n667), .E(n628), .CP(ChipClock), .Q(
        \Storage[9][0] ) );
  EDFQD1 \Storage_reg[6][10]  ( .D(n697), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][10] ) );
  EDFQD1 \Storage_reg[6][9]  ( .D(n694), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][9] ) );
  EDFQD1 \Storage_reg[6][8]  ( .D(n691), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][8] ) );
  EDFQD1 \Storage_reg[6][7]  ( .D(n688), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][7] ) );
  EDFQD1 \Storage_reg[6][6]  ( .D(n685), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][6] ) );
  EDFQD1 \Storage_reg[6][5]  ( .D(n682), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][5] ) );
  EDFQD1 \Storage_reg[6][4]  ( .D(n679), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][4] ) );
  EDFQD1 \Storage_reg[6][3]  ( .D(n676), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][3] ) );
  EDFQD1 \Storage_reg[6][2]  ( .D(n673), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][2] ) );
  EDFQD1 \Storage_reg[6][1]  ( .D(n670), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][1] ) );
  EDFQD1 \Storage_reg[6][0]  ( .D(n667), .E(n637), .CP(ChipClock), .Q(
        \Storage[6][0] ) );
  EDFQD1 \Storage_reg[5][10]  ( .D(n697), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][10] ) );
  EDFQD1 \Storage_reg[5][9]  ( .D(n694), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][9] ) );
  EDFQD1 \Storage_reg[5][8]  ( .D(n691), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][8] ) );
  EDFQD1 \Storage_reg[5][7]  ( .D(n688), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][7] ) );
  EDFQD1 \Storage_reg[5][6]  ( .D(n685), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][6] ) );
  EDFQD1 \Storage_reg[5][5]  ( .D(n682), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][5] ) );
  EDFQD1 \Storage_reg[5][4]  ( .D(n679), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][4] ) );
  EDFQD1 \Storage_reg[5][3]  ( .D(n676), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][3] ) );
  EDFQD1 \Storage_reg[5][2]  ( .D(n673), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][2] ) );
  EDFQD1 \Storage_reg[5][1]  ( .D(n670), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][1] ) );
  EDFQD1 \Storage_reg[5][0]  ( .D(n667), .E(n640), .CP(ChipClock), .Q(
        \Storage[5][0] ) );
  EDFQD1 \Storage_reg[2][10]  ( .D(n697), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][10] ) );
  EDFQD1 \Storage_reg[2][9]  ( .D(n694), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][9] ) );
  EDFQD1 \Storage_reg[2][8]  ( .D(n691), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][8] ) );
  EDFQD1 \Storage_reg[2][7]  ( .D(n688), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][7] ) );
  EDFQD1 \Storage_reg[2][6]  ( .D(n685), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][6] ) );
  EDFQD1 \Storage_reg[2][5]  ( .D(n682), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][5] ) );
  EDFQD1 \Storage_reg[2][4]  ( .D(n679), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][4] ) );
  EDFQD1 \Storage_reg[2][3]  ( .D(n676), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][3] ) );
  EDFQD1 \Storage_reg[2][2]  ( .D(n673), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][2] ) );
  EDFQD1 \Storage_reg[2][1]  ( .D(n670), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][1] ) );
  EDFQD1 \Storage_reg[2][0]  ( .D(n667), .E(n649), .CP(ChipClock), .Q(
        \Storage[2][0] ) );
  EDFQD1 \Storage_reg[1][10]  ( .D(n697), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][10] ) );
  EDFQD1 \Storage_reg[1][9]  ( .D(n694), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][9] ) );
  EDFQD1 \Storage_reg[1][8]  ( .D(n691), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][8] ) );
  EDFQD1 \Storage_reg[1][7]  ( .D(n688), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][7] ) );
  EDFQD1 \Storage_reg[1][6]  ( .D(n685), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][6] ) );
  EDFQD1 \Storage_reg[1][5]  ( .D(n682), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][5] ) );
  EDFQD1 \Storage_reg[1][4]  ( .D(n679), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][4] ) );
  EDFQD1 \Storage_reg[1][3]  ( .D(n676), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][3] ) );
  EDFQD1 \Storage_reg[1][2]  ( .D(n673), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][2] ) );
  EDFQD1 \Storage_reg[1][1]  ( .D(n670), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][1] ) );
  EDFQD1 \Storage_reg[1][0]  ( .D(n667), .E(n652), .CP(ChipClock), .Q(
        \Storage[1][0] ) );
  EDFQD1 \Storage_reg[23][10]  ( .D(n698), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][10] ) );
  EDFQD1 \Storage_reg[23][9]  ( .D(n695), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][9] ) );
  EDFQD1 \Storage_reg[23][8]  ( .D(n692), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][8] ) );
  EDFQD1 \Storage_reg[23][7]  ( .D(n689), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][7] ) );
  EDFQD1 \Storage_reg[23][6]  ( .D(n686), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][6] ) );
  EDFQD1 \Storage_reg[23][5]  ( .D(n683), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][5] ) );
  EDFQD1 \Storage_reg[23][4]  ( .D(n680), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][4] ) );
  EDFQD1 \Storage_reg[23][3]  ( .D(n677), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][3] ) );
  EDFQD1 \Storage_reg[23][2]  ( .D(n674), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][2] ) );
  EDFQD1 \Storage_reg[23][1]  ( .D(n671), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][1] ) );
  EDFQD1 \Storage_reg[23][0]  ( .D(n668), .E(n586), .CP(ChipClock), .Q(
        \Storage[23][0] ) );
  EDFQD1 \Storage_reg[20][10]  ( .D(n698), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][10] ) );
  EDFQD1 \Storage_reg[20][9]  ( .D(n695), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][9] ) );
  EDFQD1 \Storage_reg[20][8]  ( .D(n692), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][8] ) );
  EDFQD1 \Storage_reg[20][7]  ( .D(n689), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][7] ) );
  EDFQD1 \Storage_reg[20][6]  ( .D(n686), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][6] ) );
  EDFQD1 \Storage_reg[20][5]  ( .D(n683), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][5] ) );
  EDFQD1 \Storage_reg[20][4]  ( .D(n680), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][4] ) );
  EDFQD1 \Storage_reg[20][3]  ( .D(n677), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][3] ) );
  EDFQD1 \Storage_reg[20][2]  ( .D(n674), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][2] ) );
  EDFQD1 \Storage_reg[20][1]  ( .D(n671), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][1] ) );
  EDFQD1 \Storage_reg[20][0]  ( .D(n668), .E(n595), .CP(ChipClock), .Q(
        \Storage[20][0] ) );
  EDFQD1 \Storage_reg[19][10]  ( .D(n698), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][10] ) );
  EDFQD1 \Storage_reg[19][9]  ( .D(n695), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][9] ) );
  EDFQD1 \Storage_reg[19][8]  ( .D(n692), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][8] ) );
  EDFQD1 \Storage_reg[19][7]  ( .D(n689), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][7] ) );
  EDFQD1 \Storage_reg[19][6]  ( .D(n686), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][6] ) );
  EDFQD1 \Storage_reg[19][5]  ( .D(n683), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][5] ) );
  EDFQD1 \Storage_reg[19][4]  ( .D(n680), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][4] ) );
  EDFQD1 \Storage_reg[19][3]  ( .D(n677), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][3] ) );
  EDFQD1 \Storage_reg[19][2]  ( .D(n674), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][2] ) );
  EDFQD1 \Storage_reg[19][1]  ( .D(n671), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][1] ) );
  EDFQD1 \Storage_reg[19][0]  ( .D(n668), .E(n598), .CP(ChipClock), .Q(
        \Storage[19][0] ) );
  EDFQD1 \Storage_reg[16][10]  ( .D(n698), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][10] ) );
  EDFQD1 \Storage_reg[16][9]  ( .D(n695), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][9] ) );
  EDFQD1 \Storage_reg[16][8]  ( .D(n692), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][8] ) );
  EDFQD1 \Storage_reg[16][7]  ( .D(n689), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][7] ) );
  EDFQD1 \Storage_reg[16][6]  ( .D(n686), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][6] ) );
  EDFQD1 \Storage_reg[16][5]  ( .D(n683), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][5] ) );
  EDFQD1 \Storage_reg[16][4]  ( .D(n680), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][4] ) );
  EDFQD1 \Storage_reg[16][3]  ( .D(n677), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][3] ) );
  EDFQD1 \Storage_reg[16][2]  ( .D(n674), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][2] ) );
  EDFQD1 \Storage_reg[16][1]  ( .D(n671), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][1] ) );
  EDFQD1 \Storage_reg[16][0]  ( .D(n668), .E(n607), .CP(ChipClock), .Q(
        \Storage[16][0] ) );
  EDFQD1 \Storage_reg[15][10]  ( .D(n698), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][10] ) );
  EDFQD1 \Storage_reg[15][9]  ( .D(n695), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][9] ) );
  EDFQD1 \Storage_reg[15][8]  ( .D(n692), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][8] ) );
  EDFQD1 \Storage_reg[15][7]  ( .D(n689), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][7] ) );
  EDFQD1 \Storage_reg[15][6]  ( .D(n686), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][6] ) );
  EDFQD1 \Storage_reg[15][5]  ( .D(n683), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][5] ) );
  EDFQD1 \Storage_reg[15][4]  ( .D(n680), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][4] ) );
  EDFQD1 \Storage_reg[15][3]  ( .D(n677), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][3] ) );
  EDFQD1 \Storage_reg[15][2]  ( .D(n674), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][2] ) );
  EDFQD1 \Storage_reg[15][1]  ( .D(n671), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][1] ) );
  EDFQD1 \Storage_reg[15][0]  ( .D(n668), .E(n610), .CP(ChipClock), .Q(
        \Storage[15][0] ) );
  EDFQD1 \Storage_reg[12][10]  ( .D(n697), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][10] ) );
  EDFQD1 \Storage_reg[12][9]  ( .D(n695), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][9] ) );
  EDFQD1 \Storage_reg[12][8]  ( .D(n691), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][8] ) );
  EDFQD1 \Storage_reg[12][7]  ( .D(n688), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][7] ) );
  EDFQD1 \Storage_reg[12][6]  ( .D(n686), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][6] ) );
  EDFQD1 \Storage_reg[12][5]  ( .D(n683), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][5] ) );
  EDFQD1 \Storage_reg[12][4]  ( .D(n679), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][4] ) );
  EDFQD1 \Storage_reg[12][3]  ( .D(n676), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][3] ) );
  EDFQD1 \Storage_reg[12][2]  ( .D(n674), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][2] ) );
  EDFQD1 \Storage_reg[12][1]  ( .D(n670), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][1] ) );
  EDFQD1 \Storage_reg[12][0]  ( .D(n668), .E(n619), .CP(ChipClock), .Q(
        \Storage[12][0] ) );
  EDFQD1 \Storage_reg[11][10]  ( .D(n697), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][10] ) );
  EDFQD1 \Storage_reg[11][9]  ( .D(n694), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][9] ) );
  EDFQD1 \Storage_reg[11][8]  ( .D(n691), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][8] ) );
  EDFQD1 \Storage_reg[11][7]  ( .D(n688), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][7] ) );
  EDFQD1 \Storage_reg[11][6]  ( .D(n685), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][6] ) );
  EDFQD1 \Storage_reg[11][5]  ( .D(n682), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][5] ) );
  EDFQD1 \Storage_reg[11][4]  ( .D(n679), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][4] ) );
  EDFQD1 \Storage_reg[11][3]  ( .D(n676), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][3] ) );
  EDFQD1 \Storage_reg[11][2]  ( .D(n673), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][2] ) );
  EDFQD1 \Storage_reg[11][1]  ( .D(n670), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][1] ) );
  EDFQD1 \Storage_reg[11][0]  ( .D(n667), .E(n622), .CP(ChipClock), .Q(
        \Storage[11][0] ) );
  EDFQD1 \Storage_reg[8][10]  ( .D(n697), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][10] ) );
  EDFQD1 \Storage_reg[8][9]  ( .D(n694), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][9] ) );
  EDFQD1 \Storage_reg[8][8]  ( .D(n691), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][8] ) );
  EDFQD1 \Storage_reg[8][7]  ( .D(n688), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][7] ) );
  EDFQD1 \Storage_reg[8][6]  ( .D(n685), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][6] ) );
  EDFQD1 \Storage_reg[8][5]  ( .D(n682), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][5] ) );
  EDFQD1 \Storage_reg[8][4]  ( .D(n679), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][4] ) );
  EDFQD1 \Storage_reg[8][3]  ( .D(n676), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][3] ) );
  EDFQD1 \Storage_reg[8][2]  ( .D(n673), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][2] ) );
  EDFQD1 \Storage_reg[8][1]  ( .D(n670), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][1] ) );
  EDFQD1 \Storage_reg[8][0]  ( .D(n667), .E(n631), .CP(ChipClock), .Q(
        \Storage[8][0] ) );
  EDFQD1 \Storage_reg[7][10]  ( .D(n697), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][10] ) );
  EDFQD1 \Storage_reg[7][9]  ( .D(n694), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][9] ) );
  EDFQD1 \Storage_reg[7][8]  ( .D(n691), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][8] ) );
  EDFQD1 \Storage_reg[7][7]  ( .D(n688), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][7] ) );
  EDFQD1 \Storage_reg[7][6]  ( .D(n685), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][6] ) );
  EDFQD1 \Storage_reg[7][5]  ( .D(n682), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][5] ) );
  EDFQD1 \Storage_reg[7][4]  ( .D(n679), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][4] ) );
  EDFQD1 \Storage_reg[7][3]  ( .D(n676), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][3] ) );
  EDFQD1 \Storage_reg[7][2]  ( .D(n673), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][2] ) );
  EDFQD1 \Storage_reg[7][1]  ( .D(n670), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][1] ) );
  EDFQD1 \Storage_reg[7][0]  ( .D(n667), .E(n634), .CP(ChipClock), .Q(
        \Storage[7][0] ) );
  EDFQD1 \Storage_reg[4][10]  ( .D(n697), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][10] ) );
  EDFQD1 \Storage_reg[4][9]  ( .D(n694), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][9] ) );
  EDFQD1 \Storage_reg[4][8]  ( .D(n691), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][8] ) );
  EDFQD1 \Storage_reg[4][7]  ( .D(n688), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][7] ) );
  EDFQD1 \Storage_reg[4][6]  ( .D(n685), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][6] ) );
  EDFQD1 \Storage_reg[4][5]  ( .D(n682), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][5] ) );
  EDFQD1 \Storage_reg[4][4]  ( .D(n679), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][4] ) );
  EDFQD1 \Storage_reg[4][3]  ( .D(n676), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][3] ) );
  EDFQD1 \Storage_reg[4][2]  ( .D(n673), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][2] ) );
  EDFQD1 \Storage_reg[4][1]  ( .D(n670), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][1] ) );
  EDFQD1 \Storage_reg[4][0]  ( .D(n667), .E(n643), .CP(ChipClock), .Q(
        \Storage[4][0] ) );
  EDFQD1 \Storage_reg[3][10]  ( .D(n697), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][10] ) );
  EDFQD1 \Storage_reg[3][9]  ( .D(n694), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][9] ) );
  EDFQD1 \Storage_reg[3][8]  ( .D(n691), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][8] ) );
  EDFQD1 \Storage_reg[3][7]  ( .D(n688), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][7] ) );
  EDFQD1 \Storage_reg[3][6]  ( .D(n685), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][6] ) );
  EDFQD1 \Storage_reg[3][5]  ( .D(n682), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][5] ) );
  EDFQD1 \Storage_reg[3][4]  ( .D(n679), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][4] ) );
  EDFQD1 \Storage_reg[3][3]  ( .D(n676), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][3] ) );
  EDFQD1 \Storage_reg[3][2]  ( .D(n673), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][2] ) );
  EDFQD1 \Storage_reg[3][1]  ( .D(n670), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][1] ) );
  EDFQD1 \Storage_reg[3][0]  ( .D(n667), .E(n646), .CP(ChipClock), .Q(
        \Storage[3][0] ) );
  EDFQD1 \Storage_reg[0][10]  ( .D(n697), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][10] ) );
  EDFQD1 \Storage_reg[0][9]  ( .D(n694), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][9] ) );
  EDFQD1 \Storage_reg[0][8]  ( .D(n691), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][8] ) );
  EDFQD1 \Storage_reg[0][7]  ( .D(n688), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][7] ) );
  EDFQD1 \Storage_reg[0][6]  ( .D(n685), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][6] ) );
  EDFQD1 \Storage_reg[0][5]  ( .D(n682), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][5] ) );
  EDFQD1 \Storage_reg[0][4]  ( .D(n679), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][4] ) );
  EDFQD1 \Storage_reg[0][3]  ( .D(n676), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][3] ) );
  EDFQD1 \Storage_reg[0][2]  ( .D(n673), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][2] ) );
  EDFQD1 \Storage_reg[0][1]  ( .D(n670), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][1] ) );
  EDFQD1 \Storage_reg[0][0]  ( .D(n667), .E(n655), .CP(ChipClock), .Q(
        \Storage[0][0] ) );
  EDFQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][10] ) );
  EDFQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][9] ) );
  EDFQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][8] ) );
  EDFQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][7] ) );
  EDFQD1 \Storage_reg[31][6]  ( .D(DataI[6]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][6] ) );
  EDFQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][5] ) );
  EDFQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][4] ) );
  EDFQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][3] ) );
  EDFQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][2] ) );
  EDFQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][1] ) );
  EDFQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(n562), .CP(ChipClock), .Q(
        \Storage[31][0] ) );
  EDFQD1 \Storage_reg[26][32]  ( .D(n656), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][32] ) );
  EDFQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][31] ) );
  EDFQD1 \Storage_reg[26][30]  ( .D(n758), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][30] ) );
  EDFQD1 \Storage_reg[26][29]  ( .D(n755), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][29] ) );
  EDFQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][28] ) );
  EDFQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][27] ) );
  EDFQD1 \Storage_reg[26][26]  ( .D(n746), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][26] ) );
  EDFQD1 \Storage_reg[26][25]  ( .D(n743), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][25] ) );
  EDFQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][24] ) );
  EDFQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][23] ) );
  EDFQD1 \Storage_reg[26][22]  ( .D(n734), .E(n575), .CP(ChipClock), .Q(
        \Storage[26][22] ) );
  EDFQD1 \Storage_reg[26][21]  ( .D(n731), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][21] ) );
  EDFQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][20] ) );
  EDFQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][19] ) );
  EDFQD1 \Storage_reg[26][18]  ( .D(n722), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][18] ) );
  EDFQD1 \Storage_reg[26][17]  ( .D(n719), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][17] ) );
  EDFQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][16] ) );
  EDFQD1 \Storage_reg[26][15]  ( .D(n713), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][15] ) );
  EDFQD1 \Storage_reg[26][14]  ( .D(n710), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][14] ) );
  EDFQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][13] ) );
  EDFQD1 \Storage_reg[26][12]  ( .D(DataI[12]), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][12] ) );
  EDFQD1 \Storage_reg[26][11]  ( .D(n701), .E(n576), .CP(ChipClock), .Q(
        \Storage[26][11] ) );
  EDFQD1 \Storage_reg[24][32]  ( .D(n656), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][32] ) );
  EDFQD1 \Storage_reg[24][31]  ( .D(n761), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][31] ) );
  EDFQD1 \Storage_reg[24][30]  ( .D(n758), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][30] ) );
  EDFQD1 \Storage_reg[24][29]  ( .D(n755), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][29] ) );
  EDFQD1 \Storage_reg[24][28]  ( .D(n752), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][28] ) );
  EDFQD1 \Storage_reg[24][27]  ( .D(n749), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][27] ) );
  EDFQD1 \Storage_reg[24][26]  ( .D(n746), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][26] ) );
  EDFQD1 \Storage_reg[24][25]  ( .D(n743), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][25] ) );
  EDFQD1 \Storage_reg[24][24]  ( .D(n740), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][24] ) );
  EDFQD1 \Storage_reg[24][23]  ( .D(n737), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][23] ) );
  EDFQD1 \Storage_reg[24][22]  ( .D(n734), .E(n581), .CP(ChipClock), .Q(
        \Storage[24][22] ) );
  EDFQD1 \Storage_reg[24][21]  ( .D(n731), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][21] ) );
  EDFQD1 \Storage_reg[24][20]  ( .D(n728), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][20] ) );
  EDFQD1 \Storage_reg[24][19]  ( .D(n725), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][19] ) );
  EDFQD1 \Storage_reg[24][18]  ( .D(n722), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][18] ) );
  EDFQD1 \Storage_reg[24][17]  ( .D(n719), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][17] ) );
  EDFQD1 \Storage_reg[24][16]  ( .D(n716), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][16] ) );
  EDFQD1 \Storage_reg[24][15]  ( .D(n713), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][15] ) );
  EDFQD1 \Storage_reg[24][14]  ( .D(n710), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][14] ) );
  EDFQD1 \Storage_reg[24][13]  ( .D(n707), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][13] ) );
  EDFQD1 \Storage_reg[24][12]  ( .D(n704), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][12] ) );
  EDFQD1 \Storage_reg[24][11]  ( .D(n701), .E(n582), .CP(ChipClock), .Q(
        \Storage[24][11] ) );
  EDFQD1 \Storage_reg[30][32]  ( .D(n656), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][32] ) );
  EDFQD1 \Storage_reg[30][31]  ( .D(n761), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][31] ) );
  EDFQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][30] ) );
  EDFQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][29] ) );
  EDFQD1 \Storage_reg[30][28]  ( .D(n752), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][28] ) );
  EDFQD1 \Storage_reg[30][27]  ( .D(n749), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][27] ) );
  EDFQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][26] ) );
  EDFQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][25] ) );
  EDFQD1 \Storage_reg[30][24]  ( .D(n740), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][24] ) );
  EDFQD1 \Storage_reg[30][23]  ( .D(n737), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][23] ) );
  EDFQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(n563), .CP(ChipClock), .Q(
        \Storage[30][22] ) );
  EDFQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][21] ) );
  EDFQD1 \Storage_reg[30][20]  ( .D(n728), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][20] ) );
  EDFQD1 \Storage_reg[30][19]  ( .D(n725), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][19] ) );
  EDFQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][18] ) );
  EDFQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][17] ) );
  EDFQD1 \Storage_reg[30][16]  ( .D(n716), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][16] ) );
  EDFQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][15] ) );
  EDFQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][14] ) );
  EDFQD1 \Storage_reg[30][13]  ( .D(n707), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][13] ) );
  EDFQD1 \Storage_reg[30][12]  ( .D(n704), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][12] ) );
  EDFQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n564), .CP(ChipClock), .Q(
        \Storage[30][11] ) );
  EDFQD1 \Storage_reg[29][32]  ( .D(n656), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][32] ) );
  EDFQD1 \Storage_reg[29][31]  ( .D(n761), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][31] ) );
  EDFQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][30] ) );
  EDFQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][29] ) );
  EDFQD1 \Storage_reg[29][28]  ( .D(n752), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][28] ) );
  EDFQD1 \Storage_reg[29][27]  ( .D(n749), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][27] ) );
  EDFQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][26] ) );
  EDFQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][25] ) );
  EDFQD1 \Storage_reg[29][24]  ( .D(n740), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][24] ) );
  EDFQD1 \Storage_reg[29][23]  ( .D(n737), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][23] ) );
  EDFQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(n566), .CP(ChipClock), .Q(
        \Storage[29][22] ) );
  EDFQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][21] ) );
  EDFQD1 \Storage_reg[29][20]  ( .D(n728), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][20] ) );
  EDFQD1 \Storage_reg[29][19]  ( .D(n725), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][19] ) );
  EDFQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][18] ) );
  EDFQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][17] ) );
  EDFQD1 \Storage_reg[29][16]  ( .D(n716), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][16] ) );
  EDFQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][15] ) );
  EDFQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][14] ) );
  EDFQD1 \Storage_reg[29][13]  ( .D(n707), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][13] ) );
  EDFQD1 \Storage_reg[29][12]  ( .D(n704), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][12] ) );
  EDFQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(n567), .CP(ChipClock), .Q(
        \Storage[29][11] ) );
  EDFQD1 \Storage_reg[28][32]  ( .D(n656), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][32] ) );
  EDFQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][31] ) );
  EDFQD1 \Storage_reg[28][30]  ( .D(n758), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][30] ) );
  EDFQD1 \Storage_reg[28][29]  ( .D(n755), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][29] ) );
  EDFQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][28] ) );
  EDFQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][27] ) );
  EDFQD1 \Storage_reg[28][26]  ( .D(n746), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][26] ) );
  EDFQD1 \Storage_reg[28][25]  ( .D(n743), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][25] ) );
  EDFQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][24] ) );
  EDFQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][23] ) );
  EDFQD1 \Storage_reg[28][22]  ( .D(n734), .E(n569), .CP(ChipClock), .Q(
        \Storage[28][22] ) );
  EDFQD1 \Storage_reg[28][21]  ( .D(n731), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][21] ) );
  EDFQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][20] ) );
  EDFQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][19] ) );
  EDFQD1 \Storage_reg[28][18]  ( .D(n722), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][18] ) );
  EDFQD1 \Storage_reg[28][17]  ( .D(n719), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][17] ) );
  EDFQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][16] ) );
  EDFQD1 \Storage_reg[28][15]  ( .D(n713), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][15] ) );
  EDFQD1 \Storage_reg[28][14]  ( .D(n710), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][14] ) );
  EDFQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][13] ) );
  EDFQD1 \Storage_reg[28][12]  ( .D(DataI[12]), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][12] ) );
  EDFQD1 \Storage_reg[28][11]  ( .D(n701), .E(n570), .CP(ChipClock), .Q(
        \Storage[28][11] ) );
  EDFQD1 \Storage_reg[27][32]  ( .D(n656), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][32] ) );
  EDFQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][31] ) );
  EDFQD1 \Storage_reg[27][30]  ( .D(n758), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][30] ) );
  EDFQD1 \Storage_reg[27][29]  ( .D(n755), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][29] ) );
  EDFQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][28] ) );
  EDFQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][27] ) );
  EDFQD1 \Storage_reg[27][26]  ( .D(n746), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][26] ) );
  EDFQD1 \Storage_reg[27][25]  ( .D(n743), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][25] ) );
  EDFQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][24] ) );
  EDFQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][23] ) );
  EDFQD1 \Storage_reg[27][22]  ( .D(n734), .E(n572), .CP(ChipClock), .Q(
        \Storage[27][22] ) );
  EDFQD1 \Storage_reg[27][21]  ( .D(n731), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][21] ) );
  EDFQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][20] ) );
  EDFQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][19] ) );
  EDFQD1 \Storage_reg[27][18]  ( .D(n722), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][18] ) );
  EDFQD1 \Storage_reg[27][17]  ( .D(n719), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][17] ) );
  EDFQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][16] ) );
  EDFQD1 \Storage_reg[27][15]  ( .D(n713), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][15] ) );
  EDFQD1 \Storage_reg[27][14]  ( .D(n710), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][14] ) );
  EDFQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][13] ) );
  EDFQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][12] ) );
  EDFQD1 \Storage_reg[27][11]  ( .D(n701), .E(n573), .CP(ChipClock), .Q(
        \Storage[27][11] ) );
  EDFQD1 \Storage_reg[25][32]  ( .D(n656), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][32] ) );
  EDFQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][31] ) );
  EDFQD1 \Storage_reg[25][30]  ( .D(n758), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][30] ) );
  EDFQD1 \Storage_reg[25][29]  ( .D(n755), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][29] ) );
  EDFQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][28] ) );
  EDFQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][27] ) );
  EDFQD1 \Storage_reg[25][26]  ( .D(n746), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][26] ) );
  EDFQD1 \Storage_reg[25][25]  ( .D(n743), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][25] ) );
  EDFQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][24] ) );
  EDFQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][23] ) );
  EDFQD1 \Storage_reg[25][22]  ( .D(n734), .E(n578), .CP(ChipClock), .Q(
        \Storage[25][22] ) );
  EDFQD1 \Storage_reg[25][21]  ( .D(n731), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][21] ) );
  EDFQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][20] ) );
  EDFQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][19] ) );
  EDFQD1 \Storage_reg[25][18]  ( .D(n722), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][18] ) );
  EDFQD1 \Storage_reg[25][17]  ( .D(n719), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][17] ) );
  EDFQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][16] ) );
  EDFQD1 \Storage_reg[25][15]  ( .D(n713), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][15] ) );
  EDFQD1 \Storage_reg[25][14]  ( .D(n710), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][14] ) );
  EDFQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][13] ) );
  EDFQD1 \Storage_reg[25][12]  ( .D(DataI[12]), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][12] ) );
  EDFQD1 \Storage_reg[25][11]  ( .D(n701), .E(n579), .CP(ChipClock), .Q(
        \Storage[25][11] ) );
  EDFQD1 \Storage_reg[22][32]  ( .D(n656), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][32] ) );
  EDFQD1 \Storage_reg[22][31]  ( .D(n761), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][31] ) );
  EDFQD1 \Storage_reg[22][30]  ( .D(n758), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][30] ) );
  EDFQD1 \Storage_reg[22][29]  ( .D(n755), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][29] ) );
  EDFQD1 \Storage_reg[22][28]  ( .D(n752), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][28] ) );
  EDFQD1 \Storage_reg[22][27]  ( .D(n749), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][27] ) );
  EDFQD1 \Storage_reg[22][26]  ( .D(n746), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][26] ) );
  EDFQD1 \Storage_reg[22][25]  ( .D(n743), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][25] ) );
  EDFQD1 \Storage_reg[22][24]  ( .D(n740), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][24] ) );
  EDFQD1 \Storage_reg[22][23]  ( .D(n737), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][23] ) );
  EDFQD1 \Storage_reg[22][22]  ( .D(n734), .E(n587), .CP(ChipClock), .Q(
        \Storage[22][22] ) );
  EDFQD1 \Storage_reg[22][21]  ( .D(n731), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][21] ) );
  EDFQD1 \Storage_reg[22][20]  ( .D(n728), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][20] ) );
  EDFQD1 \Storage_reg[22][19]  ( .D(n725), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][19] ) );
  EDFQD1 \Storage_reg[22][18]  ( .D(n722), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][18] ) );
  EDFQD1 \Storage_reg[22][17]  ( .D(n719), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][17] ) );
  EDFQD1 \Storage_reg[22][16]  ( .D(n716), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][16] ) );
  EDFQD1 \Storage_reg[22][15]  ( .D(n713), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][15] ) );
  EDFQD1 \Storage_reg[22][14]  ( .D(n710), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][14] ) );
  EDFQD1 \Storage_reg[22][13]  ( .D(n707), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][13] ) );
  EDFQD1 \Storage_reg[22][12]  ( .D(n704), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][12] ) );
  EDFQD1 \Storage_reg[22][11]  ( .D(n701), .E(n588), .CP(ChipClock), .Q(
        \Storage[22][11] ) );
  EDFQD1 \Storage_reg[21][32]  ( .D(n656), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][32] ) );
  EDFQD1 \Storage_reg[21][31]  ( .D(n761), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][31] ) );
  EDFQD1 \Storage_reg[21][30]  ( .D(n758), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][30] ) );
  EDFQD1 \Storage_reg[21][29]  ( .D(n755), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][29] ) );
  EDFQD1 \Storage_reg[21][28]  ( .D(n752), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][28] ) );
  EDFQD1 \Storage_reg[21][27]  ( .D(n749), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][27] ) );
  EDFQD1 \Storage_reg[21][26]  ( .D(n746), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][26] ) );
  EDFQD1 \Storage_reg[21][25]  ( .D(n743), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][25] ) );
  EDFQD1 \Storage_reg[21][24]  ( .D(n740), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][24] ) );
  EDFQD1 \Storage_reg[21][23]  ( .D(n737), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][23] ) );
  EDFQD1 \Storage_reg[21][22]  ( .D(n734), .E(n590), .CP(ChipClock), .Q(
        \Storage[21][22] ) );
  EDFQD1 \Storage_reg[21][21]  ( .D(n731), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][21] ) );
  EDFQD1 \Storage_reg[21][20]  ( .D(n728), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][20] ) );
  EDFQD1 \Storage_reg[21][19]  ( .D(n725), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][19] ) );
  EDFQD1 \Storage_reg[21][18]  ( .D(n722), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][18] ) );
  EDFQD1 \Storage_reg[21][17]  ( .D(n719), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][17] ) );
  EDFQD1 \Storage_reg[21][16]  ( .D(n716), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][16] ) );
  EDFQD1 \Storage_reg[21][15]  ( .D(n713), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][15] ) );
  EDFQD1 \Storage_reg[21][14]  ( .D(n710), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][14] ) );
  EDFQD1 \Storage_reg[21][13]  ( .D(n707), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][13] ) );
  EDFQD1 \Storage_reg[21][12]  ( .D(n704), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][12] ) );
  EDFQD1 \Storage_reg[21][11]  ( .D(n701), .E(n591), .CP(ChipClock), .Q(
        \Storage[21][11] ) );
  EDFQD1 \Storage_reg[18][32]  ( .D(n657), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][32] ) );
  EDFQD1 \Storage_reg[18][31]  ( .D(n761), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][31] ) );
  EDFQD1 \Storage_reg[18][30]  ( .D(n758), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][30] ) );
  EDFQD1 \Storage_reg[18][29]  ( .D(n755), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][29] ) );
  EDFQD1 \Storage_reg[18][28]  ( .D(n752), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][28] ) );
  EDFQD1 \Storage_reg[18][27]  ( .D(n749), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][27] ) );
  EDFQD1 \Storage_reg[18][26]  ( .D(n746), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][26] ) );
  EDFQD1 \Storage_reg[18][25]  ( .D(n743), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][25] ) );
  EDFQD1 \Storage_reg[18][24]  ( .D(n740), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][24] ) );
  EDFQD1 \Storage_reg[18][23]  ( .D(n737), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][23] ) );
  EDFQD1 \Storage_reg[18][22]  ( .D(n734), .E(n599), .CP(ChipClock), .Q(
        \Storage[18][22] ) );
  EDFQD1 \Storage_reg[18][21]  ( .D(n731), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][21] ) );
  EDFQD1 \Storage_reg[18][20]  ( .D(n728), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][20] ) );
  EDFQD1 \Storage_reg[18][19]  ( .D(n725), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][19] ) );
  EDFQD1 \Storage_reg[18][18]  ( .D(n722), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][18] ) );
  EDFQD1 \Storage_reg[18][17]  ( .D(n719), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][17] ) );
  EDFQD1 \Storage_reg[18][16]  ( .D(n716), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][16] ) );
  EDFQD1 \Storage_reg[18][15]  ( .D(n713), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][15] ) );
  EDFQD1 \Storage_reg[18][14]  ( .D(n710), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][14] ) );
  EDFQD1 \Storage_reg[18][13]  ( .D(n707), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][13] ) );
  EDFQD1 \Storage_reg[18][12]  ( .D(n704), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][12] ) );
  EDFQD1 \Storage_reg[18][11]  ( .D(n701), .E(n600), .CP(ChipClock), .Q(
        \Storage[18][11] ) );
  EDFQD1 \Storage_reg[17][32]  ( .D(n657), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][32] ) );
  EDFQD1 \Storage_reg[17][31]  ( .D(n761), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][31] ) );
  EDFQD1 \Storage_reg[17][30]  ( .D(n758), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][30] ) );
  EDFQD1 \Storage_reg[17][29]  ( .D(n755), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][29] ) );
  EDFQD1 \Storage_reg[17][28]  ( .D(n752), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][28] ) );
  EDFQD1 \Storage_reg[17][27]  ( .D(n749), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][27] ) );
  EDFQD1 \Storage_reg[17][26]  ( .D(n746), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][26] ) );
  EDFQD1 \Storage_reg[17][25]  ( .D(n743), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][25] ) );
  EDFQD1 \Storage_reg[17][24]  ( .D(n740), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][24] ) );
  EDFQD1 \Storage_reg[17][23]  ( .D(n737), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][23] ) );
  EDFQD1 \Storage_reg[17][22]  ( .D(n734), .E(n602), .CP(ChipClock), .Q(
        \Storage[17][22] ) );
  EDFQD1 \Storage_reg[17][21]  ( .D(n731), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][21] ) );
  EDFQD1 \Storage_reg[17][20]  ( .D(n728), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][20] ) );
  EDFQD1 \Storage_reg[17][19]  ( .D(n725), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][19] ) );
  EDFQD1 \Storage_reg[17][18]  ( .D(n722), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][18] ) );
  EDFQD1 \Storage_reg[17][17]  ( .D(n719), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][17] ) );
  EDFQD1 \Storage_reg[17][16]  ( .D(n716), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][16] ) );
  EDFQD1 \Storage_reg[17][15]  ( .D(n713), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][15] ) );
  EDFQD1 \Storage_reg[17][14]  ( .D(n710), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][14] ) );
  EDFQD1 \Storage_reg[17][13]  ( .D(n707), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][13] ) );
  EDFQD1 \Storage_reg[17][12]  ( .D(n704), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][12] ) );
  EDFQD1 \Storage_reg[17][11]  ( .D(n701), .E(n603), .CP(ChipClock), .Q(
        \Storage[17][11] ) );
  EDFQD1 \Storage_reg[14][32]  ( .D(n657), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][32] ) );
  EDFQD1 \Storage_reg[14][31]  ( .D(n761), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][31] ) );
  EDFQD1 \Storage_reg[14][30]  ( .D(n758), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][30] ) );
  EDFQD1 \Storage_reg[14][29]  ( .D(n755), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][29] ) );
  EDFQD1 \Storage_reg[14][28]  ( .D(n752), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][28] ) );
  EDFQD1 \Storage_reg[14][27]  ( .D(n749), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][27] ) );
  EDFQD1 \Storage_reg[14][26]  ( .D(n746), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][26] ) );
  EDFQD1 \Storage_reg[14][25]  ( .D(n743), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][25] ) );
  EDFQD1 \Storage_reg[14][24]  ( .D(n740), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][24] ) );
  EDFQD1 \Storage_reg[14][23]  ( .D(n737), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][23] ) );
  EDFQD1 \Storage_reg[14][22]  ( .D(n734), .E(n611), .CP(ChipClock), .Q(
        \Storage[14][22] ) );
  EDFQD1 \Storage_reg[14][21]  ( .D(n731), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][21] ) );
  EDFQD1 \Storage_reg[14][20]  ( .D(n728), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][20] ) );
  EDFQD1 \Storage_reg[14][19]  ( .D(n725), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][19] ) );
  EDFQD1 \Storage_reg[14][18]  ( .D(n722), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][18] ) );
  EDFQD1 \Storage_reg[14][17]  ( .D(n719), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][17] ) );
  EDFQD1 \Storage_reg[14][16]  ( .D(n716), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][16] ) );
  EDFQD1 \Storage_reg[14][15]  ( .D(n713), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][15] ) );
  EDFQD1 \Storage_reg[14][14]  ( .D(n710), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][14] ) );
  EDFQD1 \Storage_reg[14][13]  ( .D(n707), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][13] ) );
  EDFQD1 \Storage_reg[14][12]  ( .D(n704), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][12] ) );
  EDFQD1 \Storage_reg[14][11]  ( .D(n701), .E(n612), .CP(ChipClock), .Q(
        \Storage[14][11] ) );
  EDFQD1 \Storage_reg[13][32]  ( .D(n657), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][32] ) );
  EDFQD1 \Storage_reg[13][31]  ( .D(n761), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][31] ) );
  EDFQD1 \Storage_reg[13][30]  ( .D(n757), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][30] ) );
  EDFQD1 \Storage_reg[13][29]  ( .D(n754), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][29] ) );
  EDFQD1 \Storage_reg[13][28]  ( .D(n752), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][28] ) );
  EDFQD1 \Storage_reg[13][27]  ( .D(n749), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][27] ) );
  EDFQD1 \Storage_reg[13][26]  ( .D(n745), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][26] ) );
  EDFQD1 \Storage_reg[13][25]  ( .D(n742), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][25] ) );
  EDFQD1 \Storage_reg[13][24]  ( .D(n740), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][24] ) );
  EDFQD1 \Storage_reg[13][23]  ( .D(n737), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][23] ) );
  EDFQD1 \Storage_reg[13][22]  ( .D(n733), .E(n614), .CP(ChipClock), .Q(
        \Storage[13][22] ) );
  EDFQD1 \Storage_reg[13][21]  ( .D(n730), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][21] ) );
  EDFQD1 \Storage_reg[13][20]  ( .D(n728), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][20] ) );
  EDFQD1 \Storage_reg[13][19]  ( .D(n725), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][19] ) );
  EDFQD1 \Storage_reg[13][18]  ( .D(n721), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][18] ) );
  EDFQD1 \Storage_reg[13][17]  ( .D(n718), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][17] ) );
  EDFQD1 \Storage_reg[13][16]  ( .D(n716), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][16] ) );
  EDFQD1 \Storage_reg[13][15]  ( .D(n712), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][15] ) );
  EDFQD1 \Storage_reg[13][14]  ( .D(n709), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][14] ) );
  EDFQD1 \Storage_reg[13][13]  ( .D(n707), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][13] ) );
  EDFQD1 \Storage_reg[13][12]  ( .D(n704), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][12] ) );
  EDFQD1 \Storage_reg[13][11]  ( .D(n700), .E(n615), .CP(ChipClock), .Q(
        \Storage[13][11] ) );
  EDFQD1 \Storage_reg[10][32]  ( .D(n657), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][32] ) );
  EDFQD1 \Storage_reg[10][31]  ( .D(n760), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][31] ) );
  EDFQD1 \Storage_reg[10][30]  ( .D(n757), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][30] ) );
  EDFQD1 \Storage_reg[10][29]  ( .D(n754), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][29] ) );
  EDFQD1 \Storage_reg[10][28]  ( .D(n751), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][28] ) );
  EDFQD1 \Storage_reg[10][27]  ( .D(n748), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][27] ) );
  EDFQD1 \Storage_reg[10][26]  ( .D(n745), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][26] ) );
  EDFQD1 \Storage_reg[10][25]  ( .D(n742), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][25] ) );
  EDFQD1 \Storage_reg[10][24]  ( .D(n739), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][24] ) );
  EDFQD1 \Storage_reg[10][23]  ( .D(n736), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][23] ) );
  EDFQD1 \Storage_reg[10][22]  ( .D(n733), .E(n623), .CP(ChipClock), .Q(
        \Storage[10][22] ) );
  EDFQD1 \Storage_reg[10][21]  ( .D(n730), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][21] ) );
  EDFQD1 \Storage_reg[10][20]  ( .D(n727), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][20] ) );
  EDFQD1 \Storage_reg[10][19]  ( .D(n724), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][19] ) );
  EDFQD1 \Storage_reg[10][18]  ( .D(n721), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][18] ) );
  EDFQD1 \Storage_reg[10][17]  ( .D(n718), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][17] ) );
  EDFQD1 \Storage_reg[10][16]  ( .D(n715), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][16] ) );
  EDFQD1 \Storage_reg[10][15]  ( .D(n712), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][15] ) );
  EDFQD1 \Storage_reg[10][14]  ( .D(n709), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][14] ) );
  EDFQD1 \Storage_reg[10][13]  ( .D(n706), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][13] ) );
  EDFQD1 \Storage_reg[10][12]  ( .D(n703), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][12] ) );
  EDFQD1 \Storage_reg[10][11]  ( .D(n700), .E(n624), .CP(ChipClock), .Q(
        \Storage[10][11] ) );
  EDFQD1 \Storage_reg[9][32]  ( .D(n658), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][32] ) );
  EDFQD1 \Storage_reg[9][31]  ( .D(n760), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][31] ) );
  EDFQD1 \Storage_reg[9][30]  ( .D(n757), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][30] ) );
  EDFQD1 \Storage_reg[9][29]  ( .D(n754), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][29] ) );
  EDFQD1 \Storage_reg[9][28]  ( .D(n751), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][28] ) );
  EDFQD1 \Storage_reg[9][27]  ( .D(n748), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][27] ) );
  EDFQD1 \Storage_reg[9][26]  ( .D(n745), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][26] ) );
  EDFQD1 \Storage_reg[9][25]  ( .D(n742), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][25] ) );
  EDFQD1 \Storage_reg[9][24]  ( .D(n739), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][24] ) );
  EDFQD1 \Storage_reg[9][23]  ( .D(n736), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][23] ) );
  EDFQD1 \Storage_reg[9][22]  ( .D(n733), .E(n626), .CP(ChipClock), .Q(
        \Storage[9][22] ) );
  EDFQD1 \Storage_reg[9][21]  ( .D(n730), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][21] ) );
  EDFQD1 \Storage_reg[9][20]  ( .D(n727), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][20] ) );
  EDFQD1 \Storage_reg[9][19]  ( .D(n724), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][19] ) );
  EDFQD1 \Storage_reg[9][18]  ( .D(n721), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][18] ) );
  EDFQD1 \Storage_reg[9][17]  ( .D(n718), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][17] ) );
  EDFQD1 \Storage_reg[9][16]  ( .D(n715), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][16] ) );
  EDFQD1 \Storage_reg[9][15]  ( .D(n712), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][15] ) );
  EDFQD1 \Storage_reg[9][14]  ( .D(n709), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][14] ) );
  EDFQD1 \Storage_reg[9][13]  ( .D(n706), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][13] ) );
  EDFQD1 \Storage_reg[9][12]  ( .D(n703), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][12] ) );
  EDFQD1 \Storage_reg[9][11]  ( .D(n700), .E(n627), .CP(ChipClock), .Q(
        \Storage[9][11] ) );
  EDFQD1 \Storage_reg[6][32]  ( .D(n658), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][32] ) );
  EDFQD1 \Storage_reg[6][31]  ( .D(n760), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][31] ) );
  EDFQD1 \Storage_reg[6][30]  ( .D(n757), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][30] ) );
  EDFQD1 \Storage_reg[6][29]  ( .D(n754), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][29] ) );
  EDFQD1 \Storage_reg[6][28]  ( .D(n751), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][28] ) );
  EDFQD1 \Storage_reg[6][27]  ( .D(n748), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][27] ) );
  EDFQD1 \Storage_reg[6][26]  ( .D(n745), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][26] ) );
  EDFQD1 \Storage_reg[6][25]  ( .D(n742), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][25] ) );
  EDFQD1 \Storage_reg[6][24]  ( .D(n739), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][24] ) );
  EDFQD1 \Storage_reg[6][23]  ( .D(n736), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][23] ) );
  EDFQD1 \Storage_reg[6][22]  ( .D(n733), .E(n635), .CP(ChipClock), .Q(
        \Storage[6][22] ) );
  EDFQD1 \Storage_reg[6][21]  ( .D(n730), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][21] ) );
  EDFQD1 \Storage_reg[6][20]  ( .D(n727), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][20] ) );
  EDFQD1 \Storage_reg[6][19]  ( .D(n724), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][19] ) );
  EDFQD1 \Storage_reg[6][18]  ( .D(n721), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][18] ) );
  EDFQD1 \Storage_reg[6][17]  ( .D(n718), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][17] ) );
  EDFQD1 \Storage_reg[6][16]  ( .D(n715), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][16] ) );
  EDFQD1 \Storage_reg[6][15]  ( .D(n712), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][15] ) );
  EDFQD1 \Storage_reg[6][14]  ( .D(n709), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][14] ) );
  EDFQD1 \Storage_reg[6][13]  ( .D(n706), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][13] ) );
  EDFQD1 \Storage_reg[6][12]  ( .D(n703), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][12] ) );
  EDFQD1 \Storage_reg[6][11]  ( .D(n700), .E(n636), .CP(ChipClock), .Q(
        \Storage[6][11] ) );
  EDFQD1 \Storage_reg[5][32]  ( .D(n658), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][32] ) );
  EDFQD1 \Storage_reg[5][31]  ( .D(n760), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][31] ) );
  EDFQD1 \Storage_reg[5][30]  ( .D(n757), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][30] ) );
  EDFQD1 \Storage_reg[5][29]  ( .D(n754), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][29] ) );
  EDFQD1 \Storage_reg[5][28]  ( .D(n751), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][28] ) );
  EDFQD1 \Storage_reg[5][27]  ( .D(n748), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][27] ) );
  EDFQD1 \Storage_reg[5][26]  ( .D(n745), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][26] ) );
  EDFQD1 \Storage_reg[5][25]  ( .D(n742), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][25] ) );
  EDFQD1 \Storage_reg[5][24]  ( .D(n739), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][24] ) );
  EDFQD1 \Storage_reg[5][23]  ( .D(n736), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][23] ) );
  EDFQD1 \Storage_reg[5][22]  ( .D(n733), .E(n638), .CP(ChipClock), .Q(
        \Storage[5][22] ) );
  EDFQD1 \Storage_reg[5][21]  ( .D(n730), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][21] ) );
  EDFQD1 \Storage_reg[5][20]  ( .D(n727), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][20] ) );
  EDFQD1 \Storage_reg[5][19]  ( .D(n724), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][19] ) );
  EDFQD1 \Storage_reg[5][18]  ( .D(n721), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][18] ) );
  EDFQD1 \Storage_reg[5][17]  ( .D(n718), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][17] ) );
  EDFQD1 \Storage_reg[5][16]  ( .D(n715), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][16] ) );
  EDFQD1 \Storage_reg[5][15]  ( .D(n712), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][15] ) );
  EDFQD1 \Storage_reg[5][14]  ( .D(n709), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][14] ) );
  EDFQD1 \Storage_reg[5][13]  ( .D(n706), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][13] ) );
  EDFQD1 \Storage_reg[5][12]  ( .D(n703), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][12] ) );
  EDFQD1 \Storage_reg[5][11]  ( .D(n700), .E(n639), .CP(ChipClock), .Q(
        \Storage[5][11] ) );
  EDFQD1 \Storage_reg[2][32]  ( .D(n658), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][32] ) );
  EDFQD1 \Storage_reg[2][31]  ( .D(n760), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][31] ) );
  EDFQD1 \Storage_reg[2][30]  ( .D(n757), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][30] ) );
  EDFQD1 \Storage_reg[2][29]  ( .D(n754), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][29] ) );
  EDFQD1 \Storage_reg[2][28]  ( .D(n751), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][28] ) );
  EDFQD1 \Storage_reg[2][27]  ( .D(n748), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][27] ) );
  EDFQD1 \Storage_reg[2][26]  ( .D(n745), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][26] ) );
  EDFQD1 \Storage_reg[2][25]  ( .D(n742), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][25] ) );
  EDFQD1 \Storage_reg[2][24]  ( .D(n739), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][24] ) );
  EDFQD1 \Storage_reg[2][23]  ( .D(n736), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][23] ) );
  EDFQD1 \Storage_reg[2][22]  ( .D(n733), .E(n647), .CP(ChipClock), .Q(
        \Storage[2][22] ) );
  EDFQD1 \Storage_reg[2][21]  ( .D(n730), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][21] ) );
  EDFQD1 \Storage_reg[2][20]  ( .D(n727), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][20] ) );
  EDFQD1 \Storage_reg[2][19]  ( .D(n724), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][19] ) );
  EDFQD1 \Storage_reg[2][18]  ( .D(n721), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][18] ) );
  EDFQD1 \Storage_reg[2][17]  ( .D(n718), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][17] ) );
  EDFQD1 \Storage_reg[2][16]  ( .D(n715), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][16] ) );
  EDFQD1 \Storage_reg[2][15]  ( .D(n712), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][15] ) );
  EDFQD1 \Storage_reg[2][14]  ( .D(n709), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][14] ) );
  EDFQD1 \Storage_reg[2][13]  ( .D(n706), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][13] ) );
  EDFQD1 \Storage_reg[2][12]  ( .D(n703), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][12] ) );
  EDFQD1 \Storage_reg[2][11]  ( .D(n700), .E(n648), .CP(ChipClock), .Q(
        \Storage[2][11] ) );
  EDFQD1 \Storage_reg[1][32]  ( .D(n658), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][32] ) );
  EDFQD1 \Storage_reg[1][31]  ( .D(n760), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][31] ) );
  EDFQD1 \Storage_reg[1][30]  ( .D(n757), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][30] ) );
  EDFQD1 \Storage_reg[1][29]  ( .D(n754), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][29] ) );
  EDFQD1 \Storage_reg[1][28]  ( .D(n751), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][28] ) );
  EDFQD1 \Storage_reg[1][27]  ( .D(n748), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][27] ) );
  EDFQD1 \Storage_reg[1][26]  ( .D(n745), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][26] ) );
  EDFQD1 \Storage_reg[1][25]  ( .D(n742), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][25] ) );
  EDFQD1 \Storage_reg[1][24]  ( .D(n739), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][24] ) );
  EDFQD1 \Storage_reg[1][23]  ( .D(n736), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][23] ) );
  EDFQD1 \Storage_reg[1][22]  ( .D(n733), .E(n650), .CP(ChipClock), .Q(
        \Storage[1][22] ) );
  EDFQD1 \Storage_reg[1][21]  ( .D(n730), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][21] ) );
  EDFQD1 \Storage_reg[1][20]  ( .D(n727), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][20] ) );
  EDFQD1 \Storage_reg[1][19]  ( .D(n724), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][19] ) );
  EDFQD1 \Storage_reg[1][18]  ( .D(n721), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][18] ) );
  EDFQD1 \Storage_reg[1][17]  ( .D(n718), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][17] ) );
  EDFQD1 \Storage_reg[1][16]  ( .D(n715), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][16] ) );
  EDFQD1 \Storage_reg[1][15]  ( .D(n712), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][15] ) );
  EDFQD1 \Storage_reg[1][14]  ( .D(n709), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][14] ) );
  EDFQD1 \Storage_reg[1][13]  ( .D(n706), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][13] ) );
  EDFQD1 \Storage_reg[1][12]  ( .D(n703), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][12] ) );
  EDFQD1 \Storage_reg[1][11]  ( .D(n700), .E(n651), .CP(ChipClock), .Q(
        \Storage[1][11] ) );
  EDFQD1 \Storage_reg[23][32]  ( .D(n656), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][32] ) );
  EDFQD1 \Storage_reg[23][31]  ( .D(n761), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][31] ) );
  EDFQD1 \Storage_reg[23][30]  ( .D(n758), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][30] ) );
  EDFQD1 \Storage_reg[23][29]  ( .D(n755), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][29] ) );
  EDFQD1 \Storage_reg[23][28]  ( .D(n752), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][28] ) );
  EDFQD1 \Storage_reg[23][27]  ( .D(n749), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][27] ) );
  EDFQD1 \Storage_reg[23][26]  ( .D(n746), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][26] ) );
  EDFQD1 \Storage_reg[23][25]  ( .D(n743), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][25] ) );
  EDFQD1 \Storage_reg[23][24]  ( .D(n740), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][24] ) );
  EDFQD1 \Storage_reg[23][23]  ( .D(n737), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][23] ) );
  EDFQD1 \Storage_reg[23][22]  ( .D(n734), .E(n584), .CP(ChipClock), .Q(
        \Storage[23][22] ) );
  EDFQD1 \Storage_reg[23][21]  ( .D(n731), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][21] ) );
  EDFQD1 \Storage_reg[23][20]  ( .D(n728), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][20] ) );
  EDFQD1 \Storage_reg[23][19]  ( .D(n725), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][19] ) );
  EDFQD1 \Storage_reg[23][18]  ( .D(n722), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][18] ) );
  EDFQD1 \Storage_reg[23][17]  ( .D(n719), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][17] ) );
  EDFQD1 \Storage_reg[23][16]  ( .D(n716), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][16] ) );
  EDFQD1 \Storage_reg[23][15]  ( .D(n713), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][15] ) );
  EDFQD1 \Storage_reg[23][14]  ( .D(n710), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][14] ) );
  EDFQD1 \Storage_reg[23][13]  ( .D(n707), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][13] ) );
  EDFQD1 \Storage_reg[23][12]  ( .D(n704), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][12] ) );
  EDFQD1 \Storage_reg[23][11]  ( .D(n701), .E(n585), .CP(ChipClock), .Q(
        \Storage[23][11] ) );
  EDFQD1 \Storage_reg[20][32]  ( .D(n657), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][32] ) );
  EDFQD1 \Storage_reg[20][31]  ( .D(n761), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][31] ) );
  EDFQD1 \Storage_reg[20][30]  ( .D(n758), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][30] ) );
  EDFQD1 \Storage_reg[20][29]  ( .D(n755), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][29] ) );
  EDFQD1 \Storage_reg[20][28]  ( .D(n752), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][28] ) );
  EDFQD1 \Storage_reg[20][27]  ( .D(n749), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][27] ) );
  EDFQD1 \Storage_reg[20][26]  ( .D(n746), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][26] ) );
  EDFQD1 \Storage_reg[20][25]  ( .D(n743), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][25] ) );
  EDFQD1 \Storage_reg[20][24]  ( .D(n740), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][24] ) );
  EDFQD1 \Storage_reg[20][23]  ( .D(n737), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][23] ) );
  EDFQD1 \Storage_reg[20][22]  ( .D(n734), .E(n593), .CP(ChipClock), .Q(
        \Storage[20][22] ) );
  EDFQD1 \Storage_reg[20][21]  ( .D(n731), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][21] ) );
  EDFQD1 \Storage_reg[20][20]  ( .D(n728), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][20] ) );
  EDFQD1 \Storage_reg[20][19]  ( .D(n725), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][19] ) );
  EDFQD1 \Storage_reg[20][18]  ( .D(n722), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][18] ) );
  EDFQD1 \Storage_reg[20][17]  ( .D(n719), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][17] ) );
  EDFQD1 \Storage_reg[20][16]  ( .D(n716), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][16] ) );
  EDFQD1 \Storage_reg[20][15]  ( .D(n713), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][15] ) );
  EDFQD1 \Storage_reg[20][14]  ( .D(n710), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][14] ) );
  EDFQD1 \Storage_reg[20][13]  ( .D(n707), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][13] ) );
  EDFQD1 \Storage_reg[20][12]  ( .D(n704), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][12] ) );
  EDFQD1 \Storage_reg[20][11]  ( .D(n701), .E(n594), .CP(ChipClock), .Q(
        \Storage[20][11] ) );
  EDFQD1 \Storage_reg[19][32]  ( .D(n657), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][32] ) );
  EDFQD1 \Storage_reg[19][31]  ( .D(n761), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][31] ) );
  EDFQD1 \Storage_reg[19][30]  ( .D(n758), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][30] ) );
  EDFQD1 \Storage_reg[19][29]  ( .D(n755), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][29] ) );
  EDFQD1 \Storage_reg[19][28]  ( .D(n752), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][28] ) );
  EDFQD1 \Storage_reg[19][27]  ( .D(n749), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][27] ) );
  EDFQD1 \Storage_reg[19][26]  ( .D(n746), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][26] ) );
  EDFQD1 \Storage_reg[19][25]  ( .D(n743), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][25] ) );
  EDFQD1 \Storage_reg[19][24]  ( .D(n740), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][24] ) );
  EDFQD1 \Storage_reg[19][23]  ( .D(n737), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][23] ) );
  EDFQD1 \Storage_reg[19][22]  ( .D(n734), .E(n596), .CP(ChipClock), .Q(
        \Storage[19][22] ) );
  EDFQD1 \Storage_reg[19][21]  ( .D(n731), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][21] ) );
  EDFQD1 \Storage_reg[19][20]  ( .D(n728), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][20] ) );
  EDFQD1 \Storage_reg[19][19]  ( .D(n725), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][19] ) );
  EDFQD1 \Storage_reg[19][18]  ( .D(n722), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][18] ) );
  EDFQD1 \Storage_reg[19][17]  ( .D(n719), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][17] ) );
  EDFQD1 \Storage_reg[19][16]  ( .D(n716), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][16] ) );
  EDFQD1 \Storage_reg[19][15]  ( .D(n713), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][15] ) );
  EDFQD1 \Storage_reg[19][14]  ( .D(n710), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][14] ) );
  EDFQD1 \Storage_reg[19][13]  ( .D(n707), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][13] ) );
  EDFQD1 \Storage_reg[19][12]  ( .D(n704), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][12] ) );
  EDFQD1 \Storage_reg[19][11]  ( .D(n701), .E(n597), .CP(ChipClock), .Q(
        \Storage[19][11] ) );
  EDFQD1 \Storage_reg[16][32]  ( .D(n657), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][32] ) );
  EDFQD1 \Storage_reg[16][31]  ( .D(n761), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][31] ) );
  EDFQD1 \Storage_reg[16][30]  ( .D(n758), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][30] ) );
  EDFQD1 \Storage_reg[16][29]  ( .D(n755), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][29] ) );
  EDFQD1 \Storage_reg[16][28]  ( .D(n752), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][28] ) );
  EDFQD1 \Storage_reg[16][27]  ( .D(n749), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][27] ) );
  EDFQD1 \Storage_reg[16][26]  ( .D(n746), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][26] ) );
  EDFQD1 \Storage_reg[16][25]  ( .D(n743), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][25] ) );
  EDFQD1 \Storage_reg[16][24]  ( .D(n740), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][24] ) );
  EDFQD1 \Storage_reg[16][23]  ( .D(n737), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][23] ) );
  EDFQD1 \Storage_reg[16][22]  ( .D(n734), .E(n605), .CP(ChipClock), .Q(
        \Storage[16][22] ) );
  EDFQD1 \Storage_reg[16][21]  ( .D(n731), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][21] ) );
  EDFQD1 \Storage_reg[16][20]  ( .D(n728), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][20] ) );
  EDFQD1 \Storage_reg[16][19]  ( .D(n725), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][19] ) );
  EDFQD1 \Storage_reg[16][18]  ( .D(n722), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][18] ) );
  EDFQD1 \Storage_reg[16][17]  ( .D(n719), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][17] ) );
  EDFQD1 \Storage_reg[16][16]  ( .D(n716), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][16] ) );
  EDFQD1 \Storage_reg[16][15]  ( .D(n713), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][15] ) );
  EDFQD1 \Storage_reg[16][14]  ( .D(n710), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][14] ) );
  EDFQD1 \Storage_reg[16][13]  ( .D(n707), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][13] ) );
  EDFQD1 \Storage_reg[16][12]  ( .D(n704), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][12] ) );
  EDFQD1 \Storage_reg[16][11]  ( .D(n701), .E(n606), .CP(ChipClock), .Q(
        \Storage[16][11] ) );
  EDFQD1 \Storage_reg[15][32]  ( .D(n657), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][32] ) );
  EDFQD1 \Storage_reg[15][31]  ( .D(n761), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][31] ) );
  EDFQD1 \Storage_reg[15][30]  ( .D(n758), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][30] ) );
  EDFQD1 \Storage_reg[15][29]  ( .D(n755), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][29] ) );
  EDFQD1 \Storage_reg[15][28]  ( .D(n752), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][28] ) );
  EDFQD1 \Storage_reg[15][27]  ( .D(n749), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][27] ) );
  EDFQD1 \Storage_reg[15][26]  ( .D(n746), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][26] ) );
  EDFQD1 \Storage_reg[15][25]  ( .D(n743), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][25] ) );
  EDFQD1 \Storage_reg[15][24]  ( .D(n740), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][24] ) );
  EDFQD1 \Storage_reg[15][23]  ( .D(n737), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][23] ) );
  EDFQD1 \Storage_reg[15][22]  ( .D(n734), .E(n608), .CP(ChipClock), .Q(
        \Storage[15][22] ) );
  EDFQD1 \Storage_reg[15][21]  ( .D(n731), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][21] ) );
  EDFQD1 \Storage_reg[15][20]  ( .D(n728), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][20] ) );
  EDFQD1 \Storage_reg[15][19]  ( .D(n725), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][19] ) );
  EDFQD1 \Storage_reg[15][18]  ( .D(n722), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][18] ) );
  EDFQD1 \Storage_reg[15][17]  ( .D(n719), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][17] ) );
  EDFQD1 \Storage_reg[15][16]  ( .D(n716), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][16] ) );
  EDFQD1 \Storage_reg[15][15]  ( .D(n713), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][15] ) );
  EDFQD1 \Storage_reg[15][14]  ( .D(n710), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][14] ) );
  EDFQD1 \Storage_reg[15][13]  ( .D(n707), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][13] ) );
  EDFQD1 \Storage_reg[15][12]  ( .D(n704), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][12] ) );
  EDFQD1 \Storage_reg[15][11]  ( .D(n701), .E(n609), .CP(ChipClock), .Q(
        \Storage[15][11] ) );
  EDFQD1 \Storage_reg[12][32]  ( .D(n657), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][32] ) );
  EDFQD1 \Storage_reg[12][31]  ( .D(n761), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][31] ) );
  EDFQD1 \Storage_reg[12][30]  ( .D(n757), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][30] ) );
  EDFQD1 \Storage_reg[12][29]  ( .D(n754), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][29] ) );
  EDFQD1 \Storage_reg[12][28]  ( .D(n752), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][28] ) );
  EDFQD1 \Storage_reg[12][27]  ( .D(n749), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][27] ) );
  EDFQD1 \Storage_reg[12][26]  ( .D(n745), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][26] ) );
  EDFQD1 \Storage_reg[12][25]  ( .D(n742), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][25] ) );
  EDFQD1 \Storage_reg[12][24]  ( .D(n740), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][24] ) );
  EDFQD1 \Storage_reg[12][23]  ( .D(n737), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][23] ) );
  EDFQD1 \Storage_reg[12][22]  ( .D(n733), .E(n617), .CP(ChipClock), .Q(
        \Storage[12][22] ) );
  EDFQD1 \Storage_reg[12][21]  ( .D(n730), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][21] ) );
  EDFQD1 \Storage_reg[12][20]  ( .D(n728), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][20] ) );
  EDFQD1 \Storage_reg[12][19]  ( .D(n725), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][19] ) );
  EDFQD1 \Storage_reg[12][18]  ( .D(n721), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][18] ) );
  EDFQD1 \Storage_reg[12][17]  ( .D(n718), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][17] ) );
  EDFQD1 \Storage_reg[12][16]  ( .D(n716), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][16] ) );
  EDFQD1 \Storage_reg[12][15]  ( .D(n712), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][15] ) );
  EDFQD1 \Storage_reg[12][14]  ( .D(n709), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][14] ) );
  EDFQD1 \Storage_reg[12][13]  ( .D(n707), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][13] ) );
  EDFQD1 \Storage_reg[12][12]  ( .D(n704), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][12] ) );
  EDFQD1 \Storage_reg[12][11]  ( .D(n700), .E(n618), .CP(ChipClock), .Q(
        \Storage[12][11] ) );
  EDFQD1 \Storage_reg[11][32]  ( .D(n657), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][32] ) );
  EDFQD1 \Storage_reg[11][31]  ( .D(n760), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][31] ) );
  EDFQD1 \Storage_reg[11][30]  ( .D(n757), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][30] ) );
  EDFQD1 \Storage_reg[11][29]  ( .D(n754), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][29] ) );
  EDFQD1 \Storage_reg[11][28]  ( .D(n751), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][28] ) );
  EDFQD1 \Storage_reg[11][27]  ( .D(n748), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][27] ) );
  EDFQD1 \Storage_reg[11][26]  ( .D(n745), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][26] ) );
  EDFQD1 \Storage_reg[11][25]  ( .D(n742), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][25] ) );
  EDFQD1 \Storage_reg[11][24]  ( .D(n739), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][24] ) );
  EDFQD1 \Storage_reg[11][23]  ( .D(n736), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][23] ) );
  EDFQD1 \Storage_reg[11][22]  ( .D(n733), .E(n620), .CP(ChipClock), .Q(
        \Storage[11][22] ) );
  EDFQD1 \Storage_reg[11][21]  ( .D(n730), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][21] ) );
  EDFQD1 \Storage_reg[11][20]  ( .D(n727), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][20] ) );
  EDFQD1 \Storage_reg[11][19]  ( .D(n724), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][19] ) );
  EDFQD1 \Storage_reg[11][18]  ( .D(n721), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][18] ) );
  EDFQD1 \Storage_reg[11][17]  ( .D(n718), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][17] ) );
  EDFQD1 \Storage_reg[11][16]  ( .D(n715), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][16] ) );
  EDFQD1 \Storage_reg[11][15]  ( .D(n712), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][15] ) );
  EDFQD1 \Storage_reg[11][14]  ( .D(n709), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][14] ) );
  EDFQD1 \Storage_reg[11][13]  ( .D(n706), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][13] ) );
  EDFQD1 \Storage_reg[11][12]  ( .D(n703), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][12] ) );
  EDFQD1 \Storage_reg[11][11]  ( .D(n700), .E(n621), .CP(ChipClock), .Q(
        \Storage[11][11] ) );
  EDFQD1 \Storage_reg[8][32]  ( .D(n658), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][32] ) );
  EDFQD1 \Storage_reg[8][31]  ( .D(n760), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][31] ) );
  EDFQD1 \Storage_reg[8][30]  ( .D(n757), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][30] ) );
  EDFQD1 \Storage_reg[8][29]  ( .D(n754), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][29] ) );
  EDFQD1 \Storage_reg[8][28]  ( .D(n751), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][28] ) );
  EDFQD1 \Storage_reg[8][27]  ( .D(n748), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][27] ) );
  EDFQD1 \Storage_reg[8][26]  ( .D(n745), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][26] ) );
  EDFQD1 \Storage_reg[8][25]  ( .D(n742), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][25] ) );
  EDFQD1 \Storage_reg[8][24]  ( .D(n739), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][24] ) );
  EDFQD1 \Storage_reg[8][23]  ( .D(n736), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][23] ) );
  EDFQD1 \Storage_reg[8][22]  ( .D(n733), .E(n629), .CP(ChipClock), .Q(
        \Storage[8][22] ) );
  EDFQD1 \Storage_reg[8][21]  ( .D(n730), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][21] ) );
  EDFQD1 \Storage_reg[8][20]  ( .D(n727), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][20] ) );
  EDFQD1 \Storage_reg[8][19]  ( .D(n724), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][19] ) );
  EDFQD1 \Storage_reg[8][18]  ( .D(n721), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][18] ) );
  EDFQD1 \Storage_reg[8][17]  ( .D(n718), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][17] ) );
  EDFQD1 \Storage_reg[8][16]  ( .D(n715), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][16] ) );
  EDFQD1 \Storage_reg[8][15]  ( .D(n712), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][15] ) );
  EDFQD1 \Storage_reg[8][14]  ( .D(n709), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][14] ) );
  EDFQD1 \Storage_reg[8][13]  ( .D(n706), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][13] ) );
  EDFQD1 \Storage_reg[8][12]  ( .D(n703), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][12] ) );
  EDFQD1 \Storage_reg[8][11]  ( .D(n700), .E(n630), .CP(ChipClock), .Q(
        \Storage[8][11] ) );
  EDFQD1 \Storage_reg[7][32]  ( .D(n658), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][32] ) );
  EDFQD1 \Storage_reg[7][31]  ( .D(n760), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][31] ) );
  EDFQD1 \Storage_reg[7][30]  ( .D(n757), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][30] ) );
  EDFQD1 \Storage_reg[7][29]  ( .D(n754), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][29] ) );
  EDFQD1 \Storage_reg[7][28]  ( .D(n751), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][28] ) );
  EDFQD1 \Storage_reg[7][27]  ( .D(n748), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][27] ) );
  EDFQD1 \Storage_reg[7][26]  ( .D(n745), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][26] ) );
  EDFQD1 \Storage_reg[7][25]  ( .D(n742), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][25] ) );
  EDFQD1 \Storage_reg[7][24]  ( .D(n739), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][24] ) );
  EDFQD1 \Storage_reg[7][23]  ( .D(n736), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][23] ) );
  EDFQD1 \Storage_reg[7][22]  ( .D(n733), .E(n632), .CP(ChipClock), .Q(
        \Storage[7][22] ) );
  EDFQD1 \Storage_reg[7][21]  ( .D(n730), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][21] ) );
  EDFQD1 \Storage_reg[7][20]  ( .D(n727), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][20] ) );
  EDFQD1 \Storage_reg[7][19]  ( .D(n724), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][19] ) );
  EDFQD1 \Storage_reg[7][18]  ( .D(n721), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][18] ) );
  EDFQD1 \Storage_reg[7][17]  ( .D(n718), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][17] ) );
  EDFQD1 \Storage_reg[7][16]  ( .D(n715), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][16] ) );
  EDFQD1 \Storage_reg[7][15]  ( .D(n712), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][15] ) );
  EDFQD1 \Storage_reg[7][14]  ( .D(n709), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][14] ) );
  EDFQD1 \Storage_reg[7][13]  ( .D(n706), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][13] ) );
  EDFQD1 \Storage_reg[7][12]  ( .D(n703), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][12] ) );
  EDFQD1 \Storage_reg[7][11]  ( .D(n700), .E(n633), .CP(ChipClock), .Q(
        \Storage[7][11] ) );
  EDFQD1 \Storage_reg[4][32]  ( .D(n658), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][32] ) );
  EDFQD1 \Storage_reg[4][31]  ( .D(n760), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][31] ) );
  EDFQD1 \Storage_reg[4][30]  ( .D(n757), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][30] ) );
  EDFQD1 \Storage_reg[4][29]  ( .D(n754), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][29] ) );
  EDFQD1 \Storage_reg[4][28]  ( .D(n751), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][28] ) );
  EDFQD1 \Storage_reg[4][27]  ( .D(n748), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][27] ) );
  EDFQD1 \Storage_reg[4][26]  ( .D(n745), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][26] ) );
  EDFQD1 \Storage_reg[4][25]  ( .D(n742), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][25] ) );
  EDFQD1 \Storage_reg[4][24]  ( .D(n739), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][24] ) );
  EDFQD1 \Storage_reg[4][23]  ( .D(n736), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][23] ) );
  EDFQD1 \Storage_reg[4][22]  ( .D(n733), .E(n641), .CP(ChipClock), .Q(
        \Storage[4][22] ) );
  EDFQD1 \Storage_reg[4][21]  ( .D(n730), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][21] ) );
  EDFQD1 \Storage_reg[4][20]  ( .D(n727), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][20] ) );
  EDFQD1 \Storage_reg[4][19]  ( .D(n724), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][19] ) );
  EDFQD1 \Storage_reg[4][18]  ( .D(n721), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][18] ) );
  EDFQD1 \Storage_reg[4][17]  ( .D(n718), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][17] ) );
  EDFQD1 \Storage_reg[4][16]  ( .D(n715), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][16] ) );
  EDFQD1 \Storage_reg[4][15]  ( .D(n712), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][15] ) );
  EDFQD1 \Storage_reg[4][14]  ( .D(n709), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][14] ) );
  EDFQD1 \Storage_reg[4][13]  ( .D(n706), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][13] ) );
  EDFQD1 \Storage_reg[4][12]  ( .D(n703), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][12] ) );
  EDFQD1 \Storage_reg[4][11]  ( .D(n700), .E(n642), .CP(ChipClock), .Q(
        \Storage[4][11] ) );
  EDFQD1 \Storage_reg[3][32]  ( .D(n658), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][32] ) );
  EDFQD1 \Storage_reg[3][31]  ( .D(n760), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][31] ) );
  EDFQD1 \Storage_reg[3][30]  ( .D(n757), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][30] ) );
  EDFQD1 \Storage_reg[3][29]  ( .D(n754), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][29] ) );
  EDFQD1 \Storage_reg[3][28]  ( .D(n751), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][28] ) );
  EDFQD1 \Storage_reg[3][27]  ( .D(n748), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][27] ) );
  EDFQD1 \Storage_reg[3][26]  ( .D(n745), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][26] ) );
  EDFQD1 \Storage_reg[3][25]  ( .D(n742), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][25] ) );
  EDFQD1 \Storage_reg[3][24]  ( .D(n739), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][24] ) );
  EDFQD1 \Storage_reg[3][23]  ( .D(n736), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][23] ) );
  EDFQD1 \Storage_reg[3][22]  ( .D(n733), .E(n644), .CP(ChipClock), .Q(
        \Storage[3][22] ) );
  EDFQD1 \Storage_reg[3][21]  ( .D(n730), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][21] ) );
  EDFQD1 \Storage_reg[3][20]  ( .D(n727), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][20] ) );
  EDFQD1 \Storage_reg[3][19]  ( .D(n724), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][19] ) );
  EDFQD1 \Storage_reg[3][18]  ( .D(n721), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][18] ) );
  EDFQD1 \Storage_reg[3][17]  ( .D(n718), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][17] ) );
  EDFQD1 \Storage_reg[3][16]  ( .D(n715), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][16] ) );
  EDFQD1 \Storage_reg[3][15]  ( .D(n712), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][15] ) );
  EDFQD1 \Storage_reg[3][14]  ( .D(n709), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][14] ) );
  EDFQD1 \Storage_reg[3][13]  ( .D(n706), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][13] ) );
  EDFQD1 \Storage_reg[3][12]  ( .D(n703), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][12] ) );
  EDFQD1 \Storage_reg[3][11]  ( .D(n700), .E(n645), .CP(ChipClock), .Q(
        \Storage[3][11] ) );
  EDFQD1 \Storage_reg[0][32]  ( .D(n658), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][32] ) );
  EDFQD1 \Storage_reg[0][31]  ( .D(n760), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][31] ) );
  EDFQD1 \Storage_reg[0][30]  ( .D(n757), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][30] ) );
  EDFQD1 \Storage_reg[0][29]  ( .D(n754), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][29] ) );
  EDFQD1 \Storage_reg[0][28]  ( .D(n751), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][28] ) );
  EDFQD1 \Storage_reg[0][27]  ( .D(n748), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][27] ) );
  EDFQD1 \Storage_reg[0][26]  ( .D(n745), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][26] ) );
  EDFQD1 \Storage_reg[0][25]  ( .D(n742), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][25] ) );
  EDFQD1 \Storage_reg[0][24]  ( .D(n739), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][24] ) );
  EDFQD1 \Storage_reg[0][23]  ( .D(n736), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][23] ) );
  EDFQD1 \Storage_reg[0][22]  ( .D(n733), .E(n653), .CP(ChipClock), .Q(
        \Storage[0][22] ) );
  EDFQD1 \Storage_reg[0][21]  ( .D(n730), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][21] ) );
  EDFQD1 \Storage_reg[0][20]  ( .D(n727), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][20] ) );
  EDFQD1 \Storage_reg[0][19]  ( .D(n724), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][19] ) );
  EDFQD1 \Storage_reg[0][18]  ( .D(n721), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][18] ) );
  EDFQD1 \Storage_reg[0][17]  ( .D(n718), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][17] ) );
  EDFQD1 \Storage_reg[0][16]  ( .D(n715), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][16] ) );
  EDFQD1 \Storage_reg[0][15]  ( .D(n712), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][15] ) );
  EDFQD1 \Storage_reg[0][14]  ( .D(n709), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][14] ) );
  EDFQD1 \Storage_reg[0][13]  ( .D(n706), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][13] ) );
  EDFQD1 \Storage_reg[0][12]  ( .D(n703), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][12] ) );
  EDFQD1 \Storage_reg[0][11]  ( .D(n700), .E(n654), .CP(ChipClock), .Q(
        \Storage[0][11] ) );
  EDFQD1 \Storage_reg[31][32]  ( .D(n656), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][32] ) );
  EDFQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][31] ) );
  EDFQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][30] ) );
  EDFQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][29] ) );
  EDFQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][28] ) );
  EDFQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][27] ) );
  EDFQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][26] ) );
  EDFQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][25] ) );
  EDFQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][24] ) );
  EDFQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][23] ) );
  EDFQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(n560), .CP(ChipClock), .Q(
        \Storage[31][22] ) );
  EDFQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][21] ) );
  EDFQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][20] ) );
  EDFQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][19] ) );
  EDFQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][18] ) );
  EDFQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][17] ) );
  EDFQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][16] ) );
  EDFQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][15] ) );
  EDFQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][14] ) );
  EDFQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][13] ) );
  EDFQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][12] ) );
  EDFQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(n561), .CP(ChipClock), .Q(
        \Storage[31][11] ) );
  EDFQD1 ParityReg_reg ( .D(N84), .E(n558), .CP(ChipClock), .Q(ParityErr) );
  EDFQD1 \DataOreg_reg[21]  ( .D(N60), .E(n557), .CP(ChipClock), .Q(
        DataOreg[21]) );
  EDFQD1 \DataOreg_reg[20]  ( .D(N61), .E(n558), .CP(ChipClock), .Q(
        DataOreg[20]) );
  EDFQD1 \DataOreg_reg[5]  ( .D(N76), .E(n557), .CP(ChipClock), .Q(DataOreg[5]) );
  EDFQD1 \DataOreg_reg[1]  ( .D(N80), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[1]) );
  EDFQD1 \DataOreg_reg[31]  ( .D(N50), .E(n557), .CP(ChipClock), .Q(
        DataOreg[31]) );
  EDFQD1 \DataOreg_reg[30]  ( .D(N51), .E(n557), .CP(ChipClock), .Q(
        DataOreg[30]) );
  EDFQD1 \DataOreg_reg[29]  ( .D(N52), .E(n557), .CP(ChipClock), .Q(
        DataOreg[29]) );
  EDFQD1 \DataOreg_reg[28]  ( .D(N53), .E(n557), .CP(ChipClock), .Q(
        DataOreg[28]) );
  EDFQD1 \DataOreg_reg[27]  ( .D(N54), .E(n557), .CP(ChipClock), .Q(
        DataOreg[27]) );
  EDFQD1 \DataOreg_reg[26]  ( .D(N55), .E(n557), .CP(ChipClock), .Q(
        DataOreg[26]) );
  EDFQD1 \DataOreg_reg[25]  ( .D(N56), .E(n557), .CP(ChipClock), .Q(
        DataOreg[25]) );
  EDFQD1 \DataOreg_reg[24]  ( .D(N57), .E(n557), .CP(ChipClock), .Q(
        DataOreg[24]) );
  EDFQD1 \DataOreg_reg[23]  ( .D(N58), .E(n557), .CP(ChipClock), .Q(
        DataOreg[23]) );
  EDFQD1 \DataOreg_reg[22]  ( .D(N59), .E(n557), .CP(ChipClock), .Q(
        DataOreg[22]) );
  EDFQD1 \DataOreg_reg[19]  ( .D(N62), .E(n558), .CP(ChipClock), .Q(
        DataOreg[19]) );
  EDFQD1 \DataOreg_reg[18]  ( .D(N63), .E(n558), .CP(ChipClock), .Q(
        DataOreg[18]) );
  EDFQD1 \DataOreg_reg[17]  ( .D(N64), .E(n558), .CP(ChipClock), .Q(
        DataOreg[17]) );
  EDFQD1 \DataOreg_reg[16]  ( .D(N65), .E(n558), .CP(ChipClock), .Q(
        DataOreg[16]) );
  EDFQD1 \DataOreg_reg[15]  ( .D(N66), .E(n558), .CP(ChipClock), .Q(
        DataOreg[15]) );
  EDFQD1 \DataOreg_reg[14]  ( .D(N67), .E(n558), .CP(ChipClock), .Q(
        DataOreg[14]) );
  EDFQD1 \DataOreg_reg[13]  ( .D(N68), .E(n558), .CP(ChipClock), .Q(
        DataOreg[13]) );
  EDFQD1 \DataOreg_reg[12]  ( .D(N69), .E(n558), .CP(ChipClock), .Q(
        DataOreg[12]) );
  EDFQD1 \DataOreg_reg[11]  ( .D(N70), .E(n558), .CP(ChipClock), .Q(
        DataOreg[11]) );
  EDFQD1 \DataOreg_reg[10]  ( .D(N71), .E(n558), .CP(ChipClock), .Q(
        DataOreg[10]) );
  EDFQD1 \DataOreg_reg[8]  ( .D(N73), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[8]) );
  EDFQD1 \DataOreg_reg[7]  ( .D(N74), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[7]) );
  EDFQD1 \DataOreg_reg[6]  ( .D(N75), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[6]) );
  EDFQD1 \DataOreg_reg[4]  ( .D(N77), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[4]) );
  EDFQD1 \DataOreg_reg[3]  ( .D(N78), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[3]) );
  EDFQD1 \DataOreg_reg[2]  ( .D(N79), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[2]) );
  EDFQD1 \DataOreg_reg[0]  ( .D(N81), .E(N2262), .CP(ChipClock), .Q(
        DataOreg[0]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOreg[10]), .OE(n1), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOreg[31]), .OE(n1), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOreg[0]), .OE(n1), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOreg[30]), .OE(n1), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOreg[6]), .OE(n1), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOreg[8]), .OE(n659), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOreg[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOreg[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOreg[2]), .OE(n1), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOreg[29]), .OE(n1), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOreg[3]), .OE(n1), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOreg[28]), .OE(n1), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOreg[4]), .OE(n1), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOreg[27]), .OE(n1), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOreg[11]), .OE(n659), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOreg[26]), .OE(n1), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOreg[12]), .OE(n659), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOreg[25]), .OE(n659), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOreg[13]), .OE(n659), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOreg[24]), .OE(n1), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOreg[14]), .OE(n659), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOreg[23]), .OE(n1), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOreg[15]), .OE(n659), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOreg[22]), .OE(n1), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOreg[16]), .OE(n659), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOreg[19]), .OE(n659), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOreg[17]), .OE(n659), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOreg[18]), .OE(n659), .Z(DataO[18]) );
  BUFFD0 U2 ( .I(N43), .Z(n535) );
  BUFFD0 U3 ( .I(N43), .Z(n536) );
  BUFFD0 U4 ( .I(N46), .Z(n506) );
  INVD0 U5 ( .I(ChipEna), .ZN(n660) );
  INVD1 U6 ( .I(n660), .ZN(n659) );
  INVD1 U7 ( .I(n660), .ZN(n1) );
  INVD1 U8 ( .I(N2262), .ZN(n559) );
  INVD1 U9 ( .I(DataI[3]), .ZN(n678) );
  INVD1 U15 ( .I(DataI[7]), .ZN(n690) );
  INVD1 U16 ( .I(DataI[8]), .ZN(n693) );
  INVD1 U17 ( .I(DataI[10]), .ZN(n699) );
  INVD1 U20 ( .I(DataI[11]), .ZN(n702) );
  INVD1 U21 ( .I(DataI[12]), .ZN(n705) );
  INVD1 U22 ( .I(DataI[13]), .ZN(n708) );
  INVD1 U23 ( .I(DataI[14]), .ZN(n711) );
  INVD1 U28 ( .I(DataI[15]), .ZN(n714) );
  INVD1 U29 ( .I(DataI[16]), .ZN(n717) );
  INVD1 U30 ( .I(DataI[17]), .ZN(n720) );
  INVD1 U31 ( .I(DataI[18]), .ZN(n723) );
  INVD1 U32 ( .I(DataI[19]), .ZN(n726) );
  INVD1 U33 ( .I(DataI[20]), .ZN(n729) );
  INVD1 U34 ( .I(DataI[21]), .ZN(n732) );
  INVD1 U35 ( .I(DataI[22]), .ZN(n735) );
  INVD1 U36 ( .I(DataI[23]), .ZN(n738) );
  INVD1 U37 ( .I(DataI[24]), .ZN(n741) );
  INVD1 U38 ( .I(DataI[25]), .ZN(n744) );
  INVD1 U39 ( .I(DataI[26]), .ZN(n747) );
  INVD1 U40 ( .I(DataI[27]), .ZN(n750) );
  INVD1 U41 ( .I(DataI[28]), .ZN(n753) );
  INVD1 U42 ( .I(DataI[29]), .ZN(n756) );
  INVD1 U43 ( .I(DataI[30]), .ZN(n759) );
  INVD1 U44 ( .I(DataI[31]), .ZN(n762) );
  INVD1 U45 ( .I(DataI[0]), .ZN(n669) );
  INVD1 U46 ( .I(DataI[1]), .ZN(n672) );
  INVD1 U47 ( .I(DataI[2]), .ZN(n675) );
  INVD1 U48 ( .I(DataI[4]), .ZN(n681) );
  INVD1 U49 ( .I(DataI[5]), .ZN(n684) );
  INVD1 U50 ( .I(DataI[6]), .ZN(n687) );
  INVD1 U51 ( .I(DataI[9]), .ZN(n696) );
  BUFFD1 U52 ( .I(n540), .Z(n546) );
  BUFFD1 U53 ( .I(n540), .Z(n545) );
  BUFFD1 U54 ( .I(n541), .Z(n544) );
  BUFFD1 U55 ( .I(n541), .Z(n543) );
  BUFFD1 U56 ( .I(n519), .Z(n529) );
  BUFFD1 U57 ( .I(n520), .Z(n525) );
  BUFFD1 U58 ( .I(n520), .Z(n526) );
  BUFFD1 U59 ( .I(n520), .Z(n527) );
  BUFFD1 U60 ( .I(n519), .Z(n528) );
  BUFFD1 U61 ( .I(n541), .Z(n542) );
  BUFFD1 U62 ( .I(n540), .Z(n547) );
  BUFFD1 U63 ( .I(n537), .Z(n548) );
  BUFFD1 U64 ( .I(n538), .Z(n549) );
  BUFFD1 U65 ( .I(n541), .Z(n550) );
  BUFFD1 U66 ( .I(n539), .Z(n551) );
  BUFFD1 U67 ( .I(n539), .Z(n552) );
  BUFFD1 U68 ( .I(n539), .Z(n553) );
  BUFFD1 U69 ( .I(n538), .Z(n554) );
  BUFFD1 U70 ( .I(n538), .Z(n555) );
  BUFFD1 U71 ( .I(n538), .Z(n556) );
  BUFFD1 U72 ( .I(n519), .Z(n530) );
  BUFFD1 U73 ( .I(n518), .Z(n531) );
  BUFFD1 U74 ( .I(n518), .Z(n532) );
  BUFFD1 U75 ( .I(n517), .Z(n534) );
  BUFFD1 U76 ( .I(n518), .Z(n533) );
  BUFFD1 U77 ( .I(n521), .Z(n523) );
  BUFFD1 U78 ( .I(n521), .Z(n524) );
  BUFFD1 U79 ( .I(n521), .Z(n522) );
  INVD1 U80 ( .I(n2), .ZN(n657) );
  INVD1 U82 ( .I(n2), .ZN(n656) );
  INVD1 U83 ( .I(n2), .ZN(n658) );
  BUFFD1 U84 ( .I(n663), .Z(n514) );
  BUFFD1 U85 ( .I(n663), .Z(n515) );
  BUFFD1 U86 ( .I(n506), .Z(n504) );
  BUFFD1 U87 ( .I(n536), .Z(n537) );
  BUFFD1 U88 ( .I(n516), .Z(n520) );
  BUFFD1 U89 ( .I(n516), .Z(n519) );
  BUFFD1 U90 ( .I(n535), .Z(n540) );
  BUFFD1 U91 ( .I(n535), .Z(n541) );
  BUFFD1 U92 ( .I(n508), .Z(n513) );
  BUFFD1 U93 ( .I(n508), .Z(n512) );
  BUFFD1 U94 ( .I(n508), .Z(n511) );
  BUFFD1 U95 ( .I(n506), .Z(n505) );
  BUFFD1 U96 ( .I(n536), .Z(n539) );
  BUFFD1 U97 ( .I(n516), .Z(n518) );
  BUFFD1 U98 ( .I(n520), .Z(n517) );
  BUFFD1 U99 ( .I(n536), .Z(n538) );
  BUFFD1 U100 ( .I(n516), .Z(n521) );
  INVD1 U101 ( .I(n4), .ZN(n583) );
  INVD1 U102 ( .I(n4), .ZN(n582) );
  INVD1 U103 ( .I(n4), .ZN(n581) );
  INVD1 U104 ( .I(n5), .ZN(n580) );
  INVD1 U105 ( .I(n5), .ZN(n579) );
  INVD1 U106 ( .I(n5), .ZN(n578) );
  INVD1 U107 ( .I(n6), .ZN(n577) );
  INVD1 U108 ( .I(n6), .ZN(n576) );
  INVD1 U109 ( .I(n6), .ZN(n575) );
  INVD1 U110 ( .I(n7), .ZN(n574) );
  INVD1 U111 ( .I(n7), .ZN(n573) );
  INVD1 U112 ( .I(n7), .ZN(n572) );
  INVD1 U113 ( .I(n8), .ZN(n571) );
  INVD1 U114 ( .I(n8), .ZN(n570) );
  INVD1 U115 ( .I(n8), .ZN(n569) );
  INVD1 U116 ( .I(n9), .ZN(n568) );
  INVD1 U117 ( .I(n9), .ZN(n567) );
  INVD1 U118 ( .I(n9), .ZN(n566) );
  INVD1 U119 ( .I(n10), .ZN(n565) );
  INVD1 U120 ( .I(n10), .ZN(n564) );
  INVD1 U121 ( .I(n10), .ZN(n563) );
  INVD1 U122 ( .I(n11), .ZN(n562) );
  INVD1 U123 ( .I(n11), .ZN(n561) );
  INVD1 U124 ( .I(n11), .ZN(n560) );
  INVD1 U125 ( .I(n12), .ZN(n655) );
  INVD1 U126 ( .I(n12), .ZN(n654) );
  INVD1 U127 ( .I(n12), .ZN(n653) );
  INVD1 U128 ( .I(n13), .ZN(n652) );
  INVD1 U129 ( .I(n13), .ZN(n651) );
  INVD1 U130 ( .I(n13), .ZN(n650) );
  INVD1 U131 ( .I(n14), .ZN(n649) );
  INVD1 U132 ( .I(n14), .ZN(n648) );
  INVD1 U133 ( .I(n14), .ZN(n647) );
  INVD1 U134 ( .I(n15), .ZN(n646) );
  INVD1 U135 ( .I(n15), .ZN(n645) );
  INVD1 U136 ( .I(n15), .ZN(n644) );
  INVD1 U137 ( .I(n16), .ZN(n643) );
  INVD1 U138 ( .I(n16), .ZN(n642) );
  INVD1 U139 ( .I(n16), .ZN(n641) );
  INVD1 U140 ( .I(n17), .ZN(n640) );
  INVD1 U141 ( .I(n17), .ZN(n639) );
  INVD1 U142 ( .I(n17), .ZN(n638) );
  INVD1 U143 ( .I(n18), .ZN(n637) );
  INVD1 U144 ( .I(n18), .ZN(n636) );
  INVD1 U145 ( .I(n18), .ZN(n635) );
  INVD1 U146 ( .I(n19), .ZN(n634) );
  INVD1 U147 ( .I(n19), .ZN(n633) );
  INVD1 U148 ( .I(n19), .ZN(n632) );
  INVD1 U149 ( .I(n20), .ZN(n631) );
  INVD1 U150 ( .I(n20), .ZN(n630) );
  INVD1 U151 ( .I(n20), .ZN(n629) );
  INVD1 U152 ( .I(n21), .ZN(n628) );
  INVD1 U153 ( .I(n21), .ZN(n627) );
  INVD1 U154 ( .I(n21), .ZN(n626) );
  INVD1 U155 ( .I(n22), .ZN(n625) );
  INVD1 U156 ( .I(n22), .ZN(n624) );
  INVD1 U157 ( .I(n22), .ZN(n623) );
  INVD1 U158 ( .I(n23), .ZN(n622) );
  INVD1 U159 ( .I(n23), .ZN(n621) );
  INVD1 U160 ( .I(n23), .ZN(n620) );
  INVD1 U161 ( .I(n24), .ZN(n619) );
  INVD1 U162 ( .I(n24), .ZN(n618) );
  INVD1 U163 ( .I(n24), .ZN(n617) );
  INVD1 U164 ( .I(n25), .ZN(n616) );
  INVD1 U165 ( .I(n25), .ZN(n615) );
  INVD1 U166 ( .I(n25), .ZN(n614) );
  INVD1 U167 ( .I(n26), .ZN(n613) );
  INVD1 U168 ( .I(n26), .ZN(n612) );
  INVD1 U169 ( .I(n26), .ZN(n611) );
  INVD1 U170 ( .I(n27), .ZN(n610) );
  INVD1 U171 ( .I(n27), .ZN(n609) );
  INVD1 U172 ( .I(n27), .ZN(n608) );
  INVD1 U173 ( .I(n28), .ZN(n607) );
  INVD1 U174 ( .I(n28), .ZN(n606) );
  INVD1 U175 ( .I(n28), .ZN(n605) );
  INVD1 U176 ( .I(n29), .ZN(n604) );
  INVD1 U177 ( .I(n29), .ZN(n603) );
  INVD1 U178 ( .I(n29), .ZN(n602) );
  INVD1 U179 ( .I(n30), .ZN(n601) );
  INVD1 U180 ( .I(n30), .ZN(n600) );
  INVD1 U181 ( .I(n30), .ZN(n599) );
  INVD1 U182 ( .I(n31), .ZN(n598) );
  INVD1 U183 ( .I(n31), .ZN(n597) );
  INVD1 U184 ( .I(n31), .ZN(n596) );
  INVD1 U185 ( .I(n32), .ZN(n595) );
  INVD1 U186 ( .I(n32), .ZN(n594) );
  INVD1 U187 ( .I(n32), .ZN(n593) );
  INVD1 U188 ( .I(n33), .ZN(n592) );
  INVD1 U189 ( .I(n33), .ZN(n591) );
  INVD1 U190 ( .I(n33), .ZN(n590) );
  INVD1 U191 ( .I(n34), .ZN(n589) );
  INVD1 U192 ( .I(n34), .ZN(n588) );
  INVD1 U193 ( .I(n34), .ZN(n587) );
  INVD1 U194 ( .I(n35), .ZN(n586) );
  INVD1 U195 ( .I(n35), .ZN(n585) );
  INVD1 U196 ( .I(n35), .ZN(n584) );
  INVD1 U197 ( .I(n666), .ZN(n502) );
  INVD1 U198 ( .I(n666), .ZN(n503) );
  XOR3D1 U199 ( .A1(n673), .A2(n670), .A3(n3), .Z(n2) );
  XNR3D1 U200 ( .A1(n667), .A2(n67), .A3(n68), .ZN(n3) );
  XOR3D1 U201 ( .A1(n73), .A2(n697), .A3(n74), .Z(n72) );
  XOR3D1 U202 ( .A1(n724), .A2(n721), .A3(n75), .Z(n74) );
  XOR3D1 U203 ( .A1(n76), .A2(n718), .A3(n77), .Z(n75) );
  XOR3D1 U204 ( .A1(n682), .A2(n679), .A3(n69), .Z(n68) );
  XOR3D1 U205 ( .A1(n70), .A2(n676), .A3(n71), .Z(n69) );
  XOR3D1 U206 ( .A1(n703), .A2(n700), .A3(n72), .Z(n71) );
  XOR3D1 U207 ( .A1(N59), .A2(N58), .A3(n87), .Z(n86) );
  XOR3D1 U208 ( .A1(n88), .A2(N57), .A3(n89), .Z(n87) );
  XOR3D1 U209 ( .A1(N78), .A2(N73), .A3(n78), .Z(N84) );
  XOR3D1 U210 ( .A1(N72), .A2(n79), .A3(n80), .Z(n78) );
  XOR3D1 U211 ( .A1(N76), .A2(N75), .A3(n81), .Z(n80) );
  XOR3D1 U212 ( .A1(N66), .A2(N65), .A3(n84), .Z(n82) );
  XOR3D1 U213 ( .A1(N64), .A2(n85), .A3(n86), .Z(n84) );
  BUFFD1 U214 ( .I(n663), .Z(n509) );
  BUFFD1 U215 ( .I(N46), .Z(n507) );
  BUFFD1 U216 ( .I(n663), .Z(n510) );
  BUFFD1 U217 ( .I(N44), .Z(n516) );
  OR2D1 U218 ( .A1(n91), .A2(n99), .Z(n4) );
  OR2D1 U219 ( .A1(n91), .A2(n98), .Z(n5) );
  OR2D1 U220 ( .A1(n91), .A2(n97), .Z(n6) );
  OR2D1 U221 ( .A1(n91), .A2(n96), .Z(n7) );
  OR2D1 U222 ( .A1(n91), .A2(n95), .Z(n8) );
  OR2D1 U223 ( .A1(n91), .A2(n94), .Z(n9) );
  OR2D1 U224 ( .A1(n91), .A2(n93), .Z(n10) );
  OR2D1 U225 ( .A1(n91), .A2(n92), .Z(n11) );
  OR2D1 U226 ( .A1(n99), .A2(n105), .Z(n12) );
  OR2D1 U227 ( .A1(n98), .A2(n105), .Z(n13) );
  OR2D1 U228 ( .A1(n97), .A2(n105), .Z(n14) );
  OR2D1 U229 ( .A1(n96), .A2(n105), .Z(n15) );
  OR2D1 U230 ( .A1(n95), .A2(n105), .Z(n16) );
  OR2D1 U231 ( .A1(n94), .A2(n105), .Z(n17) );
  OR2D1 U232 ( .A1(n93), .A2(n105), .Z(n18) );
  OR2D1 U233 ( .A1(n92), .A2(n105), .Z(n19) );
  OR2D1 U234 ( .A1(n99), .A2(n103), .Z(n20) );
  OR2D1 U235 ( .A1(n98), .A2(n103), .Z(n21) );
  OR2D1 U236 ( .A1(n97), .A2(n103), .Z(n22) );
  OR2D1 U237 ( .A1(n96), .A2(n103), .Z(n23) );
  OR2D1 U238 ( .A1(n95), .A2(n103), .Z(n24) );
  OR2D1 U239 ( .A1(n94), .A2(n103), .Z(n25) );
  OR2D1 U240 ( .A1(n93), .A2(n103), .Z(n26) );
  OR2D1 U241 ( .A1(n92), .A2(n103), .Z(n27) );
  OR2D1 U242 ( .A1(n99), .A2(n101), .Z(n28) );
  OR2D1 U243 ( .A1(n98), .A2(n101), .Z(n29) );
  OR2D1 U244 ( .A1(n97), .A2(n101), .Z(n30) );
  OR2D1 U245 ( .A1(n96), .A2(n101), .Z(n31) );
  OR2D1 U246 ( .A1(n95), .A2(n101), .Z(n32) );
  OR2D1 U247 ( .A1(n94), .A2(n101), .Z(n33) );
  OR2D1 U248 ( .A1(n93), .A2(n101), .Z(n34) );
  OR2D1 U249 ( .A1(n92), .A2(n101), .Z(n35) );
  BUFFD1 U250 ( .I(n663), .Z(n508) );
  ND3D1 U251 ( .A1(N44), .A2(N43), .A3(n663), .ZN(n92) );
  INVD1 U252 ( .I(n559), .ZN(n558) );
  INVD1 U253 ( .I(n559), .ZN(n557) );
  CKAN2D0 U254 ( .A1(DreadyReg), .A2(ChipEna), .Z(Dready) );
  INVD1 U255 ( .I(n711), .ZN(n709) );
  INVD1 U256 ( .I(n714), .ZN(n712) );
  INVD1 U257 ( .I(n732), .ZN(n730) );
  INVD1 U258 ( .I(n735), .ZN(n733) );
  INVD1 U259 ( .I(n744), .ZN(n742) );
  INVD1 U260 ( .I(n747), .ZN(n745) );
  INVD1 U261 ( .I(n756), .ZN(n754) );
  INVD1 U262 ( .I(n759), .ZN(n757) );
  INVD1 U263 ( .I(n699), .ZN(n697) );
  INVD1 U264 ( .I(n702), .ZN(n700) );
  INVD1 U265 ( .I(n720), .ZN(n718) );
  INVD1 U266 ( .I(n723), .ZN(n721) );
  INVD1 U267 ( .I(n708), .ZN(n706) );
  INVD1 U268 ( .I(n717), .ZN(n715) );
  INVD1 U269 ( .I(n729), .ZN(n727) );
  INVD1 U270 ( .I(n738), .ZN(n736) );
  INVD1 U271 ( .I(n741), .ZN(n739) );
  INVD1 U272 ( .I(n750), .ZN(n748) );
  INVD1 U273 ( .I(n753), .ZN(n751) );
  INVD1 U274 ( .I(n762), .ZN(n760) );
  INVD1 U275 ( .I(n705), .ZN(n703) );
  INVD1 U276 ( .I(n726), .ZN(n724) );
  INVD1 U277 ( .I(n690), .ZN(n688) );
  INVD1 U278 ( .I(n693), .ZN(n691) );
  INVD1 U279 ( .I(n672), .ZN(n670) );
  INVD1 U280 ( .I(n678), .ZN(n676) );
  INVD1 U281 ( .I(n681), .ZN(n679) );
  INVD1 U282 ( .I(n672), .ZN(n671) );
  INVD1 U283 ( .I(n678), .ZN(n677) );
  INVD1 U284 ( .I(n681), .ZN(n680) );
  INVD1 U285 ( .I(n690), .ZN(n689) );
  INVD1 U286 ( .I(n693), .ZN(n692) );
  INVD1 U287 ( .I(n699), .ZN(n698) );
  INVD1 U288 ( .I(n702), .ZN(n701) );
  INVD1 U289 ( .I(n711), .ZN(n710) );
  INVD1 U290 ( .I(n714), .ZN(n713) );
  INVD1 U291 ( .I(n720), .ZN(n719) );
  INVD1 U292 ( .I(n723), .ZN(n722) );
  INVD1 U293 ( .I(n732), .ZN(n731) );
  INVD1 U294 ( .I(n735), .ZN(n734) );
  INVD1 U295 ( .I(n744), .ZN(n743) );
  INVD1 U296 ( .I(n747), .ZN(n746) );
  INVD1 U297 ( .I(n756), .ZN(n755) );
  INVD1 U298 ( .I(n759), .ZN(n758) );
  INVD1 U299 ( .I(n687), .ZN(n685) );
  INVD1 U300 ( .I(n696), .ZN(n694) );
  INVD1 U301 ( .I(n669), .ZN(n667) );
  INVD1 U302 ( .I(n675), .ZN(n673) );
  INVD1 U303 ( .I(n684), .ZN(n682) );
  INVD1 U304 ( .I(n669), .ZN(n668) );
  INVD1 U305 ( .I(n675), .ZN(n674) );
  INVD1 U306 ( .I(n684), .ZN(n683) );
  INVD1 U307 ( .I(n687), .ZN(n686) );
  INVD1 U308 ( .I(n696), .ZN(n695) );
  INVD1 U309 ( .I(n705), .ZN(n704) );
  INVD1 U310 ( .I(n708), .ZN(n707) );
  INVD1 U311 ( .I(n717), .ZN(n716) );
  INVD1 U312 ( .I(n726), .ZN(n725) );
  INVD1 U313 ( .I(n729), .ZN(n728) );
  INVD1 U314 ( .I(n738), .ZN(n737) );
  INVD1 U315 ( .I(n741), .ZN(n740) );
  INVD1 U316 ( .I(n750), .ZN(n749) );
  INVD1 U317 ( .I(n753), .ZN(n752) );
  INVD1 U318 ( .I(n762), .ZN(n761) );
  INVD1 U319 ( .I(n664), .ZN(n663) );
  ND3D1 U320 ( .A1(n100), .A2(n666), .A3(N46), .ZN(n103) );
  ND3D1 U321 ( .A1(n665), .A2(n666), .A3(n100), .ZN(n105) );
  ND3D1 U322 ( .A1(n100), .A2(n665), .A3(N47), .ZN(n101) );
  ND3D1 U323 ( .A1(N46), .A2(n100), .A3(N47), .ZN(n91) );
  ND3D1 U324 ( .A1(n662), .A2(n664), .A3(N43), .ZN(n98) );
  ND3D1 U325 ( .A1(n661), .A2(n664), .A3(N44), .ZN(n97) );
  ND3D1 U326 ( .A1(N43), .A2(n664), .A3(N44), .ZN(n96) );
  ND3D1 U327 ( .A1(n661), .A2(n662), .A3(n663), .ZN(n95) );
  ND3D1 U328 ( .A1(N43), .A2(n662), .A3(n663), .ZN(n94) );
  ND3D1 U329 ( .A1(N44), .A2(n661), .A3(n663), .ZN(n93) );
  ND3D1 U330 ( .A1(n662), .A2(n664), .A3(n661), .ZN(n99) );
  INR2D1 U331 ( .A1(ChipEna), .B1(n90), .ZN(N2262) );
  MUX4ND0 U332 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n536), .S1(n518), .ZN(
        n492) );
  MUX4ND0 U333 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n550), .S1(n522), .ZN(
        n310) );
  MUX4ND0 U334 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n537), .S1(n517), .ZN(
        n323) );
  MUX4ND0 U335 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n537), .S1(n524), .ZN(
        n336) );
  MUX4ND0 U336 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n539), .S1(n518), .ZN(
        n349) );
  MUX4ND0 U337 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n535), .S1(n521), .ZN(
        n388) );
  MUX4ND0 U338 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n535), .S1(n521), .ZN(
        n401) );
  MUX4ND0 U339 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n537), .S1(n521), .ZN(
        n414) );
  MUX4ND0 U340 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n538), .S1(n518), .ZN(
        n427) );
  MUX4ND0 U341 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n540), .S1(n517), .ZN(
        n440) );
  MUX4ND0 U342 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n539), .S1(n517), .ZN(
        n453) );
  MUX4ND0 U343 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n535), .S1(n518), .ZN(
        n466) );
  MUX4ND0 U344 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n537), .S1(n517), .ZN(
        n479) );
  MUX4D0 U345 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n535), .S1(n528), .Z(
        n493) );
  MUX4D0 U346 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n537), .S1(n525), .Z(
        n389) );
  MUX4D0 U347 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n542), .S1(n525), .Z(
        n402) );
  MUX4D0 U348 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n536), .S1(n526), .Z(
        n415) );
  MUX4D0 U349 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n542), .S1(n526), .Z(
        n428) );
  MUX4D0 U350 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n539), .S1(n527), .Z(
        n441) );
  MUX4D0 U351 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n539), .S1(n527), .Z(
        n454) );
  MUX4D0 U352 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n542), .S1(n527), .Z(
        n467) );
  MUX4D0 U353 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(N43), .S1(n528), .Z(
        n480) );
  MUX4D0 U354 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n535), .S1(n529), .Z(
        n497) );
  MUX4D0 U355 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n536), .S1(n529), .Z(
        n495) );
  MUX4D0 U356 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n539), .S1(n525), .Z(
        n393) );
  MUX4D0 U357 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n540), .S1(n525), .Z(
        n391) );
  MUX4D0 U358 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n538), .S1(n525), .Z(
        n406) );
  MUX4D0 U359 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(N43), .S1(n525), .Z(
        n404) );
  MUX4D0 U360 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n536), .S1(n526), .Z(
        n419) );
  MUX4D0 U361 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n536), .S1(n526), .Z(
        n417) );
  MUX4D0 U362 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n539), .S1(n526), .Z(
        n432) );
  MUX4D0 U363 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n542), .S1(n526), .Z(
        n430) );
  MUX4D0 U364 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n536), .S1(n527), .Z(
        n445) );
  MUX4D0 U365 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n539), .S1(n527), .Z(
        n443) );
  MUX4D0 U366 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n542), .S1(n527), .Z(
        n458) );
  MUX4D0 U367 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n542), .S1(n527), .Z(
        n456) );
  MUX4D0 U368 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n540), .S1(n528), .Z(
        n471) );
  MUX4D0 U369 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n538), .S1(n528), .Z(
        n469) );
  MUX4D0 U370 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n542), .S1(n528), .Z(
        n484) );
  MUX4D0 U371 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n537), .S1(n528), .Z(
        n482) );
  MUX4D0 U372 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(N43), .S1(n528), .Z(
        n494) );
  MUX4D0 U373 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n541), .S1(n525), .Z(
        n390) );
  MUX4D0 U374 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n542), .S1(n525), .Z(
        n403) );
  MUX4D0 U375 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n540), .S1(n526), .Z(
        n416) );
  MUX4D0 U376 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n540), .S1(n526), .Z(
        n429) );
  MUX4D0 U377 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(N43), .S1(n527), .Z(
        n442) );
  MUX4D0 U378 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n539), .S1(n527), .Z(
        n455) );
  MUX4D0 U379 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n536), .S1(n528), .Z(
        n468) );
  MUX4D0 U380 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n540), .S1(n528), .Z(
        n481) );
  MUX4D0 U381 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n536), .S1(n529), .Z(
        n498) );
  MUX4D0 U382 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n535), .S1(n529), .Z(
        n496) );
  MUX4D0 U383 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n537), .S1(n522), .Z(
        n316) );
  MUX4D0 U384 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n539), .S1(n523), .Z(
        n342) );
  MUX4D0 U385 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n556), .S1(n524), .Z(
        n355) );
  MUX4D0 U386 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n537), .S1(n525), .Z(
        n394) );
  MUX4D0 U387 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n540), .S1(n525), .Z(
        n392) );
  MUX4D0 U388 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n541), .S1(n526), .Z(
        n407) );
  MUX4D0 U389 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n539), .S1(n525), .Z(
        n405) );
  MUX4D0 U390 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n538), .S1(n526), .Z(
        n420) );
  MUX4D0 U391 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n535), .S1(n526), .Z(
        n418) );
  MUX4D0 U392 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n536), .S1(n526), .Z(
        n433) );
  MUX4D0 U393 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(N43), .S1(n526), .Z(
        n431) );
  MUX4D0 U394 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n539), .S1(n527), .Z(
        n446) );
  MUX4D0 U395 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(N43), .S1(n527), .Z(
        n444) );
  MUX4D0 U396 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n542), .S1(n527), .Z(
        n459) );
  MUX4D0 U397 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n538), .S1(n527), .Z(
        n457) );
  MUX4D0 U398 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n538), .S1(n528), .Z(
        n472) );
  MUX4D0 U399 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n538), .S1(n528), .Z(
        n470) );
  MUX4D0 U400 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n540), .S1(n528), .Z(
        n485) );
  MUX4D0 U401 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n539), .S1(n528), .Z(
        n483) );
  INVD1 U402 ( .I(N43), .ZN(n661) );
  INVD1 U403 ( .I(N45), .ZN(n664) );
  INVD1 U404 ( .I(N44), .ZN(n662) );
  INVD1 U405 ( .I(N46), .ZN(n665) );
  MUX4ND0 U406 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n547), .S1(n517), .ZN(
        n193) );
  MUX4ND0 U407 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n548), .S1(n522), .ZN(
        n39) );
  MUX4ND0 U408 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n547), .S1(n522), .ZN(
        n52) );
  MUX4ND0 U409 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n547), .S1(n522), .ZN(
        n65) );
  MUX4ND0 U410 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n547), .S1(n517), .ZN(
        n115) );
  MUX4ND0 U411 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n547), .S1(n534), .ZN(
        n128) );
  MUX4ND0 U412 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n547), .S1(n516), .ZN(
        n141) );
  MUX4ND0 U413 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n547), .S1(n518), .ZN(
        n154) );
  MUX4ND0 U414 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n547), .S1(n531), .ZN(
        n167) );
  MUX4ND0 U415 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n547), .S1(n518), .ZN(
        n180) );
  MUX4ND0 U416 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n547), .S1(n532), .ZN(
        n206) );
  MUX4ND0 U417 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n547), .S1(n530), .ZN(
        n219) );
  MUX4ND0 U418 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n547), .S1(n531), .ZN(
        n232) );
  MUX4ND0 U419 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n554), .S1(n534), .ZN(
        n245) );
  MUX4ND0 U420 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n555), .S1(n532), .ZN(
        n258) );
  MUX4ND0 U421 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n549), .S1(n530), .ZN(
        n271) );
  MUX4ND0 U422 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n548), .S1(n533), .ZN(
        n284) );
  MUX4ND0 U423 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n550), .S1(n518), .ZN(
        n297) );
  MUX4ND0 U424 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n555), .S1(n533), .ZN(
        n362) );
  MUX4ND0 U425 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n554), .S1(n519), .ZN(
        n375) );
  MUX4D0 U426 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n552), .S1(n533), .Z(
        n194) );
  MUX4D0 U427 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n553), .S1(n521), .Z(n40) );
  MUX4D0 U428 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n548), .S1(n529), .Z(n53) );
  MUX4D0 U429 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n548), .S1(n530), .Z(n66) );
  MUX4D0 U430 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n549), .S1(n530), .Z(
        n116) );
  MUX4D0 U431 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n549), .S1(n531), .Z(
        n129) );
  MUX4D0 U432 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n550), .S1(n531), .Z(
        n142) );
  MUX4D0 U433 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n550), .S1(n532), .Z(
        n155) );
  MUX4D0 U434 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n551), .S1(n532), .Z(
        n168) );
  MUX4D0 U435 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n551), .S1(n532), .Z(
        n181) );
  MUX4D0 U436 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n552), .S1(n533), .Z(
        n207) );
  MUX4D0 U437 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n553), .S1(n516), .Z(
        n220) );
  MUX4D0 U438 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n553), .S1(n534), .Z(
        n233) );
  MUX4D0 U439 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n554), .S1(n534), .Z(
        n246) );
  MUX4D0 U440 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n554), .S1(n534), .Z(
        n259) );
  MUX4D0 U441 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n555), .S1(n516), .Z(
        n272) );
  MUX4D0 U442 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n555), .S1(N44), .Z(
        n285) );
  MUX4D0 U443 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n556), .S1(n517), .Z(
        n298) );
  MUX4D0 U444 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n556), .S1(n522), .Z(
        n311) );
  MUX4D0 U445 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n538), .S1(n522), .Z(
        n324) );
  MUX4D0 U446 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n535), .S1(n523), .Z(
        n337) );
  MUX4D0 U447 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n554), .S1(n523), .Z(
        n350) );
  MUX4D0 U448 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n541), .S1(n524), .Z(
        n363) );
  MUX4D0 U449 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n553), .S1(n524), .Z(
        n376) );
  MUX4D0 U450 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n552), .S1(n533), .Z(n198)
         );
  MUX4D0 U451 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n552), .S1(n525), .Z(
        n196) );
  MUX4D0 U452 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n548), .S1(n529), .Z(n44)
         );
  MUX4D0 U453 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n549), .S1(n529), .Z(n42) );
  MUX4D0 U454 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n548), .S1(n530), .Z(n57)
         );
  MUX4D0 U455 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n548), .S1(n529), .Z(n55) );
  MUX4D0 U456 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n548), .S1(n530), .Z(n107)
         );
  MUX4D0 U457 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n548), .S1(n530), .Z(
        n104) );
  MUX4D0 U458 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n549), .S1(n530), .Z(n120)
         );
  MUX4D0 U459 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n549), .S1(n530), .Z(
        n118) );
  MUX4D0 U460 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n549), .S1(n531), .Z(n133)
         );
  MUX4D0 U461 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n549), .S1(n531), .Z(
        n131) );
  MUX4D0 U462 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n550), .S1(n531), .Z(n146)
         );
  MUX4D0 U463 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n550), .S1(n531), .Z(
        n144) );
  MUX4D0 U464 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n550), .S1(n532), .Z(n159)
         );
  MUX4D0 U465 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n550), .S1(n532), .Z(
        n157) );
  MUX4D0 U466 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n551), .S1(n532), .Z(n172)
         );
  MUX4D0 U467 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n551), .S1(n532), .Z(
        n170) );
  MUX4D0 U468 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n551), .S1(n533), .Z(n185)
         );
  MUX4D0 U469 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n551), .S1(n533), .Z(
        n183) );
  MUX4D0 U470 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n552), .S1(n520), .Z(
        n211) );
  MUX4D0 U471 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n552), .S1(n520), .Z(
        n209) );
  MUX4D0 U472 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n553), .S1(n517), .Z(
        n224) );
  MUX4D0 U473 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n553), .S1(n516), .Z(
        n222) );
  MUX4D0 U474 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n553), .S1(n534), .Z(
        n237) );
  MUX4D0 U475 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n553), .S1(n534), .Z(
        n235) );
  MUX4D0 U476 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n554), .S1(n526), .Z(
        n250) );
  MUX4D0 U477 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n554), .S1(n534), .Z(
        n248) );
  MUX4D0 U478 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n554), .S1(n534), .Z(
        n263) );
  MUX4D0 U479 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n554), .S1(n534), .Z(
        n261) );
  MUX4D0 U480 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n555), .S1(n516), .Z(
        n276) );
  MUX4D0 U481 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n555), .S1(N44), .Z(
        n274) );
  MUX4D0 U482 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n555), .S1(n521), .Z(
        n289) );
  MUX4D0 U483 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n555), .S1(n517), .Z(
        n287) );
  MUX4D0 U484 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n556), .S1(n533), .Z(
        n302) );
  MUX4D0 U485 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n556), .S1(n517), .Z(
        n300) );
  MUX4D0 U486 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n556), .S1(n522), .Z(
        n315) );
  MUX4D0 U487 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n556), .S1(n522), .Z(
        n313) );
  MUX4D0 U488 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n537), .S1(n523), .Z(
        n328) );
  MUX4D0 U489 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n541), .S1(n522), .Z(
        n326) );
  MUX4D0 U490 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n537), .S1(n523), .Z(
        n341) );
  MUX4D0 U491 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n540), .S1(n523), .Z(
        n339) );
  MUX4D0 U492 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n537), .S1(n524), .Z(
        n354) );
  MUX4D0 U493 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n537), .S1(n523), .Z(
        n352) );
  MUX4D0 U494 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n551), .S1(n524), .Z(
        n367) );
  MUX4D0 U495 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n552), .S1(n524), .Z(
        n365) );
  MUX4D0 U496 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n540), .S1(n524), .Z(
        n380) );
  MUX4D0 U497 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n535), .S1(n524), .Z(
        n378) );
  MUX4D0 U498 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n552), .S1(n533), .Z(
        n195) );
  MUX4D0 U499 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n552), .S1(n529), .Z(n41) );
  MUX4D0 U500 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n548), .S1(n529), .Z(n54) );
  MUX4D0 U501 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n548), .S1(n530), .Z(
        n102) );
  MUX4D0 U502 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n549), .S1(n530), .Z(
        n117) );
  MUX4D0 U503 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n549), .S1(n531), .Z(
        n130) );
  MUX4D0 U504 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n550), .S1(n531), .Z(
        n143) );
  MUX4D0 U505 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n550), .S1(n532), .Z(
        n156) );
  MUX4D0 U506 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n551), .S1(n532), .Z(
        n169) );
  MUX4D0 U507 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n551), .S1(n533), .Z(
        n182) );
  MUX4D0 U508 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n552), .S1(n533), .Z(
        n208) );
  MUX4D0 U509 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n553), .S1(n516), .Z(
        n221) );
  MUX4D0 U510 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n553), .S1(n516), .Z(
        n234) );
  MUX4D0 U511 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n554), .S1(n534), .Z(
        n247) );
  MUX4D0 U512 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n554), .S1(n520), .Z(
        n260) );
  MUX4D0 U513 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n555), .S1(n534), .Z(
        n273) );
  MUX4D0 U514 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n555), .S1(n518), .Z(
        n286) );
  MUX4D0 U515 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n556), .S1(n519), .Z(
        n299) );
  MUX4D0 U516 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n556), .S1(n522), .Z(
        n312) );
  MUX4D0 U517 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n540), .S1(n522), .Z(
        n325) );
  MUX4D0 U518 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n541), .S1(n523), .Z(
        n338) );
  MUX4D0 U519 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n540), .S1(n523), .Z(
        n351) );
  MUX4D0 U520 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n551), .S1(n524), .Z(
        n364) );
  MUX4D0 U521 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n538), .S1(n524), .Z(
        n377) );
  MUX4D0 U522 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n552), .S1(n533), .Z(n199)
         );
  MUX4D0 U523 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n552), .S1(n533), .Z(
        n197) );
  MUX4D0 U524 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n550), .S1(n529), .Z(n45)
         );
  MUX4D0 U525 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n549), .S1(n529), .Z(n43) );
  MUX4D0 U526 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n548), .S1(n530), .Z(n58)
         );
  MUX4D0 U527 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n548), .S1(n529), .Z(n56) );
  MUX4D0 U528 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n548), .S1(n530), .Z(n108)
         );
  MUX4D0 U529 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n548), .S1(n530), .Z(
        n106) );
  MUX4D0 U530 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n549), .S1(n531), .Z(n121)
         );
  MUX4D0 U531 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n549), .S1(n530), .Z(
        n119) );
  MUX4D0 U532 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n549), .S1(n531), .Z(n134)
         );
  MUX4D0 U533 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n549), .S1(n531), .Z(
        n132) );
  MUX4D0 U534 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n550), .S1(n531), .Z(n147)
         );
  MUX4D0 U535 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n550), .S1(n531), .Z(
        n145) );
  MUX4D0 U536 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n550), .S1(n532), .Z(n160)
         );
  MUX4D0 U537 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n550), .S1(n532), .Z(
        n158) );
  MUX4D0 U538 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n551), .S1(n532), .Z(n173)
         );
  MUX4D0 U539 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n551), .S1(n532), .Z(
        n171) );
  MUX4D0 U540 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n551), .S1(n533), .Z(n186)
         );
  MUX4D0 U541 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n551), .S1(n533), .Z(
        n184) );
  MUX4D0 U542 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n552), .S1(n519), .Z(
        n212) );
  MUX4D0 U543 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n552), .S1(n519), .Z(
        n210) );
  MUX4D0 U544 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n553), .S1(n526), .Z(
        n225) );
  MUX4D0 U545 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n553), .S1(n516), .Z(
        n223) );
  MUX4D0 U546 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n554), .S1(n534), .Z(
        n238) );
  MUX4D0 U547 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n553), .S1(n534), .Z(
        n236) );
  MUX4D0 U548 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n554), .S1(n534), .Z(
        n251) );
  MUX4D0 U549 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n554), .S1(n517), .Z(
        n249) );
  MUX4D0 U550 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n555), .S1(n528), .Z(
        n264) );
  MUX4D0 U551 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n554), .S1(n527), .Z(
        n262) );
  MUX4D0 U552 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n555), .S1(n520), .Z(
        n277) );
  MUX4D0 U553 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n555), .S1(N44), .Z(
        n275) );
  MUX4D0 U554 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n556), .S1(n522), .Z(
        n290) );
  MUX4D0 U555 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n555), .S1(n516), .Z(
        n288) );
  MUX4D0 U556 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n556), .S1(n522), .Z(
        n303) );
  MUX4D0 U557 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n556), .S1(n525), .Z(
        n301) );
  MUX4D0 U558 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n556), .S1(n522), .Z(
        n314) );
  MUX4D0 U559 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n537), .S1(n523), .Z(
        n329) );
  MUX4D0 U560 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n538), .S1(n523), .Z(
        n327) );
  MUX4D0 U561 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n556), .S1(n523), .Z(
        n340) );
  MUX4D0 U562 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n538), .S1(n523), .Z(
        n353) );
  MUX4D0 U563 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n555), .S1(n524), .Z(
        n368) );
  MUX4D0 U564 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n553), .S1(n524), .Z(
        n366) );
  MUX4D0 U565 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n537), .S1(n525), .Z(
        n381) );
  MUX4D0 U566 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n541), .S1(n524), .Z(
        n379) );
  INVD1 U567 ( .I(N47), .ZN(n666) );
  AN3D1 U568 ( .A1(n90), .A2(n659), .A3(Write), .Z(n100) );
  MUX3ND0 U569 ( .I0(n37), .I1(n38), .I2(n39), .S0(n517), .S1(n512), .ZN(n36)
         );
  MUX3ND0 U570 ( .I0(n46), .I1(n47), .I2(n48), .S0(n506), .S1(N47), .ZN(N81)
         );
  MUX3ND0 U571 ( .I0(n50), .I1(n51), .I2(n52), .S0(n519), .S1(n508), .ZN(n49)
         );
  MUX3ND0 U572 ( .I0(n59), .I1(n60), .I2(n61), .S0(N46), .S1(n502), .ZN(N80)
         );
  MUX3ND0 U573 ( .I0(n63), .I1(n64), .I2(n65), .S0(N44), .S1(n508), .ZN(n62)
         );
  MUX3ND0 U574 ( .I0(n109), .I1(n110), .I2(n111), .S0(N46), .S1(n502), .ZN(N79) );
  MUX3ND0 U575 ( .I0(n113), .I1(n114), .I2(n115), .S0(N44), .S1(n510), .ZN(
        n112) );
  MUX3ND0 U576 ( .I0(n122), .I1(n123), .I2(n124), .S0(n507), .S1(N47), .ZN(N78) );
  MUX3ND0 U577 ( .I0(n126), .I1(n127), .I2(n128), .S0(n516), .S1(n508), .ZN(
        n125) );
  MUX3ND0 U578 ( .I0(n135), .I1(n136), .I2(n137), .S0(n507), .S1(N47), .ZN(N77) );
  MUX3ND0 U579 ( .I0(n139), .I1(n140), .I2(n141), .S0(n521), .S1(n508), .ZN(
        n138) );
  MUX3ND0 U580 ( .I0(n148), .I1(n149), .I2(n150), .S0(n506), .S1(N47), .ZN(N76) );
  MUX3ND0 U581 ( .I0(n152), .I1(n153), .I2(n154), .S0(n519), .S1(n508), .ZN(
        n151) );
  MUX3ND0 U582 ( .I0(n161), .I1(n162), .I2(n163), .S0(n507), .S1(N47), .ZN(N75) );
  MUX3ND0 U583 ( .I0(n165), .I1(n166), .I2(n167), .S0(n521), .S1(N45), .ZN(
        n164) );
  MUX3ND0 U584 ( .I0(n174), .I1(n175), .I2(n176), .S0(n507), .S1(n502), .ZN(
        N74) );
  MUX3ND0 U585 ( .I0(n178), .I1(n179), .I2(n180), .S0(n521), .S1(n508), .ZN(
        n177) );
  MUX3ND0 U586 ( .I0(n187), .I1(n188), .I2(n189), .S0(n506), .S1(n502), .ZN(
        N73) );
  MUX3ND0 U587 ( .I0(n191), .I1(n192), .I2(n193), .S0(n518), .S1(n514), .ZN(
        n190) );
  MUX3ND0 U588 ( .I0(n200), .I1(n201), .I2(n202), .S0(n507), .S1(n502), .ZN(
        N72) );
  MUX3ND0 U589 ( .I0(n204), .I1(n205), .I2(n206), .S0(N44), .S1(n508), .ZN(
        n203) );
  MUX3ND0 U590 ( .I0(n213), .I1(n214), .I2(n215), .S0(n506), .S1(n502), .ZN(
        N71) );
  MUX3ND0 U591 ( .I0(n217), .I1(n218), .I2(n219), .S0(n524), .S1(N45), .ZN(
        n216) );
  MUX3ND0 U592 ( .I0(n226), .I1(n227), .I2(n228), .S0(n506), .S1(n502), .ZN(
        N70) );
  MUX3ND0 U593 ( .I0(n230), .I1(n231), .I2(n232), .S0(n529), .S1(n513), .ZN(
        n229) );
  MUX3ND0 U594 ( .I0(n239), .I1(n240), .I2(n241), .S0(n507), .S1(n502), .ZN(
        N69) );
  MUX3ND0 U595 ( .I0(n243), .I1(n244), .I2(n245), .S0(n521), .S1(n512), .ZN(
        n242) );
  MUX3ND0 U596 ( .I0(n252), .I1(n253), .I2(n254), .S0(N46), .S1(n502), .ZN(N68) );
  MUX3ND0 U597 ( .I0(n256), .I1(n257), .I2(n258), .S0(N44), .S1(n513), .ZN(
        n255) );
  MUX3ND0 U598 ( .I0(n265), .I1(n266), .I2(n267), .S0(N46), .S1(n502), .ZN(N67) );
  MUX3ND0 U599 ( .I0(n269), .I1(n270), .I2(n271), .S0(n523), .S1(n510), .ZN(
        n268) );
  MUX3ND0 U600 ( .I0(n278), .I1(n279), .I2(n280), .S0(N46), .S1(n502), .ZN(N66) );
  MUX3ND0 U601 ( .I0(n282), .I1(n283), .I2(n284), .S0(n525), .S1(n510), .ZN(
        n281) );
  MUX3ND0 U602 ( .I0(n291), .I1(n292), .I2(n293), .S0(N46), .S1(n502), .ZN(N65) );
  MUX3ND0 U603 ( .I0(n295), .I1(n296), .I2(n297), .S0(n527), .S1(n510), .ZN(
        n294) );
  MUX3ND0 U604 ( .I0(n304), .I1(n305), .I2(n306), .S0(N46), .S1(n502), .ZN(N64) );
  MUX3ND0 U605 ( .I0(n308), .I1(n309), .I2(n310), .S0(n516), .S1(n510), .ZN(
        n307) );
  MUX3ND0 U606 ( .I0(n317), .I1(n318), .I2(n319), .S0(n506), .S1(n502), .ZN(
        N63) );
  MUX3ND0 U607 ( .I0(n321), .I1(n322), .I2(n323), .S0(n521), .S1(n510), .ZN(
        n320) );
  MUX3ND0 U608 ( .I0(n330), .I1(n331), .I2(n332), .S0(n507), .S1(n502), .ZN(
        N62) );
  MUX3ND0 U609 ( .I0(n334), .I1(n335), .I2(n336), .S0(n518), .S1(n510), .ZN(
        n333) );
  MUX3ND0 U610 ( .I0(n343), .I1(n344), .I2(n345), .S0(n506), .S1(n503), .ZN(
        N61) );
  MUX3ND0 U611 ( .I0(n347), .I1(n348), .I2(n349), .S0(n519), .S1(n510), .ZN(
        n346) );
  MUX3ND0 U612 ( .I0(n356), .I1(n357), .I2(n358), .S0(n507), .S1(n503), .ZN(
        N60) );
  MUX3ND0 U613 ( .I0(n360), .I1(n361), .I2(n362), .S0(N44), .S1(n510), .ZN(
        n359) );
  MUX3ND0 U614 ( .I0(n369), .I1(n370), .I2(n371), .S0(N46), .S1(n503), .ZN(N59) );
  MUX3ND0 U615 ( .I0(n373), .I1(n374), .I2(n375), .S0(n517), .S1(n510), .ZN(
        n372) );
  MUX3ND0 U616 ( .I0(n382), .I1(n383), .I2(n384), .S0(N46), .S1(n503), .ZN(N58) );
  MUX3ND0 U617 ( .I0(n386), .I1(n387), .I2(n388), .S0(n523), .S1(n510), .ZN(
        n385) );
  MUX3ND0 U618 ( .I0(n395), .I1(n396), .I2(n397), .S0(n505), .S1(n503), .ZN(
        N57) );
  MUX3ND0 U619 ( .I0(n399), .I1(n400), .I2(n401), .S0(n519), .S1(n510), .ZN(
        n398) );
  MUX3ND0 U620 ( .I0(n408), .I1(n409), .I2(n410), .S0(n507), .S1(n503), .ZN(
        N56) );
  MUX3ND0 U621 ( .I0(n412), .I1(n413), .I2(n414), .S0(n521), .S1(n510), .ZN(
        n411) );
  MUX3ND0 U622 ( .I0(n421), .I1(n422), .I2(n423), .S0(n507), .S1(n503), .ZN(
        N55) );
  MUX3ND0 U623 ( .I0(n425), .I1(n426), .I2(n427), .S0(n517), .S1(n510), .ZN(
        n424) );
  MUX3ND0 U624 ( .I0(n434), .I1(n435), .I2(n436), .S0(n507), .S1(n503), .ZN(
        N54) );
  MUX3ND0 U625 ( .I0(n438), .I1(n439), .I2(n440), .S0(n518), .S1(n508), .ZN(
        n437) );
  MUX3ND0 U626 ( .I0(n447), .I1(n448), .I2(n449), .S0(n507), .S1(n503), .ZN(
        N53) );
  MUX3ND0 U627 ( .I0(n451), .I1(n452), .I2(n453), .S0(n518), .S1(n663), .ZN(
        n450) );
  MUX3ND0 U628 ( .I0(n460), .I1(n461), .I2(n462), .S0(n506), .S1(n503), .ZN(
        N52) );
  MUX3ND0 U629 ( .I0(n464), .I1(n465), .I2(n466), .S0(n521), .S1(n508), .ZN(
        n463) );
  MUX3ND0 U630 ( .I0(n473), .I1(n474), .I2(n475), .S0(n507), .S1(n503), .ZN(
        N51) );
  MUX3ND0 U631 ( .I0(n477), .I1(n478), .I2(n479), .S0(n529), .S1(n663), .ZN(
        n476) );
  MUX3ND0 U632 ( .I0(n486), .I1(n487), .I2(n488), .S0(n504), .S1(n503), .ZN(
        N50) );
  MUX3ND0 U633 ( .I0(n490), .I1(n491), .I2(n492), .S0(n519), .S1(N45), .ZN(
        n489) );
  MUX3ND0 U634 ( .I0(n499), .I1(n500), .I2(n501), .S0(n506), .S1(n503), .ZN(
        N49) );
  MUX2ND0 U635 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n542), .ZN(
        n38) );
  MUX2ND0 U636 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n542), .ZN(
        n37) );
  MUX3ND0 U637 ( .I0(n41), .I1(n40), .I2(n36), .S0(n515), .S1(n504), .ZN(n48)
         );
  MUX2ND0 U638 ( .I0(n43), .I1(n42), .S(n513), .ZN(n47) );
  MUX2ND0 U639 ( .I0(n45), .I1(n44), .S(n512), .ZN(n46) );
  MUX2ND0 U640 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n543), .ZN(
        n51) );
  MUX2ND0 U641 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n543), .ZN(
        n50) );
  MUX3ND0 U642 ( .I0(n54), .I1(n53), .I2(n49), .S0(n515), .S1(n506), .ZN(n61)
         );
  MUX2ND0 U643 ( .I0(n56), .I1(n55), .S(n511), .ZN(n60) );
  MUX2ND0 U644 ( .I0(n58), .I1(n57), .S(n513), .ZN(n59) );
  MUX2ND0 U645 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n543), .ZN(
        n64) );
  MUX2ND0 U646 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n543), .ZN(
        n63) );
  MUX3ND0 U647 ( .I0(n102), .I1(n66), .I2(n62), .S0(n515), .S1(n506), .ZN(n111) );
  MUX2ND0 U648 ( .I0(n106), .I1(n104), .S(n513), .ZN(n110) );
  MUX2ND0 U649 ( .I0(n108), .I1(n107), .S(n512), .ZN(n109) );
  MUX2ND0 U650 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n544), .ZN(
        n114) );
  MUX2ND0 U651 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n544), .ZN(
        n113) );
  MUX3ND0 U652 ( .I0(n117), .I1(n116), .I2(n112), .S0(n515), .S1(n507), .ZN(
        n124) );
  MUX2ND0 U653 ( .I0(n119), .I1(n118), .S(n513), .ZN(n123) );
  MUX2ND0 U654 ( .I0(n121), .I1(n120), .S(n512), .ZN(n122) );
  MUX2ND0 U655 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n545), .ZN(
        n127) );
  MUX2ND0 U656 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n544), .ZN(
        n126) );
  MUX3ND0 U657 ( .I0(n130), .I1(n129), .I2(n125), .S0(n515), .S1(n506), .ZN(
        n137) );
  MUX2ND0 U658 ( .I0(n132), .I1(n131), .S(n513), .ZN(n136) );
  MUX2ND0 U659 ( .I0(n134), .I1(n133), .S(n513), .ZN(n135) );
  MUX2ND0 U660 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n545), .ZN(
        n140) );
  MUX2ND0 U661 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n545), .ZN(
        n139) );
  MUX3ND0 U662 ( .I0(n143), .I1(n142), .I2(n138), .S0(n514), .S1(n507), .ZN(
        n150) );
  MUX2ND0 U663 ( .I0(n145), .I1(n144), .S(n512), .ZN(n149) );
  MUX2ND0 U664 ( .I0(n147), .I1(n146), .S(n512), .ZN(n148) );
  MUX2ND0 U665 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n546), .ZN(
        n153) );
  MUX2ND0 U666 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n545), .ZN(
        n152) );
  MUX3ND0 U667 ( .I0(n156), .I1(n155), .I2(n151), .S0(n514), .S1(n505), .ZN(
        n163) );
  MUX2ND0 U668 ( .I0(n158), .I1(n157), .S(n512), .ZN(n162) );
  MUX2ND0 U669 ( .I0(n160), .I1(n159), .S(n512), .ZN(n161) );
  MUX2ND0 U670 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n546), .ZN(
        n166) );
  MUX2ND0 U671 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n546), .ZN(
        n165) );
  MUX3ND0 U672 ( .I0(n169), .I1(n168), .I2(n164), .S0(n513), .S1(n505), .ZN(
        n176) );
  MUX2ND0 U673 ( .I0(n171), .I1(n170), .S(n512), .ZN(n175) );
  MUX2ND0 U674 ( .I0(n173), .I1(n172), .S(n512), .ZN(n174) );
  MUX2ND0 U675 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n547), .ZN(
        n179) );
  MUX2ND0 U676 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n546), .ZN(
        n178) );
  MUX3ND0 U677 ( .I0(n182), .I1(n181), .I2(n177), .S0(n515), .S1(n505), .ZN(
        n189) );
  MUX2ND0 U678 ( .I0(n184), .I1(n183), .S(n512), .ZN(n188) );
  MUX2ND0 U679 ( .I0(n186), .I1(n185), .S(n512), .ZN(n187) );
  MUX2ND0 U680 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n546), .ZN(
        n192) );
  MUX2ND0 U681 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n547), .ZN(
        n191) );
  MUX3ND0 U682 ( .I0(n195), .I1(n194), .I2(n190), .S0(n514), .S1(n505), .ZN(
        n202) );
  MUX2ND0 U683 ( .I0(n197), .I1(n196), .S(n512), .ZN(n201) );
  MUX2ND0 U684 ( .I0(n199), .I1(n198), .S(n511), .ZN(n200) );
  MUX2ND0 U685 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n547), 
        .ZN(n205) );
  MUX2ND0 U686 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n546), 
        .ZN(n204) );
  MUX3ND0 U687 ( .I0(n208), .I1(n207), .I2(n203), .S0(n513), .S1(n505), .ZN(
        n215) );
  MUX2ND0 U688 ( .I0(n210), .I1(n209), .S(n511), .ZN(n214) );
  MUX2ND0 U689 ( .I0(n212), .I1(n211), .S(n511), .ZN(n213) );
  MUX2ND0 U690 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n546), 
        .ZN(n218) );
  MUX2ND0 U691 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n546), 
        .ZN(n217) );
  MUX3ND0 U692 ( .I0(n221), .I1(n220), .I2(n216), .S0(n513), .S1(n505), .ZN(
        n228) );
  MUX2ND0 U693 ( .I0(n223), .I1(n222), .S(n512), .ZN(n227) );
  MUX2ND0 U694 ( .I0(n225), .I1(n224), .S(n511), .ZN(n226) );
  MUX2ND0 U695 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n546), 
        .ZN(n231) );
  MUX2ND0 U696 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n546), 
        .ZN(n230) );
  MUX3ND0 U697 ( .I0(n234), .I1(n233), .I2(n229), .S0(n514), .S1(n505), .ZN(
        n241) );
  MUX2ND0 U698 ( .I0(n236), .I1(n235), .S(n511), .ZN(n240) );
  MUX2ND0 U699 ( .I0(n238), .I1(n237), .S(n511), .ZN(n239) );
  MUX2ND0 U700 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n546), 
        .ZN(n244) );
  MUX2ND0 U701 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n546), 
        .ZN(n243) );
  MUX3ND0 U702 ( .I0(n247), .I1(n246), .I2(n242), .S0(n514), .S1(n505), .ZN(
        n254) );
  MUX2ND0 U703 ( .I0(n249), .I1(n248), .S(n511), .ZN(n253) );
  MUX2ND0 U704 ( .I0(n251), .I1(n250), .S(n511), .ZN(n252) );
  MUX2ND0 U705 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n546), 
        .ZN(n257) );
  MUX2ND0 U706 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n545), 
        .ZN(n256) );
  MUX3ND0 U707 ( .I0(n260), .I1(n259), .I2(n255), .S0(n513), .S1(n505), .ZN(
        n267) );
  MUX2ND0 U708 ( .I0(n262), .I1(n261), .S(n511), .ZN(n266) );
  MUX2ND0 U709 ( .I0(n264), .I1(n263), .S(n511), .ZN(n265) );
  MUX2ND0 U710 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n545), 
        .ZN(n270) );
  MUX2ND0 U711 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n546), 
        .ZN(n269) );
  MUX3ND0 U712 ( .I0(n273), .I1(n272), .I2(n268), .S0(n513), .S1(n505), .ZN(
        n280) );
  MUX2ND0 U713 ( .I0(n275), .I1(n274), .S(n511), .ZN(n279) );
  MUX2ND0 U714 ( .I0(n277), .I1(n276), .S(N45), .ZN(n278) );
  MUX2ND0 U715 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n545), 
        .ZN(n283) );
  MUX2ND0 U716 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n545), 
        .ZN(n282) );
  MUX3ND0 U717 ( .I0(n286), .I1(n285), .I2(n281), .S0(n514), .S1(n505), .ZN(
        n293) );
  MUX2ND0 U718 ( .I0(n288), .I1(n287), .S(N45), .ZN(n292) );
  MUX2ND0 U719 ( .I0(n290), .I1(n289), .S(N45), .ZN(n291) );
  MUX2ND0 U720 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n545), 
        .ZN(n296) );
  MUX2ND0 U721 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n545), 
        .ZN(n295) );
  MUX3ND0 U722 ( .I0(n299), .I1(n298), .I2(n294), .S0(n514), .S1(n505), .ZN(
        n306) );
  MUX2ND0 U723 ( .I0(n301), .I1(n300), .S(N45), .ZN(n305) );
  MUX2ND0 U724 ( .I0(n303), .I1(n302), .S(n663), .ZN(n304) );
  MUX2ND0 U725 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n545), 
        .ZN(n309) );
  MUX2ND0 U726 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n545), 
        .ZN(n308) );
  MUX3ND0 U727 ( .I0(n312), .I1(n311), .I2(n307), .S0(n514), .S1(n505), .ZN(
        n319) );
  MUX2ND0 U728 ( .I0(n314), .I1(n313), .S(n663), .ZN(n318) );
  MUX2ND0 U729 ( .I0(n316), .I1(n315), .S(n508), .ZN(n317) );
  MUX2ND0 U730 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n545), 
        .ZN(n322) );
  MUX2ND0 U731 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n545), 
        .ZN(n321) );
  MUX3ND0 U732 ( .I0(n325), .I1(n324), .I2(n320), .S0(n513), .S1(n504), .ZN(
        n332) );
  MUX2ND0 U733 ( .I0(n327), .I1(n326), .S(n663), .ZN(n331) );
  MUX2ND0 U734 ( .I0(n329), .I1(n328), .S(n510), .ZN(n330) );
  MUX2ND0 U735 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n545), 
        .ZN(n335) );
  MUX2ND0 U736 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n544), 
        .ZN(n334) );
  MUX3ND0 U737 ( .I0(n338), .I1(n337), .I2(n333), .S0(n514), .S1(n504), .ZN(
        n345) );
  MUX2ND0 U738 ( .I0(n340), .I1(n339), .S(n509), .ZN(n344) );
  MUX2ND0 U739 ( .I0(n342), .I1(n341), .S(N45), .ZN(n343) );
  MUX2ND0 U740 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n544), 
        .ZN(n348) );
  MUX2ND0 U741 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n544), 
        .ZN(n347) );
  MUX3ND0 U742 ( .I0(n351), .I1(n350), .I2(n346), .S0(n513), .S1(n504), .ZN(
        n358) );
  MUX2ND0 U743 ( .I0(n353), .I1(n352), .S(n508), .ZN(n357) );
  MUX2ND0 U744 ( .I0(n355), .I1(n354), .S(n515), .ZN(n356) );
  MUX2ND0 U745 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n544), 
        .ZN(n361) );
  MUX2ND0 U746 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n544), 
        .ZN(n360) );
  MUX3ND0 U747 ( .I0(n364), .I1(n363), .I2(n359), .S0(n515), .S1(n504), .ZN(
        n371) );
  MUX2ND0 U748 ( .I0(n366), .I1(n365), .S(n508), .ZN(n370) );
  MUX2ND0 U749 ( .I0(n368), .I1(n367), .S(n509), .ZN(n369) );
  MUX2ND0 U750 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n544), 
        .ZN(n374) );
  MUX2ND0 U751 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n544), 
        .ZN(n373) );
  MUX3ND0 U752 ( .I0(n377), .I1(n376), .I2(n372), .S0(n514), .S1(n504), .ZN(
        n384) );
  MUX2ND0 U753 ( .I0(n379), .I1(n378), .S(n509), .ZN(n383) );
  MUX2ND0 U754 ( .I0(n381), .I1(n380), .S(n509), .ZN(n382) );
  MUX2ND0 U755 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n544), 
        .ZN(n387) );
  MUX2ND0 U756 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n544), 
        .ZN(n386) );
  MUX3ND0 U757 ( .I0(n390), .I1(n389), .I2(n385), .S0(n514), .S1(n504), .ZN(
        n397) );
  MUX2ND0 U758 ( .I0(n392), .I1(n391), .S(n509), .ZN(n396) );
  MUX2ND0 U759 ( .I0(n394), .I1(n393), .S(n509), .ZN(n395) );
  MUX2ND0 U760 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n544), 
        .ZN(n400) );
  MUX2ND0 U761 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n544), 
        .ZN(n399) );
  MUX3ND0 U762 ( .I0(n403), .I1(n402), .I2(n398), .S0(n514), .S1(n504), .ZN(
        n410) );
  MUX2ND0 U763 ( .I0(n405), .I1(n404), .S(n509), .ZN(n409) );
  MUX2ND0 U764 ( .I0(n407), .I1(n406), .S(n509), .ZN(n408) );
  MUX2ND0 U765 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n544), 
        .ZN(n413) );
  MUX2ND0 U766 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n543), 
        .ZN(n412) );
  MUX3ND0 U767 ( .I0(n416), .I1(n415), .I2(n411), .S0(n515), .S1(n504), .ZN(
        n423) );
  MUX2ND0 U768 ( .I0(n418), .I1(n417), .S(n509), .ZN(n422) );
  MUX2ND0 U769 ( .I0(n420), .I1(n419), .S(n509), .ZN(n421) );
  MUX2ND0 U770 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n543), 
        .ZN(n426) );
  MUX2ND0 U771 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n543), 
        .ZN(n425) );
  MUX3ND0 U772 ( .I0(n429), .I1(n428), .I2(n424), .S0(n514), .S1(n504), .ZN(
        n436) );
  MUX2ND0 U773 ( .I0(n431), .I1(n430), .S(n509), .ZN(n435) );
  MUX2ND0 U774 ( .I0(n433), .I1(n432), .S(n509), .ZN(n434) );
  MUX2ND0 U775 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n543), 
        .ZN(n439) );
  MUX2ND0 U776 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n543), 
        .ZN(n438) );
  MUX3ND0 U777 ( .I0(n442), .I1(n441), .I2(n437), .S0(n515), .S1(n504), .ZN(
        n449) );
  MUX2ND0 U778 ( .I0(n444), .I1(n443), .S(n509), .ZN(n448) );
  MUX2ND0 U779 ( .I0(n446), .I1(n445), .S(n509), .ZN(n447) );
  MUX2ND0 U780 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n543), 
        .ZN(n452) );
  MUX2ND0 U781 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n543), 
        .ZN(n451) );
  MUX3ND0 U782 ( .I0(n455), .I1(n454), .I2(n450), .S0(n515), .S1(n504), .ZN(
        n462) );
  MUX2ND0 U783 ( .I0(n457), .I1(n456), .S(N45), .ZN(n461) );
  MUX2ND0 U784 ( .I0(n459), .I1(n458), .S(n663), .ZN(n460) );
  MUX2ND0 U785 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n543), 
        .ZN(n465) );
  MUX2ND0 U786 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n543), 
        .ZN(n464) );
  MUX3ND0 U787 ( .I0(n468), .I1(n467), .I2(n463), .S0(n515), .S1(n504), .ZN(
        n475) );
  MUX2ND0 U788 ( .I0(n470), .I1(n469), .S(N45), .ZN(n474) );
  MUX2ND0 U789 ( .I0(n472), .I1(n471), .S(n509), .ZN(n473) );
  MUX2ND0 U790 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n543), 
        .ZN(n478) );
  MUX2ND0 U791 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n543), 
        .ZN(n477) );
  MUX3ND0 U792 ( .I0(n481), .I1(n480), .I2(n476), .S0(n515), .S1(n504), .ZN(
        n488) );
  MUX2ND0 U793 ( .I0(n483), .I1(n482), .S(N45), .ZN(n487) );
  MUX2ND0 U794 ( .I0(n485), .I1(n484), .S(n514), .ZN(n486) );
  MUX2ND0 U795 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n542), 
        .ZN(n491) );
  MUX2ND0 U796 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n546), 
        .ZN(n490) );
  MUX3ND0 U797 ( .I0(n494), .I1(n493), .I2(n489), .S0(n515), .S1(n505), .ZN(
        n501) );
  MUX2ND0 U798 ( .I0(n496), .I1(n495), .S(N45), .ZN(n500) );
  MUX2ND0 U799 ( .I0(n498), .I1(n497), .S(n511), .ZN(n499) );
  INVD0 U800 ( .I(Read), .ZN(n90) );
endmodule


module FIFOStateM_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(SUM[5]), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKND0 U1 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_DW01_inc_4 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

