��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5�h��%��Xcbp��'����Q4KҲ��r�D� �m�'�t�חEʭ�3�Jld��q�G�~��Z2��˝1~OT������oPY̅���c�PƐt
׫�J��q{�f��a�:&�>��s�z+/�c�Z�J
_䆼�\�v�����{�{\J�yG����y��\�vť���ҧ`�S�*H������=t����w���@�|��].��'���Xwd�n]Nِ����_H;a(􆿳���A�b,�my$�N���Uە��GV��y�&_3#ڸZ鎬����D�OBp�b}��BB϶q��{l�f|�ό���.Ӳ�[O�"���Ig`i�ҋX����@�ڗe'��E4�Mʸ|��].��'���Xw�-X��-���Ig`i�ҋX����@�ڗe'�@.�>�ȼ�|��].��'���Xw����UA����Ig`i7G#+���[H�����2��~��o�b�x�'�6LE�EYZ/���)֨9 >�j��O0E>�������fHa��!A{�H]�%�Iߎn?�e"�2ao
r��FE���r#�9l$���޸�����C�O"I��MjX��k���`���F(ĕL2	X�vb�)�S�����]�c.��'1����1\���k�e1i��Q,�&d���ݚev3Y�IkT˱ ��O�������]�U�����8�o��@�<�qؚ��L�NG�>)�����7������7�� �����R=�;@R��Ω�dBj#/����@$˺/tw�ԝD=��٭@�FϟQ�-i�`�g``FD�e3>�ƙ�Ǘ���mC��XH�����wI�d��`���1�E��)֨9 E3����=E�EYZ/�@�L0�6#����"'W�9�p��y��9��L����Lo�I��'��恭�h�I��'�%�e���Ĕ^ֻ��X�x%}�����
D�5tm�c�oL�~j�F},M�5����`K�����svfY������;5B5Y+���o�(�)��;U��tm�c�oL�������FTVP��b�M:�8U(�d�٣��c�A�L'��y�!�;&����˚�T�\ �����j�|�z#:rQ��q�X�G[��;ۂ���cY�~�"���ʷ��1�(ʌ�N�M8�U����t��h~��J����^Mf���9���q���U�pzl��a��i��؂ۃ�y�wjאﻋ-�����S8�l��`�_gi�.�!����Wy����`y����s��d�\��MN����!I/�������A��X�@�5��6�l��sХ+�:R 8*!Ē\��c�PƐt
�20)�_�5�e��a)�m�d�so�}a�C�ub;�;���A���g?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��LC6���i��y�L*���8�^�.eO��q��S��;�(e)��v��=����'�$��u,��y�"���Չ-d��r�b+��/6!��Ei�gz�����n�|W;"V7��evwJ���&�o�\,9o$aϛ`!�A���
+,I�2Sj�	�$ɜ�\�۟�-?�d���&����{ԕ�h7�{`��������* -��ed.:E������ƄH����[��2����s�Z�. |�����D�U(�	~nU�L���႔}��xq)�:"ɽ�gW��t_!0h��(Z+�<Vo�eo[߽�M�b�_gi�.�!6PJAzs�U�R�X��3){]�8�~�G4PN��g��U-�eJ+*H�)��>J�p����Q��x�$��J����^�%�[�:V�SƠ��b��7��e�A*"v%)��2������K��A7����C �v��Z�	�і��>Y!���b"��6[�F/��d�>q��,E��n
V~$����[����J����^<���Hn
V~$�E��<^�_�;+�}�pPo��z�#�>B���nF���<�W�.�P��Dbgo���M�ܚp:���fM��X��WG ���}�h�b�B~fQ0�u]9�#�I�X��WG ����7��� �24���W��\v�9�i	A��Z���Ӗ��x�?�+��d��MT�+	�}.�A��R�ߋQ"���_ޓ�@�Ԕ�LS���W)��/807���>�V�T۳�͕���ƒtJ�Ʌ�X�G[�cGK��W�X�G[�����5Orw�&�z<a��r�����K�J�����s��qs����>�C�;��,��V�.o)�\���&%�_1�/�hA��R�ߋ\5�/ X���͖n��r)��"�l���n�2�����t;�i��؂����p���m��Jc�}���F��靤�}O�"L?���H��+��g&)�6�=�#��-���g��U-�e7sQ��4����+9�:�m(��a(􆿳�^~>��m+�����Ur�K�f�AjHt��t��Q��rw�&�z<aSm�6��`4�04�jf�5ߧE4��Fi��|�3;c�<𷜏���'�֔�"�we����e�fke��.���E.t�