
module BIST_AWid5_DWid32_DW01_inc_5 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_4 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module BIST_AWid5_DWid32 ( DataO, Addr, ReadCmd, WriteCmd, Testing, TestOK, 
        DataI, DoSelfTest, ParityErr, Clk, Reset );
  output [31:0] DataO;
  output [4:0] Addr;
  input [31:0] DataI;
  input DoSelfTest, ParityErr, Clk, Reset;
  output ReadCmd, WriteCmd, Testing, TestOK;
  wire   n294, TDone5, TDone3, TDone1, TRes5, TRes3, TRes1, AllDoner, N132,
         N138, N145, N151, N158, N165, N170, N172, N184, N185, N186, N203,
         N204, N205, N206, N208, N210, N211, N212, N214, N216, N217, N218,
         N219, N220, N226, N227, N228, N229, N230, N233, N272, N284, N285,
         N286, N287, N288, N319, N320, N321, N322, N323, N326, N364, N370,
         N371, N372, N373, N374, N404, N405, N406, N407, N408, N411, N449,
         N455, N456, N457, N458, N459, n204, n206, n208, n210, n212, n216,
         n218, n220, n222, n224, n228, n230, n232, n234, n237, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n205, n207, n209, n211, n213, n214, n215,
         n217, n219, n221, n223, n225, n226, n227, n229, n231, n233, n235,
         n236, n238, n239, n240, n287, n288, n289, n290, n291, n292, n293;
  wire   [6:1] TestDone;
  wire   [2:0] TestNo;
  wire   [4:0] Addr1;
  wire   [4:0] Addr3;
  wire   [4:0] Addr5;
  wire   [31:0] DataO1;
  wire   [2:0] State;
  wire   [4:0] i1;
  wire   [4:0] i2;
  wire   [4:0] i3;
  wire   [4:0] i4;
  wire   [4:0] i5;
  wire   [4:0] i6;
  assign DataO[31] = N364;

  DFND1 \Addr2_reg[3]  ( .D(n283), .CPN(Clk), .Q(n239), .QN(n22) );
  DFND1 \Addr2_reg[0]  ( .D(n281), .CPN(Clk), .Q(n291), .QN(n18) );
  DFND1 \Addr2_reg[1]  ( .D(n279), .CPN(Clk), .Q(n289), .QN(n19) );
  DFND1 \Addr2_reg[2]  ( .D(n277), .CPN(Clk), .Q(n287), .QN(n20) );
  DFND1 \Addr2_reg[4]  ( .D(n275), .CPN(Clk), .Q(n236), .QN(n21) );
  DFND1 \Addr4_reg[3]  ( .D(n270), .CPN(Clk), .Q(n240), .QN(n23) );
  DFND1 \Addr4_reg[0]  ( .D(n268), .CPN(Clk), .Q(n292), .QN(n14) );
  DFND1 \Addr4_reg[1]  ( .D(n266), .CPN(Clk), .Q(n290), .QN(n15) );
  DFND1 \Addr4_reg[2]  ( .D(n264), .CPN(Clk), .Q(n288), .QN(n16) );
  DFND1 \Addr4_reg[4]  ( .D(n262), .CPN(Clk), .Q(n238), .QN(n17) );
  DFND1 \Addr6_reg[3]  ( .D(n251), .CPN(Clk), .QN(n10) );
  DFND1 \Addr6_reg[0]  ( .D(n249), .CPN(Clk), .QN(n9) );
  DFND1 \Addr6_reg[1]  ( .D(n247), .CPN(Clk), .QN(n8) );
  DFND1 \Addr6_reg[2]  ( .D(n245), .CPN(Clk), .QN(n7) );
  DFND1 \Addr6_reg[4]  ( .D(n243), .CPN(Clk), .QN(n6) );
  BIST_AWid5_DWid32_DW01_inc_0 \TestPhase06/DelayedSample/add_544  ( .A(i6), 
        .SUM({N459, N458, N457, N456, N455}) );
  BIST_AWid5_DWid32_DW01_inc_1 \TestPhase05/add_506  ( .A(i5), .SUM({N408, 
        N407, N406, N405, N404}) );
  BIST_AWid5_DWid32_DW01_inc_2 \TestPhase04/DelayedSample/add_476  ( .A(i4), 
        .SUM({N374, N373, N372, N371, N370}) );
  BIST_AWid5_DWid32_DW01_inc_3 \TestPhase03/add_438  ( .A(i3), .SUM({N323, 
        N322, N321, N320, N319}) );
  BIST_AWid5_DWid32_DW01_inc_4 \TestPhase02/DelayedSample/add_408  ( .A(i2), 
        .SUM({N288, N287, N286, N285, N284}) );
  BIST_AWid5_DWid32_DW01_inc_5 \TestPhase01/add_366  ( .A(i1), .SUM({N230, 
        N229, N228, N227, N226}) );
  DFNSND1 Wait2_reg ( .D(n274), .CPN(Clk), .SDN(n286), .Q(n3), .QN(n227) );
  DFNSND1 Wait4_reg ( .D(n272), .CPN(Clk), .SDN(n286), .Q(n1), .QN(n226) );
  DFNSND1 Wait6_reg ( .D(n253), .CPN(Clk), .SDN(n286), .Q(n2), .QN(n229) );
  EDFQD1 \DataO1_reg[27]  ( .D(i1[3]), .E(N272), .CP(Clk), .Q(DataO1[27]) );
  EDFQD1 \DataO1_reg[25]  ( .D(i1[1]), .E(N272), .CP(Clk), .Q(DataO1[25]) );
  EDFQD1 \DataO1_reg[19]  ( .D(i1[3]), .E(N272), .CP(Clk), .Q(DataO1[19]) );
  EDFQD1 \DataO1_reg[17]  ( .D(i1[1]), .E(N272), .CP(Clk), .Q(DataO1[17]) );
  EDFQD1 \DataO1_reg[11]  ( .D(i1[3]), .E(N272), .CP(Clk), .Q(DataO1[11]) );
  EDFQD1 \DataO1_reg[9]  ( .D(i1[1]), .E(N272), .CP(Clk), .Q(DataO1[9]) );
  EDFQD1 \DataO1_reg[3]  ( .D(i1[3]), .E(N272), .CP(Clk), .Q(DataO1[3]) );
  EDFQD1 \DataO1_reg[1]  ( .D(i1[1]), .E(N272), .CP(Clk), .Q(DataO1[1]) );
  EDFQD1 \DataO1_reg[0]  ( .D(i1[0]), .E(N272), .CP(Clk), .Q(DataO1[0]) );
  EDFQD1 \DataO1_reg[2]  ( .D(i1[2]), .E(N272), .CP(Clk), .Q(DataO1[2]) );
  EDFQD1 \DataO1_reg[4]  ( .D(i1[4]), .E(N272), .CP(Clk), .Q(DataO1[4]) );
  EDFQD1 \DataO1_reg[8]  ( .D(i1[0]), .E(N272), .CP(Clk), .Q(DataO1[8]) );
  EDFQD1 \DataO1_reg[10]  ( .D(i1[2]), .E(N272), .CP(Clk), .Q(DataO1[10]) );
  EDFQD1 \DataO1_reg[12]  ( .D(i1[4]), .E(N272), .CP(Clk), .Q(DataO1[12]) );
  EDFQD1 \DataO1_reg[16]  ( .D(i1[0]), .E(N272), .CP(Clk), .Q(DataO1[16]) );
  EDFQD1 \DataO1_reg[18]  ( .D(i1[2]), .E(N272), .CP(Clk), .Q(DataO1[18]) );
  EDFQD1 \DataO1_reg[20]  ( .D(i1[4]), .E(N272), .CP(Clk), .Q(DataO1[20]) );
  EDFQD1 \DataO1_reg[24]  ( .D(i1[0]), .E(N272), .CP(Clk), .Q(DataO1[24]) );
  EDFQD1 \DataO1_reg[26]  ( .D(i1[2]), .E(N272), .CP(Clk), .Q(DataO1[26]) );
  EDFQD1 \DataO1_reg[28]  ( .D(i1[4]), .E(N272), .CP(Clk), .Q(DataO1[28]) );
  EDFQD1 \Addr1_reg[4]  ( .D(i1[4]), .E(N272), .CP(Clk), .Q(Addr1[4]) );
  EDFQD1 \Addr1_reg[2]  ( .D(i1[2]), .E(N272), .CP(Clk), .Q(Addr1[2]) );
  EDFQD1 \Addr1_reg[0]  ( .D(i1[0]), .E(N272), .CP(Clk), .Q(Addr1[0]) );
  EDFQD1 \Addr1_reg[1]  ( .D(i1[1]), .E(N272), .CP(Clk), .Q(Addr1[1]) );
  EDFQD1 \Addr1_reg[3]  ( .D(i1[3]), .E(N272), .CP(Clk), .Q(Addr1[3]) );
  EDFQD1 \Addr3_reg[4]  ( .D(i3[4]), .E(N364), .CP(Clk), .Q(Addr3[4]) );
  EDFQD1 \Addr3_reg[2]  ( .D(i3[2]), .E(N364), .CP(Clk), .Q(Addr3[2]) );
  EDFQD1 \Addr3_reg[0]  ( .D(i3[0]), .E(N364), .CP(Clk), .Q(Addr3[0]) );
  EDFQD1 \Addr3_reg[1]  ( .D(i3[1]), .E(N364), .CP(Clk), .Q(Addr3[1]) );
  EDFQD1 \Addr3_reg[3]  ( .D(i3[3]), .E(N364), .CP(Clk), .Q(Addr3[3]) );
  EDFQD1 \Addr5_reg[4]  ( .D(i5[4]), .E(N449), .CP(Clk), .Q(Addr5[4]) );
  EDFQD1 \Addr5_reg[2]  ( .D(i5[2]), .E(N449), .CP(Clk), .Q(Addr5[2]) );
  EDFQD1 \Addr5_reg[0]  ( .D(i5[0]), .E(N449), .CP(Clk), .Q(Addr5[0]) );
  EDFQD1 \Addr5_reg[1]  ( .D(i5[1]), .E(N449), .CP(Clk), .Q(Addr5[1]) );
  EDFQD1 \Addr5_reg[3]  ( .D(i5[3]), .E(N449), .CP(Clk), .Q(Addr5[3]) );
  DFNCND1 \i2_reg[4]  ( .D(n276), .CPN(Clk), .CDN(n286), .Q(i2[4]), .QN(n228)
         );
  DFNCND1 \i4_reg[4]  ( .D(n263), .CPN(Clk), .CDN(n286), .Q(i4[4]), .QN(n216)
         );
  DFNCND1 \i6_reg[4]  ( .D(n244), .CPN(Clk), .CDN(n286), .Q(i6[4]), .QN(n204)
         );
  DFNCND1 TDone6_reg ( .D(n285), .CPN(Clk), .CDN(n286), .QN(n11) );
  DFNCND1 TDone4_reg ( .D(n260), .CPN(Clk), .CDN(n286), .QN(n12) );
  DFNCND1 TDone2_reg ( .D(n241), .CPN(Clk), .CDN(n286), .QN(n13) );
  EDFCNQD1 WriteCmdr_reg ( .D(N186), .E(n4), .CP(Clk), .CDN(n286), .Q(WriteCmd) );
  EDFCNQD1 ReadCmdr_reg ( .D(N185), .E(n4), .CP(Clk), .CDN(n286), .Q(ReadCmd)
         );
  DFCNQD1 TRes1_reg ( .D(n259), .CP(Clk), .CDN(n286), .Q(TRes1) );
  DFCNQD1 TDone1_reg ( .D(n258), .CP(Clk), .CDN(n286), .Q(TDone1) );
  DFCNQD1 TRes5_reg ( .D(n255), .CP(Clk), .CDN(n286), .Q(TRes5) );
  DFCNQD1 TDone3_reg ( .D(n256), .CP(Clk), .CDN(n286), .Q(TDone3) );
  DFCNQD1 TDone5_reg ( .D(n254), .CP(Clk), .CDN(n286), .Q(TDone5) );
  EDFCNQD1 AllDoner_reg ( .D(N206), .E(N205), .CP(Clk), .CDN(n286), .Q(
        AllDoner) );
  EDFCNQD1 \i3_reg[4]  ( .D(N323), .E(N326), .CP(Clk), .CDN(n286), .Q(i3[4])
         );
  EDFCNQD1 \i5_reg[4]  ( .D(N408), .E(N411), .CP(Clk), .CDN(n286), .Q(i5[4])
         );
  DFNCND1 \i2_reg[3]  ( .D(n284), .CPN(Clk), .CDN(n286), .Q(i2[3]), .QN(n237)
         );
  DFNCND1 \i2_reg[1]  ( .D(n280), .CPN(Clk), .CDN(n286), .Q(i2[1]), .QN(n232)
         );
  DFNCND1 \i2_reg[2]  ( .D(n278), .CPN(Clk), .CDN(n286), .Q(i2[2]), .QN(n230)
         );
  DFNCND1 \i4_reg[3]  ( .D(n271), .CPN(Clk), .CDN(n286), .Q(i4[3]), .QN(n224)
         );
  DFNCND1 \i4_reg[1]  ( .D(n267), .CPN(Clk), .CDN(n286), .Q(i4[1]), .QN(n220)
         );
  DFNCND1 \i4_reg[2]  ( .D(n265), .CPN(Clk), .CDN(n286), .Q(i4[2]), .QN(n218)
         );
  DFNCND1 \i6_reg[3]  ( .D(n252), .CPN(Clk), .CDN(n286), .Q(i6[3]), .QN(n212)
         );
  DFNCND1 \i6_reg[1]  ( .D(n248), .CPN(Clk), .CDN(n286), .Q(i6[1]), .QN(n208)
         );
  DFNCND1 \i6_reg[2]  ( .D(n246), .CPN(Clk), .CDN(n286), .Q(i6[2]), .QN(n206)
         );
  DFNCND1 \i2_reg[0]  ( .D(n282), .CPN(Clk), .CDN(n286), .Q(i2[0]), .QN(n234)
         );
  DFNCND1 \i4_reg[0]  ( .D(n269), .CPN(Clk), .CDN(n286), .Q(i4[0]), .QN(n222)
         );
  DFNCND1 \i6_reg[0]  ( .D(n250), .CPN(Clk), .CDN(n286), .Q(i6[0]), .QN(n210)
         );
  DFNCND1 TRes6_reg ( .D(n242), .CPN(Clk), .CDN(n286), .Q(n231) );
  DFCNQD1 TRes3_reg ( .D(n257), .CP(Clk), .CDN(n286), .Q(TRes3) );
  EDFCNQD1 \TestNo_reg[2]  ( .D(N212), .E(N211), .CP(Clk), .CDN(n286), .Q(
        TestNo[2]) );
  EDFCND1 \TestNo_reg[1]  ( .D(N210), .E(N211), .CP(Clk), .CDN(n286), .Q(n293), 
        .QN(n5) );
  EDFCNQD1 \i3_reg[1]  ( .D(N320), .E(N326), .CP(Clk), .CDN(n286), .Q(i3[1])
         );
  EDFCNQD1 \i3_reg[2]  ( .D(N321), .E(N326), .CP(Clk), .CDN(n286), .Q(i3[2])
         );
  EDFCNQD1 \i3_reg[3]  ( .D(N322), .E(N326), .CP(Clk), .CDN(n286), .Q(i3[3])
         );
  EDFCNQD1 \i5_reg[1]  ( .D(N405), .E(N411), .CP(Clk), .CDN(n286), .Q(i5[1])
         );
  EDFCNQD1 \i5_reg[2]  ( .D(N406), .E(N411), .CP(Clk), .CDN(n286), .Q(i5[2])
         );
  EDFCNQD1 \i5_reg[3]  ( .D(N407), .E(N411), .CP(Clk), .CDN(n286), .Q(i5[3])
         );
  EDFCNQD1 \i3_reg[0]  ( .D(N319), .E(N326), .CP(Clk), .CDN(n286), .Q(i3[0])
         );
  EDFCNQD1 \i5_reg[0]  ( .D(N404), .E(N411), .CP(Clk), .CDN(n286), .Q(i5[0])
         );
  DFNCND1 TRes2_reg ( .D(n273), .CPN(Clk), .CDN(n286), .Q(n235) );
  DFNCND1 TRes4_reg ( .D(n261), .CPN(Clk), .CDN(n286), .Q(n233) );
  EDFCNQD1 \TestNo_reg[0]  ( .D(N208), .E(N211), .CP(Clk), .CDN(n286), .Q(
        TestNo[0]) );
  EDFCNQD1 \i1_reg[4]  ( .D(N230), .E(N233), .CP(Clk), .CDN(n286), .Q(i1[4])
         );
  EDFCNQD1 \i1_reg[1]  ( .D(N227), .E(N233), .CP(Clk), .CDN(n286), .Q(i1[1])
         );
  EDFCNQD1 \i1_reg[2]  ( .D(N228), .E(N233), .CP(Clk), .CDN(n286), .Q(i1[2])
         );
  EDFCNQD1 \i1_reg[3]  ( .D(N229), .E(N233), .CP(Clk), .CDN(n286), .Q(i1[3])
         );
  EDFCNQD1 \i1_reg[0]  ( .D(N226), .E(N233), .CP(Clk), .CDN(n286), .Q(i1[0])
         );
  EDFCNQD1 \State_reg[1]  ( .D(N216), .E(N217), .CP(Clk), .CDN(n286), .Q(
        State[1]) );
  EDFCNQD1 \State_reg[2]  ( .D(N218), .E(N217), .CP(Clk), .CDN(n286), .Q(
        State[2]) );
  EDFCNQD1 \State_reg[0]  ( .D(N214), .E(N217), .CP(Clk), .CDN(n286), .Q(
        State[0]) );
  EDFCNQD1 Testingr_reg ( .D(N204), .E(N203), .CP(Clk), .CDN(n286), .Q(Testing) );
  EDFCNQD1 TestOKr_reg ( .D(N220), .E(N219), .CP(Clk), .CDN(n286), .Q(n294) );
  ND2D1 U3 ( .A1(N326), .A2(n286), .ZN(n205) );
  NR3D0 U4 ( .A1(AllDoner), .A2(ParityErr), .A3(n201), .ZN(n4) );
  AN2D2 U5 ( .A1(N233), .A2(n286), .Z(N272) );
  CKBD0 U6 ( .CLK(n26), .C(n24) );
  CKNXD16 U7 ( .I(n24), .ZN(TestOK) );
  CKND0 U8 ( .CLK(n294), .CN(n26) );
  INVD3 U9 ( .I(Reset), .ZN(n286) );
  CKND0 U10 ( .CLK(Testing), .CN(n27) );
  NR2XD0 U11 ( .A1(n27), .A2(n198), .ZN(n166) );
  INVD0 U12 ( .I(n200), .ZN(n165) );
  CKAN2D0 U13 ( .A1(N411), .A2(n286), .Z(N449) );
  NR2D1 U14 ( .A1(n74), .A2(Reset), .ZN(n65) );
  NR2D1 U15 ( .A1(n86), .A2(Reset), .ZN(n78) );
  CKAN2D0 U16 ( .A1(TDone3), .A2(n286), .Z(TestDone[3]) );
  CKAN2D0 U17 ( .A1(TDone5), .A2(n286), .Z(TestDone[5]) );
  INR2D1 U18 ( .A1(State[0]), .B1(TestDone[1]), .ZN(n43) );
  ND2D1 U19 ( .A1(State[0]), .A2(N132), .ZN(n47) );
  INR2D1 U20 ( .A1(State[0]), .B1(N132), .ZN(n44) );
  INR2D1 U21 ( .A1(State[0]), .B1(N132), .ZN(n45) );
  MUX3ND0 U22 ( .I0(n43), .I1(n58), .I2(n57), .S0(State[2]), .S1(State[1]), 
        .ZN(n28) );
  AN2D1 U23 ( .A1(TestDone[6]), .A2(n161), .Z(n50) );
  INVD1 U24 ( .I(n205), .ZN(DataO[30]) );
  INVD1 U25 ( .I(n205), .ZN(DataO[29]) );
  INVD1 U26 ( .I(n205), .ZN(DataO[23]) );
  INVD1 U27 ( .I(n205), .ZN(DataO[22]) );
  INVD1 U28 ( .I(n205), .ZN(DataO[21]) );
  INVD1 U29 ( .I(n205), .ZN(DataO[15]) );
  INVD1 U30 ( .I(n205), .ZN(DataO[14]) );
  INVD1 U31 ( .I(n205), .ZN(DataO[13]) );
  INVD1 U32 ( .I(n205), .ZN(DataO[7]) );
  INVD1 U33 ( .I(n205), .ZN(DataO[6]) );
  INVD1 U34 ( .I(n205), .ZN(DataO[5]) );
  OR2D1 U35 ( .A1(N165), .A2(State[0]), .Z(n46) );
  MUX3ND0 U36 ( .I0(n47), .I1(n48), .I2(n49), .S0(State[2]), .S1(State[1]), 
        .ZN(N184) );
  OR2D1 U37 ( .A1(N165), .A2(State[0]), .Z(n51) );
  MUX3ND0 U38 ( .I0(n44), .I1(n52), .I2(n53), .S0(State[2]), .S1(State[1]), 
        .ZN(N172) );
  OR2D1 U39 ( .A1(N165), .A2(State[0]), .Z(n54) );
  MUX3ND0 U40 ( .I0(n45), .I1(n55), .I2(n56), .S0(State[2]), .S1(State[1]), 
        .ZN(N170) );
  MUX3ND0 U41 ( .I0(N138), .I1(N145), .I2(n46), .S0(State[0]), .S1(State[2]), 
        .ZN(n49) );
  MUX2ND0 U42 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n48) );
  MUX3ND0 U43 ( .I0(TestDone[2]), .I1(TestDone[3]), .I2(n50), .S0(State[0]), 
        .S1(State[2]), .ZN(n57) );
  MUX2ND0 U44 ( .I0(TestDone[4]), .I1(TestDone[5]), .S(State[0]), .ZN(n58) );
  MUX3ND0 U45 ( .I0(N138), .I1(N145), .I2(n51), .S0(State[0]), .S1(State[2]), 
        .ZN(n53) );
  MUX2ND0 U46 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n52) );
  MUX3ND0 U47 ( .I0(N138), .I1(N145), .I2(n54), .S0(State[0]), .S1(State[2]), 
        .ZN(n56) );
  MUX2ND0 U48 ( .I0(N151), .I1(N158), .S(State[0]), .ZN(n55) );
  OAI31D0 U49 ( .A1(n2), .A2(n59), .A3(n60), .B(n11), .ZN(n285) );
  AN2D0 U50 ( .A1(n61), .A2(n62), .Z(n59) );
  MUX2ND0 U51 ( .I0(n63), .I1(n237), .S(n64), .ZN(n284) );
  MUX2ND0 U52 ( .I0(n22), .I1(n237), .S(n65), .ZN(n283) );
  MUX2ND0 U53 ( .I0(n66), .I1(n234), .S(n64), .ZN(n282) );
  MUX2ND0 U54 ( .I0(n18), .I1(n234), .S(n65), .ZN(n281) );
  MUX2ND0 U55 ( .I0(n67), .I1(n232), .S(n64), .ZN(n280) );
  MUX2ND0 U56 ( .I0(n19), .I1(n232), .S(n65), .ZN(n279) );
  MUX2ND0 U57 ( .I0(n68), .I1(n230), .S(n64), .ZN(n278) );
  CKND0 U58 ( .CLK(N286), .CN(n68) );
  MUX2ND0 U59 ( .I0(n20), .I1(n230), .S(n65), .ZN(n277) );
  MUX2ND0 U60 ( .I0(n69), .I1(n228), .S(n64), .ZN(n276) );
  CKND0 U61 ( .CLK(N288), .CN(n69) );
  MUX2ND0 U62 ( .I0(n21), .I1(n228), .S(n65), .ZN(n275) );
  OAI21D0 U63 ( .A1(n227), .A2(n70), .B(n64), .ZN(n274) );
  OAI21D0 U64 ( .A1(n64), .A2(n71), .B(n72), .ZN(n273) );
  OAI31D0 U65 ( .A1(n3), .A2(n73), .A3(n74), .B(n235), .ZN(n72) );
  ND3D0 U66 ( .A1(n73), .A2(n70), .A3(n227), .ZN(n64) );
  OAI21D0 U67 ( .A1(n226), .A2(n75), .B(n76), .ZN(n272) );
  MUX2ND0 U68 ( .I0(n77), .I1(n224), .S(n76), .ZN(n271) );
  MUX2ND0 U69 ( .I0(n23), .I1(n224), .S(n78), .ZN(n270) );
  MUX2ND0 U70 ( .I0(n79), .I1(n222), .S(n76), .ZN(n269) );
  MUX2ND0 U71 ( .I0(n14), .I1(n222), .S(n78), .ZN(n268) );
  MUX2ND0 U72 ( .I0(n80), .I1(n220), .S(n76), .ZN(n267) );
  MUX2ND0 U73 ( .I0(n15), .I1(n220), .S(n78), .ZN(n266) );
  MUX2ND0 U74 ( .I0(n81), .I1(n218), .S(n76), .ZN(n265) );
  CKND0 U75 ( .CLK(N372), .CN(n81) );
  MUX2ND0 U76 ( .I0(n16), .I1(n218), .S(n78), .ZN(n264) );
  MUX2ND0 U77 ( .I0(n82), .I1(n216), .S(n76), .ZN(n263) );
  CKND0 U78 ( .CLK(N374), .CN(n82) );
  MUX2ND0 U79 ( .I0(n17), .I1(n216), .S(n78), .ZN(n262) );
  OAI21D0 U80 ( .A1(n76), .A2(n83), .B(n84), .ZN(n261) );
  OAI31D0 U81 ( .A1(n1), .A2(n85), .A3(n86), .B(n233), .ZN(n84) );
  ND3D0 U82 ( .A1(n85), .A2(n75), .A3(n226), .ZN(n76) );
  OAI31D0 U83 ( .A1(n1), .A2(n87), .A3(n86), .B(n12), .ZN(n260) );
  AN2D0 U84 ( .A1(n83), .A2(n85), .Z(n87) );
  AN2D0 U85 ( .A1(n88), .A2(n89), .Z(n85) );
  NR4D0 U86 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(n89) );
  ND4D0 U87 ( .A1(DataI[10]), .A2(DataI[4]), .A3(DataI[2]), .A4(DataI[1]), 
        .ZN(n93) );
  ND4D0 U88 ( .A1(DataI[3]), .A2(DataI[0]), .A3(DataI[28]), .A4(DataI[26]), 
        .ZN(n92) );
  ND4D0 U89 ( .A1(DataI[25]), .A2(DataI[27]), .A3(DataI[20]), .A4(DataI[19]), 
        .ZN(n91) );
  ND4D0 U90 ( .A1(DataI[24]), .A2(DataI[17]), .A3(DataI[16]), .A4(DataI[18]), 
        .ZN(n90) );
  NR4D0 U91 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n88) );
  ND4D0 U92 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[5]), .A4(DataI[31]), 
        .ZN(n97) );
  ND4D0 U93 ( .A1(DataI[30]), .A2(DataI[29]), .A3(DataI[23]), .A4(DataI[22]), 
        .ZN(n96) );
  ND4D0 U94 ( .A1(DataI[21]), .A2(DataI[15]), .A3(DataI[14]), .A4(DataI[13]), 
        .ZN(n95) );
  ND4D0 U95 ( .A1(DataI[9]), .A2(DataI[12]), .A3(DataI[11]), .A4(DataI[8]), 
        .ZN(n94) );
  ND3D0 U96 ( .A1(N374), .A2(N372), .A3(n98), .ZN(n83) );
  NR3D0 U97 ( .A1(n80), .A2(n77), .A3(n79), .ZN(n98) );
  CKND0 U98 ( .CLK(N370), .CN(n79) );
  CKND0 U99 ( .CLK(N373), .CN(n77) );
  CKND0 U100 ( .CLK(N371), .CN(n80) );
  IND2D0 U101 ( .A1(TRes1), .B1(n99), .ZN(n259) );
  IND2D0 U102 ( .A1(TDone1), .B1(n99), .ZN(n258) );
  ND4D0 U103 ( .A1(N226), .A2(N233), .A3(N227), .A4(n100), .ZN(n99) );
  AN3D0 U104 ( .A1(N229), .A2(N228), .A3(N230), .Z(n100) );
  CKND2D0 U105 ( .A1(n101), .A2(n102), .ZN(n257) );
  IND2D0 U106 ( .A1(TDone3), .B1(n102), .ZN(n256) );
  ND4D0 U107 ( .A1(N319), .A2(N326), .A3(N320), .A4(n103), .ZN(n102) );
  AN3D0 U108 ( .A1(N322), .A2(N321), .A3(N323), .Z(n103) );
  IND2D0 U109 ( .A1(TRes5), .B1(n104), .ZN(n255) );
  IND2D0 U110 ( .A1(TDone5), .B1(n104), .ZN(n254) );
  ND4D0 U111 ( .A1(N404), .A2(N411), .A3(N405), .A4(n105), .ZN(n104) );
  AN3D0 U112 ( .A1(N407), .A2(N406), .A3(N408), .Z(n105) );
  OAI21D0 U113 ( .A1(n229), .A2(n106), .B(n107), .ZN(n253) );
  MUX2ND0 U114 ( .I0(n108), .I1(n212), .S(n107), .ZN(n252) );
  CKND0 U115 ( .CLK(N458), .CN(n108) );
  MUX2ND0 U116 ( .I0(n212), .I1(n10), .S(n109), .ZN(n251) );
  MUX2ND0 U117 ( .I0(n110), .I1(n210), .S(n107), .ZN(n250) );
  MUX2ND0 U118 ( .I0(n210), .I1(n9), .S(n109), .ZN(n249) );
  MUX2ND0 U119 ( .I0(n111), .I1(n208), .S(n107), .ZN(n248) );
  MUX2ND0 U120 ( .I0(n208), .I1(n8), .S(n109), .ZN(n247) );
  MUX2ND0 U121 ( .I0(n112), .I1(n206), .S(n107), .ZN(n246) );
  MUX2ND0 U122 ( .I0(n206), .I1(n7), .S(n109), .ZN(n245) );
  MUX2ND0 U123 ( .I0(n113), .I1(n204), .S(n107), .ZN(n244) );
  CKND0 U124 ( .CLK(N459), .CN(n113) );
  MUX2ND0 U125 ( .I0(n204), .I1(n6), .S(n109), .ZN(n243) );
  OAI21D0 U126 ( .A1(n107), .A2(n61), .B(n114), .ZN(n242) );
  OAI31D0 U127 ( .A1(n2), .A2(n62), .A3(n60), .B(n231), .ZN(n114) );
  CKND0 U128 ( .CLK(n106), .CN(n60) );
  ND3D0 U129 ( .A1(N459), .A2(N458), .A3(n115), .ZN(n61) );
  NR3D0 U130 ( .A1(n112), .A2(n110), .A3(n111), .ZN(n115) );
  CKND0 U131 ( .CLK(N456), .CN(n111) );
  CKND0 U132 ( .CLK(N455), .CN(n110) );
  CKND0 U133 ( .CLK(N457), .CN(n112) );
  ND3D0 U134 ( .A1(n106), .A2(n62), .A3(n229), .ZN(n107) );
  AN3D0 U135 ( .A1(n116), .A2(n117), .A3(n118), .Z(n62) );
  INR4D0 U136 ( .A1(n119), .B1(n120), .B2(DataI[24]), .B3(DataI[20]), .ZN(n118) );
  OR3D0 U137 ( .A1(DataI[26]), .A2(DataI[27]), .A3(DataI[25]), .Z(n120) );
  INR4D0 U138 ( .A1(n121), .B1(DataI[2]), .B2(DataI[3]), .B3(DataI[28]), .ZN(
        n119) );
  NR3D0 U139 ( .A1(DataI[4]), .A2(DataI[9]), .A3(DataI[8]), .ZN(n121) );
  NR3D0 U140 ( .A1(n122), .A2(DataI[17]), .A3(DataI[16]), .ZN(n117) );
  OR3D0 U141 ( .A1(DataI[19]), .A2(DataI[1]), .A3(DataI[18]), .Z(n122) );
  NR3D0 U142 ( .A1(n123), .A2(DataI[0]), .A3(n124), .ZN(n116) );
  OR3D0 U143 ( .A1(DataI[11]), .A2(DataI[12]), .A3(DataI[10]), .Z(n123) );
  OAI31D0 U144 ( .A1(n3), .A2(n125), .A3(n74), .B(n13), .ZN(n241) );
  AN2D0 U145 ( .A1(n71), .A2(n73), .Z(n125) );
  AN4D0 U146 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .Z(n73) );
  NR4D0 U147 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .ZN(n129) );
  XNR2D0 U148 ( .A1(n237), .A2(DataI[19]), .ZN(n133) );
  XNR2D0 U149 ( .A1(n234), .A2(DataI[24]), .ZN(n132) );
  XNR2D0 U150 ( .A1(n228), .A2(DataI[20]), .ZN(n131) );
  ND3D0 U151 ( .A1(n134), .A2(n135), .A3(n136), .ZN(n130) );
  CKXOR2D0 U152 ( .A1(n232), .A2(DataI[17]), .Z(n136) );
  CKXOR2D0 U153 ( .A1(n230), .A2(DataI[18]), .Z(n135) );
  CKXOR2D0 U154 ( .A1(n234), .A2(DataI[16]), .Z(n134) );
  NR3D0 U155 ( .A1(n137), .A2(n138), .A3(n139), .ZN(n128) );
  XNR2D0 U156 ( .A1(n234), .A2(DataI[0]), .ZN(n139) );
  XNR2D0 U157 ( .A1(n228), .A2(DataI[28]), .ZN(n138) );
  ND3D0 U158 ( .A1(n140), .A2(n141), .A3(n142), .ZN(n137) );
  CKXOR2D0 U159 ( .A1(n230), .A2(DataI[26]), .Z(n142) );
  CKXOR2D0 U160 ( .A1(n237), .A2(DataI[27]), .Z(n141) );
  CKXOR2D0 U161 ( .A1(n232), .A2(DataI[25]), .Z(n140) );
  NR3D0 U162 ( .A1(n143), .A2(n144), .A3(n145), .ZN(n127) );
  XNR2D0 U163 ( .A1(n230), .A2(DataI[10]), .ZN(n145) );
  XNR2D0 U164 ( .A1(n228), .A2(DataI[4]), .ZN(n144) );
  ND3D0 U165 ( .A1(n146), .A2(n147), .A3(n148), .ZN(n143) );
  CKXOR2D0 U166 ( .A1(n230), .A2(DataI[2]), .Z(n148) );
  CKXOR2D0 U167 ( .A1(n237), .A2(DataI[3]), .Z(n147) );
  CKXOR2D0 U168 ( .A1(n232), .A2(DataI[1]), .Z(n146) );
  NR3D0 U169 ( .A1(n149), .A2(n150), .A3(n124), .ZN(n126) );
  ND4D0 U170 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(n124) );
  NR3D0 U171 ( .A1(DataI[5]), .A2(DataI[7]), .A3(DataI[6]), .ZN(n154) );
  NR3D0 U172 ( .A1(DataI[29]), .A2(DataI[31]), .A3(DataI[30]), .ZN(n153) );
  NR3D0 U173 ( .A1(DataI[21]), .A2(DataI[23]), .A3(DataI[22]), .ZN(n152) );
  NR3D0 U174 ( .A1(DataI[13]), .A2(DataI[15]), .A3(DataI[14]), .ZN(n151) );
  XNR2D0 U175 ( .A1(n232), .A2(DataI[9]), .ZN(n150) );
  ND3D0 U176 ( .A1(n155), .A2(n156), .A3(n157), .ZN(n149) );
  CKXOR2D0 U177 ( .A1(n228), .A2(DataI[12]), .Z(n157) );
  CKXOR2D0 U178 ( .A1(n234), .A2(DataI[8]), .Z(n156) );
  CKXOR2D0 U179 ( .A1(n237), .A2(DataI[11]), .Z(n155) );
  ND3D0 U180 ( .A1(N288), .A2(N286), .A3(n158), .ZN(n71) );
  NR3D0 U181 ( .A1(n67), .A2(n63), .A3(n66), .ZN(n158) );
  CKND0 U182 ( .CLK(N284), .CN(n66) );
  CKND0 U183 ( .CLK(N287), .CN(n63) );
  CKND0 U184 ( .CLK(N285), .CN(n67) );
  NR4D0 U185 ( .A1(n159), .A2(n160), .A3(n161), .A4(n101), .ZN(N220) );
  CKND2D0 U186 ( .A1(n162), .A2(n163), .ZN(n160) );
  ND4D0 U187 ( .A1(n164), .A2(n231), .A3(n233), .A4(n235), .ZN(n159) );
  AO22D0 U188 ( .A1(n165), .A2(ParityErr), .B1(N170), .B2(n166), .Z(N219) );
  AOI31D0 U189 ( .A1(n167), .A2(n168), .A3(n169), .B(n170), .ZN(N218) );
  OA21D0 U190 ( .A1(n171), .A2(n163), .B(n172), .Z(n169) );
  AO21D0 U191 ( .A1(n286), .A2(n235), .B(n173), .Z(n167) );
  IOA21D0 U192 ( .A1(n28), .A2(n4), .B(n174), .ZN(N217) );
  AOI31D0 U193 ( .A1(n171), .A2(n175), .A3(n176), .B(n170), .ZN(N216) );
  AOI21D0 U194 ( .A1(n177), .A2(n178), .B(n179), .ZN(n176) );
  CKND2D0 U195 ( .A1(n233), .A2(n286), .ZN(n178) );
  AOI31D0 U196 ( .A1(n180), .A2(State[0]), .A3(n181), .B(n170), .ZN(N214) );
  AOI22D0 U197 ( .A1(n182), .A2(n183), .B1(n184), .B2(n185), .ZN(n181) );
  CKND0 U198 ( .CLK(n179), .CN(n180) );
  OAI211D0 U199 ( .A1(n186), .A2(n187), .B(n168), .C(n173), .ZN(n179) );
  NR2D0 U200 ( .A1(Reset), .A2(n101), .ZN(n186) );
  CKND0 U201 ( .CLK(TRes3), .CN(n101) );
  NR2D0 U202 ( .A1(n188), .A2(n170), .ZN(N212) );
  OA222D0 U203 ( .A1(n189), .A2(N151), .B1(n175), .B2(N158), .C1(n168), .C2(
        N165), .Z(n188) );
  CKND2D0 U204 ( .A1(n174), .A2(n190), .ZN(N211) );
  OAI21D0 U205 ( .A1(n161), .A2(n191), .B(n4), .ZN(n190) );
  NR2D0 U206 ( .A1(n192), .A2(n170), .ZN(N210) );
  OA222D0 U207 ( .A1(n173), .A2(N138), .B1(n187), .B2(N145), .C1(n168), .C2(
        N165), .Z(n192) );
  AOI21D0 U208 ( .A1(n193), .A2(n194), .B(n170), .ZN(N208) );
  CKND0 U209 ( .CLK(n166), .CN(n170) );
  AOI22D0 U210 ( .A1(n195), .A2(TRes3), .B1(n182), .B2(n163), .ZN(n194) );
  AOI21D0 U211 ( .A1(n184), .A2(n164), .B(n196), .ZN(n193) );
  CKND0 U212 ( .CLK(n185), .CN(n164) );
  AO211D0 U213 ( .A1(n191), .A2(n4), .B(n165), .C(n162), .Z(N206) );
  NR3D0 U214 ( .A1(n197), .A2(n198), .A3(n199), .ZN(n162) );
  ND3D0 U215 ( .A1(n171), .A2(n173), .A3(n172), .ZN(n191) );
  NR3D0 U216 ( .A1(n184), .A2(n177), .A3(n195), .ZN(n172) );
  CKND0 U217 ( .CLK(n189), .CN(n177) );
  AO211D0 U218 ( .A1(N172), .A2(n166), .B(ParityErr), .C(n201), .Z(N205) );
  IND3D0 U219 ( .A1(N184), .B1(n200), .B2(n174), .ZN(N203) );
  NR2D0 U220 ( .A1(n201), .A2(N204), .ZN(n174) );
  NR2D0 U221 ( .A1(n198), .A2(Testing), .ZN(N204) );
  CKND0 U222 ( .CLK(n4), .CN(n198) );
  CKND0 U223 ( .CLK(DoSelfTest), .CN(n201) );
  OAI21D0 U224 ( .A1(ParityErr), .A2(AllDoner), .B(DoSelfTest), .ZN(n200) );
  AN2D0 U225 ( .A1(n196), .A2(Testing), .Z(N186) );
  OAI222D0 U226 ( .A1(TestDone[1]), .A2(n171), .B1(TestDone[3]), .B2(n187), 
        .C1(TestDone[5]), .C2(n175), .ZN(n196) );
  CKND0 U227 ( .CLK(n184), .CN(n175) );
  NR3D0 U228 ( .A1(n199), .A2(State[1]), .A3(n161), .ZN(n184) );
  CKND0 U229 ( .CLK(n195), .CN(n187) );
  NR3D0 U230 ( .A1(n197), .A2(State[2]), .A3(n161), .ZN(n195) );
  CKND0 U231 ( .CLK(n182), .CN(n171) );
  NR3D0 U232 ( .A1(State[1]), .A2(State[2]), .A3(n161), .ZN(n182) );
  CKND0 U233 ( .CLK(n202), .CN(TestDone[1]) );
  NR2D0 U234 ( .A1(n203), .A2(n27), .ZN(N185) );
  OA222D0 U235 ( .A1(n173), .A2(TestDone[2]), .B1(n168), .B2(TestDone[6]), 
        .C1(n189), .C2(TestDone[4]), .Z(n203) );
  ND3D0 U236 ( .A1(n161), .A2(n197), .A3(State[2]), .ZN(n189) );
  CKND0 U237 ( .CLK(State[1]), .CN(n197) );
  ND3D0 U238 ( .A1(State[1]), .A2(n161), .A3(State[2]), .ZN(n168) );
  ND3D0 U239 ( .A1(n161), .A2(n199), .A3(State[1]), .ZN(n173) );
  CKND0 U240 ( .CLK(State[2]), .CN(n199) );
  CKND0 U241 ( .CLK(State[0]), .CN(n161) );
  INR2D0 U242 ( .A1(TestDone[6]), .B1(n231), .ZN(N165) );
  NR2D0 U243 ( .A1(n11), .A2(Reset), .ZN(TestDone[6]) );
  AN2D0 U244 ( .A1(TestDone[5]), .A2(n185), .Z(N158) );
  CKND2D0 U245 ( .A1(TRes5), .A2(n286), .ZN(n185) );
  INR2D0 U246 ( .A1(TestDone[4]), .B1(n233), .ZN(N151) );
  NR2D0 U247 ( .A1(n12), .A2(Reset), .ZN(TestDone[4]) );
  INR2D0 U248 ( .A1(TestDone[3]), .B1(TRes3), .ZN(N145) );
  INR2D0 U249 ( .A1(TestDone[2]), .B1(n235), .ZN(N138) );
  NR2D0 U250 ( .A1(n13), .A2(Reset), .ZN(TestDone[2]) );
  NR2D0 U251 ( .A1(n163), .A2(n202), .ZN(N132) );
  CKND2D0 U252 ( .A1(TDone1), .A2(n286), .ZN(n202) );
  CKND0 U253 ( .CLK(n183), .CN(n163) );
  CKND2D0 U254 ( .A1(TRes1), .A2(n286), .ZN(n183) );
  IOA21D0 U255 ( .A1(DataO1[9]), .A2(N272), .B(n205), .ZN(DataO[9]) );
  IOA21D0 U256 ( .A1(DataO1[8]), .A2(N272), .B(n205), .ZN(DataO[8]) );
  IOA21D0 U257 ( .A1(DataO1[4]), .A2(N272), .B(n205), .ZN(DataO[4]) );
  IOA21D0 U258 ( .A1(DataO1[3]), .A2(N272), .B(n205), .ZN(DataO[3]) );
  IOA21D0 U259 ( .A1(DataO1[2]), .A2(N272), .B(n205), .ZN(DataO[2]) );
  IOA21D0 U260 ( .A1(DataO1[28]), .A2(N272), .B(n205), .ZN(DataO[28]) );
  IOA21D0 U261 ( .A1(DataO1[27]), .A2(N272), .B(n205), .ZN(DataO[27]) );
  IOA21D0 U262 ( .A1(DataO1[26]), .A2(N272), .B(n205), .ZN(DataO[26]) );
  IOA21D0 U263 ( .A1(DataO1[25]), .A2(N272), .B(n205), .ZN(DataO[25]) );
  IOA21D0 U264 ( .A1(DataO1[24]), .A2(N272), .B(n205), .ZN(DataO[24]) );
  IOA21D0 U265 ( .A1(DataO1[20]), .A2(N272), .B(n205), .ZN(DataO[20]) );
  IOA21D0 U266 ( .A1(DataO1[1]), .A2(N272), .B(n205), .ZN(DataO[1]) );
  IOA21D0 U267 ( .A1(DataO1[19]), .A2(N272), .B(n205), .ZN(DataO[19]) );
  IOA21D0 U268 ( .A1(DataO1[18]), .A2(N272), .B(n205), .ZN(DataO[18]) );
  IOA21D0 U269 ( .A1(DataO1[17]), .A2(N272), .B(n205), .ZN(DataO[17]) );
  IOA21D0 U270 ( .A1(DataO1[16]), .A2(N272), .B(n205), .ZN(DataO[16]) );
  IOA21D0 U271 ( .A1(DataO1[12]), .A2(N272), .B(n205), .ZN(DataO[12]) );
  IOA21D0 U272 ( .A1(DataO1[11]), .A2(N272), .B(n205), .ZN(DataO[11]) );
  IOA21D0 U273 ( .A1(DataO1[10]), .A2(N272), .B(n205), .ZN(DataO[10]) );
  IOA21D0 U274 ( .A1(DataO1[0]), .A2(N272), .B(n205), .ZN(DataO[0]) );
  OAI211D0 U275 ( .A1(n109), .A2(n6), .B(n207), .C(n209), .ZN(Addr[4]) );
  AOI222D0 U276 ( .A1(Addr3[4]), .A2(N364), .B1(Addr1[4]), .B2(N272), .C1(
        Addr5[4]), .C2(N449), .ZN(n209) );
  AOI22D0 U277 ( .A1(n236), .A2(n65), .B1(n238), .B2(n78), .ZN(n207) );
  OAI211D0 U278 ( .A1(n10), .A2(n109), .B(n211), .C(n213), .ZN(Addr[3]) );
  AOI222D0 U279 ( .A1(Addr3[3]), .A2(N364), .B1(Addr1[3]), .B2(N272), .C1(
        Addr5[3]), .C2(N449), .ZN(n213) );
  AOI22D0 U280 ( .A1(n65), .A2(n239), .B1(n78), .B2(n240), .ZN(n211) );
  OAI211D0 U281 ( .A1(n109), .A2(n7), .B(n214), .C(n215), .ZN(Addr[2]) );
  AOI222D0 U282 ( .A1(Addr3[2]), .A2(N364), .B1(Addr1[2]), .B2(N272), .C1(
        Addr5[2]), .C2(N449), .ZN(n215) );
  AOI22D0 U283 ( .A1(n287), .A2(n65), .B1(n288), .B2(n78), .ZN(n214) );
  OAI211D0 U284 ( .A1(n109), .A2(n8), .B(n217), .C(n219), .ZN(Addr[1]) );
  AOI222D0 U285 ( .A1(Addr3[1]), .A2(N364), .B1(Addr1[1]), .B2(N272), .C1(
        Addr5[1]), .C2(N449), .ZN(n219) );
  AOI22D0 U286 ( .A1(n289), .A2(n65), .B1(n290), .B2(n78), .ZN(n217) );
  OAI211D0 U287 ( .A1(n109), .A2(n9), .B(n221), .C(n223), .ZN(Addr[0]) );
  AOI222D0 U288 ( .A1(Addr3[0]), .A2(N364), .B1(Addr1[0]), .B2(N272), .C1(
        Addr5[0]), .C2(N449), .ZN(n223) );
  AN3D0 U289 ( .A1(TestNo[0]), .A2(TestNo[2]), .A3(n5), .Z(N411) );
  AN3D0 U290 ( .A1(TestNo[0]), .A2(n225), .A3(n5), .Z(N233) );
  CKND0 U291 ( .CLK(n205), .CN(N364) );
  AN3D0 U292 ( .A1(TestNo[0]), .A2(n293), .A3(n225), .Z(N326) );
  AOI22D0 U293 ( .A1(n291), .A2(n65), .B1(n292), .B2(n78), .ZN(n221) );
  CKND0 U294 ( .CLK(n75), .CN(n86) );
  NR3D0 U295 ( .A1(TestNo[0]), .A2(n293), .A3(n225), .ZN(n75) );
  CKND0 U296 ( .CLK(n70), .CN(n74) );
  NR3D0 U297 ( .A1(TestNo[0]), .A2(TestNo[2]), .A3(n5), .ZN(n70) );
  CKND2D0 U298 ( .A1(n106), .A2(n286), .ZN(n109) );
  NR3D0 U299 ( .A1(n225), .A2(TestNo[0]), .A3(n5), .ZN(n106) );
  CKND0 U300 ( .CLK(TestNo[2]), .CN(n225) );
endmodule


module Mem_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, ClkR, 
        ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, n572, ClockR, ClockW, Dreadyr,
         \Storage[31][32] , \Storage[31][31] , \Storage[31][30] ,
         \Storage[31][29] , \Storage[31][28] , \Storage[31][27] ,
         \Storage[31][26] , \Storage[31][25] , \Storage[31][24] ,
         \Storage[31][23] , \Storage[31][22] , \Storage[31][21] ,
         \Storage[31][20] , \Storage[31][19] , \Storage[31][18] ,
         \Storage[31][17] , \Storage[31][16] , \Storage[31][15] ,
         \Storage[31][14] , \Storage[31][13] , \Storage[31][12] ,
         \Storage[31][11] , \Storage[31][10] , \Storage[31][9] ,
         \Storage[31][8] , \Storage[31][7] , \Storage[31][6] ,
         \Storage[31][5] , \Storage[31][4] , \Storage[31][3] ,
         \Storage[31][2] , \Storage[31][1] , \Storage[31][0] ,
         \Storage[30][32] , \Storage[30][31] , \Storage[30][30] ,
         \Storage[30][29] , \Storage[30][28] , \Storage[30][27] ,
         \Storage[30][26] , \Storage[30][25] , \Storage[30][24] ,
         \Storage[30][23] , \Storage[30][22] , \Storage[30][21] ,
         \Storage[30][20] , \Storage[30][19] , \Storage[30][18] ,
         \Storage[30][17] , \Storage[30][16] , \Storage[30][15] ,
         \Storage[30][14] , \Storage[30][13] , \Storage[30][12] ,
         \Storage[30][11] , \Storage[30][10] , \Storage[30][9] ,
         \Storage[30][8] , \Storage[30][7] , \Storage[30][6] ,
         \Storage[30][5] , \Storage[30][4] , \Storage[30][3] ,
         \Storage[30][2] , \Storage[30][1] , \Storage[30][0] ,
         \Storage[29][32] , \Storage[29][31] , \Storage[29][30] ,
         \Storage[29][29] , \Storage[29][28] , \Storage[29][27] ,
         \Storage[29][26] , \Storage[29][25] , \Storage[29][24] ,
         \Storage[29][23] , \Storage[29][22] , \Storage[29][21] ,
         \Storage[29][20] , \Storage[29][19] , \Storage[29][18] ,
         \Storage[29][17] , \Storage[29][16] , \Storage[29][15] ,
         \Storage[29][14] , \Storage[29][13] , \Storage[29][12] ,
         \Storage[29][11] , \Storage[29][10] , \Storage[29][9] ,
         \Storage[29][8] , \Storage[29][7] , \Storage[29][6] ,
         \Storage[29][5] , \Storage[29][4] , \Storage[29][3] ,
         \Storage[29][2] , \Storage[29][1] , \Storage[29][0] ,
         \Storage[28][32] , \Storage[28][31] , \Storage[28][30] ,
         \Storage[28][29] , \Storage[28][28] , \Storage[28][27] ,
         \Storage[28][26] , \Storage[28][25] , \Storage[28][24] ,
         \Storage[28][23] , \Storage[28][22] , \Storage[28][21] ,
         \Storage[28][20] , \Storage[28][19] , \Storage[28][18] ,
         \Storage[28][17] , \Storage[28][16] , \Storage[28][15] ,
         \Storage[28][14] , \Storage[28][13] , \Storage[28][12] ,
         \Storage[28][11] , \Storage[28][10] , \Storage[28][9] ,
         \Storage[28][8] , \Storage[28][7] , \Storage[28][6] ,
         \Storage[28][5] , \Storage[28][4] , \Storage[28][3] ,
         \Storage[28][2] , \Storage[28][1] , \Storage[28][0] ,
         \Storage[27][32] , \Storage[27][31] , \Storage[27][30] ,
         \Storage[27][29] , \Storage[27][28] , \Storage[27][27] ,
         \Storage[27][26] , \Storage[27][25] , \Storage[27][24] ,
         \Storage[27][23] , \Storage[27][22] , \Storage[27][21] ,
         \Storage[27][20] , \Storage[27][19] , \Storage[27][18] ,
         \Storage[27][17] , \Storage[27][16] , \Storage[27][15] ,
         \Storage[27][14] , \Storage[27][13] , \Storage[27][12] ,
         \Storage[27][11] , \Storage[27][10] , \Storage[27][9] ,
         \Storage[27][8] , \Storage[27][7] , \Storage[27][6] ,
         \Storage[27][5] , \Storage[27][4] , \Storage[27][3] ,
         \Storage[27][2] , \Storage[27][1] , \Storage[27][0] ,
         \Storage[26][32] , \Storage[26][31] , \Storage[26][30] ,
         \Storage[26][29] , \Storage[26][28] , \Storage[26][27] ,
         \Storage[26][26] , \Storage[26][25] , \Storage[26][24] ,
         \Storage[26][23] , \Storage[26][22] , \Storage[26][21] ,
         \Storage[26][20] , \Storage[26][19] , \Storage[26][18] ,
         \Storage[26][17] , \Storage[26][16] , \Storage[26][15] ,
         \Storage[26][14] , \Storage[26][13] , \Storage[26][12] ,
         \Storage[26][11] , \Storage[26][10] , \Storage[26][9] ,
         \Storage[26][8] , \Storage[26][7] , \Storage[26][6] ,
         \Storage[26][5] , \Storage[26][4] , \Storage[26][3] ,
         \Storage[26][2] , \Storage[26][1] , \Storage[26][0] ,
         \Storage[25][32] , \Storage[25][31] , \Storage[25][30] ,
         \Storage[25][29] , \Storage[25][28] , \Storage[25][27] ,
         \Storage[25][26] , \Storage[25][25] , \Storage[25][24] ,
         \Storage[25][23] , \Storage[25][22] , \Storage[25][21] ,
         \Storage[25][20] , \Storage[25][19] , \Storage[25][18] ,
         \Storage[25][17] , \Storage[25][16] , \Storage[25][15] ,
         \Storage[25][14] , \Storage[25][13] , \Storage[25][12] ,
         \Storage[25][11] , \Storage[25][10] , \Storage[25][9] ,
         \Storage[25][8] , \Storage[25][7] , \Storage[25][6] ,
         \Storage[25][5] , \Storage[25][4] , \Storage[25][3] ,
         \Storage[25][2] , \Storage[25][1] , \Storage[25][0] ,
         \Storage[24][32] , \Storage[24][31] , \Storage[24][30] ,
         \Storage[24][29] , \Storage[24][28] , \Storage[24][27] ,
         \Storage[24][26] , \Storage[24][25] , \Storage[24][24] ,
         \Storage[24][23] , \Storage[24][22] , \Storage[24][21] ,
         \Storage[24][20] , \Storage[24][19] , \Storage[24][18] ,
         \Storage[24][17] , \Storage[24][16] , \Storage[24][15] ,
         \Storage[24][14] , \Storage[24][13] , \Storage[24][12] ,
         \Storage[24][11] , \Storage[24][10] , \Storage[24][9] ,
         \Storage[24][8] , \Storage[24][7] , \Storage[24][6] ,
         \Storage[24][5] , \Storage[24][4] , \Storage[24][3] ,
         \Storage[24][2] , \Storage[24][1] , \Storage[24][0] ,
         \Storage[23][32] , \Storage[23][31] , \Storage[23][30] ,
         \Storage[23][29] , \Storage[23][28] , \Storage[23][27] ,
         \Storage[23][26] , \Storage[23][25] , \Storage[23][24] ,
         \Storage[23][23] , \Storage[23][22] , \Storage[23][21] ,
         \Storage[23][20] , \Storage[23][19] , \Storage[23][18] ,
         \Storage[23][17] , \Storage[23][16] , \Storage[23][15] ,
         \Storage[23][14] , \Storage[23][13] , \Storage[23][12] ,
         \Storage[23][11] , \Storage[23][10] , \Storage[23][9] ,
         \Storage[23][8] , \Storage[23][7] , \Storage[23][6] ,
         \Storage[23][5] , \Storage[23][4] , \Storage[23][3] ,
         \Storage[23][2] , \Storage[23][1] , \Storage[23][0] ,
         \Storage[22][32] , \Storage[22][31] , \Storage[22][30] ,
         \Storage[22][29] , \Storage[22][28] , \Storage[22][27] ,
         \Storage[22][26] , \Storage[22][25] , \Storage[22][24] ,
         \Storage[22][23] , \Storage[22][22] , \Storage[22][21] ,
         \Storage[22][20] , \Storage[22][19] , \Storage[22][18] ,
         \Storage[22][17] , \Storage[22][16] , \Storage[22][15] ,
         \Storage[22][14] , \Storage[22][13] , \Storage[22][12] ,
         \Storage[22][11] , \Storage[22][10] , \Storage[22][9] ,
         \Storage[22][8] , \Storage[22][7] , \Storage[22][6] ,
         \Storage[22][5] , \Storage[22][4] , \Storage[22][3] ,
         \Storage[22][2] , \Storage[22][1] , \Storage[22][0] ,
         \Storage[21][32] , \Storage[21][31] , \Storage[21][30] ,
         \Storage[21][29] , \Storage[21][28] , \Storage[21][27] ,
         \Storage[21][26] , \Storage[21][25] , \Storage[21][24] ,
         \Storage[21][23] , \Storage[21][22] , \Storage[21][21] ,
         \Storage[21][20] , \Storage[21][19] , \Storage[21][18] ,
         \Storage[21][17] , \Storage[21][16] , \Storage[21][15] ,
         \Storage[21][14] , \Storage[21][13] , \Storage[21][12] ,
         \Storage[21][11] , \Storage[21][10] , \Storage[21][9] ,
         \Storage[21][8] , \Storage[21][7] , \Storage[21][6] ,
         \Storage[21][5] , \Storage[21][4] , \Storage[21][3] ,
         \Storage[21][2] , \Storage[21][1] , \Storage[21][0] ,
         \Storage[20][32] , \Storage[20][31] , \Storage[20][30] ,
         \Storage[20][29] , \Storage[20][28] , \Storage[20][27] ,
         \Storage[20][26] , \Storage[20][25] , \Storage[20][24] ,
         \Storage[20][23] , \Storage[20][22] , \Storage[20][21] ,
         \Storage[20][20] , \Storage[20][19] , \Storage[20][18] ,
         \Storage[20][17] , \Storage[20][16] , \Storage[20][15] ,
         \Storage[20][14] , \Storage[20][13] , \Storage[20][12] ,
         \Storage[20][11] , \Storage[20][10] , \Storage[20][9] ,
         \Storage[20][8] , \Storage[20][7] , \Storage[20][6] ,
         \Storage[20][5] , \Storage[20][4] , \Storage[20][3] ,
         \Storage[20][2] , \Storage[20][1] , \Storage[20][0] ,
         \Storage[19][32] , \Storage[19][31] , \Storage[19][30] ,
         \Storage[19][29] , \Storage[19][28] , \Storage[19][27] ,
         \Storage[19][26] , \Storage[19][25] , \Storage[19][24] ,
         \Storage[19][23] , \Storage[19][22] , \Storage[19][21] ,
         \Storage[19][20] , \Storage[19][19] , \Storage[19][18] ,
         \Storage[19][17] , \Storage[19][16] , \Storage[19][15] ,
         \Storage[19][14] , \Storage[19][13] , \Storage[19][12] ,
         \Storage[19][11] , \Storage[19][10] , \Storage[19][9] ,
         \Storage[19][8] , \Storage[19][7] , \Storage[19][6] ,
         \Storage[19][5] , \Storage[19][4] , \Storage[19][3] ,
         \Storage[19][2] , \Storage[19][1] , \Storage[19][0] ,
         \Storage[18][32] , \Storage[18][31] , \Storage[18][30] ,
         \Storage[18][29] , \Storage[18][28] , \Storage[18][27] ,
         \Storage[18][26] , \Storage[18][25] , \Storage[18][24] ,
         \Storage[18][23] , \Storage[18][22] , \Storage[18][21] ,
         \Storage[18][20] , \Storage[18][19] , \Storage[18][18] ,
         \Storage[18][17] , \Storage[18][16] , \Storage[18][15] ,
         \Storage[18][14] , \Storage[18][13] , \Storage[18][12] ,
         \Storage[18][11] , \Storage[18][10] , \Storage[18][9] ,
         \Storage[18][8] , \Storage[18][7] , \Storage[18][6] ,
         \Storage[18][5] , \Storage[18][4] , \Storage[18][3] ,
         \Storage[18][2] , \Storage[18][1] , \Storage[18][0] ,
         \Storage[17][32] , \Storage[17][31] , \Storage[17][30] ,
         \Storage[17][29] , \Storage[17][28] , \Storage[17][27] ,
         \Storage[17][26] , \Storage[17][25] , \Storage[17][24] ,
         \Storage[17][23] , \Storage[17][22] , \Storage[17][21] ,
         \Storage[17][20] , \Storage[17][19] , \Storage[17][18] ,
         \Storage[17][17] , \Storage[17][16] , \Storage[17][15] ,
         \Storage[17][14] , \Storage[17][13] , \Storage[17][12] ,
         \Storage[17][11] , \Storage[17][10] , \Storage[17][9] ,
         \Storage[17][8] , \Storage[17][7] , \Storage[17][6] ,
         \Storage[17][5] , \Storage[17][4] , \Storage[17][3] ,
         \Storage[17][2] , \Storage[17][1] , \Storage[17][0] ,
         \Storage[16][32] , \Storage[16][31] , \Storage[16][30] ,
         \Storage[16][29] , \Storage[16][28] , \Storage[16][27] ,
         \Storage[16][26] , \Storage[16][25] , \Storage[16][24] ,
         \Storage[16][23] , \Storage[16][22] , \Storage[16][21] ,
         \Storage[16][20] , \Storage[16][19] , \Storage[16][18] ,
         \Storage[16][17] , \Storage[16][16] , \Storage[16][15] ,
         \Storage[16][14] , \Storage[16][13] , \Storage[16][12] ,
         \Storage[16][11] , \Storage[16][10] , \Storage[16][9] ,
         \Storage[16][8] , \Storage[16][7] , \Storage[16][6] ,
         \Storage[16][5] , \Storage[16][4] , \Storage[16][3] ,
         \Storage[16][2] , \Storage[16][1] , \Storage[16][0] ,
         \Storage[15][32] , \Storage[15][31] , \Storage[15][30] ,
         \Storage[15][29] , \Storage[15][28] , \Storage[15][27] ,
         \Storage[15][26] , \Storage[15][25] , \Storage[15][24] ,
         \Storage[15][23] , \Storage[15][22] , \Storage[15][21] ,
         \Storage[15][20] , \Storage[15][19] , \Storage[15][18] ,
         \Storage[15][17] , \Storage[15][16] , \Storage[15][15] ,
         \Storage[15][14] , \Storage[15][13] , \Storage[15][12] ,
         \Storage[15][11] , \Storage[15][10] , \Storage[15][9] ,
         \Storage[15][8] , \Storage[15][7] , \Storage[15][6] ,
         \Storage[15][5] , \Storage[15][4] , \Storage[15][3] ,
         \Storage[15][2] , \Storage[15][1] , \Storage[15][0] ,
         \Storage[14][32] , \Storage[14][31] , \Storage[14][30] ,
         \Storage[14][29] , \Storage[14][28] , \Storage[14][27] ,
         \Storage[14][26] , \Storage[14][25] , \Storage[14][24] ,
         \Storage[14][23] , \Storage[14][22] , \Storage[14][21] ,
         \Storage[14][20] , \Storage[14][19] , \Storage[14][18] ,
         \Storage[14][17] , \Storage[14][16] , \Storage[14][15] ,
         \Storage[14][14] , \Storage[14][13] , \Storage[14][12] ,
         \Storage[14][11] , \Storage[14][10] , \Storage[14][9] ,
         \Storage[14][8] , \Storage[14][7] , \Storage[14][6] ,
         \Storage[14][5] , \Storage[14][4] , \Storage[14][3] ,
         \Storage[14][2] , \Storage[14][1] , \Storage[14][0] ,
         \Storage[13][32] , \Storage[13][31] , \Storage[13][30] ,
         \Storage[13][29] , \Storage[13][28] , \Storage[13][27] ,
         \Storage[13][26] , \Storage[13][25] , \Storage[13][24] ,
         \Storage[13][23] , \Storage[13][22] , \Storage[13][21] ,
         \Storage[13][20] , \Storage[13][19] , \Storage[13][18] ,
         \Storage[13][17] , \Storage[13][16] , \Storage[13][15] ,
         \Storage[13][14] , \Storage[13][13] , \Storage[13][12] ,
         \Storage[13][11] , \Storage[13][10] , \Storage[13][9] ,
         \Storage[13][8] , \Storage[13][7] , \Storage[13][6] ,
         \Storage[13][5] , \Storage[13][4] , \Storage[13][3] ,
         \Storage[13][2] , \Storage[13][1] , \Storage[13][0] ,
         \Storage[12][32] , \Storage[12][31] , \Storage[12][30] ,
         \Storage[12][29] , \Storage[12][28] , \Storage[12][27] ,
         \Storage[12][26] , \Storage[12][25] , \Storage[12][24] ,
         \Storage[12][23] , \Storage[12][22] , \Storage[12][21] ,
         \Storage[12][20] , \Storage[12][19] , \Storage[12][18] ,
         \Storage[12][17] , \Storage[12][16] , \Storage[12][15] ,
         \Storage[12][14] , \Storage[12][13] , \Storage[12][12] ,
         \Storage[12][11] , \Storage[12][10] , \Storage[12][9] ,
         \Storage[12][8] , \Storage[12][7] , \Storage[12][6] ,
         \Storage[12][5] , \Storage[12][4] , \Storage[12][3] ,
         \Storage[12][2] , \Storage[12][1] , \Storage[12][0] ,
         \Storage[11][32] , \Storage[11][31] , \Storage[11][30] ,
         \Storage[11][29] , \Storage[11][28] , \Storage[11][27] ,
         \Storage[11][26] , \Storage[11][25] , \Storage[11][24] ,
         \Storage[11][23] , \Storage[11][22] , \Storage[11][21] ,
         \Storage[11][20] , \Storage[11][19] , \Storage[11][18] ,
         \Storage[11][17] , \Storage[11][16] , \Storage[11][15] ,
         \Storage[11][14] , \Storage[11][13] , \Storage[11][12] ,
         \Storage[11][11] , \Storage[11][10] , \Storage[11][9] ,
         \Storage[11][8] , \Storage[11][7] , \Storage[11][6] ,
         \Storage[11][5] , \Storage[11][4] , \Storage[11][3] ,
         \Storage[11][2] , \Storage[11][1] , \Storage[11][0] ,
         \Storage[10][32] , \Storage[10][31] , \Storage[10][30] ,
         \Storage[10][29] , \Storage[10][28] , \Storage[10][27] ,
         \Storage[10][26] , \Storage[10][25] , \Storage[10][24] ,
         \Storage[10][23] , \Storage[10][22] , \Storage[10][21] ,
         \Storage[10][20] , \Storage[10][19] , \Storage[10][18] ,
         \Storage[10][17] , \Storage[10][16] , \Storage[10][15] ,
         \Storage[10][14] , \Storage[10][13] , \Storage[10][12] ,
         \Storage[10][11] , \Storage[10][10] , \Storage[10][9] ,
         \Storage[10][8] , \Storage[10][7] , \Storage[10][6] ,
         \Storage[10][5] , \Storage[10][4] , \Storage[10][3] ,
         \Storage[10][2] , \Storage[10][1] , \Storage[10][0] ,
         \Storage[9][32] , \Storage[9][31] , \Storage[9][30] ,
         \Storage[9][29] , \Storage[9][28] , \Storage[9][27] ,
         \Storage[9][26] , \Storage[9][25] , \Storage[9][24] ,
         \Storage[9][23] , \Storage[9][22] , \Storage[9][21] ,
         \Storage[9][20] , \Storage[9][19] , \Storage[9][18] ,
         \Storage[9][17] , \Storage[9][16] , \Storage[9][15] ,
         \Storage[9][14] , \Storage[9][13] , \Storage[9][12] ,
         \Storage[9][11] , \Storage[9][10] , \Storage[9][9] , \Storage[9][8] ,
         \Storage[9][7] , \Storage[9][6] , \Storage[9][5] , \Storage[9][4] ,
         \Storage[9][3] , \Storage[9][2] , \Storage[9][1] , \Storage[9][0] ,
         \Storage[8][32] , \Storage[8][31] , \Storage[8][30] ,
         \Storage[8][29] , \Storage[8][28] , \Storage[8][27] ,
         \Storage[8][26] , \Storage[8][25] , \Storage[8][24] ,
         \Storage[8][23] , \Storage[8][22] , \Storage[8][21] ,
         \Storage[8][20] , \Storage[8][19] , \Storage[8][18] ,
         \Storage[8][17] , \Storage[8][16] , \Storage[8][15] ,
         \Storage[8][14] , \Storage[8][13] , \Storage[8][12] ,
         \Storage[8][11] , \Storage[8][10] , \Storage[8][9] , \Storage[8][8] ,
         \Storage[8][7] , \Storage[8][6] , \Storage[8][5] , \Storage[8][4] ,
         \Storage[8][3] , \Storage[8][2] , \Storage[8][1] , \Storage[8][0] ,
         \Storage[7][32] , \Storage[7][31] , \Storage[7][30] ,
         \Storage[7][29] , \Storage[7][28] , \Storage[7][27] ,
         \Storage[7][26] , \Storage[7][25] , \Storage[7][24] ,
         \Storage[7][23] , \Storage[7][22] , \Storage[7][21] ,
         \Storage[7][20] , \Storage[7][19] , \Storage[7][18] ,
         \Storage[7][17] , \Storage[7][16] , \Storage[7][15] ,
         \Storage[7][14] , \Storage[7][13] , \Storage[7][12] ,
         \Storage[7][11] , \Storage[7][10] , \Storage[7][9] , \Storage[7][8] ,
         \Storage[7][7] , \Storage[7][6] , \Storage[7][5] , \Storage[7][4] ,
         \Storage[7][3] , \Storage[7][2] , \Storage[7][1] , \Storage[7][0] ,
         \Storage[6][32] , \Storage[6][31] , \Storage[6][30] ,
         \Storage[6][29] , \Storage[6][28] , \Storage[6][27] ,
         \Storage[6][26] , \Storage[6][25] , \Storage[6][24] ,
         \Storage[6][23] , \Storage[6][22] , \Storage[6][21] ,
         \Storage[6][20] , \Storage[6][19] , \Storage[6][18] ,
         \Storage[6][17] , \Storage[6][16] , \Storage[6][15] ,
         \Storage[6][14] , \Storage[6][13] , \Storage[6][12] ,
         \Storage[6][11] , \Storage[6][10] , \Storage[6][9] , \Storage[6][8] ,
         \Storage[6][7] , \Storage[6][6] , \Storage[6][5] , \Storage[6][4] ,
         \Storage[6][3] , \Storage[6][2] , \Storage[6][1] , \Storage[6][0] ,
         \Storage[5][32] , \Storage[5][31] , \Storage[5][30] ,
         \Storage[5][29] , \Storage[5][28] , \Storage[5][27] ,
         \Storage[5][26] , \Storage[5][25] , \Storage[5][24] ,
         \Storage[5][23] , \Storage[5][22] , \Storage[5][21] ,
         \Storage[5][20] , \Storage[5][19] , \Storage[5][18] ,
         \Storage[5][17] , \Storage[5][16] , \Storage[5][15] ,
         \Storage[5][14] , \Storage[5][13] , \Storage[5][12] ,
         \Storage[5][11] , \Storage[5][10] , \Storage[5][9] , \Storage[5][8] ,
         \Storage[5][7] , \Storage[5][6] , \Storage[5][5] , \Storage[5][4] ,
         \Storage[5][3] , \Storage[5][2] , \Storage[5][1] , \Storage[5][0] ,
         \Storage[4][32] , \Storage[4][31] , \Storage[4][30] ,
         \Storage[4][29] , \Storage[4][28] , \Storage[4][27] ,
         \Storage[4][26] , \Storage[4][25] , \Storage[4][24] ,
         \Storage[4][23] , \Storage[4][22] , \Storage[4][21] ,
         \Storage[4][20] , \Storage[4][19] , \Storage[4][18] ,
         \Storage[4][17] , \Storage[4][16] , \Storage[4][15] ,
         \Storage[4][14] , \Storage[4][13] , \Storage[4][12] ,
         \Storage[4][11] , \Storage[4][10] , \Storage[4][9] , \Storage[4][8] ,
         \Storage[4][7] , \Storage[4][6] , \Storage[4][5] , \Storage[4][4] ,
         \Storage[4][3] , \Storage[4][2] , \Storage[4][1] , \Storage[4][0] ,
         \Storage[3][32] , \Storage[3][31] , \Storage[3][30] ,
         \Storage[3][29] , \Storage[3][28] , \Storage[3][27] ,
         \Storage[3][26] , \Storage[3][25] , \Storage[3][24] ,
         \Storage[3][23] , \Storage[3][22] , \Storage[3][21] ,
         \Storage[3][20] , \Storage[3][19] , \Storage[3][18] ,
         \Storage[3][17] , \Storage[3][16] , \Storage[3][15] ,
         \Storage[3][14] , \Storage[3][13] , \Storage[3][12] ,
         \Storage[3][11] , \Storage[3][10] , \Storage[3][9] , \Storage[3][8] ,
         \Storage[3][7] , \Storage[3][6] , \Storage[3][5] , \Storage[3][4] ,
         \Storage[3][3] , \Storage[3][2] , \Storage[3][1] , \Storage[3][0] ,
         \Storage[2][32] , \Storage[2][31] , \Storage[2][30] ,
         \Storage[2][29] , \Storage[2][28] , \Storage[2][27] ,
         \Storage[2][26] , \Storage[2][25] , \Storage[2][24] ,
         \Storage[2][23] , \Storage[2][22] , \Storage[2][21] ,
         \Storage[2][20] , \Storage[2][19] , \Storage[2][18] ,
         \Storage[2][17] , \Storage[2][16] , \Storage[2][15] ,
         \Storage[2][14] , \Storage[2][13] , \Storage[2][12] ,
         \Storage[2][11] , \Storage[2][10] , \Storage[2][9] , \Storage[2][8] ,
         \Storage[2][7] , \Storage[2][6] , \Storage[2][5] , \Storage[2][4] ,
         \Storage[2][3] , \Storage[2][2] , \Storage[2][1] , \Storage[2][0] ,
         \Storage[1][32] , \Storage[1][31] , \Storage[1][30] ,
         \Storage[1][29] , \Storage[1][28] , \Storage[1][27] ,
         \Storage[1][26] , \Storage[1][25] , \Storage[1][24] ,
         \Storage[1][23] , \Storage[1][22] , \Storage[1][21] ,
         \Storage[1][20] , \Storage[1][19] , \Storage[1][18] ,
         \Storage[1][17] , \Storage[1][16] , \Storage[1][15] ,
         \Storage[1][14] , \Storage[1][13] , \Storage[1][12] ,
         \Storage[1][11] , \Storage[1][10] , \Storage[1][9] , \Storage[1][8] ,
         \Storage[1][7] , \Storage[1][6] , \Storage[1][5] , \Storage[1][4] ,
         \Storage[1][3] , \Storage[1][2] , \Storage[1][1] , \Storage[1][0] ,
         \Storage[0][32] , \Storage[0][31] , \Storage[0][30] ,
         \Storage[0][29] , \Storage[0][28] , \Storage[0][27] ,
         \Storage[0][26] , \Storage[0][25] , \Storage[0][24] ,
         \Storage[0][23] , \Storage[0][22] , \Storage[0][21] ,
         \Storage[0][20] , \Storage[0][19] , \Storage[0][18] ,
         \Storage[0][17] , \Storage[0][16] , \Storage[0][15] ,
         \Storage[0][14] , \Storage[0][13] , \Storage[0][12] ,
         \Storage[0][11] , \Storage[0][10] , \Storage[0][9] , \Storage[0][8] ,
         \Storage[0][7] , \Storage[0][6] , \Storage[0][5] , \Storage[0][4] ,
         \Storage[0][3] , \Storage[0][2] , \Storage[0][1] , \Storage[0][0] ,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N85, N150, N183, N216, N249, N282, N315,
         N348, N381, N414, N447, N480, N513, N546, N579, N612, N645, N678,
         N711, N744, N777, N810, N843, N876, N909, N942, N975, N999, N1041,
         N1074, N1107, N1140, N1173, n107, n108, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  BUFTD1 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD1 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD1 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD1 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD1 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD1 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD1 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD1 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD1 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD1 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD1 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD1 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD1 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD1 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD1 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD1 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD1 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD1 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD1 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD1 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD1 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD1 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD1 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD1 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD1 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD1 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD1 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD1 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD1 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD1 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD1 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD1 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(N85), .E(N999), .CP(n61), .CDN(n8), .Q(
        \Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(DataI[31]), .E(N999), .CP(n66), .CDN(n8), 
        .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(DataI[30]), .E(N999), .CP(n67), .CDN(n8), 
        .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(DataI[29]), .E(N999), .CP(n69), .CDN(n8), 
        .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(DataI[28]), .E(N999), .CP(n63), .CDN(n8), 
        .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(DataI[27]), .E(N999), .CP(n60), .CDN(n8), 
        .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(DataI[26]), .E(N999), .CP(n62), .CDN(n8), 
        .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(DataI[25]), .E(N999), .CP(n61), .CDN(n8), 
        .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(DataI[24]), .E(N999), .CP(n67), .CDN(n7), 
        .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(DataI[23]), .E(N999), .CP(n66), .CDN(n7), 
        .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(DataI[22]), .E(N999), .CP(n65), .CDN(n7), 
        .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(DataI[21]), .E(N999), .CP(n59), .CDN(n7), 
        .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(DataI[20]), .E(N999), .CP(n45), .CDN(n7), 
        .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(DataI[19]), .E(N999), .CP(n50), .CDN(n7), 
        .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(DataI[18]), .E(N999), .CP(n70), .CDN(n7), 
        .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(DataI[17]), .E(N999), .CP(n62), .CDN(n7), 
        .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(DataI[16]), .E(N999), .CP(n55), .CDN(n7), 
        .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(DataI[15]), .E(N999), .CP(n68), .CDN(n7), 
        .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(DataI[14]), .E(N999), .CP(n61), .CDN(n7), 
        .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(DataI[13]), .E(N999), .CP(n65), .CDN(n6), 
        .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(DataI[12]), .E(N999), .CP(n64), .CDN(n6), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(DataI[11]), .E(N999), .CP(n61), .CDN(n6), 
        .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(DataI[10]), .E(N999), .CP(n59), .CDN(n6), 
        .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(DataI[9]), .E(N999), .CP(n44), .CDN(n6), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(DataI[8]), .E(N999), .CP(n46), .CDN(n6), 
        .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(DataI[7]), .E(N999), .CP(n52), .CDN(n6), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(DataI[6]), .E(N999), .CP(n53), .CDN(n6), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(DataI[5]), .E(N999), .CP(n41), .CDN(n6), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(DataI[4]), .E(N999), .CP(n69), .CDN(n6), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(DataI[3]), .E(N999), .CP(n63), .CDN(n6), 
        .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(DataI[2]), .E(N999), .CP(n68), .CDN(n5), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(DataI[1]), .E(N999), .CP(n66), .CDN(n5), 
        .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(DataI[0]), .E(N999), .CP(n69), .CDN(n5), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(N85), .E(N942), .CP(n45), .CDN(n34), .Q(
        \Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(DataI[31]), .E(N942), .CP(n45), .CDN(n31), .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(DataI[30]), .E(N942), .CP(n45), .CDN(n3), 
        .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(DataI[29]), .E(N942), .CP(n45), .CDN(n39), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(DataI[28]), .E(N942), .CP(n45), .CDN(n29), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(DataI[27]), .E(N942), .CP(n45), .CDN(n33), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(DataI[26]), .E(N942), .CP(n45), .CDN(n35), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(DataI[25]), .E(N942), .CP(n45), .CDN(n37), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(DataI[24]), .E(N942), .CP(n45), .CDN(n20), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(DataI[23]), .E(N942), .CP(n44), .CDN(n5), 
        .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(DataI[22]), .E(N942), .CP(n44), .CDN(n4), 
        .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(DataI[21]), .E(N942), .CP(n44), .CDN(n11), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(DataI[20]), .E(N942), .CP(n44), .CDN(n9), 
        .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(DataI[19]), .E(N942), .CP(n44), .CDN(n10), .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(DataI[18]), .E(N942), .CP(n44), .CDN(n7), 
        .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(DataI[17]), .E(N942), .CP(n44), .CDN(n8), 
        .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(DataI[16]), .E(N942), .CP(n44), .CDN(n31), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(DataI[15]), .E(N942), .CP(n44), .CDN(n3), 
        .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(DataI[14]), .E(N942), .CP(n44), .CDN(n29), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(DataI[13]), .E(N942), .CP(n43), .CDN(n30), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(DataI[12]), .E(N942), .CP(n43), .CDN(n36), .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(DataI[11]), .E(N942), .CP(n43), .CDN(n12), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(DataI[10]), .E(N942), .CP(n43), .CDN(n13), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(DataI[9]), .E(N942), .CP(n43), .CDN(n21), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(DataI[8]), .E(N942), .CP(n43), .CDN(n24), 
        .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(DataI[7]), .E(N942), .CP(n43), .CDN(n23), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(DataI[6]), .E(N942), .CP(n43), .CDN(n22), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(DataI[5]), .E(N942), .CP(n43), .CDN(n5), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(DataI[4]), .E(N942), .CP(n43), .CDN(n4), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(DataI[3]), .E(N942), .CP(n42), .CDN(n11), 
        .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(DataI[2]), .E(N942), .CP(n42), .CDN(n28), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(DataI[1]), .E(N942), .CP(n42), .CDN(n27), 
        .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(DataI[0]), .E(N942), .CP(n42), .CDN(n26), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(N85), .E(N1140), .CP(n52), .CDN(n27), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(N1140), .CP(n52), .CDN(
        n24), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(N1140), .CP(n52), .CDN(
        n38), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(N1140), .CP(n52), .CDN(
        n22), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(N1140), .CP(n52), .CDN(
        n34), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(N1140), .CP(n51), .CDN(
        n21), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(N1140), .CP(n51), .CDN(n6), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(N1140), .CP(n51), .CDN(
        n33), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(N1140), .CP(n51), .CDN(
        n40), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(N1140), .CP(n51), .CDN(
        n24), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(N1140), .CP(n51), .CDN(
        n14), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(N1140), .CP(n51), .CDN(
        n34), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(N1140), .CP(n51), .CDN(n4), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(N1140), .CP(n51), .CDN(
        n25), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(N1140), .CP(n51), .CDN(
        n21), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(N1140), .CP(n50), .CDN(
        n31), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(N1140), .CP(n50), .CDN(
        n31), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(N1140), .CP(n50), .CDN(
        n24), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(N1140), .CP(n50), .CDN(n3), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(N1140), .CP(n50), .CDN(
        n12), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(DataI[12]), .E(N1140), .CP(n50), .CDN(
        n12), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(N1140), .CP(n50), .CDN(
        n12), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(N1140), .CP(n50), .CDN(
        n12), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(DataI[9]), .E(N1140), .CP(n50), .CDN(n12), 
        .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(N1140), .CP(n50), .CDN(n12), 
        .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(N1140), .CP(n49), .CDN(n12), 
        .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(DataI[6]), .E(N1140), .CP(n49), .CDN(n12), 
        .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(DataI[5]), .E(N1140), .CP(n49), .CDN(n12), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(N1140), .CP(n49), .CDN(n12), 
        .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(N1140), .CP(n49), .CDN(n12), 
        .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(DataI[2]), .E(N1140), .CP(n49), .CDN(n11), 
        .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(N1140), .CP(n49), .CDN(n11), 
        .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(DataI[0]), .E(N1140), .CP(n49), .CDN(n11), 
        .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(N85), .E(N1107), .CP(n55), .CDN(n8), .Q(
        \Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(N1107), .CP(n55), .CDN(
        n39), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(N1107), .CP(n55), .CDN(
        n28), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(N1107), .CP(n55), .CDN(
        n35), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(N1107), .CP(n55), .CDN(
        n16), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(DataI[27]), .E(N1107), .CP(n55), .CDN(
        n23), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(N1107), .CP(n55), .CDN(
        n27), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(N1107), .CP(n55), .CDN(
        n34), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(N1107), .CP(n54), .CDN(
        n12), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(DataI[23]), .E(N1107), .CP(n54), .CDN(
        n30), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(N1107), .CP(n54), .CDN(
        n32), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(N1107), .CP(n54), .CDN(
        n33), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(N1107), .CP(n54), .CDN(n8), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(N1107), .CP(n54), .CDN(
        n38), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(N1107), .CP(n54), .CDN(
        n40), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(N1107), .CP(n54), .CDN(
        n36), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(N1107), .CP(n54), .CDN(
        n35), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(N1107), .CP(n54), .CDN(
        n37), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(N1107), .CP(n53), .CDN(
        n29), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(DataI[13]), .E(N1107), .CP(n53), .CDN(
        n37), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(N1107), .CP(n53), .CDN(
        n30), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(N1107), .CP(n53), .CDN(
        n23), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(N1107), .CP(n53), .CDN(
        n28), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(N1107), .CP(n53), .CDN(n29), 
        .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(N1107), .CP(n53), .CDN(n3), 
        .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(N1107), .CP(n53), .CDN(n39), 
        .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(DataI[6]), .E(N1107), .CP(n53), .CDN(n29), 
        .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(DataI[5]), .E(N1107), .CP(n53), .CDN(n12), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(N1107), .CP(n52), .CDN(n40), 
        .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(N1107), .CP(n52), .CDN(n35), 
        .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(N1107), .CP(n52), .CDN(n25), 
        .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(N1107), .CP(n52), .CDN(n4), 
        .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(DataI[0]), .E(N1107), .CP(n52), .CDN(n5), 
        .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(N85), .E(N1074), .CP(n59), .CDN(n10), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(DataI[31]), .E(N1074), .CP(n58), .CDN(n4), .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(DataI[30]), .E(N1074), .CP(n58), .CDN(n5), .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(DataI[29]), .E(N1074), .CP(n58), .CDN(n6), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(DataI[28]), .E(N1074), .CP(n58), .CDN(
        n11), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(DataI[27]), .E(N1074), .CP(n58), .CDN(
        n23), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(DataI[26]), .E(N1074), .CP(n58), .CDN(
        n30), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(DataI[25]), .E(N1074), .CP(n58), .CDN(
        n27), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(DataI[24]), .E(N1074), .CP(n58), .CDN(
        n37), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(DataI[23]), .E(N1074), .CP(n58), .CDN(
        n21), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(DataI[22]), .E(N1074), .CP(n58), .CDN(
        n38), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(DataI[21]), .E(N1074), .CP(n57), .CDN(
        n25), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(DataI[20]), .E(N1074), .CP(n57), .CDN(
        n24), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(DataI[19]), .E(N1074), .CP(n57), .CDN(
        n21), .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(DataI[18]), .E(N1074), .CP(n57), .CDN(
        n22), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(DataI[17]), .E(N1074), .CP(n57), .CDN(
        n36), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(DataI[16]), .E(N1074), .CP(n57), .CDN(
        n34), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(DataI[15]), .E(N1074), .CP(n57), .CDN(
        n32), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(DataI[14]), .E(N1074), .CP(n57), .CDN(
        n12), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(DataI[13]), .E(N1074), .CP(n57), .CDN(n8), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(DataI[12]), .E(N1074), .CP(n57), .CDN(
        n32), .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(DataI[11]), .E(N1074), .CP(n56), .CDN(
        n28), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(DataI[10]), .E(N1074), .CP(n56), .CDN(
        n14), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(DataI[9]), .E(N1074), .CP(n56), .CDN(n15), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(DataI[8]), .E(N1074), .CP(n56), .CDN(n16), 
        .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(DataI[7]), .E(N1074), .CP(n56), .CDN(n13), 
        .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(DataI[6]), .E(N1074), .CP(n56), .CDN(n20), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(DataI[5]), .E(N1074), .CP(n56), .CDN(n17), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(DataI[4]), .E(N1074), .CP(n56), .CDN(n18), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(DataI[3]), .E(N1074), .CP(n56), .CDN(n19), 
        .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(DataI[2]), .E(N1074), .CP(n56), .CDN(n6), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(DataI[1]), .E(N1074), .CP(n55), .CDN(n25), 
        .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(DataI[0]), .E(N1074), .CP(n55), .CDN(n40), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(N85), .E(N1041), .CP(n61), .CDN(n31), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(DataI[31]), .E(N1041), .CP(n55), .CDN(
        n11), .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(DataI[30]), .E(N1041), .CP(n47), .CDN(n7), .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(DataI[29]), .E(N1041), .CP(n56), .CDN(
        n27), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(DataI[28]), .E(N1041), .CP(n70), .CDN(
        n12), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(DataI[27]), .E(N1041), .CP(n65), .CDN(
        n29), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(DataI[26]), .E(N1041), .CP(n64), .CDN(
        n12), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(DataI[25]), .E(N1041), .CP(n62), .CDN(
        n22), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(DataI[24]), .E(N1041), .CP(n60), .CDN(n5), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(DataI[23]), .E(N1041), .CP(n61), .CDN(n6), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(DataI[22]), .E(N1041), .CP(n66), .CDN(
        n19), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(DataI[21]), .E(N1041), .CP(n54), .CDN(
        n18), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(DataI[20]), .E(N1041), .CP(n62), .CDN(
        n17), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(DataI[19]), .E(N1041), .CP(n46), .CDN(
        n20), .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(DataI[18]), .E(N1041), .CP(n57), .CDN(
        n13), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(DataI[17]), .E(N1041), .CP(n57), .CDN(
        n16), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(DataI[16]), .E(N1041), .CP(n56), .CDN(
        n15), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(DataI[15]), .E(N1041), .CP(n58), .CDN(
        n14), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(DataI[14]), .E(N1041), .CP(n44), .CDN(
        n26), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(DataI[13]), .E(N1041), .CP(n49), .CDN(
        n19), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(DataI[12]), .E(N1041), .CP(n55), .CDN(
        n33), .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(DataI[11]), .E(N1041), .CP(n41), .CDN(n4), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(DataI[10]), .E(N1041), .CP(n65), .CDN(n5), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(DataI[9]), .E(N1041), .CP(n42), .CDN(n6), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(DataI[8]), .E(N1041), .CP(n59), .CDN(n8), 
        .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(DataI[7]), .E(N1041), .CP(n59), .CDN(n7), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(DataI[6]), .E(N1041), .CP(n59), .CDN(n10), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(DataI[5]), .E(N1041), .CP(n59), .CDN(n9), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(DataI[4]), .E(N1041), .CP(n59), .CDN(n28), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(DataI[3]), .E(N1041), .CP(n59), .CDN(n27), 
        .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(DataI[2]), .E(N1041), .CP(n59), .CDN(n33), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(DataI[1]), .E(N1041), .CP(n59), .CDN(n32), 
        .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(DataI[0]), .E(N1041), .CP(n59), .CDN(n31), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(N85), .E(N975), .CP(n42), .CDN(n16), .Q(
        \Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(DataI[31]), .E(N975), .CP(n42), .CDN(n29), .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(DataI[30]), .E(N975), .CP(n42), .CDN(n9), 
        .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(DataI[29]), .E(N975), .CP(n42), .CDN(n25), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(DataI[28]), .E(N975), .CP(n42), .CDN(n6), 
        .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(DataI[27]), .E(N975), .CP(n42), .CDN(n20), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(DataI[26]), .E(N975), .CP(n66), .CDN(n17), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(DataI[25]), .E(N975), .CP(n49), .CDN(n18), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(DataI[24]), .E(N975), .CP(n48), .CDN(n10), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(DataI[23]), .E(N975), .CP(n41), .CDN(n10), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(DataI[22]), .E(N975), .CP(n52), .CDN(n10), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(DataI[21]), .E(N975), .CP(n53), .CDN(n10), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(DataI[20]), .E(N975), .CP(n51), .CDN(n10), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(DataI[19]), .E(N975), .CP(n50), .CDN(n10), .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(DataI[18]), .E(N975), .CP(n64), .CDN(n10), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(DataI[17]), .E(N975), .CP(n42), .CDN(n10), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(DataI[16]), .E(N975), .CP(n41), .CDN(n10), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(DataI[15]), .E(N975), .CP(n41), .CDN(n10), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(DataI[14]), .E(N975), .CP(n41), .CDN(n10), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(DataI[13]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(DataI[12]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(DataI[11]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(DataI[10]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(DataI[9]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(DataI[8]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(DataI[7]), .E(N975), .CP(n41), .CDN(n9), 
        .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(DataI[6]), .E(N975), .CP(n65), .CDN(n9), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(DataI[5]), .E(N975), .CP(n47), .CDN(n9), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(DataI[4]), .E(N975), .CP(n59), .CDN(n9), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(DataI[3]), .E(N975), .CP(n67), .CDN(n9), 
        .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(DataI[2]), .E(N975), .CP(n42), .CDN(n8), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(DataI[1]), .E(N975), .CP(n49), .CDN(n8), 
        .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(DataI[0]), .E(N975), .CP(n48), .CDN(n8), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(N85), .E(N876), .CP(n68), .CDN(n35), .Q(
        \Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(DataI[31]), .E(N876), .CP(n53), .CDN(n15), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(DataI[30]), .E(N876), .CP(n52), .CDN(n21), .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(DataI[29]), .E(N876), .CP(n48), .CDN(n7), 
        .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(DataI[28]), .E(N876), .CP(n49), .CDN(n39), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(DataI[27]), .E(N876), .CP(n41), .CDN(n11), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(DataI[26]), .E(N876), .CP(n44), .CDN(n28), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(DataI[25]), .E(N876), .CP(n55), .CDN(n40), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(DataI[24]), .E(N876), .CP(n42), .CDN(n25), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(DataI[23]), .E(N876), .CP(n65), .CDN(n29), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(DataI[22]), .E(N876), .CP(n64), .CDN(n11), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(DataI[21]), .E(N876), .CP(n57), .CDN(n28), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(DataI[20]), .E(N876), .CP(n59), .CDN(n27), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(DataI[19]), .E(N876), .CP(n60), .CDN(n26), .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(DataI[18]), .E(N876), .CP(n61), .CDN(n19), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(DataI[17]), .E(N876), .CP(n66), .CDN(n14), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(DataI[16]), .E(N876), .CP(n67), .CDN(n15), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(DataI[15]), .E(N876), .CP(n43), .CDN(n16), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(DataI[14]), .E(N876), .CP(n42), .CDN(n13), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(DataI[13]), .E(N876), .CP(n41), .CDN(n24), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(DataI[12]), .E(N876), .CP(n54), .CDN(n34), .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(DataI[11]), .E(N876), .CP(n58), .CDN(n31), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(DataI[10]), .E(N876), .CP(n63), .CDN(n19), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(DataI[9]), .E(N876), .CP(n66), .CDN(n40), 
        .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(DataI[8]), .E(N876), .CP(n51), .CDN(n13), 
        .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(DataI[7]), .E(N876), .CP(n50), .CDN(n32), 
        .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(DataI[6]), .E(N876), .CP(n55), .CDN(n12), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(DataI[5]), .E(N876), .CP(n54), .CDN(n25), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(DataI[4]), .E(N876), .CP(n58), .CDN(n30), 
        .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(DataI[3]), .E(N876), .CP(n59), .CDN(n11), 
        .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(DataI[2]), .E(N876), .CP(n66), .CDN(n6), 
        .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(DataI[1]), .E(N876), .CP(n67), .CDN(n25), 
        .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(DataI[0]), .E(N876), .CP(n66), .CDN(n30), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(N85), .E(N843), .CP(n55), .CDN(n31), .Q(
        \Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(DataI[31]), .E(N843), .CP(n62), .CDN(n30), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(DataI[30]), .E(N843), .CP(n62), .CDN(n22), .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(DataI[29]), .E(N843), .CP(n44), .CDN(n13), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(DataI[28]), .E(N843), .CP(n42), .CDN(n18), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(DataI[27]), .E(N843), .CP(n43), .CDN(n17), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(DataI[26]), .E(N843), .CP(n55), .CDN(n33), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(DataI[25]), .E(N843), .CP(n54), .CDN(n18), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(DataI[24]), .E(N843), .CP(n58), .CDN(n37), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(DataI[23]), .E(N843), .CP(n59), .CDN(n27), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(DataI[22]), .E(N843), .CP(n56), .CDN(n30), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(DataI[21]), .E(N843), .CP(n57), .CDN(n22), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(DataI[20]), .E(N843), .CP(n60), .CDN(n3), 
        .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(DataI[19]), .E(N843), .CP(n48), .CDN(n29), .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(DataI[18]), .E(N843), .CP(n42), .CDN(n39), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(DataI[17]), .E(N843), .CP(n69), .CDN(
        n108), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(DataI[16]), .E(N843), .CP(n51), .CDN(n10), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(DataI[15]), .E(N843), .CP(ClockW), .CDN(
        n30), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(DataI[14]), .E(N843), .CP(n68), .CDN(n24), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(DataI[13]), .E(N843), .CP(n44), .CDN(n4), 
        .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(DataI[12]), .E(N843), .CP(n60), .CDN(n36), .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(DataI[11]), .E(N843), .CP(n66), .CDN(n27), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(DataI[10]), .E(N843), .CP(n64), .CDN(n38), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(DataI[9]), .E(N843), .CP(n62), .CDN(n40), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(DataI[8]), .E(N843), .CP(n59), .CDN(n28), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(DataI[7]), .E(N843), .CP(n62), .CDN(n24), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(DataI[6]), .E(N843), .CP(n68), .CDN(n29), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(DataI[5]), .E(N843), .CP(n54), .CDN(n12), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(DataI[4]), .E(N843), .CP(n50), .CDN(n10), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(DataI[3]), .E(N843), .CP(n51), .CDN(n22), 
        .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(DataI[2]), .E(N843), .CP(n54), .CDN(n36), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(DataI[1]), .E(N843), .CP(n55), .CDN(n16), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(DataI[0]), .E(N843), .CP(n59), .CDN(n11), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N85), .E(N744), .CP(n56), .CDN(n32), .Q(
        \Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(DataI[31]), .E(N744), .CP(n42), .CDN(n30), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(DataI[30]), .E(N744), .CP(n70), .CDN(n31), .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(DataI[29]), .E(N744), .CP(n70), .CDN(n35), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(DataI[28]), .E(N744), .CP(n63), .CDN(n33), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(DataI[27]), .E(N744), .CP(n58), .CDN(n3), 
        .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(DataI[26]), .E(N744), .CP(n43), .CDN(n39), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(DataI[25]), .E(N744), .CP(n46), .CDN(
        n108), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(DataI[24]), .E(N744), .CP(n70), .CDN(n24), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(DataI[23]), .E(N744), .CP(n55), .CDN(n36), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(DataI[22]), .E(N744), .CP(n64), .CDN(n30), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(DataI[21]), .E(N744), .CP(n54), .CDN(n3), 
        .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(DataI[20]), .E(N744), .CP(n60), .CDN(n37), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(DataI[19]), .E(N744), .CP(n65), .CDN(n7), 
        .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(DataI[18]), .E(N744), .CP(n49), .CDN(n3), 
        .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(DataI[17]), .E(N744), .CP(ClockW), .CDN(
        n28), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(DataI[16]), .E(N744), .CP(n68), .CDN(n27), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(DataI[15]), .E(N744), .CP(n69), .CDN(n26), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(DataI[14]), .E(N744), .CP(n52), .CDN(n22), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(DataI[13]), .E(N744), .CP(n52), .CDN(n24), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(DataI[12]), .E(N744), .CP(n61), .CDN(n36), .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(DataI[11]), .E(N744), .CP(n69), .CDN(n23), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(DataI[10]), .E(N744), .CP(n62), .CDN(n25), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(DataI[9]), .E(N744), .CP(n44), .CDN(n40), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(DataI[8]), .E(N744), .CP(n57), .CDN(n21), 
        .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(DataI[7]), .E(N744), .CP(n43), .CDN(n26), 
        .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(DataI[6]), .E(N744), .CP(n46), .CDN(n40), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(DataI[5]), .E(N744), .CP(n47), .CDN(n13), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(DataI[4]), .E(N744), .CP(n59), .CDN(n16), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(DataI[3]), .E(N744), .CP(n45), .CDN(n15), 
        .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(DataI[2]), .E(N744), .CP(n41), .CDN(n17), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(DataI[1]), .E(N744), .CP(n69), .CDN(n4), 
        .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(DataI[0]), .E(N744), .CP(n55), .CDN(n5), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(N85), .E(N711), .CP(n50), .CDN(n19), .Q(
        \Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(DataI[31]), .E(N711), .CP(n69), .CDN(n18), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(DataI[30]), .E(N711), .CP(n56), .CDN(n17), .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(DataI[29]), .E(N711), .CP(n57), .CDN(n20), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(DataI[28]), .E(N711), .CP(n58), .CDN(n21), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(DataI[27]), .E(N711), .CP(n46), .CDN(n19), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(DataI[26]), .E(N711), .CP(n41), .CDN(n34), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(DataI[25]), .E(N711), .CP(n43), .CDN(n23), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(DataI[24]), .E(N711), .CP(n52), .CDN(n36), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(DataI[23]), .E(N711), .CP(n46), .CDN(n8), 
        .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(DataI[22]), .E(N711), .CP(n60), .CDN(n7), 
        .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(DataI[21]), .E(N711), .CP(n47), .CDN(n4), 
        .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(DataI[20]), .E(N711), .CP(n46), .CDN(n5), 
        .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(DataI[19]), .E(N711), .CP(n45), .CDN(n33), .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(DataI[18]), .E(N711), .CP(n54), .CDN(n25), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(DataI[17]), .E(N711), .CP(n68), .CDN(n19), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(DataI[16]), .E(N711), .CP(n69), .CDN(n23), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(DataI[15]), .E(N711), .CP(n45), .CDN(n25), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(DataI[14]), .E(N711), .CP(n69), .CDN(n38), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(DataI[13]), .E(N711), .CP(n51), .CDN(n20), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(DataI[12]), .E(N711), .CP(n56), .CDN(n23), .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(DataI[11]), .E(N711), .CP(n64), .CDN(n4), 
        .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(DataI[10]), .E(N711), .CP(n44), .CDN(n32), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(DataI[9]), .E(N711), .CP(n62), .CDN(n36), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(DataI[8]), .E(N711), .CP(n45), .CDN(n5), 
        .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(DataI[7]), .E(N711), .CP(n70), .CDN(n26), 
        .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(DataI[6]), .E(N711), .CP(n65), .CDN(n14), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(DataI[5]), .E(N711), .CP(n63), .CDN(n15), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(DataI[4]), .E(N711), .CP(n64), .CDN(n16), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(DataI[3]), .E(N711), .CP(n62), .CDN(n13), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(DataI[2]), .E(N711), .CP(n60), .CDN(n7), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(DataI[1]), .E(N711), .CP(n61), .CDN(n29), 
        .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(DataI[0]), .E(N711), .CP(n68), .CDN(n36), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N85), .E(N612), .CP(n66), .CDN(n13), .Q(
        \Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(DataI[31]), .E(N612), .CP(n49), .CDN(n13), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(DataI[30]), .E(N612), .CP(n70), .CDN(n13), .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(DataI[29]), .E(N612), .CP(n65), .CDN(n13), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(DataI[28]), .E(N612), .CP(n63), .CDN(n13), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(DataI[27]), .E(N612), .CP(n64), .CDN(n13), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(DataI[26]), .E(N612), .CP(n62), .CDN(n13), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(DataI[25]), .E(N612), .CP(n68), .CDN(n38), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(DataI[24]), .E(N612), .CP(n45), .CDN(n32), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(DataI[23]), .E(N612), .CP(n66), .CDN(n8), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(DataI[22]), .E(N612), .CP(n56), .CDN(n4), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(DataI[21]), .E(N612), .CP(n46), .CDN(n29), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(DataI[20]), .E(N612), .CP(n60), .CDN(n35), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(DataI[19]), .E(N612), .CP(n67), .CDN(n28), .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(DataI[18]), .E(N612), .CP(n64), .CDN(n39), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(DataI[17]), .E(N612), .CP(n56), .CDN(n37), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(DataI[16]), .E(N612), .CP(n67), .CDN(n36), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(DataI[15]), .E(N612), .CP(n62), .CDN(n40), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(DataI[14]), .E(N612), .CP(n46), .CDN(n14), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(DataI[13]), .E(N612), .CP(ClockW), .CDN(
        n28), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(DataI[12]), .E(N612), .CP(n70), .CDN(n31), .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(DataI[11]), .E(N612), .CP(n65), .CDN(n14), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(DataI[10]), .E(N612), .CP(n63), .CDN(
        n108), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(DataI[9]), .E(N612), .CP(n64), .CDN(n14), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(DataI[8]), .E(N612), .CP(n62), .CDN(n34), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(DataI[7]), .E(N612), .CP(n60), .CDN(n20), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(DataI[6]), .E(N612), .CP(n61), .CDN(n3), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(DataI[5]), .E(N612), .CP(n62), .CDN(n30), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(DataI[4]), .E(N612), .CP(n45), .CDN(n3), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(DataI[3]), .E(N612), .CP(ClockW), .CDN(
        n30), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(DataI[2]), .E(N612), .CP(n61), .CDN(n30), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(DataI[1]), .E(N612), .CP(n70), .CDN(n32), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(DataI[0]), .E(N612), .CP(n64), .CDN(n33), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N85), .E(N579), .CP(n70), .CDN(n16), .Q(
        \Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(DataI[31]), .E(N579), .CP(n47), .CDN(n16), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(DataI[30]), .E(N579), .CP(n55), .CDN(n16), .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(DataI[29]), .E(N579), .CP(n52), .CDN(n16), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(DataI[28]), .E(N579), .CP(n41), .CDN(n16), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(DataI[27]), .E(N579), .CP(n64), .CDN(n16), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(DataI[26]), .E(N579), .CP(n57), .CDN(n16), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(DataI[25]), .E(N579), .CP(n54), .CDN(n15), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(DataI[24]), .E(N579), .CP(n65), .CDN(n15), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(DataI[23]), .E(N579), .CP(n67), .CDN(n15), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(DataI[22]), .E(N579), .CP(n62), .CDN(n15), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(DataI[21]), .E(N579), .CP(n65), .CDN(n15), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(DataI[20]), .E(N579), .CP(n67), .CDN(n15), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(DataI[19]), .E(N579), .CP(ClockW), .CDN(
        n15), .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(DataI[18]), .E(N579), .CP(n69), .CDN(n15), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(DataI[17]), .E(N579), .CP(n56), .CDN(n15), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(DataI[16]), .E(N579), .CP(n57), .CDN(n15), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(DataI[15]), .E(N579), .CP(n69), .CDN(n15), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(DataI[14]), .E(N579), .CP(n49), .CDN(n14), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(DataI[13]), .E(N579), .CP(n60), .CDN(n14), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(DataI[12]), .E(N579), .CP(n45), .CDN(n14), .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(DataI[11]), .E(N579), .CP(n67), .CDN(n14), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(DataI[10]), .E(N579), .CP(n66), .CDN(n14), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(DataI[9]), .E(N579), .CP(n44), .CDN(n14), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(DataI[8]), .E(N579), .CP(n49), .CDN(n14), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(DataI[7]), .E(N579), .CP(n68), .CDN(n14), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(DataI[6]), .E(N579), .CP(ClockW), .CDN(
        n14), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(DataI[5]), .E(N579), .CP(n61), .CDN(n14), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(DataI[4]), .E(N579), .CP(n68), .CDN(n14), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(DataI[3]), .E(N579), .CP(n47), .CDN(n13), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(DataI[2]), .E(N579), .CP(n60), .CDN(n13), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(DataI[1]), .E(N579), .CP(n61), .CDN(n13), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(DataI[0]), .E(N579), .CP(n65), .CDN(n13), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N85), .E(N480), .CP(n68), .CDN(n25), .Q(
        \Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(DataI[31]), .E(N480), .CP(n51), .CDN(n25), .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(DataI[30]), .E(N480), .CP(n65), .CDN(n25), .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(DataI[29]), .E(N480), .CP(n68), .CDN(n25), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(DataI[28]), .E(N480), .CP(n41), .CDN(n25), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(DataI[27]), .E(N480), .CP(n56), .CDN(n25), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(DataI[26]), .E(N480), .CP(n54), .CDN(n25), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(DataI[25]), .E(N480), .CP(n54), .CDN(n24), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(DataI[24]), .E(N480), .CP(n43), .CDN(n24), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(DataI[23]), .E(N480), .CP(n66), .CDN(n24), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(DataI[22]), .E(N480), .CP(n56), .CDN(n24), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(DataI[21]), .E(N480), .CP(n42), .CDN(n24), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(DataI[20]), .E(N480), .CP(n46), .CDN(n24), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(DataI[19]), .E(N480), .CP(n60), .CDN(n24), .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(DataI[18]), .E(N480), .CP(n59), .CDN(n24), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(DataI[17]), .E(N480), .CP(n65), .CDN(n24), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(DataI[16]), .E(N480), .CP(n62), .CDN(n24), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(DataI[15]), .E(N480), .CP(n42), .CDN(n24), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(DataI[14]), .E(N480), .CP(n60), .CDN(n23), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(DataI[13]), .E(N480), .CP(n46), .CDN(n23), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(DataI[12]), .E(N480), .CP(n59), .CDN(n23), .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(DataI[11]), .E(N480), .CP(n62), .CDN(n23), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(DataI[10]), .E(N480), .CP(n60), .CDN(n23), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(DataI[9]), .E(N480), .CP(n61), .CDN(n23), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(DataI[8]), .E(N480), .CP(n65), .CDN(n23), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(DataI[7]), .E(N480), .CP(n63), .CDN(n23), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(DataI[6]), .E(N480), .CP(n64), .CDN(n23), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(DataI[5]), .E(N480), .CP(n67), .CDN(n23), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(DataI[4]), .E(N480), .CP(n69), .CDN(n23), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(DataI[3]), .E(N480), .CP(n56), .CDN(n22), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(DataI[2]), .E(N480), .CP(n48), .CDN(n22), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(DataI[1]), .E(N480), .CP(n46), .CDN(n22), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(DataI[0]), .E(N480), .CP(n66), .CDN(n22), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N85), .E(N447), .CP(n69), .CDN(n17), .Q(
        \Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(DataI[31]), .E(N447), .CP(n58), .CDN(n20), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(DataI[30]), .E(N447), .CP(n41), .CDN(n34), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(DataI[29]), .E(N447), .CP(n58), .CDN(n32), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(DataI[28]), .E(N447), .CP(n61), .CDN(n31), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(DataI[27]), .E(N447), .CP(n63), .CDN(n30), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(DataI[26]), .E(N447), .CP(n51), .CDN(n3), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(DataI[25]), .E(N447), .CP(n67), .CDN(n30), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(DataI[24]), .E(N447), .CP(n53), .CDN(n17), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(DataI[23]), .E(N447), .CP(n57), .CDN(n20), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(DataI[22]), .E(N447), .CP(n49), .CDN(n26), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(DataI[21]), .E(N447), .CP(n59), .CDN(n13), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(DataI[20]), .E(N447), .CP(n57), .CDN(n16), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(DataI[19]), .E(N447), .CP(n66), .CDN(n15), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(DataI[18]), .E(N447), .CP(n50), .CDN(n14), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(DataI[17]), .E(N447), .CP(n55), .CDN(n12), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(DataI[16]), .E(N447), .CP(n47), .CDN(n18), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(DataI[15]), .E(N447), .CP(n68), .CDN(n19), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(DataI[14]), .E(N447), .CP(n43), .CDN(n36), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(DataI[13]), .E(N447), .CP(n45), .CDN(n30), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(DataI[12]), .E(N447), .CP(n48), .CDN(n40), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(DataI[11]), .E(N447), .CP(n44), .CDN(n38), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(DataI[10]), .E(N447), .CP(n66), .CDN(n10), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(DataI[9]), .E(N447), .CP(n64), .CDN(n33), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(DataI[8]), .E(N447), .CP(ClockW), .CDN(n17), .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(DataI[7]), .E(N447), .CP(n54), .CDN(n20), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(DataI[6]), .E(N447), .CP(n55), .CDN(n4), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(DataI[5]), .E(N447), .CP(n70), .CDN(n5), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(DataI[4]), .E(N447), .CP(n47), .CDN(n6), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(DataI[3]), .E(N447), .CP(n58), .CDN(n25), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(DataI[2]), .E(N447), .CP(n62), .CDN(n25), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(DataI[1]), .E(N447), .CP(n67), .CDN(n25), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(DataI[0]), .E(N447), .CP(n53), .CDN(n25), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N85), .E(N348), .CP(n59), .CDN(n15), .Q(
        \Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(N348), .CP(n69), .CDN(n9), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(N348), .CP(n53), .CDN(n8), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(N348), .CP(n66), .CDN(n40), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(N348), .CP(n64), .CDN(n38), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(N348), .CP(n45), .CDN(n30), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(N348), .CP(n56), .CDN(n13), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(N348), .CP(n68), .CDN(n34), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(N348), .CP(n49), .CDN(n26), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(N348), .CP(n46), .CDN(n11), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(N348), .CP(n43), .CDN(n18), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(N348), .CP(n52), .CDN(n4), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(N348), .CP(n68), .CDN(n40), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(N348), .CP(n68), .CDN(n6), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(N348), .CP(n69), .CDN(n39), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(N348), .CP(n48), .CDN(n13), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(N348), .CP(ClockW), .CDN(
        n28), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(N348), .CP(n45), .CDN(n34), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(N348), .CP(n53), .CDN(n27), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(N348), .CP(n47), .CDN(n29), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(N348), .CP(n46), .CDN(n108), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(N348), .CP(n61), .CDN(n33), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(N348), .CP(ClockW), .CDN(
        n32), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(N348), .CP(n44), .CDN(n31), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(N348), .CP(n65), .CDN(n30), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(N348), .CP(n50), .CDN(n13), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(N348), .CP(n63), .CDN(n35), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(N348), .CP(n41), .CDN(n16), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(N348), .CP(n44), .CDN(n23), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(N348), .CP(n68), .CDN(n33), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(N348), .CP(n67), .CDN(n6), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(N348), .CP(n66), .CDN(n30), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(N348), .CP(n60), .CDN(n33), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N85), .E(N315), .CP(n52), .CDN(n32), .Q(
        \Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(N315), .CP(n55), .CDN(n6), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(N315), .CP(n42), .CDN(n15), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(N315), .CP(n60), .CDN(n13), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(N315), .CP(n45), .CDN(n10), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(N315), .CP(n49), .CDN(n36), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(N315), .CP(n45), .CDN(n15), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(N315), .CP(ClockW), .CDN(
        n35), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(N315), .CP(n44), .CDN(n6), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(N315), .CP(n52), .CDN(n16), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(N315), .CP(n50), .CDN(n33), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(N315), .CP(n62), .CDN(n31), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(N315), .CP(n63), .CDN(n108), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(N315), .CP(n67), .CDN(n29), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(N315), .CP(n47), .CDN(n40), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(N315), .CP(n62), .CDN(n39), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(N315), .CP(n45), .CDN(n13), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(N315), .CP(n53), .CDN(n20), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(N315), .CP(n51), .CDN(n36), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(N315), .CP(ClockW), .CDN(
        n30), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(N315), .CP(n45), .CDN(n34), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(N315), .CP(n66), .CDN(n37), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(N315), .CP(n67), .CDN(n35), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(N315), .CP(n45), .CDN(n108), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(N315), .CP(n47), .CDN(n19), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(N315), .CP(n44), .CDN(n9), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(N315), .CP(n68), .CDN(n36), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(N315), .CP(n46), .CDN(n38), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(N315), .CP(n42), .CDN(n40), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(N315), .CP(n43), .CDN(n30), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(N315), .CP(n51), .CDN(n12), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(N315), .CP(n41), .CDN(n9), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(N315), .CP(n51), .CDN(n37), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(N216), .CP(n68), .CDN(n35), .Q(
        \Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(N216), .CP(n48), .CDN(n38), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(N216), .CP(n69), .CDN(n18), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(N216), .CP(n70), .CDN(n14), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(N216), .CP(n62), .CDN(n35), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(N216), .CP(n41), .CDN(n18), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(N216), .CP(n66), .CDN(n8), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(N216), .CP(n42), .CDN(n3), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(N216), .CP(n61), .CDN(n33), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(N216), .CP(n66), .CDN(n11), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(N216), .CP(n67), .CDN(n38), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(N216), .CP(n44), .CDN(n108), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(N216), .CP(n50), .CDN(n38), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(N216), .CP(n43), .CDN(n15), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(N216), .CP(n64), .CDN(n32), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(N216), .CP(n61), .CDN(n29), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(N216), .CP(n63), .CDN(n20), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(N216), .CP(n61), .CDN(n9), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(N216), .CP(n68), .CDN(n34), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(N216), .CP(ClockW), .CDN(
        n18), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(N216), .CP(n51), .CDN(n40), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(N216), .CP(n61), .CDN(n108), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(N216), .CP(n43), .CDN(n33), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(N216), .CP(n44), .CDN(n32), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(N216), .CP(n41), .CDN(n21), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(N216), .CP(ClockW), .CDN(n29), .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(N216), .CP(n51), .CDN(n39), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(N216), .CP(n63), .CDN(n29), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(N216), .CP(n43), .CDN(n36), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(N216), .CP(n49), .CDN(n40), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(N216), .CP(n50), .CDN(n36), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(N216), .CP(n66), .CDN(n35), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(N216), .CP(n46), .CDN(n19), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N85), .E(N183), .CP(n50), .CDN(n21), .Q(
        \Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(N183), .CP(n64), .CDN(n31), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(N183), .CP(n54), .CDN(n38), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(N183), .CP(n45), .CDN(n7), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(N183), .CP(n58), .CDN(n26), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(N183), .CP(n48), .CDN(n27), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(N183), .CP(n53), .CDN(n39), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(N183), .CP(n52), .CDN(n29), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(N183), .CP(n63), .CDN(n38), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(N183), .CP(n68), .CDN(n16), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(N183), .CP(n46), .CDN(n37), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(N183), .CP(n47), .CDN(n36), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(N183), .CP(n62), .CDN(n37), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(N183), .CP(n58), .CDN(n8), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(N183), .CP(n52), .CDN(n32), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(N183), .CP(n69), .CDN(n7), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(N183), .CP(n52), .CDN(n19), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(N183), .CP(ClockW), .CDN(
        n34), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(N183), .CP(n68), .CDN(n38), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(N183), .CP(n43), .CDN(n28), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(N183), .CP(n58), .CDN(n7), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(N183), .CP(n63), .CDN(n26), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(N183), .CP(n64), .CDN(n34), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(N183), .CP(n62), .CDN(n15), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(N183), .CP(n60), .CDN(n30), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(N183), .CP(n61), .CDN(n31), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(N183), .CP(n66), .CDN(n32), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(N183), .CP(n67), .CDN(n33), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(N183), .CP(n63), .CDN(n14), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(N183), .CP(n53), .CDN(n37), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(N183), .CP(n47), .CDN(n36), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(N183), .CP(n43), .CDN(n37), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(N183), .CP(n50), .CDN(n31), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(N414), .CP(n57), .CDN(n28), .Q(
        \Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(DataI[31]), .E(N414), .CP(n63), .CDN(n28), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(DataI[30]), .E(N414), .CP(n44), .CDN(n28), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(DataI[29]), .E(N414), .CP(n47), .CDN(n28), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(DataI[28]), .E(N414), .CP(n68), .CDN(n28), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(N150), .CP(n58), .CDN(n28), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(N85), .E(N909), .CP(n63), .CDN(n12), .Q(
        \Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(DataI[31]), .E(N909), .CP(n44), .CDN(n39), .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(DataI[30]), .E(N909), .CP(n70), .CDN(n29), .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(DataI[29]), .E(N909), .CP(n42), .CDN(n35), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(DataI[28]), .E(N909), .CP(n43), .CDN(n36), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(DataI[27]), .E(N909), .CP(n46), .CDN(n37), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(DataI[26]), .E(N909), .CP(n47), .CDN(n13), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(DataI[25]), .E(N909), .CP(n63), .CDN(n13), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(DataI[24]), .E(N909), .CP(n54), .CDN(n21), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(DataI[23]), .E(N909), .CP(n58), .CDN(n23), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(DataI[22]), .E(N909), .CP(n43), .CDN(n7), 
        .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(DataI[21]), .E(N909), .CP(n42), .CDN(n10), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(DataI[20]), .E(N909), .CP(n44), .CDN(n9), 
        .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(DataI[19]), .E(N909), .CP(n45), .CDN(n32), .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(DataI[18]), .E(N909), .CP(n46), .CDN(n23), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(DataI[17]), .E(N909), .CP(n47), .CDN(n20), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(DataI[16]), .E(N909), .CP(n52), .CDN(n17), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(DataI[15]), .E(N909), .CP(n56), .CDN(n18), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(DataI[14]), .E(N909), .CP(n66), .CDN(n24), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(DataI[13]), .E(N909), .CP(n63), .CDN(n5), 
        .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(DataI[12]), .E(N909), .CP(n69), .CDN(n22), .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(DataI[11]), .E(N909), .CP(n67), .CDN(n18), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(DataI[10]), .E(N909), .CP(n41), .CDN(n17), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(DataI[9]), .E(N909), .CP(n61), .CDN(n20), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(DataI[8]), .E(N909), .CP(n47), .CDN(n24), 
        .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(DataI[7]), .E(N909), .CP(n46), .CDN(n23), 
        .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(DataI[6]), .E(N909), .CP(n57), .CDN(n33), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(DataI[5]), .E(N909), .CP(n58), .CDN(n25), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(DataI[4]), .E(N909), .CP(n57), .CDN(n11), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(DataI[3]), .E(N909), .CP(n60), .CDN(n38), 
        .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(DataI[2]), .E(N909), .CP(n64), .CDN(n18), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(DataI[1]), .E(N909), .CP(n57), .CDN(n5), 
        .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(DataI[0]), .E(N909), .CP(n63), .CDN(n37), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N85), .E(N810), .CP(n49), .CDN(n24), .Q(
        \Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(DataI[31]), .E(N810), .CP(n48), .CDN(n21), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(DataI[30]), .E(N810), .CP(n52), .CDN(n10), .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(DataI[29]), .E(N810), .CP(n53), .CDN(n15), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(DataI[28]), .E(N810), .CP(n50), .CDN(n38), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(DataI[27]), .E(N810), .CP(n51), .CDN(n3), 
        .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(DataI[26]), .E(N810), .CP(n55), .CDN(n31), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(DataI[25]), .E(N810), .CP(n50), .CDN(n25), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(DataI[24]), .E(N810), .CP(n63), .CDN(n26), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(DataI[23]), .E(N810), .CP(n47), .CDN(n10), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(DataI[22]), .E(N810), .CP(n67), .CDN(n21), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(DataI[21]), .E(N810), .CP(n69), .CDN(n25), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(DataI[20]), .E(N810), .CP(n69), .CDN(n35), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(DataI[19]), .E(N810), .CP(n50), .CDN(n23), .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(DataI[18]), .E(N810), .CP(n52), .CDN(n13), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(DataI[17]), .E(N810), .CP(n57), .CDN(n16), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(DataI[16]), .E(N810), .CP(n69), .CDN(n15), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(DataI[15]), .E(N810), .CP(n41), .CDN(n14), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(DataI[14]), .E(N810), .CP(n43), .CDN(n19), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(DataI[13]), .E(N810), .CP(n65), .CDN(n32), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(DataI[12]), .E(N810), .CP(n56), .CDN(n23), .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(DataI[11]), .E(N810), .CP(n64), .CDN(n33), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(DataI[10]), .E(N810), .CP(n63), .CDN(n17), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(DataI[9]), .E(N810), .CP(n65), .CDN(n31), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(DataI[8]), .E(N810), .CP(n61), .CDN(n20), 
        .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(DataI[7]), .E(N810), .CP(n60), .CDN(n38), 
        .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(DataI[6]), .E(N810), .CP(n51), .CDN(n33), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(DataI[5]), .E(N810), .CP(n68), .CDN(n22), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(DataI[4]), .E(N810), .CP(n70), .CDN(n30), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(DataI[3]), .E(N810), .CP(n52), .CDN(n7), 
        .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(DataI[2]), .E(N810), .CP(n66), .CDN(n34), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(DataI[1]), .E(N810), .CP(n67), .CDN(n10), 
        .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(DataI[0]), .E(N810), .CP(n60), .CDN(n21), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(N85), .E(N777), .CP(n68), .CDN(n8), .Q(
        \Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(DataI[31]), .E(N777), .CP(n60), .CDN(n7), 
        .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(DataI[30]), .E(N777), .CP(n61), .CDN(n10), .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(DataI[29]), .E(N777), .CP(n64), .CDN(n9), 
        .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(DataI[28]), .E(N777), .CP(n63), .CDN(n5), 
        .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(DataI[27]), .E(N777), .CP(n55), .CDN(n33), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(DataI[26]), .E(N777), .CP(n70), .CDN(n17), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(DataI[25]), .E(N777), .CP(n59), .CDN(n6), 
        .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(DataI[24]), .E(N777), .CP(n59), .CDN(n8), 
        .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(DataI[23]), .E(N777), .CP(n58), .CDN(n32), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(DataI[22]), .E(N777), .CP(n69), .CDN(n31), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(DataI[21]), .E(N777), .CP(n70), .CDN(n3), 
        .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(DataI[20]), .E(N777), .CP(n43), .CDN(n11), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(DataI[19]), .E(N777), .CP(n70), .CDN(n35), .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(DataI[18]), .E(N777), .CP(n64), .CDN(n22), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(DataI[17]), .E(N777), .CP(n41), .CDN(n12), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(DataI[16]), .E(N777), .CP(n53), .CDN(n40), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(DataI[15]), .E(N777), .CP(n51), .CDN(n15), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(DataI[14]), .E(N777), .CP(n67), .CDN(n35), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(DataI[13]), .E(N777), .CP(n64), .CDN(n40), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(DataI[12]), .E(N777), .CP(n57), .CDN(n38), .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(DataI[11]), .E(N777), .CP(n56), .CDN(n28), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(DataI[10]), .E(N777), .CP(n48), .CDN(n36), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(DataI[9]), .E(N777), .CP(n49), .CDN(n35), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(DataI[8]), .E(N777), .CP(n53), .CDN(n20), 
        .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(DataI[7]), .E(N777), .CP(n52), .CDN(n38), 
        .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(DataI[6]), .E(N777), .CP(n50), .CDN(n19), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(DataI[5]), .E(N777), .CP(n51), .CDN(n37), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(DataI[4]), .E(N777), .CP(n60), .CDN(n14), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(DataI[3]), .E(N777), .CP(n65), .CDN(n39), 
        .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(DataI[2]), .E(N777), .CP(n57), .CDN(n32), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(DataI[1]), .E(N777), .CP(n56), .CDN(n8), 
        .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(DataI[0]), .E(N777), .CP(n59), .CDN(n7), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(N678), .CP(n43), .CDN(n35), .Q(
        \Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(DataI[31]), .E(N678), .CP(n42), .CDN(n6), 
        .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(DataI[30]), .E(N678), .CP(n45), .CDN(n4), 
        .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(DataI[29]), .E(N678), .CP(n45), .CDN(n5), 
        .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(DataI[28]), .E(N678), .CP(n67), .CDN(n6), 
        .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(DataI[27]), .E(N678), .CP(n58), .CDN(n8), 
        .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(DataI[26]), .E(N678), .CP(n56), .CDN(n7), 
        .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(DataI[25]), .E(N678), .CP(n70), .CDN(n10), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(DataI[24]), .E(N678), .CP(n50), .CDN(n12), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(DataI[23]), .E(N678), .CP(n51), .CDN(n4), 
        .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(DataI[22]), .E(N678), .CP(n53), .CDN(n9), 
        .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(DataI[21]), .E(N678), .CP(n44), .CDN(n10), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(DataI[20]), .E(N678), .CP(n42), .CDN(n18), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(DataI[19]), .E(N678), .CP(n54), .CDN(n34), .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(DataI[18]), .E(N678), .CP(n48), .CDN(n29), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(DataI[17]), .E(N678), .CP(n55), .CDN(n35), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(DataI[16]), .E(N678), .CP(n53), .CDN(n11), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(DataI[15]), .E(N678), .CP(n63), .CDN(n37), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(DataI[14]), .E(N678), .CP(n53), .CDN(n26), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(DataI[13]), .E(N678), .CP(n49), .CDN(n8), 
        .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(DataI[12]), .E(N678), .CP(ClockW), .CDN(
        n18), .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(DataI[11]), .E(N678), .CP(ClockW), .CDN(
        n38), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(DataI[10]), .E(N678), .CP(n41), .CDN(n19), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(DataI[9]), .E(N678), .CP(n53), .CDN(n39), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(DataI[8]), .E(N678), .CP(n49), .CDN(n9), 
        .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(DataI[7]), .E(N678), .CP(n54), .CDN(n12), 
        .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(DataI[6]), .E(N678), .CP(n61), .CDN(n6), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(DataI[5]), .E(N678), .CP(n42), .CDN(n33), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(DataI[4]), .E(N678), .CP(n59), .CDN(n39), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(DataI[3]), .E(N678), .CP(n54), .CDN(n40), 
        .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(DataI[2]), .E(N678), .CP(n55), .CDN(n19), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(DataI[1]), .E(N678), .CP(n51), .CDN(n18), 
        .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(DataI[0]), .E(N678), .CP(n50), .CDN(n32), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N85), .E(N645), .CP(n63), .CDN(n34), .Q(
        \Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(DataI[31]), .E(N645), .CP(n65), .CDN(n34), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(DataI[30]), .E(N645), .CP(n61), .CDN(n9), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(DataI[29]), .E(N645), .CP(n60), .CDN(n16), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(DataI[28]), .E(N645), .CP(n54), .CDN(n34), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(DataI[27]), .E(N645), .CP(n63), .CDN(n36), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(DataI[26]), .E(N645), .CP(n54), .CDN(n14), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(DataI[25]), .E(N645), .CP(n48), .CDN(n39), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(DataI[24]), .E(N645), .CP(n55), .CDN(n33), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(DataI[23]), .E(N645), .CP(n64), .CDN(n30), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(DataI[22]), .E(N645), .CP(n52), .CDN(n39), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(DataI[21]), .E(N645), .CP(n66), .CDN(n16), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(DataI[20]), .E(N645), .CP(n66), .CDN(n39), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(DataI[19]), .E(N645), .CP(n45), .CDN(n4), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(DataI[18]), .E(N645), .CP(ClockW), .CDN(
        n15), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(DataI[17]), .E(N645), .CP(n53), .CDN(n26), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(DataI[16]), .E(N645), .CP(ClockW), .CDN(
        n12), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(DataI[15]), .E(N645), .CP(n69), .CDN(
        n108), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(DataI[14]), .E(N645), .CP(n54), .CDN(n21), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(DataI[13]), .E(N645), .CP(n59), .CDN(n17), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(DataI[12]), .E(N645), .CP(n67), .CDN(n29), .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(DataI[11]), .E(N645), .CP(n53), .CDN(n38), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(DataI[10]), .E(N645), .CP(n48), .CDN(n31), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(DataI[9]), .E(N645), .CP(n70), .CDN(n37), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(DataI[8]), .E(N645), .CP(n70), .CDN(n31), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(DataI[7]), .E(N645), .CP(n42), .CDN(n24), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(DataI[6]), .E(N645), .CP(n70), .CDN(n24), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(DataI[5]), .E(N645), .CP(ClockW), .CDN(n9), .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(DataI[4]), .E(N645), .CP(n61), .CDN(n14), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(DataI[3]), .E(N645), .CP(n60), .CDN(n40), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(DataI[2]), .E(N645), .CP(n62), .CDN(n23), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(DataI[1]), .E(N645), .CP(n63), .CDN(n15), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(DataI[0]), .E(N645), .CP(n65), .CDN(n35), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(N546), .CP(n45), .CDN(n19), .Q(
        \Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(DataI[31]), .E(N546), .CP(n54), .CDN(n19), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(DataI[30]), .E(N546), .CP(n42), .CDN(n19), .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(DataI[29]), .E(N546), .CP(n53), .CDN(n19), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(DataI[28]), .E(N546), .CP(n47), .CDN(n19), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(DataI[27]), .E(N546), .CP(n66), .CDN(n19), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(DataI[26]), .E(N546), .CP(n57), .CDN(n19), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(DataI[25]), .E(N546), .CP(n50), .CDN(n18), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(DataI[24]), .E(N546), .CP(n47), .CDN(n18), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(DataI[23]), .E(N546), .CP(ClockW), .CDN(
        n18), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(DataI[22]), .E(N546), .CP(n67), .CDN(n18), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(DataI[21]), .E(N546), .CP(n47), .CDN(n18), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(DataI[20]), .E(N546), .CP(n43), .CDN(n18), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(DataI[19]), .E(N546), .CP(n44), .CDN(n18), .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(DataI[18]), .E(N546), .CP(n59), .CDN(n18), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(DataI[17]), .E(N546), .CP(n56), .CDN(n18), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(DataI[16]), .E(N546), .CP(n59), .CDN(n18), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(DataI[15]), .E(N546), .CP(n65), .CDN(n18), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(DataI[14]), .E(N546), .CP(n57), .CDN(n17), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(DataI[13]), .E(N546), .CP(n48), .CDN(n17), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(DataI[12]), .E(N546), .CP(n50), .CDN(n17), .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(DataI[11]), .E(N546), .CP(n47), .CDN(n17), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(DataI[10]), .E(N546), .CP(ClockW), .CDN(
        n17), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(DataI[9]), .E(N546), .CP(n48), .CDN(n17), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(DataI[8]), .E(N546), .CP(n41), .CDN(n17), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(DataI[7]), .E(N546), .CP(n51), .CDN(n17), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(DataI[6]), .E(N546), .CP(ClockW), .CDN(
        n17), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(DataI[5]), .E(N546), .CP(n66), .CDN(n17), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(DataI[4]), .E(N546), .CP(n49), .CDN(n17), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(DataI[3]), .E(N546), .CP(n60), .CDN(n16), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(DataI[2]), .E(N546), .CP(n64), .CDN(n16), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(DataI[1]), .E(N546), .CP(n47), .CDN(n16), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(DataI[0]), .E(N546), .CP(n69), .CDN(n16), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N85), .E(N513), .CP(n61), .CDN(n22), .Q(
        \Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(DataI[31]), .E(N513), .CP(n59), .CDN(n22), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(DataI[30]), .E(N513), .CP(n46), .CDN(n22), .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(DataI[29]), .E(N513), .CP(n65), .CDN(n22), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(DataI[28]), .E(N513), .CP(ClockW), .CDN(
        n22), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(DataI[27]), .E(N513), .CP(n65), .CDN(n22), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(DataI[26]), .E(N513), .CP(n45), .CDN(n22), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(DataI[25]), .E(N513), .CP(n56), .CDN(n21), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(DataI[24]), .E(N513), .CP(n57), .CDN(n21), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(DataI[23]), .E(N513), .CP(n46), .CDN(n21), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(DataI[22]), .E(N513), .CP(n69), .CDN(n21), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(DataI[21]), .E(N513), .CP(n68), .CDN(n21), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(DataI[20]), .E(N513), .CP(n44), .CDN(n21), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(DataI[19]), .E(N513), .CP(n43), .CDN(n21), .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(DataI[18]), .E(N513), .CP(n70), .CDN(n21), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(DataI[17]), .E(N513), .CP(n52), .CDN(n21), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(DataI[16]), .E(N513), .CP(n48), .CDN(n21), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(DataI[15]), .E(N513), .CP(n41), .CDN(n21), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(DataI[14]), .E(N513), .CP(n59), .CDN(n20), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(DataI[13]), .E(N513), .CP(n42), .CDN(n20), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(DataI[12]), .E(N513), .CP(n63), .CDN(n20), .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(DataI[11]), .E(N513), .CP(n47), .CDN(n20), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(DataI[10]), .E(N513), .CP(n70), .CDN(n20), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(DataI[9]), .E(N513), .CP(n41), .CDN(n20), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(DataI[8]), .E(N513), .CP(n62), .CDN(n20), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(DataI[7]), .E(N513), .CP(n49), .CDN(n20), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(DataI[6]), .E(N513), .CP(n70), .CDN(n20), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(DataI[5]), .E(N513), .CP(n49), .CDN(n20), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(DataI[4]), .E(N513), .CP(n44), .CDN(n20), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(DataI[3]), .E(N513), .CP(n48), .CDN(n19), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(DataI[2]), .E(N513), .CP(n70), .CDN(n19), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(DataI[1]), .E(N513), .CP(n58), .CDN(n19), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(DataI[0]), .E(N513), .CP(n41), .CDN(n19), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(DataI[27]), .E(N414), .CP(n70), .CDN(n28), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(DataI[26]), .E(N414), .CP(n60), .CDN(n28), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(DataI[25]), .E(N414), .CP(n57), .CDN(n27), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(DataI[24]), .E(N414), .CP(n42), .CDN(n27), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(DataI[23]), .E(N414), .CP(n42), .CDN(n27), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(DataI[22]), .E(N414), .CP(n60), .CDN(n27), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(DataI[21]), .E(N414), .CP(n51), .CDN(n27), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(DataI[20]), .E(N414), .CP(n66), .CDN(n27), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(DataI[19]), .E(N414), .CP(n54), .CDN(n27), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(DataI[18]), .E(N414), .CP(n62), .CDN(n27), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(DataI[17]), .E(N414), .CP(n64), .CDN(n27), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(DataI[16]), .E(N414), .CP(n58), .CDN(n27), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(DataI[15]), .E(N414), .CP(ClockW), .CDN(
        n27), .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(DataI[14]), .E(N414), .CP(n46), .CDN(n26), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(DataI[13]), .E(N414), .CP(ClockW), .CDN(
        n26), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(DataI[12]), .E(N414), .CP(n53), .CDN(n26), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(DataI[11]), .E(N414), .CP(n50), .CDN(n26), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(DataI[10]), .E(N414), .CP(n48), .CDN(n26), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(DataI[9]), .E(N414), .CP(n49), .CDN(n26), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(DataI[8]), .E(N414), .CP(n62), .CDN(n26), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(DataI[7]), .E(N414), .CP(n61), .CDN(n26), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(DataI[6]), .E(N414), .CP(n62), .CDN(n26), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(DataI[5]), .E(N414), .CP(n70), .CDN(n26), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(DataI[4]), .E(N414), .CP(n65), .CDN(n26), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(DataI[3]), .E(N414), .CP(n48), .CDN(n39), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(DataI[2]), .E(N414), .CP(ClockW), .CDN(n29), .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(DataI[1]), .E(N414), .CP(ClockW), .CDN(n37), .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(DataI[0]), .E(N414), .CP(n68), .CDN(n35), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N85), .E(N381), .CP(n54), .CDN(n12), .Q(
        \Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(N381), .CP(n65), .CDN(n38), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(N381), .CP(n55), .CDN(n25), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(N381), .CP(n54), .CDN(n22), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(N381), .CP(n59), .CDN(n27), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(N381), .CP(n58), .CDN(n37), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(N381), .CP(n57), .CDN(n35), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(N381), .CP(n56), .CDN(n40), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(N381), .CP(n51), .CDN(n11), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(N381), .CP(n50), .CDN(n17), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(N381), .CP(n52), .CDN(n20), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(N381), .CP(n59), .CDN(n22), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(N381), .CP(n60), .CDN(n21), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(N381), .CP(n49), .CDN(n24), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(N381), .CP(n48), .CDN(n23), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(N381), .CP(n52), .CDN(n25), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(N381), .CP(n53), .CDN(n36), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(N381), .CP(n51), .CDN(n22), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(N381), .CP(n50), .CDN(n11), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(N381), .CP(n55), .CDN(n7), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(N381), .CP(n54), .CDN(n12), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(N381), .CP(n67), .CDN(n17), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(N381), .CP(n48), .CDN(n26), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(N381), .CP(n69), .CDN(n14), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(N381), .CP(n57), .CDN(n28), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(N381), .CP(n56), .CDN(n27), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(N381), .CP(n63), .CDN(n26), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(N381), .CP(n48), .CDN(n12), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(N381), .CP(n49), .CDN(n9), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(N381), .CP(n44), .CDN(n33), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(N381), .CP(n44), .CDN(n9), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(N381), .CP(n67), .CDN(n38), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(N381), .CP(n51), .CDN(n3), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(N282), .CP(n56), .CDN(n8), .Q(
        \Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(N282), .CP(n68), .CDN(n28), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(N282), .CP(n48), .CDN(n16), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(N282), .CP(n43), .CDN(n17), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(N282), .CP(n63), .CDN(n10), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(N282), .CP(n68), .CDN(n31), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(N282), .CP(n69), .CDN(n27), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(N282), .CP(n67), .CDN(n30), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(N282), .CP(n55), .CDN(n3), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(N282), .CP(n70), .CDN(n39), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(N282), .CP(n63), .CDN(n21), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(N282), .CP(n55), .CDN(n37), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(N282), .CP(n64), .CDN(n25), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(N282), .CP(n45), .CDN(n39), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(N282), .CP(n49), .CDN(n39), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(N282), .CP(ClockW), .CDN(
        n29), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(N282), .CP(n62), .CDN(n22), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(N282), .CP(n60), .CDN(n8), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(N282), .CP(n61), .CDN(n37), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(N282), .CP(n64), .CDN(n28), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(N282), .CP(ClockW), .CDN(
        n26), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(N282), .CP(n65), .CDN(n9), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(N282), .CP(n63), .CDN(n4), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(N282), .CP(n61), .CDN(n14), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(N282), .CP(n48), .CDN(n37), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(N282), .CP(n58), .CDN(n36), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(N282), .CP(n53), .CDN(n40), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(N282), .CP(n64), .CDN(n108), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(N282), .CP(ClockW), .CDN(n38), .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(N282), .CP(n53), .CDN(n35), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(N282), .CP(n69), .CDN(n31), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(N282), .CP(n49), .CDN(n34), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(N282), .CP(n68), .CDN(n6), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N85), .E(N249), .CP(n52), .CDN(n39), .Q(
        \Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(N249), .CP(n70), .CDN(n5), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(N249), .CP(n43), .CDN(n34), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(N249), .CP(n67), .CDN(n40), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(N249), .CP(n46), .CDN(n39), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(N249), .CP(ClockW), .CDN(
        n29), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(N249), .CP(n51), .CDN(n26), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(N249), .CP(n52), .CDN(n108), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(N249), .CP(n56), .CDN(n35), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(N249), .CP(n65), .CDN(n37), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(N249), .CP(n50), .CDN(n19), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(N249), .CP(n58), .CDN(n5), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(N249), .CP(n41), .CDN(n10), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(N249), .CP(n42), .CDN(n5), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(N249), .CP(n47), .CDN(n35), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(N249), .CP(n44), .CDN(n19), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(N249), .CP(n65), .CDN(n36), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(N249), .CP(n49), .CDN(n15), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(N249), .CP(ClockW), .CDN(
        n40), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(N249), .CP(ClockW), .CDN(
        n16), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(N249), .CP(n68), .CDN(n38), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(N249), .CP(n69), .CDN(n108), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(N249), .CP(n43), .CDN(n22), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(N249), .CP(ClockW), .CDN(n11), .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(N249), .CP(n60), .CDN(n27), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(N249), .CP(n65), .CDN(n14), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(N249), .CP(n58), .CDN(n20), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(N249), .CP(n65), .CDN(n36), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(N249), .CP(n55), .CDN(n34), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(N249), .CP(n59), .CDN(n7), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(N249), .CP(n64), .CDN(n30), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(N249), .CP(n66), .CDN(n31), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(N249), .CP(n70), .CDN(n32), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(N150), .CP(n64), .CDN(n36), .Q(
        \Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(N150), .CP(n67), .CDN(n37), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(N150), .CP(n56), .CDN(n10), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(N150), .CP(n45), .CDN(n11), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(N150), .CP(n42), .CDN(n24), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(N150), .CP(n67), .CDN(n40), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(N150), .CP(n52), .CDN(n38), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(N150), .CP(n60), .CDN(n17), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(N150), .CP(n41), .CDN(n35), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(N150), .CP(n57), .CDN(n30), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(N150), .CP(n69), .CDN(n108), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(N150), .CP(n66), .CDN(n34), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(N150), .CP(n62), .CDN(n27), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(N150), .CP(n60), .CDN(n32), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(N150), .CP(n58), .CDN(n33), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(N150), .CP(n55), .CDN(n13), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(N150), .CP(n61), .CDN(n31), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(N150), .CP(n69), .CDN(n40), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(N150), .CP(n58), .CDN(n29), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(N150), .CP(n67), .CDN(n37), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(N150), .CP(n65), .CDN(n9), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(N150), .CP(n70), .CDN(n34), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(N150), .CP(n62), .CDN(n16), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(N150), .CP(n50), .CDN(n29), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(N150), .CP(n57), .CDN(n32), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(N150), .CP(n51), .CDN(n37), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(N150), .CP(n53), .CDN(n26), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(N150), .CP(n67), .CDN(n32), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(N150), .CP(n70), .CDN(n39), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(N150), .CP(n61), .CDN(n40), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(N150), .CP(n43), .CDN(n35), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(N150), .CP(n46), .CDN(n23), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(N85), .E(N1173), .CP(n49), .CDN(n11), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(N1173), .CP(n49), .CDN(
        n11), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(N1173), .CP(n48), .CDN(
        n11), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(N1173), .CP(n48), .CDN(
        n22), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(N1173), .CP(n48), .CDN(
        n21), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(N1173), .CP(n48), .CDN(
        n24), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(N1173), .CP(n48), .CDN(
        n23), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(N1173), .CP(n47), .CDN(
        n25), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(N1173), .CP(n47), .CDN(
        n34), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(N1173), .CP(n47), .CDN(
        n32), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(N1173), .CP(n47), .CDN(
        n31), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(N1173), .CP(n47), .CDN(n3), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(N1173), .CP(n47), .CDN(
        n39), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(N1173), .CP(n47), .CDN(
        n29), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(N1173), .CP(n47), .CDN(
        n18), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(N1173), .CP(n47), .CDN(n4), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(N1173), .CP(n47), .CDN(n5), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(N1173), .CP(n46), .CDN(n6), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(N1173), .CP(n46), .CDN(n11), 
        .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(N1173), .CP(n46), .CDN(n8), 
        .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(N1173), .CP(n46), .CDN(n7), 
        .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(DataI[6]), .E(N1173), .CP(n46), .CDN(n10), 
        .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(N1173), .CP(n46), .CDN(n9), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(N1173), .CP(n46), .CDN(n28), 
        .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(N1173), .CP(n46), .CDN(n27), 
        .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(N1173), .CP(n46), .CDN(n36), 
        .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(N1173), .CP(n46), .CDN(n39), 
        .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(N1173), .CP(n45), .CDN(n22), 
        .Q(\Storage[31][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n107), .CP(ClockR), .CDN(n3), .Q(Dreadyr) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N51), .E(Read), .CP(ClockR), .CDN(n38), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N52), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N53), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N54), .E(Read), .CP(ClockR), .CDN(n28), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N55), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N56), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N57), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N58), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N59), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N60), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N61), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N62), .E(Read), .CP(ClockR), .CDN(n3), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N63), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N64), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N65), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N66), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N67), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N68), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N69), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N70), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N71), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N72), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N73), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N74), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N75), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N76), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N77), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N78), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N79), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N80), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N81), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N82), .E(Read), .CP(ClockR), .CDN(n28), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N83), .E(Read), .CP(ClockR), .CDN(n28), .Q(n572)
         );
  AN2D1 U3 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  INVD1 U4 ( .I(n2), .ZN(ParityErr) );
  CKAN2D0 U5 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  CKND0 U6 ( .CLK(n572), .CN(n2) );
  NR2D2P5 U7 ( .A1(n535), .A2(n537), .ZN(N876) );
  NR2D2P5 U8 ( .A1(n531), .A2(n566), .ZN(N480) );
  NR2D2P5 U9 ( .A1(n564), .A2(n568), .ZN(N249) );
  NR2D2P5 U10 ( .A1(n532), .A2(n536), .ZN(N1173) );
  NR2D2P5 U11 ( .A1(n535), .A2(n550), .ZN(N843) );
  NR2D2P5 U12 ( .A1(n532), .A2(n533), .ZN(N975) );
  NR2D2P5 U13 ( .A1(n531), .A2(n568), .ZN(N216) );
  NR2D2P5 U14 ( .A1(n535), .A2(n563), .ZN(N810) );
  ND3D1 U15 ( .A1(AddrW[4]), .A2(n565), .A3(Write), .ZN(n535) );
  NR2D2P5 U16 ( .A1(n537), .A2(n566), .ZN(N612) );
  NR2D2P5 U17 ( .A1(n550), .A2(n566), .ZN(N579) );
  ND3D1 U18 ( .A1(AddrW[3]), .A2(n567), .A3(Write), .ZN(n566) );
  NR2D2P5 U19 ( .A1(n536), .A2(n568), .ZN(N381) );
  ND3D1 U20 ( .A1(n565), .A2(n567), .A3(Write), .ZN(n568) );
  NR2D2P5 U21 ( .A1(n532), .A2(n563), .ZN(N1074) );
  NR2D2P5 U22 ( .A1(n532), .A2(n564), .ZN(N1041) );
  ND3D1 U23 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n532) );
  NR2D2P5 U24 ( .A1(n535), .A2(n536), .ZN(N909) );
  NR2D2P5 U25 ( .A1(n533), .A2(n566), .ZN(N447) );
  NR2D2P5 U26 ( .A1(n550), .A2(n568), .ZN(N315) );
  NR2D2P5 U27 ( .A1(n532), .A2(n537), .ZN(N1140) );
  NR2D2P5 U28 ( .A1(n535), .A2(n564), .ZN(N777) );
  NR2D2P5 U29 ( .A1(n533), .A2(n568), .ZN(N183) );
  NR2D2P5 U30 ( .A1(n563), .A2(n566), .ZN(N546) );
  NR2D2P5 U31 ( .A1(n532), .A2(n534), .ZN(N942) );
  ND3D0 U32 ( .A1(n571), .A2(n570), .A3(n569), .ZN(n534) );
  NR2D2P5 U33 ( .A1(n531), .A2(n535), .ZN(N744) );
  NR2D2P5 U34 ( .A1(n536), .A2(n566), .ZN(N645) );
  NR2D2P5 U35 ( .A1(n537), .A2(n568), .ZN(N348) );
  NR2D2P5 U36 ( .A1(n532), .A2(n550), .ZN(N1107) );
  NR2D2P5 U37 ( .A1(n564), .A2(n566), .ZN(N513) );
  NR2D2P5 U38 ( .A1(n563), .A2(n568), .ZN(N282) );
  NR2D2P5 U39 ( .A1(n534), .A2(n535), .ZN(N678) );
  AN2D1 U40 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  NR2D2P5 U41 ( .A1(n531), .A2(n532), .ZN(N999) );
  NR2D2P5 U42 ( .A1(n533), .A2(n535), .ZN(N711) );
  NR2D2P5 U43 ( .A1(n534), .A2(n566), .ZN(N414) );
  NR2D2P5 U44 ( .A1(n534), .A2(n568), .ZN(N150) );
  XOR3D1 U45 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n538), .Z(N85) );
  BUFFD0 U46 ( .I(N44), .Z(n84) );
  BUFFD0 U47 ( .I(N46), .Z(n99) );
  BUFFD0 U48 ( .I(N46), .Z(n98) );
  BUFFD1 U49 ( .I(n64), .Z(n43) );
  BUFFD1 U50 ( .I(n67), .Z(n44) );
  BUFFD1 U51 ( .I(n62), .Z(n41) );
  BUFFD1 U52 ( .I(n70), .Z(n42) );
  BUFFD1 U53 ( .I(n61), .Z(n56) );
  BUFFD1 U54 ( .I(n61), .Z(n57) );
  BUFFD1 U55 ( .I(n60), .Z(n58) );
  BUFFD1 U56 ( .I(n60), .Z(n59) );
  BUFFD1 U57 ( .I(n63), .Z(n53) );
  BUFFD1 U58 ( .I(n62), .Z(n54) );
  BUFFD1 U59 ( .I(n62), .Z(n55) );
  BUFFD1 U60 ( .I(n64), .Z(n50) );
  BUFFD1 U61 ( .I(n64), .Z(n51) );
  BUFFD1 U62 ( .I(n63), .Z(n52) );
  BUFFD1 U63 ( .I(n67), .Z(n45) );
  BUFFD1 U64 ( .I(n66), .Z(n46) );
  BUFFD1 U65 ( .I(n66), .Z(n47) );
  BUFFD1 U66 ( .I(n65), .Z(n48) );
  BUFFD1 U67 ( .I(n65), .Z(n49) );
  BUFFD1 U68 ( .I(n31), .Z(n23) );
  BUFFD1 U69 ( .I(n31), .Z(n24) );
  BUFFD1 U70 ( .I(n30), .Z(n25) );
  BUFFD1 U71 ( .I(n32), .Z(n20) );
  BUFFD1 U72 ( .I(n31), .Z(n21) );
  BUFFD1 U73 ( .I(n31), .Z(n22) );
  BUFFD1 U74 ( .I(n32), .Z(n17) );
  BUFFD1 U75 ( .I(n32), .Z(n18) );
  BUFFD1 U76 ( .I(n32), .Z(n19) );
  BUFFD1 U77 ( .I(n33), .Z(n14) );
  BUFFD1 U78 ( .I(n33), .Z(n15) );
  BUFFD1 U79 ( .I(n33), .Z(n16) );
  BUFFD1 U80 ( .I(n33), .Z(n13) );
  BUFFD1 U81 ( .I(n33), .Z(n12) );
  BUFFD1 U82 ( .I(n40), .Z(n11) );
  BUFFD1 U83 ( .I(n69), .Z(n61) );
  BUFFD1 U84 ( .I(n69), .Z(n60) );
  BUFFD1 U85 ( .I(n69), .Z(n62) );
  BUFFD1 U86 ( .I(n68), .Z(n64) );
  BUFFD1 U87 ( .I(n68), .Z(n63) );
  BUFFD1 U88 ( .I(n61), .Z(n67) );
  BUFFD1 U89 ( .I(n62), .Z(n66) );
  BUFFD1 U90 ( .I(n68), .Z(n65) );
  BUFFD1 U91 ( .I(n38), .Z(n3) );
  BUFFD1 U92 ( .I(n29), .Z(n26) );
  BUFFD1 U93 ( .I(n29), .Z(n27) );
  BUFFD1 U94 ( .I(n34), .Z(n9) );
  BUFFD1 U95 ( .I(n34), .Z(n10) );
  BUFFD1 U96 ( .I(n37), .Z(n6) );
  BUFFD1 U97 ( .I(n34), .Z(n7) );
  BUFFD1 U98 ( .I(n34), .Z(n8) );
  BUFFD1 U99 ( .I(n30), .Z(n5) );
  BUFFD1 U100 ( .I(n35), .Z(n4) );
  BUFFD1 U101 ( .I(n29), .Z(n28) );
  BUFFD1 U102 ( .I(n82), .Z(n76) );
  BUFFD1 U103 ( .I(n71), .Z(n77) );
  BUFFD1 U104 ( .I(n84), .Z(n78) );
  BUFFD1 U105 ( .I(n83), .Z(n73) );
  BUFFD1 U106 ( .I(N44), .Z(n72) );
  BUFFD1 U107 ( .I(n84), .Z(n71) );
  BUFFD1 U108 ( .I(n82), .Z(n75) );
  BUFFD1 U109 ( .I(n83), .Z(n74) );
  BUFFD1 U110 ( .I(n92), .Z(n85) );
  BUFFD1 U111 ( .I(n91), .Z(n87) );
  BUFFD1 U112 ( .I(n92), .Z(n86) );
  BUFFD1 U113 ( .I(n90), .Z(n89) );
  BUFFD1 U114 ( .I(n91), .Z(n88) );
  BUFFD1 U115 ( .I(n70), .Z(n69) );
  BUFFD1 U116 ( .I(n70), .Z(n68) );
  BUFFD1 U117 ( .I(n37), .Z(n30) );
  BUFFD1 U118 ( .I(n37), .Z(n31) );
  BUFFD1 U119 ( .I(n36), .Z(n32) );
  BUFFD1 U120 ( .I(n36), .Z(n33) );
  BUFFD1 U121 ( .I(n81), .Z(n79) );
  BUFFD1 U122 ( .I(n99), .Z(n95) );
  BUFFD1 U123 ( .I(n99), .Z(n94) );
  BUFFD1 U124 ( .I(n98), .Z(n97) );
  BUFFD1 U125 ( .I(n98), .Z(n96) );
  BUFFD1 U126 ( .I(n81), .Z(n80) );
  BUFFD1 U127 ( .I(n87), .Z(n90) );
  BUFFD1 U128 ( .I(n93), .Z(n91) );
  BUFFD1 U129 ( .I(n93), .Z(n92) );
  BUFFD1 U130 ( .I(ClockW), .Z(n70) );
  BUFFD1 U131 ( .I(n39), .Z(n37) );
  BUFFD1 U132 ( .I(n39), .Z(n36) );
  BUFFD1 U133 ( .I(n84), .Z(n82) );
  BUFFD1 U134 ( .I(n84), .Z(n83) );
  BUFFD1 U135 ( .I(n35), .Z(n34) );
  BUFFD1 U136 ( .I(n38), .Z(n29) );
  BUFFD1 U137 ( .I(n39), .Z(n38) );
  BUFFD1 U138 ( .I(N45), .Z(n93) );
  BUFFD1 U139 ( .I(n108), .Z(n39) );
  BUFFD1 U140 ( .I(n40), .Z(n35) );
  BUFFD1 U141 ( .I(n108), .Z(n40) );
  BUFFD1 U142 ( .I(n71), .Z(n81) );
  MUX4ND0 U143 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n74), .S1(n92), .ZN(
        n521) );
  MUX4ND0 U144 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n76), .S1(N45), .ZN(n118) );
  MUX4ND0 U145 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n76), .S1(n86), .ZN(n131) );
  MUX4ND0 U146 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n76), .S1(n93), .ZN(n144) );
  MUX4ND0 U147 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n76), .S1(n91), .ZN(n157) );
  MUX4ND0 U148 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n76), .S1(n92), .ZN(n170) );
  MUX4ND0 U149 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n76), .S1(N45), .ZN(n183) );
  MUX4ND0 U150 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n76), .S1(n87), .ZN(n196) );
  MUX4ND0 U151 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n76), .S1(n88), .ZN(n209) );
  MUX4ND0 U152 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n76), .S1(n89), .ZN(n222) );
  MUX4ND0 U153 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n75), .S1(n88), .ZN(
        n235) );
  MUX4ND0 U154 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n75), .S1(n86), .ZN(
        n248) );
  MUX4ND0 U155 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n75), .S1(n85), .ZN(
        n261) );
  MUX4ND0 U156 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n75), .S1(n92), .ZN(
        n274) );
  MUX4ND0 U157 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n75), .S1(n91), .ZN(
        n287) );
  MUX4ND0 U158 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n75), .S1(n93), .ZN(
        n300) );
  MUX4ND0 U159 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n75), .S1(n93), .ZN(
        n313) );
  MUX4ND0 U160 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n75), .S1(n88), .ZN(
        n326) );
  MUX4ND0 U161 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n75), .S1(n90), .ZN(
        n339) );
  MUX4ND0 U162 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n75), .S1(n90), .ZN(
        n352) );
  MUX4ND0 U163 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n75), .S1(n93), .ZN(
        n365) );
  MUX4ND0 U164 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n75), .S1(N45), .ZN(
        n378) );
  MUX4ND0 U165 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n74), .S1(n89), .ZN(
        n391) );
  MUX4ND0 U166 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n74), .S1(n88), .ZN(
        n404) );
  MUX4ND0 U167 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n74), .S1(n89), .ZN(
        n417) );
  MUX4ND0 U168 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n74), .S1(n86), .ZN(
        n430) );
  MUX4ND0 U169 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n74), .S1(n90), .ZN(
        n443) );
  MUX4ND0 U170 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n74), .S1(n87), .ZN(
        n456) );
  MUX4ND0 U171 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n74), .S1(n86), .ZN(
        n469) );
  MUX4ND0 U172 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n74), .S1(n91), .ZN(n103) );
  MUX4ND0 U173 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n74), .S1(n85), .ZN(
        n482) );
  MUX4ND0 U174 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n74), .S1(n87), .ZN(
        n495) );
  MUX4ND0 U175 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n74), .S1(n89), .ZN(
        n508) );
  MUX4D0 U176 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n73), .S1(n86), .Z(
        n522) );
  MUX4D0 U177 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n81), .S1(n88), .Z(n104)
         );
  MUX4D0 U178 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n83), .S1(n87), .Z(n119)
         );
  MUX4D0 U179 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n82), .S1(n86), .Z(n132)
         );
  MUX4D0 U180 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n84), .S1(n85), .Z(n145)
         );
  MUX4D0 U181 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n84), .S1(n91), .Z(n158)
         );
  MUX4D0 U182 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n80), .S1(n90), .Z(n171)
         );
  MUX4D0 U183 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n71), .S1(n88), .Z(n184)
         );
  MUX4D0 U184 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n82), .S1(n89), .Z(n197)
         );
  MUX4D0 U185 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n82), .S1(n89), .Z(n210)
         );
  MUX4D0 U186 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(N44), .S1(n90), .Z(n223)
         );
  MUX4D0 U187 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n77), .S1(n87), .Z(
        n236) );
  MUX4D0 U188 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n81), .S1(n91), .Z(
        n249) );
  MUX4D0 U189 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n74), .S1(n88), .Z(
        n262) );
  MUX4D0 U190 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n84), .S1(n91), .Z(
        n275) );
  MUX4D0 U191 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n74), .S1(n92), .Z(
        n288) );
  MUX4D0 U192 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n73), .S1(n93), .Z(
        n301) );
  MUX4D0 U193 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n73), .S1(n90), .Z(
        n314) );
  MUX4D0 U194 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n76), .S1(n90), .Z(
        n327) );
  MUX4D0 U195 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n74), .S1(n88), .Z(
        n340) );
  MUX4D0 U196 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n73), .S1(n88), .Z(
        n353) );
  MUX4D0 U197 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n74), .S1(n92), .Z(
        n366) );
  MUX4D0 U198 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n80), .S1(n88), .Z(
        n379) );
  MUX4D0 U199 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n83), .S1(n87), .Z(
        n392) );
  MUX4D0 U200 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n73), .S1(n93), .Z(
        n405) );
  MUX4D0 U201 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n72), .S1(n91), .Z(
        n418) );
  MUX4D0 U202 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n72), .S1(n91), .Z(
        n431) );
  MUX4D0 U203 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n71), .S1(n88), .Z(
        n444) );
  MUX4D0 U204 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n71), .S1(n85), .Z(
        n457) );
  MUX4D0 U205 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n77), .S1(n91), .Z(
        n470) );
  MUX4D0 U206 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n79), .S1(n92), .Z(
        n483) );
  MUX4D0 U207 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n79), .S1(n89), .Z(
        n496) );
  MUX4D0 U208 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n76), .S1(n92), .Z(
        n509) );
  MUX4D0 U209 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n73), .S1(n88), .Z(
        n524) );
  MUX4D0 U210 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n82), .S1(n92), .Z(n526)
         );
  MUX4D0 U211 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(N44), .S1(n93), .Z(n106)
         );
  MUX4D0 U212 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n84), .S1(n85), .Z(n110)
         );
  MUX4D0 U213 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n71), .S1(n93), .Z(n121)
         );
  MUX4D0 U214 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n76), .S1(n88), .Z(n123)
         );
  MUX4D0 U215 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n83), .S1(n85), .Z(n134)
         );
  MUX4D0 U216 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n73), .S1(n88), .Z(n136)
         );
  MUX4D0 U217 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n83), .S1(n89), .Z(n147)
         );
  MUX4D0 U218 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n80), .S1(n89), .Z(n149)
         );
  MUX4D0 U219 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n81), .S1(n93), .Z(n160)
         );
  MUX4D0 U220 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n82), .S1(n93), .Z(n162)
         );
  MUX4D0 U221 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n77), .S1(n91), .Z(n173)
         );
  MUX4D0 U222 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n71), .S1(n89), .Z(n175)
         );
  MUX4D0 U223 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n82), .S1(n93), .Z(n186)
         );
  MUX4D0 U224 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n72), .S1(n93), .Z(n188)
         );
  MUX4D0 U225 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n83), .S1(n89), .Z(n199)
         );
  MUX4D0 U226 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n83), .S1(n89), .Z(n201)
         );
  MUX4D0 U227 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n72), .S1(n89), .Z(n212)
         );
  MUX4D0 U228 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n83), .S1(n89), .Z(n214)
         );
  MUX4D0 U229 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n75), .S1(n92), .Z(n225)
         );
  MUX4D0 U230 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n80), .S1(n91), .Z(n227)
         );
  MUX4D0 U231 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n80), .S1(n91), .Z(
        n238) );
  MUX4D0 U232 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n81), .S1(n87), .Z(n240)
         );
  MUX4D0 U233 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n72), .S1(n93), .Z(
        n251) );
  MUX4D0 U234 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(N44), .S1(n85), .Z(n253)
         );
  MUX4D0 U235 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n82), .S1(n87), .Z(
        n264) );
  MUX4D0 U236 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n81), .S1(n89), .Z(n266)
         );
  MUX4D0 U237 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n77), .S1(n90), .Z(
        n277) );
  MUX4D0 U238 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n82), .S1(n86), .Z(n279)
         );
  MUX4D0 U239 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(N44), .S1(n92), .Z(
        n290) );
  MUX4D0 U240 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n73), .S1(n91), .Z(n292)
         );
  MUX4D0 U241 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n73), .S1(n87), .Z(
        n303) );
  MUX4D0 U242 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n73), .S1(n92), .Z(n305)
         );
  MUX4D0 U243 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n73), .S1(n86), .Z(
        n316) );
  MUX4D0 U244 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n74), .S1(n92), .Z(n318)
         );
  MUX4D0 U245 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n73), .S1(N45), .Z(
        n329) );
  MUX4D0 U246 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n75), .S1(n90), .Z(n331)
         );
  MUX4D0 U247 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n76), .S1(n88), .Z(
        n342) );
  MUX4D0 U248 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n80), .S1(n91), .Z(n344)
         );
  MUX4D0 U249 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n79), .S1(n88), .Z(
        n355) );
  MUX4D0 U250 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n82), .S1(n90), .Z(n357)
         );
  MUX4D0 U251 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n75), .S1(n88), .Z(
        n368) );
  MUX4D0 U252 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(N44), .S1(n88), .Z(n370)
         );
  MUX4D0 U253 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n83), .S1(n93), .Z(
        n381) );
  MUX4D0 U254 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n82), .S1(n86), .Z(n383)
         );
  MUX4D0 U255 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n72), .S1(n92), .Z(
        n394) );
  MUX4D0 U256 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n81), .S1(n87), .Z(n396)
         );
  MUX4D0 U257 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n80), .S1(n85), .Z(
        n407) );
  MUX4D0 U258 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(N44), .S1(N45), .Z(n409)
         );
  MUX4D0 U259 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n72), .S1(n90), .Z(
        n420) );
  MUX4D0 U260 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n72), .S1(n86), .Z(n422)
         );
  MUX4D0 U261 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n72), .S1(N45), .Z(
        n433) );
  MUX4D0 U262 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n71), .S1(n90), .Z(n435)
         );
  MUX4D0 U263 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n71), .S1(n91), .Z(
        n446) );
  MUX4D0 U264 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n71), .S1(n92), .Z(n448)
         );
  MUX4D0 U265 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n71), .S1(N45), .Z(
        n459) );
  MUX4D0 U266 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n78), .S1(n93), .Z(n461)
         );
  MUX4D0 U267 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n82), .S1(n86), .Z(
        n472) );
  MUX4D0 U268 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n81), .S1(N45), .Z(n474)
         );
  MUX4D0 U269 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n78), .S1(n89), .Z(
        n485) );
  MUX4D0 U270 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n82), .S1(n93), .Z(n487)
         );
  MUX4D0 U271 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n83), .S1(n90), .Z(
        n498) );
  MUX4D0 U272 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n81), .S1(n92), .Z(n500)
         );
  MUX4D0 U273 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n80), .S1(n88), .Z(
        n511) );
  MUX4D0 U274 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n72), .S1(n90), .Z(n513)
         );
  MUX4D0 U275 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n75), .S1(N45), .Z(
        n523) );
  MUX4D0 U276 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(N44), .S1(n93), .Z(n105)
         );
  MUX4D0 U277 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n81), .S1(n85), .Z(n120)
         );
  MUX4D0 U278 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n75), .S1(n88), .Z(n133)
         );
  MUX4D0 U279 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n84), .S1(n92), .Z(n146)
         );
  MUX4D0 U280 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n73), .S1(n91), .Z(n159)
         );
  MUX4D0 U281 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n76), .S1(n91), .Z(n172)
         );
  MUX4D0 U282 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n81), .S1(n93), .Z(n185)
         );
  MUX4D0 U283 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n75), .S1(n89), .Z(n198)
         );
  MUX4D0 U284 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n83), .S1(n89), .Z(n211)
         );
  MUX4D0 U285 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(N44), .S1(n89), .Z(n224)
         );
  MUX4D0 U286 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n81), .S1(n88), .Z(
        n237) );
  MUX4D0 U287 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n78), .S1(n86), .Z(
        n250) );
  MUX4D0 U288 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n83), .S1(n93), .Z(
        n263) );
  MUX4D0 U289 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n82), .S1(n90), .Z(
        n276) );
  MUX4D0 U290 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n82), .S1(n90), .Z(
        n289) );
  MUX4D0 U291 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n73), .S1(n90), .Z(
        n302) );
  MUX4D0 U292 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n73), .S1(n87), .Z(
        n315) );
  MUX4D0 U293 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n73), .S1(n90), .Z(
        n328) );
  MUX4D0 U294 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n74), .S1(n85), .Z(
        n341) );
  MUX4D0 U295 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n81), .S1(n90), .Z(
        n354) );
  MUX4D0 U296 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n83), .S1(n88), .Z(
        n367) );
  MUX4D0 U297 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n78), .S1(n93), .Z(
        n380) );
  MUX4D0 U298 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n83), .S1(n85), .Z(
        n393) );
  MUX4D0 U299 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n71), .S1(n86), .Z(
        n406) );
  MUX4D0 U300 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n72), .S1(n90), .Z(
        n419) );
  MUX4D0 U301 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n72), .S1(n92), .Z(
        n432) );
  MUX4D0 U302 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n71), .S1(n91), .Z(
        n445) );
  MUX4D0 U303 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n71), .S1(n88), .Z(
        n458) );
  MUX4D0 U304 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n83), .S1(N45), .Z(
        n471) );
  MUX4D0 U305 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n83), .S1(n93), .Z(
        n484) );
  MUX4D0 U306 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n81), .S1(n86), .Z(
        n497) );
  MUX4D0 U307 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n72), .S1(n91), .Z(
        n510) );
  MUX4D0 U308 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n72), .S1(n87), .Z(
        n525) );
  MUX4D0 U309 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n71), .S1(n93), .Z(n527)
         );
  MUX4D0 U310 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n71), .S1(n91), .Z(n109)
         );
  MUX4D0 U311 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n81), .S1(n87), .Z(n111)
         );
  MUX4D0 U312 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n78), .S1(n89), .Z(n122)
         );
  MUX4D0 U313 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n76), .S1(n89), .Z(n124)
         );
  MUX4D0 U314 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n81), .S1(n89), .Z(n135)
         );
  MUX4D0 U315 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n83), .S1(n91), .Z(n137)
         );
  MUX4D0 U316 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n83), .S1(n92), .Z(n148)
         );
  MUX4D0 U317 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(N44), .S1(n90), .Z(n150)
         );
  MUX4D0 U318 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n73), .S1(n85), .Z(n161)
         );
  MUX4D0 U319 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n81), .S1(n91), .Z(n163)
         );
  MUX4D0 U320 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n75), .S1(n85), .Z(n174)
         );
  MUX4D0 U321 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n78), .S1(n89), .Z(n176)
         );
  MUX4D0 U322 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n79), .S1(n90), .Z(n187)
         );
  MUX4D0 U323 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n78), .S1(n93), .Z(n189)
         );
  MUX4D0 U324 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n84), .S1(n89), .Z(n200)
         );
  MUX4D0 U325 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n82), .S1(n89), .Z(n202)
         );
  MUX4D0 U326 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n83), .S1(n89), .Z(n213)
         );
  MUX4D0 U327 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n75), .S1(n92), .Z(n215)
         );
  MUX4D0 U328 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n79), .S1(n87), .Z(n226)
         );
  MUX4D0 U329 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n73), .S1(n90), .Z(n228)
         );
  MUX4D0 U330 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n83), .S1(n87), .Z(
        n239) );
  MUX4D0 U331 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n72), .S1(n91), .Z(n241)
         );
  MUX4D0 U332 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n74), .S1(n92), .Z(
        n252) );
  MUX4D0 U333 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n72), .S1(n90), .Z(n254)
         );
  MUX4D0 U334 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n77), .S1(n85), .Z(
        n265) );
  MUX4D0 U335 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n81), .S1(n93), .Z(n267)
         );
  MUX4D0 U336 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n81), .S1(n91), .Z(
        n278) );
  MUX4D0 U337 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n82), .S1(n92), .Z(n280)
         );
  MUX4D0 U338 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n79), .S1(N45), .Z(
        n291) );
  MUX4D0 U339 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n73), .S1(n88), .Z(n293)
         );
  MUX4D0 U340 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n73), .S1(n89), .Z(
        n304) );
  MUX4D0 U341 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n73), .S1(n85), .Z(n306)
         );
  MUX4D0 U342 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n71), .S1(n93), .Z(
        n317) );
  MUX4D0 U343 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n72), .S1(n90), .Z(n319)
         );
  MUX4D0 U344 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n80), .S1(n88), .Z(
        n330) );
  MUX4D0 U345 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n74), .S1(n92), .Z(n332)
         );
  MUX4D0 U346 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n74), .S1(n88), .Z(
        n343) );
  MUX4D0 U347 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n83), .S1(n88), .Z(n345)
         );
  MUX4D0 U348 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n79), .S1(n88), .Z(
        n356) );
  MUX4D0 U349 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n77), .S1(n89), .Z(n358)
         );
  MUX4D0 U350 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n84), .S1(n89), .Z(
        n369) );
  MUX4D0 U351 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n82), .S1(n93), .Z(n371)
         );
  MUX4D0 U352 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n84), .S1(n91), .Z(
        n382) );
  MUX4D0 U353 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n82), .S1(n92), .Z(n384)
         );
  MUX4D0 U354 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n77), .S1(n88), .Z(
        n395) );
  MUX4D0 U355 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n82), .S1(n90), .Z(n397)
         );
  MUX4D0 U356 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n75), .S1(n91), .Z(
        n408) );
  MUX4D0 U357 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n72), .S1(n92), .Z(n410)
         );
  MUX4D0 U358 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n72), .S1(N45), .Z(
        n421) );
  MUX4D0 U359 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n72), .S1(N45), .Z(n423)
         );
  MUX4D0 U360 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n72), .S1(n92), .Z(
        n434) );
  MUX4D0 U361 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n71), .S1(n90), .Z(n436)
         );
  MUX4D0 U362 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n71), .S1(n86), .Z(
        n447) );
  MUX4D0 U363 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n71), .S1(N45), .Z(n449)
         );
  MUX4D0 U364 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n80), .S1(n85), .Z(
        n460) );
  MUX4D0 U365 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n76), .S1(n91), .Z(n462)
         );
  MUX4D0 U366 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n78), .S1(n92), .Z(
        n473) );
  MUX4D0 U367 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n82), .S1(n92), .Z(n475)
         );
  MUX4D0 U368 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n80), .S1(n93), .Z(
        n486) );
  MUX4D0 U369 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n76), .S1(n92), .Z(n488)
         );
  MUX4D0 U370 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n80), .S1(n91), .Z(
        n499) );
  MUX4D0 U371 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n71), .S1(n86), .Z(n501)
         );
  MUX4D0 U372 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n71), .S1(n90), .Z(
        n512) );
  MUX4D0 U373 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n81), .S1(n93), .Z(n514)
         );
  MUX3ND0 U374 ( .I0(n101), .I1(n102), .I2(n103), .S0(n85), .S1(n94), .ZN(n100) );
  MUX3ND0 U375 ( .I0(n112), .I1(n113), .I2(n114), .S0(N47), .S1(N48), .ZN(N82)
         );
  MUX3ND0 U376 ( .I0(n116), .I1(n117), .I2(n118), .S0(n85), .S1(n99), .ZN(n115) );
  MUX3ND0 U377 ( .I0(n125), .I1(n126), .I2(n127), .S0(N47), .S1(N48), .ZN(N81)
         );
  MUX3ND0 U378 ( .I0(n129), .I1(n130), .I2(n131), .S0(n85), .S1(n94), .ZN(n128) );
  MUX3ND0 U379 ( .I0(n138), .I1(n139), .I2(n140), .S0(N47), .S1(N48), .ZN(N80)
         );
  MUX3ND0 U380 ( .I0(n142), .I1(n143), .I2(n144), .S0(n86), .S1(n98), .ZN(n141) );
  MUX3ND0 U381 ( .I0(n151), .I1(n152), .I2(n153), .S0(N47), .S1(N48), .ZN(N79)
         );
  MUX3ND0 U382 ( .I0(n155), .I1(n156), .I2(n157), .S0(n85), .S1(n96), .ZN(n154) );
  MUX3ND0 U383 ( .I0(n164), .I1(n165), .I2(n166), .S0(N47), .S1(N48), .ZN(N78)
         );
  MUX3ND0 U384 ( .I0(n168), .I1(n169), .I2(n170), .S0(n87), .S1(N46), .ZN(n167) );
  MUX3ND0 U385 ( .I0(n177), .I1(n178), .I2(n179), .S0(N47), .S1(N48), .ZN(N77)
         );
  MUX3ND0 U386 ( .I0(n181), .I1(n182), .I2(n183), .S0(n86), .S1(n99), .ZN(n180) );
  MUX3ND0 U387 ( .I0(n190), .I1(n191), .I2(n192), .S0(N47), .S1(N48), .ZN(N76)
         );
  MUX3ND0 U388 ( .I0(n194), .I1(n195), .I2(n196), .S0(n87), .S1(n97), .ZN(n193) );
  MUX3ND0 U389 ( .I0(n203), .I1(n204), .I2(n205), .S0(N47), .S1(N48), .ZN(N75)
         );
  MUX3ND0 U390 ( .I0(n207), .I1(n208), .I2(n209), .S0(n87), .S1(n98), .ZN(n206) );
  MUX3ND0 U391 ( .I0(n216), .I1(n217), .I2(n218), .S0(N47), .S1(N48), .ZN(N74)
         );
  MUX3ND0 U392 ( .I0(n220), .I1(n221), .I2(n222), .S0(n87), .S1(N46), .ZN(n219) );
  MUX3ND0 U393 ( .I0(n229), .I1(n230), .I2(n231), .S0(N47), .S1(N48), .ZN(N73)
         );
  MUX3ND0 U394 ( .I0(n233), .I1(n234), .I2(n235), .S0(n85), .S1(N46), .ZN(n232) );
  MUX3ND0 U395 ( .I0(n242), .I1(n243), .I2(n244), .S0(N47), .S1(N48), .ZN(N72)
         );
  MUX3ND0 U396 ( .I0(n246), .I1(n247), .I2(n248), .S0(n87), .S1(n95), .ZN(n245) );
  MUX3ND0 U397 ( .I0(n255), .I1(n256), .I2(n257), .S0(N47), .S1(N48), .ZN(N71)
         );
  MUX3ND0 U398 ( .I0(n259), .I1(n260), .I2(n261), .S0(n87), .S1(n99), .ZN(n258) );
  MUX3ND0 U399 ( .I0(n268), .I1(n269), .I2(n270), .S0(N47), .S1(N48), .ZN(N70)
         );
  MUX3ND0 U400 ( .I0(n272), .I1(n273), .I2(n274), .S0(n86), .S1(n97), .ZN(n271) );
  MUX3ND0 U401 ( .I0(n281), .I1(n282), .I2(n283), .S0(N47), .S1(N48), .ZN(N69)
         );
  MUX3ND0 U402 ( .I0(n285), .I1(n286), .I2(n287), .S0(n85), .S1(n98), .ZN(n284) );
  MUX3ND0 U403 ( .I0(n294), .I1(n295), .I2(n296), .S0(N47), .S1(N48), .ZN(N68)
         );
  MUX3ND0 U404 ( .I0(n298), .I1(n299), .I2(n300), .S0(n86), .S1(N46), .ZN(n297) );
  MUX3ND0 U405 ( .I0(n307), .I1(n308), .I2(n309), .S0(N47), .S1(N48), .ZN(N67)
         );
  MUX3ND0 U406 ( .I0(n311), .I1(n312), .I2(n313), .S0(n86), .S1(n95), .ZN(n310) );
  MUX3ND0 U407 ( .I0(n320), .I1(n321), .I2(n322), .S0(N47), .S1(N48), .ZN(N66)
         );
  MUX3ND0 U408 ( .I0(n324), .I1(n325), .I2(n326), .S0(n85), .S1(n99), .ZN(n323) );
  MUX3ND0 U409 ( .I0(n333), .I1(n334), .I2(n335), .S0(N47), .S1(N48), .ZN(N65)
         );
  MUX3ND0 U410 ( .I0(n337), .I1(n338), .I2(n339), .S0(n85), .S1(n96), .ZN(n336) );
  MUX3ND0 U411 ( .I0(n346), .I1(n347), .I2(n348), .S0(N47), .S1(N48), .ZN(N64)
         );
  MUX3ND0 U412 ( .I0(n350), .I1(n351), .I2(n352), .S0(n85), .S1(n98), .ZN(n349) );
  MUX3ND0 U413 ( .I0(n359), .I1(n360), .I2(n361), .S0(N47), .S1(N48), .ZN(N63)
         );
  MUX3ND0 U414 ( .I0(n363), .I1(n364), .I2(n365), .S0(n86), .S1(n97), .ZN(n362) );
  MUX3ND0 U415 ( .I0(n372), .I1(n373), .I2(n374), .S0(N47), .S1(N48), .ZN(N62)
         );
  MUX3ND0 U416 ( .I0(n376), .I1(n377), .I2(n378), .S0(n86), .S1(N46), .ZN(n375) );
  MUX3ND0 U417 ( .I0(n385), .I1(n386), .I2(n387), .S0(N47), .S1(N48), .ZN(N61)
         );
  MUX3ND0 U418 ( .I0(n389), .I1(n390), .I2(n391), .S0(n86), .S1(n98), .ZN(n388) );
  MUX3ND0 U419 ( .I0(n398), .I1(n399), .I2(n400), .S0(N47), .S1(N48), .ZN(N60)
         );
  MUX3ND0 U420 ( .I0(n402), .I1(n403), .I2(n404), .S0(n86), .S1(N46), .ZN(n401) );
  MUX3ND0 U421 ( .I0(n411), .I1(n412), .I2(n413), .S0(N47), .S1(N48), .ZN(N59)
         );
  MUX3ND0 U422 ( .I0(n415), .I1(n416), .I2(n417), .S0(n87), .S1(n99), .ZN(n414) );
  MUX3ND0 U423 ( .I0(n424), .I1(n425), .I2(n426), .S0(N47), .S1(N48), .ZN(N58)
         );
  MUX3ND0 U424 ( .I0(n428), .I1(n429), .I2(n430), .S0(n87), .S1(n99), .ZN(n427) );
  MUX3ND0 U425 ( .I0(n437), .I1(n438), .I2(n439), .S0(N47), .S1(N48), .ZN(N57)
         );
  MUX3ND0 U426 ( .I0(n441), .I1(n442), .I2(n443), .S0(n87), .S1(n95), .ZN(n440) );
  MUX3ND0 U427 ( .I0(n450), .I1(n451), .I2(n452), .S0(N47), .S1(N48), .ZN(N56)
         );
  MUX3ND0 U428 ( .I0(n454), .I1(n455), .I2(n456), .S0(n87), .S1(n98), .ZN(n453) );
  MUX3ND0 U429 ( .I0(n463), .I1(n464), .I2(n465), .S0(N47), .S1(N48), .ZN(N55)
         );
  MUX3ND0 U430 ( .I0(n467), .I1(n468), .I2(n469), .S0(n85), .S1(n99), .ZN(n466) );
  MUX3ND0 U431 ( .I0(n476), .I1(n477), .I2(n478), .S0(N47), .S1(N48), .ZN(N54)
         );
  MUX3ND0 U432 ( .I0(n480), .I1(n481), .I2(n482), .S0(n87), .S1(n99), .ZN(n479) );
  MUX3ND0 U433 ( .I0(n489), .I1(n490), .I2(n491), .S0(N47), .S1(N48), .ZN(N53)
         );
  MUX3ND0 U434 ( .I0(n493), .I1(n494), .I2(n495), .S0(n86), .S1(n98), .ZN(n492) );
  MUX3ND0 U435 ( .I0(n502), .I1(n503), .I2(n504), .S0(N47), .S1(N48), .ZN(N52)
         );
  MUX3ND0 U436 ( .I0(n506), .I1(n507), .I2(n508), .S0(n86), .S1(n96), .ZN(n505) );
  MUX3ND0 U437 ( .I0(n515), .I1(n516), .I2(n517), .S0(N47), .S1(N48), .ZN(N51)
         );
  MUX3ND0 U438 ( .I0(n519), .I1(n520), .I2(n521), .S0(n85), .S1(n95), .ZN(n518) );
  MUX3ND0 U439 ( .I0(n528), .I1(n529), .I2(n530), .S0(N47), .S1(N48), .ZN(N50)
         );
  MUX2ND0 U440 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n80), .ZN(
        n102) );
  MUX2ND0 U441 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n80), .ZN(
        n101) );
  MUX3ND0 U442 ( .I0(n105), .I1(n104), .I2(n100), .S0(n95), .S1(N47), .ZN(n114) );
  MUX2ND0 U443 ( .I0(n109), .I1(n106), .S(N46), .ZN(n113) );
  MUX2ND0 U444 ( .I0(n111), .I1(n110), .S(n99), .ZN(n112) );
  MUX2ND0 U445 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n80), .ZN(
        n117) );
  MUX2ND0 U446 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n79), .ZN(
        n116) );
  MUX3ND0 U447 ( .I0(n120), .I1(n119), .I2(n115), .S0(N46), .S1(N47), .ZN(n127) );
  MUX2ND0 U448 ( .I0(n122), .I1(n121), .S(n95), .ZN(n126) );
  MUX2ND0 U449 ( .I0(n124), .I1(n123), .S(n94), .ZN(n125) );
  MUX2ND0 U450 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n79), .ZN(
        n130) );
  MUX2ND0 U451 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n79), .ZN(
        n129) );
  MUX3ND0 U452 ( .I0(n133), .I1(n132), .I2(n128), .S0(n95), .S1(N47), .ZN(n140) );
  MUX2ND0 U453 ( .I0(n135), .I1(n134), .S(n98), .ZN(n139) );
  MUX2ND0 U454 ( .I0(n137), .I1(n136), .S(n97), .ZN(n138) );
  MUX2ND0 U455 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n79), .ZN(
        n143) );
  MUX2ND0 U456 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n78), .ZN(
        n142) );
  MUX3ND0 U457 ( .I0(n146), .I1(n145), .I2(n141), .S0(n95), .S1(N47), .ZN(n153) );
  MUX2ND0 U458 ( .I0(n148), .I1(n147), .S(N46), .ZN(n152) );
  MUX2ND0 U459 ( .I0(n150), .I1(n149), .S(n99), .ZN(n151) );
  MUX2ND0 U460 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n78), .ZN(
        n156) );
  MUX2ND0 U461 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n78), .ZN(
        n155) );
  MUX3ND0 U462 ( .I0(n159), .I1(n158), .I2(n154), .S0(n95), .S1(N47), .ZN(n166) );
  MUX2ND0 U463 ( .I0(n161), .I1(n160), .S(n98), .ZN(n165) );
  MUX2ND0 U464 ( .I0(n163), .I1(n162), .S(N46), .ZN(n164) );
  MUX2ND0 U465 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n78), .ZN(
        n169) );
  MUX2ND0 U466 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n77), .ZN(
        n168) );
  MUX3ND0 U467 ( .I0(n172), .I1(n171), .I2(n167), .S0(n98), .S1(N47), .ZN(n179) );
  MUX2ND0 U468 ( .I0(n174), .I1(n173), .S(n98), .ZN(n178) );
  MUX2ND0 U469 ( .I0(n176), .I1(n175), .S(n97), .ZN(n177) );
  MUX2ND0 U470 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n77), .ZN(
        n182) );
  MUX2ND0 U471 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n77), .ZN(
        n181) );
  MUX3ND0 U472 ( .I0(n185), .I1(n184), .I2(n180), .S0(n95), .S1(N47), .ZN(n192) );
  MUX2ND0 U473 ( .I0(n187), .I1(n186), .S(n97), .ZN(n191) );
  MUX2ND0 U474 ( .I0(n189), .I1(n188), .S(n97), .ZN(n190) );
  MUX2ND0 U475 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n77), .ZN(
        n195) );
  MUX2ND0 U476 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n76), .ZN(
        n194) );
  MUX3ND0 U477 ( .I0(n198), .I1(n197), .I2(n193), .S0(n96), .S1(N47), .ZN(n205) );
  MUX2ND0 U478 ( .I0(n200), .I1(n199), .S(n97), .ZN(n204) );
  MUX2ND0 U479 ( .I0(n202), .I1(n201), .S(n97), .ZN(n203) );
  MUX2ND0 U480 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n76), .ZN(
        n208) );
  MUX2ND0 U481 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n76), .ZN(
        n207) );
  MUX3ND0 U482 ( .I0(n211), .I1(n210), .I2(n206), .S0(n94), .S1(N47), .ZN(n218) );
  MUX2ND0 U483 ( .I0(n213), .I1(n212), .S(n97), .ZN(n217) );
  MUX2ND0 U484 ( .I0(n215), .I1(n214), .S(n97), .ZN(n216) );
  MUX2ND0 U485 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n77), .ZN(
        n221) );
  MUX2ND0 U486 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n76), .ZN(
        n220) );
  MUX3ND0 U487 ( .I0(n224), .I1(n223), .I2(n219), .S0(N46), .S1(N47), .ZN(n231) );
  MUX2ND0 U488 ( .I0(n226), .I1(n225), .S(n97), .ZN(n230) );
  MUX2ND0 U489 ( .I0(n228), .I1(n227), .S(n97), .ZN(n229) );
  MUX2ND0 U490 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n76), .ZN(
        n234) );
  MUX2ND0 U491 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n77), .ZN(
        n233) );
  MUX3ND0 U492 ( .I0(n237), .I1(n236), .I2(n232), .S0(n95), .S1(N47), .ZN(n244) );
  MUX2ND0 U493 ( .I0(n239), .I1(n238), .S(n97), .ZN(n243) );
  MUX2ND0 U494 ( .I0(n241), .I1(n240), .S(n97), .ZN(n242) );
  MUX2ND0 U495 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n77), .ZN(
        n247) );
  MUX2ND0 U496 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n77), .ZN(
        n246) );
  MUX3ND0 U497 ( .I0(n250), .I1(n249), .I2(n245), .S0(n96), .S1(N47), .ZN(n257) );
  MUX2ND0 U498 ( .I0(n252), .I1(n251), .S(n97), .ZN(n256) );
  MUX2ND0 U499 ( .I0(n254), .I1(n253), .S(n97), .ZN(n255) );
  MUX2ND0 U500 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n77), .ZN(
        n260) );
  MUX2ND0 U501 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n77), .ZN(
        n259) );
  MUX3ND0 U502 ( .I0(n263), .I1(n262), .I2(n258), .S0(n97), .S1(N47), .ZN(n270) );
  MUX2ND0 U503 ( .I0(n265), .I1(n264), .S(n96), .ZN(n269) );
  MUX2ND0 U504 ( .I0(n267), .I1(n266), .S(n95), .ZN(n268) );
  MUX2ND0 U505 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n77), .ZN(
        n273) );
  MUX2ND0 U506 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n77), .ZN(
        n272) );
  MUX3ND0 U507 ( .I0(n276), .I1(n275), .I2(n271), .S0(n94), .S1(N47), .ZN(n283) );
  MUX2ND0 U508 ( .I0(n278), .I1(n277), .S(n97), .ZN(n282) );
  MUX2ND0 U509 ( .I0(n280), .I1(n279), .S(n95), .ZN(n281) );
  MUX2ND0 U510 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n77), .ZN(
        n286) );
  MUX2ND0 U511 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n77), .ZN(
        n285) );
  MUX3ND0 U512 ( .I0(n289), .I1(n288), .I2(n284), .S0(n95), .S1(N47), .ZN(n296) );
  MUX2ND0 U513 ( .I0(n291), .I1(n290), .S(n96), .ZN(n295) );
  MUX2ND0 U514 ( .I0(n293), .I1(n292), .S(n96), .ZN(n294) );
  MUX2ND0 U515 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n78), .ZN(
        n299) );
  MUX2ND0 U516 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n77), .ZN(
        n298) );
  MUX3ND0 U517 ( .I0(n302), .I1(n301), .I2(n297), .S0(n97), .S1(N47), .ZN(n309) );
  MUX2ND0 U518 ( .I0(n304), .I1(n303), .S(n94), .ZN(n308) );
  MUX2ND0 U519 ( .I0(n306), .I1(n305), .S(n94), .ZN(n307) );
  MUX2ND0 U520 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n77), .ZN(
        n312) );
  MUX2ND0 U521 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n78), .ZN(
        n311) );
  MUX3ND0 U522 ( .I0(n315), .I1(n314), .I2(n310), .S0(n94), .S1(N47), .ZN(n322) );
  MUX2ND0 U523 ( .I0(n317), .I1(n316), .S(n94), .ZN(n321) );
  MUX2ND0 U524 ( .I0(n319), .I1(n318), .S(n96), .ZN(n320) );
  MUX2ND0 U525 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n78), .ZN(
        n325) );
  MUX2ND0 U526 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n78), .ZN(
        n324) );
  MUX3ND0 U527 ( .I0(n328), .I1(n327), .I2(n323), .S0(n94), .S1(N47), .ZN(n335) );
  MUX2ND0 U528 ( .I0(n330), .I1(n329), .S(n95), .ZN(n334) );
  MUX2ND0 U529 ( .I0(n332), .I1(n331), .S(n96), .ZN(n333) );
  MUX2ND0 U530 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n78), .ZN(
        n338) );
  MUX2ND0 U531 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n78), .ZN(
        n337) );
  MUX3ND0 U532 ( .I0(n341), .I1(n340), .I2(n336), .S0(n95), .S1(N47), .ZN(n348) );
  MUX2ND0 U533 ( .I0(n343), .I1(n342), .S(n94), .ZN(n347) );
  MUX2ND0 U534 ( .I0(n345), .I1(n344), .S(n94), .ZN(n346) );
  MUX2ND0 U535 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n78), .ZN(
        n351) );
  MUX2ND0 U536 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n78), .ZN(
        n350) );
  MUX3ND0 U537 ( .I0(n354), .I1(n353), .I2(n349), .S0(n99), .S1(N47), .ZN(n361) );
  MUX2ND0 U538 ( .I0(n356), .I1(n355), .S(n95), .ZN(n360) );
  MUX2ND0 U539 ( .I0(n358), .I1(n357), .S(n95), .ZN(n359) );
  MUX2ND0 U540 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n78), .ZN(
        n364) );
  MUX2ND0 U541 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n78), .ZN(
        n363) );
  MUX3ND0 U542 ( .I0(n367), .I1(n366), .I2(n362), .S0(n94), .S1(N47), .ZN(n374) );
  MUX2ND0 U543 ( .I0(n369), .I1(n368), .S(n96), .ZN(n373) );
  MUX2ND0 U544 ( .I0(n371), .I1(n370), .S(n97), .ZN(n372) );
  MUX2ND0 U545 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n78), .ZN(
        n377) );
  MUX2ND0 U546 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n78), .ZN(
        n376) );
  MUX3ND0 U547 ( .I0(n380), .I1(n379), .I2(n375), .S0(n94), .S1(N47), .ZN(n387) );
  MUX2ND0 U548 ( .I0(n382), .I1(n381), .S(n97), .ZN(n386) );
  MUX2ND0 U549 ( .I0(n384), .I1(n383), .S(n95), .ZN(n385) );
  MUX2ND0 U550 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n78), .ZN(
        n390) );
  MUX2ND0 U551 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n79), .ZN(
        n389) );
  MUX3ND0 U552 ( .I0(n393), .I1(n392), .I2(n388), .S0(n95), .S1(N47), .ZN(n400) );
  MUX2ND0 U553 ( .I0(n395), .I1(n394), .S(n96), .ZN(n399) );
  MUX2ND0 U554 ( .I0(n397), .I1(n396), .S(n94), .ZN(n398) );
  MUX2ND0 U555 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n79), .ZN(
        n403) );
  MUX2ND0 U556 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n79), .ZN(
        n402) );
  MUX3ND0 U557 ( .I0(n406), .I1(n405), .I2(n401), .S0(n95), .S1(N47), .ZN(n413) );
  MUX2ND0 U558 ( .I0(n408), .I1(n407), .S(n95), .ZN(n412) );
  MUX2ND0 U559 ( .I0(n410), .I1(n409), .S(n96), .ZN(n411) );
  MUX2ND0 U560 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n79), .ZN(
        n416) );
  MUX2ND0 U561 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n79), .ZN(
        n415) );
  MUX3ND0 U562 ( .I0(n419), .I1(n418), .I2(n414), .S0(n95), .S1(N47), .ZN(n426) );
  MUX2ND0 U563 ( .I0(n421), .I1(n420), .S(n96), .ZN(n425) );
  MUX2ND0 U564 ( .I0(n423), .I1(n422), .S(n94), .ZN(n424) );
  MUX2ND0 U565 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n79), .ZN(
        n429) );
  MUX2ND0 U566 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n79), .ZN(
        n428) );
  MUX3ND0 U567 ( .I0(n432), .I1(n431), .I2(n427), .S0(n95), .S1(N47), .ZN(n439) );
  MUX2ND0 U568 ( .I0(n434), .I1(n433), .S(n96), .ZN(n438) );
  MUX2ND0 U569 ( .I0(n436), .I1(n435), .S(n96), .ZN(n437) );
  MUX2ND0 U570 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n79), .ZN(
        n442) );
  MUX2ND0 U571 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n79), .ZN(
        n441) );
  MUX3ND0 U572 ( .I0(n445), .I1(n444), .I2(n440), .S0(n94), .S1(N47), .ZN(n452) );
  MUX2ND0 U573 ( .I0(n447), .I1(n446), .S(n96), .ZN(n451) );
  MUX2ND0 U574 ( .I0(n449), .I1(n448), .S(n96), .ZN(n450) );
  MUX2ND0 U575 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n79), .ZN(
        n455) );
  MUX2ND0 U576 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n79), .ZN(
        n454) );
  MUX3ND0 U577 ( .I0(n458), .I1(n457), .I2(n453), .S0(n94), .S1(N47), .ZN(n465) );
  MUX2ND0 U578 ( .I0(n460), .I1(n459), .S(n97), .ZN(n464) );
  MUX2ND0 U579 ( .I0(n462), .I1(n461), .S(n96), .ZN(n463) );
  MUX2ND0 U580 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n79), .ZN(
        n468) );
  MUX2ND0 U581 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n79), .ZN(
        n467) );
  MUX3ND0 U582 ( .I0(n471), .I1(n470), .I2(n466), .S0(n94), .S1(N47), .ZN(n478) );
  MUX2ND0 U583 ( .I0(n473), .I1(n472), .S(n96), .ZN(n477) );
  MUX2ND0 U584 ( .I0(n475), .I1(n474), .S(n94), .ZN(n476) );
  MUX2ND0 U585 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n80), .ZN(
        n481) );
  MUX2ND0 U586 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n80), .ZN(
        n480) );
  MUX3ND0 U587 ( .I0(n484), .I1(n483), .I2(n479), .S0(n94), .S1(N47), .ZN(n491) );
  MUX2ND0 U588 ( .I0(n486), .I1(n485), .S(n97), .ZN(n490) );
  MUX2ND0 U589 ( .I0(n488), .I1(n487), .S(n96), .ZN(n489) );
  MUX2ND0 U590 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n80), .ZN(
        n494) );
  MUX2ND0 U591 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n80), .ZN(
        n493) );
  MUX3ND0 U592 ( .I0(n497), .I1(n496), .I2(n492), .S0(n94), .S1(N47), .ZN(n504) );
  MUX2ND0 U593 ( .I0(n499), .I1(n498), .S(n96), .ZN(n503) );
  MUX2ND0 U594 ( .I0(n501), .I1(n500), .S(n96), .ZN(n502) );
  MUX2ND0 U595 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n80), .ZN(
        n507) );
  MUX2ND0 U596 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n80), .ZN(
        n506) );
  MUX3ND0 U597 ( .I0(n510), .I1(n509), .I2(n505), .S0(n94), .S1(N47), .ZN(n517) );
  MUX2ND0 U598 ( .I0(n512), .I1(n511), .S(n95), .ZN(n516) );
  MUX2ND0 U599 ( .I0(n514), .I1(n513), .S(n96), .ZN(n515) );
  MUX2ND0 U600 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n80), .ZN(
        n520) );
  MUX2ND0 U601 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n77), .ZN(
        n519) );
  MUX3ND0 U602 ( .I0(n523), .I1(n522), .I2(n518), .S0(n94), .S1(N47), .ZN(n530) );
  MUX2ND0 U603 ( .I0(n525), .I1(n524), .S(n96), .ZN(n529) );
  MUX2ND0 U604 ( .I0(n527), .I1(n526), .S(n97), .ZN(n528) );
  CKND0 U605 ( .CLK(Reset), .CN(n108) );
  OR2D0 U606 ( .A1(Read), .A2(Dreadyr), .Z(n107) );
  XOR3D0 U607 ( .A1(DataI[0]), .A2(n539), .A3(n540), .Z(n538) );
  XOR3D0 U608 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n541), .Z(n540) );
  XOR3D0 U609 ( .A1(n542), .A2(DataI[3]), .A3(n543), .Z(n541) );
  XOR3D0 U610 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n544), .Z(n543) );
  XOR3D0 U611 ( .A1(n545), .A2(DataI[10]), .A3(n546), .Z(n544) );
  XOR3D0 U612 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n547), .Z(n546) );
  XOR3D0 U613 ( .A1(n548), .A2(DataI[17]), .A3(n549), .Z(n547) );
  XNR4D0 U614 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n549) );
  XOR4D0 U615 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n548) );
  XOR4D0 U616 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n545) );
  XOR4D0 U617 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n542) );
  XNR4D0 U618 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n539) );
  XOR4D0 U619 ( .A1(n551), .A2(N79), .A3(n552), .A4(n553), .Z(N83) );
  XNR4D0 U620 ( .A1(N76), .A2(N75), .A3(N78), .A4(N77), .ZN(n553) );
  XNR3D0 U621 ( .A1(N82), .A2(N81), .A3(N80), .ZN(n552) );
  XOR3D0 U622 ( .A1(N74), .A2(N73), .A3(n554), .Z(n551) );
  XOR3D0 U623 ( .A1(N72), .A2(n555), .A3(n556), .Z(n554) );
  XOR3D0 U624 ( .A1(N67), .A2(N66), .A3(n557), .Z(n556) );
  XOR3D0 U625 ( .A1(n558), .A2(N65), .A3(n559), .Z(n557) );
  XOR3D0 U626 ( .A1(N60), .A2(N59), .A3(n560), .Z(n559) );
  XOR3D0 U627 ( .A1(n561), .A2(N58), .A3(n562), .Z(n560) );
  XNR4D0 U628 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n562) );
  XOR4D0 U629 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n561) );
  XOR4D0 U630 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .Z(n558) );
  XNR4D0 U631 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n555) );
  ND3D0 U632 ( .A1(n569), .A2(n570), .A3(AddrW[1]), .ZN(n531) );
  ND3D0 U633 ( .A1(n571), .A2(n570), .A3(AddrW[0]), .ZN(n533) );
  CKND0 U634 ( .CLK(AddrW[4]), .CN(n567) );
  CKND0 U635 ( .CLK(AddrW[3]), .CN(n565) );
  ND3D0 U636 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n536) );
  ND3D0 U637 ( .A1(AddrW[1]), .A2(n569), .A3(AddrW[2]), .ZN(n537) );
  ND3D0 U638 ( .A1(AddrW[0]), .A2(n571), .A3(AddrW[2]), .ZN(n550) );
  ND3D0 U639 ( .A1(n569), .A2(n571), .A3(AddrW[2]), .ZN(n563) );
  CKND0 U640 ( .CLK(AddrW[1]), .CN(n571) );
  CKND0 U641 ( .CLK(AddrW[0]), .CN(n569) );
  ND3D0 U642 ( .A1(AddrW[1]), .A2(n570), .A3(AddrW[0]), .ZN(n564) );
  CKND0 U643 ( .CLK(AddrW[2]), .CN(n570) );
endmodule


module MemBIST_Top ( Dready, ParityErr, Testing, TestOK, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, DoSelfTest, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, DoSelfTest, Read, Write, Reset;
  output Dready, ParityErr, Testing, TestOK;
  wire   N9, n145, n146, Dreadyw, ClkWw, Readw, ReadCmdBISTw, Writew,
         WriteCmdBISTw, n129, n130, n131, n133, n135, n136, n137, n138, n139,
         n140, n141, n143, n144;
  wire   [31:0] DataOw;
  wire   [31:0] DataIw;
  wire   [31:0] DataOBISTw;
  wire   [4:0] AddrRw;
  wire   [4:0] AddrBISTw;
  wire   [4:0] AddrWw;
  wire   [31:0] DataIBISTw;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10;

  BUFTD1 \DataIBISTw_tri[2]  ( .I(DataOw[2]), .OE(n137), .Z(DataIBISTw[2]) );
  BUFTD1 \DataIBISTw_tri[3]  ( .I(DataOw[3]), .OE(N9), .Z(DataIBISTw[3]) );
  BUFTD1 \DataIBISTw_tri[16]  ( .I(DataOw[16]), .OE(n138), .Z(DataIBISTw[16])
         );
  BUFTD1 \DataIBISTw_tri[17]  ( .I(DataOw[17]), .OE(n138), .Z(DataIBISTw[17])
         );
  BUFTD1 \DataIBISTw_tri[20]  ( .I(DataOw[20]), .OE(n137), .Z(DataIBISTw[20])
         );
  BUFTD1 \DataIBISTw_tri[24]  ( .I(DataOw[24]), .OE(n138), .Z(DataIBISTw[24])
         );
  Mem_AWid5_DWid32 Mem_U1 ( .Dready(Dreadyw), .ParityErr(n146), .DataO(DataOw), 
        .DataI(DataIw), .AddrR({AddrRw[4:3], n130, AddrRw[1], n131}), .AddrW(
        AddrWw), .ClkR(n140), .ClkW(ClkWw), .ChipEna(n139), .Read(Readw), 
        .Write(Writew), .Reset(Reset) );
  BIST_AWid5_DWid32 BIST_U1 ( .DataO({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, DataOBISTw[28:24], 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, DataOBISTw[20:16], SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, DataOBISTw[12:7], 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, DataOBISTw[4:0]}), 
        .Addr(AddrBISTw), .ReadCmd(ReadCmdBISTw), .WriteCmd(WriteCmdBISTw), 
        .Testing(N9), .TestOK(TestOK), .DataI(DataIBISTw), .DoSelfTest(
        DoSelfTest), .ParityErr(n136), .Clk(n140), .Reset(Reset) );
  BUFTD0 \DataIBISTw_tri[4]  ( .I(DataOw[4]), .OE(N9), .Z(DataIBISTw[4]) );
  BUFTD0 \DataIBISTw_tri[9]  ( .I(DataOw[9]), .OE(n138), .Z(DataIBISTw[9]) );
  BUFTD0 \DataIBISTw_tri[0]  ( .I(DataOw[0]), .OE(n137), .Z(DataIBISTw[0]) );
  BUFTD0 \DataIBISTw_tri[28]  ( .I(DataOw[28]), .OE(N9), .Z(DataIBISTw[28]) );
  BUFTD0 \DataIBISTw_tri[8]  ( .I(DataOw[8]), .OE(n137), .Z(DataIBISTw[8]) );
  BUFTD0 \DataIBISTw_tri[25]  ( .I(DataOw[25]), .OE(n138), .Z(DataIBISTw[25])
         );
  BUFTD0 \DataIBISTw_tri[10]  ( .I(DataOw[10]), .OE(n138), .Z(DataIBISTw[10])
         );
  BUFTD0 \DataIBISTw_tri[11]  ( .I(DataOw[11]), .OE(n138), .Z(DataIBISTw[11])
         );
  BUFTD0 \DataIBISTw_tri[18]  ( .I(DataOw[18]), .OE(N9), .Z(DataIBISTw[18]) );
  BUFTD0 \DataIBISTw_tri[26]  ( .I(DataOw[26]), .OE(n138), .Z(DataIBISTw[26])
         );
  BUFTD0 \DataIBISTw_tri[27]  ( .I(DataOw[27]), .OE(N9), .Z(DataIBISTw[27]) );
  BUFTD0 \DataIBISTw_tri[12]  ( .I(DataOw[12]), .OE(n137), .Z(DataIBISTw[12])
         );
  BUFTD0 \DataIBISTw_tri[1]  ( .I(DataOw[1]), .OE(n138), .Z(DataIBISTw[1]) );
  BUFTD0 \DataIBISTw_tri[19]  ( .I(DataOw[19]), .OE(n137), .Z(DataIBISTw[19])
         );
  BUFTD0 \DataIBISTw_tri[21]  ( .I(DataOw[21]), .OE(N9), .Z(DataIBISTw[21]) );
  BUFTD0 \DataIBISTw_tri[5]  ( .I(DataOw[5]), .OE(N9), .Z(DataIBISTw[5]) );
  BUFTD0 \DataIBISTw_tri[7]  ( .I(DataOw[7]), .OE(n138), .Z(DataIBISTw[7]) );
  BUFTD0 \DataIBISTw_tri[29]  ( .I(DataOw[29]), .OE(n137), .Z(DataIBISTw[29])
         );
  BUFTD0 \DataIBISTw_tri[23]  ( .I(DataOw[23]), .OE(N9), .Z(DataIBISTw[23]) );
  BUFTD0 \DataIBISTw_tri[30]  ( .I(DataOw[30]), .OE(n137), .Z(DataIBISTw[30])
         );
  BUFTD0 \DataIBISTw_tri[13]  ( .I(DataOw[13]), .OE(n137), .Z(DataIBISTw[13])
         );
  BUFTD0 \DataIBISTw_tri[15]  ( .I(DataOw[15]), .OE(N9), .Z(DataIBISTw[15]) );
  BUFTD0 \DataIBISTw_tri[6]  ( .I(DataOw[6]), .OE(n138), .Z(DataIBISTw[6]) );
  BUFTD0 \DataIBISTw_tri[31]  ( .I(DataOw[31]), .OE(N9), .Z(DataIBISTw[31]) );
  BUFTD0 \DataIBISTw_tri[14]  ( .I(DataOw[14]), .OE(n137), .Z(DataIBISTw[14])
         );
  BUFTD0 \DataIBISTw_tri[22]  ( .I(DataOw[22]), .OE(n138), .Z(DataIBISTw[22])
         );
  BUFTD16 \DataO_tri[0]  ( .I(DataOw[0]), .OE(n129), .Z(DataO[0]) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOw[31]), .OE(n129), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOw[1]), .OE(n129), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOw[30]), .OE(n129), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOw[2]), .OE(n129), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOw[29]), .OE(n129), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOw[3]), .OE(n129), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOw[28]), .OE(n129), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOw[4]), .OE(n129), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOw[27]), .OE(n129), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOw[5]), .OE(n129), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOw[26]), .OE(n129), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOw[6]), .OE(n129), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOw[25]), .OE(n129), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOw[7]), .OE(n129), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOw[24]), .OE(n129), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOw[23]), .OE(n129), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOw[8]), .OE(n129), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOw[22]), .OE(n129), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOw[9]), .OE(n129), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOw[21]), .OE(n129), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOw[10]), .OE(n129), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOw[20]), .OE(n129), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOw[11]), .OE(n129), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOw[19]), .OE(n129), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOw[12]), .OE(n129), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOw[18]), .OE(n129), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOw[13]), .OE(n129), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOw[17]), .OE(n129), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOw[14]), .OE(n129), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOw[16]), .OE(n129), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOw[15]), .OE(n129), .Z(DataO[15]) );
  INVD3 U49 ( .I(N9), .ZN(n129) );
  INVD1 U50 ( .I(n135), .ZN(n136) );
  MUX2D0 U51 ( .I0(AddrR[2]), .I1(AddrBISTw[2]), .S(n138), .Z(n130) );
  MUX2D0 U52 ( .I0(AddrR[0]), .I1(AddrBISTw[0]), .S(n137), .Z(n131) );
  CKNXD16 U53 ( .I(n135), .ZN(ParityErr) );
  CKBXD0 U54 ( .I(n129), .Z(n133) );
  CKNXD16 U55 ( .I(n133), .ZN(Testing) );
  INVD1 U56 ( .I(n129), .ZN(n138) );
  INVD1 U57 ( .I(n129), .ZN(n137) );
  CKND0 U58 ( .CLK(n146), .CN(n135) );
  BUFFD2 U59 ( .I(ChipEna), .Z(n139) );
  BUFFD4 U60 ( .I(ClkR), .Z(n140) );
  MUX2D1 U61 ( .I0(DataI[19]), .I1(DataOBISTw[19]), .S(N9), .Z(DataIw[19]) );
  MUX2D1 U62 ( .I0(DataI[20]), .I1(DataOBISTw[20]), .S(N9), .Z(DataIw[20]) );
  MUX2D1 U63 ( .I0(DataI[16]), .I1(DataOBISTw[16]), .S(N9), .Z(DataIw[16]) );
  MUX2D1 U64 ( .I0(DataI[24]), .I1(DataOBISTw[24]), .S(n138), .Z(DataIw[24])
         );
  MUX2D1 U65 ( .I0(DataI[12]), .I1(DataOBISTw[12]), .S(n138), .Z(DataIw[12])
         );
  MUX2D1 U66 ( .I0(DataI[27]), .I1(DataOBISTw[27]), .S(n137), .Z(DataIw[27])
         );
  MUX2D1 U67 ( .I0(DataI[9]), .I1(DataOBISTw[9]), .S(n137), .Z(DataIw[9]) );
  MUX2D1 U68 ( .I0(DataI[28]), .I1(DataOBISTw[28]), .S(n137), .Z(DataIw[28])
         );
  MUX2D1 U69 ( .I0(DataI[0]), .I1(DataOBISTw[0]), .S(n138), .Z(DataIw[0]) );
  MUX2D1 U70 ( .I0(DataI[2]), .I1(DataOBISTw[2]), .S(n138), .Z(DataIw[2]) );
  MUX2D1 U71 ( .I0(DataI[10]), .I1(DataOBISTw[10]), .S(n137), .Z(DataIw[10])
         );
  MUX2D1 U72 ( .I0(DataI[11]), .I1(DataOBISTw[11]), .S(n137), .Z(DataIw[11])
         );
  MUX2D1 U73 ( .I0(DataI[4]), .I1(DataOBISTw[4]), .S(n137), .Z(DataIw[4]) );
  MUX2D1 U74 ( .I0(DataI[17]), .I1(DataOBISTw[17]), .S(n137), .Z(DataIw[17])
         );
  MUX2D1 U75 ( .I0(DataI[3]), .I1(DataOBISTw[3]), .S(N9), .Z(DataIw[3]) );
  MUX2D1 U76 ( .I0(DataI[18]), .I1(DataOBISTw[18]), .S(n137), .Z(DataIw[18])
         );
  MUX2D1 U77 ( .I0(DataI[1]), .I1(DataOBISTw[1]), .S(n138), .Z(DataIw[1]) );
  MUX2D1 U78 ( .I0(DataI[25]), .I1(DataOBISTw[25]), .S(n138), .Z(DataIw[25])
         );
  MUX2D1 U79 ( .I0(DataI[8]), .I1(DataOBISTw[8]), .S(n138), .Z(DataIw[8]) );
  MUX2D1 U80 ( .I0(DataI[26]), .I1(DataOBISTw[26]), .S(n138), .Z(DataIw[26])
         );
  MUX2D2 U81 ( .I0(AddrR[4]), .I1(AddrBISTw[4]), .S(N9), .Z(AddrRw[4]) );
  MUX2D2 U82 ( .I0(Read), .I1(ReadCmdBISTw), .S(N9), .Z(Readw) );
  CKBXD0 U83 ( .I(n143), .Z(n141) );
  CKNXD16 U84 ( .I(n141), .ZN(Dready) );
  CKND0 U85 ( .CLK(n145), .CN(n143) );
  MUX2D4 U86 ( .I0(AddrR[3]), .I1(AddrBISTw[3]), .S(n137), .Z(AddrRw[3]) );
  IOA21D1 U87 ( .A1(DataI[7]), .A2(n129), .B(n144), .ZN(DataIw[7]) );
  IOA21D1 U88 ( .A1(DataI[21]), .A2(n129), .B(n144), .ZN(DataIw[21]) );
  IOA21D1 U89 ( .A1(DataI[22]), .A2(n129), .B(n144), .ZN(DataIw[22]) );
  IOA21D1 U90 ( .A1(DataI[14]), .A2(n129), .B(n144), .ZN(DataIw[14]) );
  IOA21D1 U91 ( .A1(DataI[15]), .A2(n129), .B(n144), .ZN(DataIw[15]) );
  IOA21D1 U92 ( .A1(DataI[29]), .A2(n129), .B(n144), .ZN(DataIw[29]) );
  IOA21D1 U93 ( .A1(DataI[30]), .A2(n129), .B(n144), .ZN(DataIw[30]) );
  IOA21D1 U94 ( .A1(DataI[5]), .A2(n129), .B(n144), .ZN(DataIw[5]) );
  IOA21D1 U95 ( .A1(DataI[6]), .A2(n129), .B(n144), .ZN(DataIw[6]) );
  IOA21D1 U96 ( .A1(DataI[23]), .A2(n129), .B(n144), .ZN(DataIw[23]) );
  IOA21D1 U97 ( .A1(DataI[13]), .A2(n129), .B(n144), .ZN(DataIw[13]) );
  IOA21D1 U98 ( .A1(DataI[31]), .A2(n129), .B(n144), .ZN(DataIw[31]) );
  MUX2D0 U99 ( .I0(Write), .I1(WriteCmdBISTw), .S(n137), .Z(Writew) );
  INR2D0 U100 ( .A1(Dreadyw), .B1(n138), .ZN(n145) );
  CKND2D0 U101 ( .A1(DataOBISTw[7]), .A2(n137), .ZN(n144) );
  MUX2D0 U102 ( .I0(ClkW), .I1(n140), .S(n138), .Z(ClkWw) );
  MUX2D0 U103 ( .I0(AddrW[4]), .I1(AddrBISTw[4]), .S(N9), .Z(AddrWw[4]) );
  MUX2D0 U104 ( .I0(AddrW[3]), .I1(AddrBISTw[3]), .S(N9), .Z(AddrWw[3]) );
  MUX2D0 U105 ( .I0(AddrW[2]), .I1(AddrBISTw[2]), .S(n137), .Z(AddrWw[2]) );
  MUX2D0 U106 ( .I0(AddrW[1]), .I1(AddrBISTw[1]), .S(n138), .Z(AddrWw[1]) );
  MUX2D0 U107 ( .I0(AddrW[0]), .I1(AddrBISTw[0]), .S(N9), .Z(AddrWw[0]) );
  MUX2D0 U108 ( .I0(AddrR[1]), .I1(AddrBISTw[1]), .S(n137), .Z(AddrRw[1]) );
endmodule

