
module FullDup ( OutParDataA, OutParDataB, InParDataA, InParDataB, InParValidA, 
        InParValidB, ClockA, ClockB, Reset );
  output [31:0] OutParDataA;
  output [31:0] OutParDataB;
  input [31:0] InParDataA;
  input [31:0] InParDataB;
  input InParValidA, InParValidB, ClockA, ClockB, Reset;
  wire   n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, \SerDes_U1/Rx_ParClk ,
         \SerDes_U1/Tx_SerClk , \SerDes_U1/SerLineValid ,
         \SerDes_U1/Des_U1/SerRxToDecode , \SerDes_U1/Des_U1/SerialClk ,
         \SerDes_U1/Des_U1/N34 , \SerDes_U1/Des_U1/N33 ,
         \SerDes_U1/Des_U1/N32 , \SerDes_U1/Des_U1/N31 ,
         \SerDes_U1/Des_U1/N30 , \SerDes_U1/Des_U1/N29 ,
         \SerDes_U1/Des_U1/N28 , \SerDes_U1/Des_U1/N27 ,
         \SerDes_U1/Des_U1/N26 , \SerDes_U1/Des_U1/N25 ,
         \SerDes_U1/Des_U1/N24 , \SerDes_U1/Des_U1/N23 ,
         \SerDes_U1/Des_U1/N22 , \SerDes_U1/Des_U1/N21 ,
         \SerDes_U1/Des_U1/N20 , \SerDes_U1/Des_U1/N19 ,
         \SerDes_U1/Des_U1/N18 , \SerDes_U1/Des_U1/N17 ,
         \SerDes_U1/Des_U1/N16 , \SerDes_U1/Des_U1/N15 ,
         \SerDes_U1/Des_U1/N14 , \SerDes_U1/Des_U1/N13 ,
         \SerDes_U1/Des_U1/N12 , \SerDes_U1/Des_U1/N11 ,
         \SerDes_U1/Des_U1/N10 , \SerDes_U1/Des_U1/N9 , \SerDes_U1/Des_U1/N8 ,
         \SerDes_U1/Des_U1/N7 , \SerDes_U1/Des_U1/N6 , \SerDes_U1/Des_U1/N5 ,
         \SerDes_U1/Des_U1/N4 , \SerDes_U1/Des_U1/N3 , \SerDes_U2/Rx_ParClk ,
         \SerDes_U2/Tx_SerClk , \SerDes_U2/SerLineValid ,
         \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ,
         \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ,
         \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N84 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N82 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N80 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N78 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N76 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N74 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N72 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N70 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N68 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N66 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N64 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N62 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N60 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N58 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N56 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N54 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N28 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N26 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N24 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ,
         \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N83 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N81 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N79 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N77 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N75 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N73 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N71 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N69 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N67 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N65 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N63 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N61 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N59 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N57 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N55 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N53 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N29 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N27 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N25 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N24 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N23 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ,
         \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 , \SerDes_U2/Des_U1/SerRxToDecode ,
         \SerDes_U2/Des_U1/SerialClk , \SerDes_U2/Des_U1/N34 ,
         \SerDes_U2/Des_U1/N33 , \SerDes_U2/Des_U1/N32 ,
         \SerDes_U2/Des_U1/N31 , \SerDes_U2/Des_U1/N30 ,
         \SerDes_U2/Des_U1/N29 , \SerDes_U2/Des_U1/N28 ,
         \SerDes_U2/Des_U1/N27 , \SerDes_U2/Des_U1/N26 ,
         \SerDes_U2/Des_U1/N25 , \SerDes_U2/Des_U1/N24 ,
         \SerDes_U2/Des_U1/N23 , \SerDes_U2/Des_U1/N22 ,
         \SerDes_U2/Des_U1/N21 , \SerDes_U2/Des_U1/N20 ,
         \SerDes_U2/Des_U1/N19 , \SerDes_U2/Des_U1/N18 ,
         \SerDes_U2/Des_U1/N17 , \SerDes_U2/Des_U1/N16 ,
         \SerDes_U2/Des_U1/N15 , \SerDes_U2/Des_U1/N14 ,
         \SerDes_U2/Des_U1/N13 , \SerDes_U2/Des_U1/N12 ,
         \SerDes_U2/Des_U1/N11 , \SerDes_U2/Des_U1/N10 , \SerDes_U2/Des_U1/N9 ,
         \SerDes_U2/Des_U1/N8 , \SerDes_U2/Des_U1/N7 , \SerDes_U2/Des_U1/N6 ,
         \SerDes_U2/Des_U1/N5 , \SerDes_U2/Des_U1/N4 , \SerDes_U2/Des_U1/N3 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ,
         \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ,
         \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ,
         \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N79 , \SerDes_U1/Des_U1/DesDec_Rx1/N47 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N43 , \SerDes_U1/Des_U1/DesDec_Rx1/N42 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N41 , \SerDes_U1/Des_U1/DesDec_Rx1/N40 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N39 , \SerDes_U1/Des_U1/DesDec_Rx1/N38 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N37 , \SerDes_U1/Des_U1/DesDec_Rx1/N34 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N33 , \SerDes_U1/Des_U1/DesDec_Rx1/N32 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/N31 , \SerDes_U1/Des_U1/DesDec_Rx1/N30 ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ,
         \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N79 , \SerDes_U2/Des_U1/DesDec_Rx1/N47 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N43 , \SerDes_U2/Des_U1/DesDec_Rx1/N42 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N41 , \SerDes_U2/Des_U1/DesDec_Rx1/N40 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N39 , \SerDes_U2/Des_U1/DesDec_Rx1/N38 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N37 , \SerDes_U2/Des_U1/DesDec_Rx1/N34 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N33 , \SerDes_U2/Des_U1/DesDec_Rx1/N32 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/N31 , \SerDes_U2/Des_U1/DesDec_Rx1/N30 ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ,
         \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ,
         \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ,
         \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ,
         \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ,
         \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 , n717, n721, n723,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n762,
         n764, n766, n768, n770, n772, n774, n776, n778, n780, n782, n784,
         n786, n788, n790, n792, n794, n796, n798, n800, n802, n804, n806,
         n808, n810, n812, n814, n816, n818, n820, n822, n837, n841, n842,
         n849, n855, n856, n858, n864, n869, n871, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n910, n912, n914, n916, n918,
         n920, n922, n924, n926, n928, n930, n932, n934, n936, n938, n940,
         n942, n944, n946, n948, n950, n952, n954, n956, n958, n960, n962,
         n964, n966, n968, n970, n985, n989, n990, n997, n1003, n1004, n1006,
         n1011, n1015, n1016, n1018, n1024, n1030, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1406, n1408, n1410,
         n1412, n1414, n1416, n1418, n1420, n1422, n1424, n1426, n1428, n1430,
         n1432, n1434, n1436, n1438, n1440, n1442, n1444, n1446, n1448, n1450,
         n1452, n1454, n1456, n1458, n1460, n1462, n1464, n1466, n1468, n1470,
         n1472, n1474, n1476, n1478, n1480, n1482, n1484, n1486, n1488, n1490,
         n1492, n1494, n1496, n1498, n1500, n1502, n1504, n1506, n1508, n1510,
         n1512, n1514, n1516, n1518, n1520, n1522, n1524, n1526, n1528, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997;
  wire   [31:0] \SerDes_U1/Ser_U1/FIFO_Out ;
  wire   [31:0] \SerDes_U1/Des_U1/DecodeToFIFO ;
  wire   [31:0] \SerDes_U2/Ser_U1/FIFO_Out ;
  wire   [3:0] \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr ;
  wire   [3:0] \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState ;
  wire   [2:0] \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState ;
  wire   [31:0] \SerDes_U2/Des_U1/DecodeToFIFO ;
  wire   [2:0] \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr ;
  wire   [2:0] \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState ;
  wire   [2:0] \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState ;
  wire   [1:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq ;
  wire   [1:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq ;
  wire   [1:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq ;
  wire   [1:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq ;
  wire   [5:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD ;
  wire   [5:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD ;
  wire   [3:0] \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr ;
  wire   [3:0] \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr ;

  DEL005 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/SM_DeGlitcher1  ( .I(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ), .Z(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleDelay1  ( .I(ClockA), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleDelay1  ( .I(
        \SerDes_U1/Rx_ParClk ), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleDelay1  ( .I(ClockB), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleDelay1  ( .I(
        \SerDes_U2/Rx_ParClk ), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [1]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[4].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[3].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [4]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[2].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [3]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[1].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [2]) );
  DEL005 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DelayLine[0].Delay85ps  ( 
        .I(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [1]) );
  CKND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/I_2  ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/I_2  ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/I_2  ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [0]) );
  CKND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/I_2  ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [0]) );
  DFND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/FullFIFOr_reg  ( .D(n1246), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(n2967) );
  DFND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/EmptyFIFOr_reg  ( .D(n1232), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(n1302), .QN(n1036) );
  DFND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/EmptyFIFOr_reg  ( .D(n1231), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(n1299), .QN(n1035) );
  DFND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/FullFIFOr_reg  ( .D(n1230), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .Q(n2962), .QN(n1401) );
  EDFCNQD2 \SerDes_U2/Des_U1/DesDec_Rx1/ParClkr_reg  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N37 ), .E(
        \SerDes_U2/Des_U1/DesDec_Rx1/N43 ), .CP(n2284), .CDN(n1247), .Q(
        \SerDes_U2/Rx_ParClk ) );
  FullDup_DW01_inc_0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/add_16  ( .A(
        {\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/add_16  ( .A(
        {\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_2 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/add_16  ( .A(
        {\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 }) );
  FullDup_DW01_inc_3 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/add_16  ( .A(
        {\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 }) );
  FullDup_DW01_dec_0 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 }) );
  FullDup_DW01_inc_4 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 }) );
  FullDup_DW01_inc_5 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 , 
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 }) );
  FullDup_DW01_dec_1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 }) );
  FullDup_DW01_inc_6 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 }) );
  FullDup_DW01_inc_7 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 , 
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 }) );
  FullDup_DW01_dec_2 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 }) );
  FullDup_DW01_inc_8 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 }) );
  FullDup_DW01_inc_9 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 , 
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 }) );
  FullDup_DW01_dec_3 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/sub_193  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 }) );
  FullDup_DW01_inc_10 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/Sampler/add_190  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 }) );
  FullDup_DW01_inc_11 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutGen/add_171  ( 
        .A({\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 , 
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 }) );
  FullDup_DW01_inc_12 \SerDes_U2/Des_U1/DesDec_Rx1/ClkGen/add_206  ( .A({
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] , 
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] }), .SUM({
        \SerDes_U2/Des_U1/DesDec_Rx1/N34 , \SerDes_U2/Des_U1/DesDec_Rx1/N33 , 
        \SerDes_U2/Des_U1/DesDec_Rx1/N32 , \SerDes_U2/Des_U1/DesDec_Rx1/N31 , 
        \SerDes_U2/Des_U1/DesDec_Rx1/N30 }) );
  FullDup_DW01_inc_13 \SerDes_U1/Des_U1/DesDec_Rx1/ClkGen/add_206  ( .A({
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] , 
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] }), .SUM({
        \SerDes_U1/Des_U1/DesDec_Rx1/N34 , \SerDes_U1/Des_U1/DesDec_Rx1/N33 , 
        \SerDes_U1/Des_U1/DesDec_Rx1/N32 , \SerDes_U1/Des_U1/DesDec_Rx1/N31 , 
        \SerDes_U1/Des_U1/DesDec_Rx1/N30 }) );
  FullDup_DW01_dec_4 \SerDes_U2/Ser_U1/SerEnc_Tx1/ShifterBlock/sub_132  ( .A({
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 }), .SUM({
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 , 
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 })
         );
  FullDup_DW01_dec_5 \SerDes_U1/Ser_U1/SerEnc_Tx1/ShifterBlock/sub_132  ( .A({
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N6 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N4 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 }), .SUM({
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 , 
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 , \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 })
         );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[31]  ( .D(\SerDes_U2/Des_U1/N34 ), .CP(
        ClockA), .CDN(n2216), .Q(n2998) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[30]  ( .D(\SerDes_U2/Des_U1/N33 ), .CP(
        ClockA), .CDN(n2215), .Q(n2999) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[29]  ( .D(\SerDes_U2/Des_U1/N32 ), .CP(
        ClockA), .CDN(n2216), .Q(n3000) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[28]  ( .D(\SerDes_U2/Des_U1/N31 ), .CP(
        ClockA), .CDN(n2215), .Q(n3001) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[27]  ( .D(\SerDes_U2/Des_U1/N30 ), .CP(
        ClockA), .CDN(n2227), .Q(n3002) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[26]  ( .D(\SerDes_U2/Des_U1/N29 ), .CP(
        ClockA), .CDN(n2232), .Q(n3003) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[25]  ( .D(\SerDes_U2/Des_U1/N28 ), .CP(
        ClockA), .CDN(n2220), .Q(n3004) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[24]  ( .D(\SerDes_U2/Des_U1/N27 ), .CP(
        ClockA), .CDN(n2215), .Q(n3005) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[23]  ( .D(\SerDes_U2/Des_U1/N26 ), .CP(
        ClockA), .CDN(n2216), .Q(n3006) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[22]  ( .D(\SerDes_U2/Des_U1/N25 ), .CP(
        ClockA), .CDN(n2215), .Q(n3007) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[21]  ( .D(\SerDes_U2/Des_U1/N24 ), .CP(
        ClockA), .CDN(n2218), .Q(n3008) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[20]  ( .D(\SerDes_U2/Des_U1/N23 ), .CP(
        ClockA), .CDN(n2215), .Q(n3009) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[19]  ( .D(\SerDes_U2/Des_U1/N22 ), .CP(
        ClockA), .CDN(n2228), .Q(n3010) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[18]  ( .D(\SerDes_U2/Des_U1/N21 ), .CP(
        ClockA), .CDN(n2215), .Q(n3011) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[17]  ( .D(\SerDes_U2/Des_U1/N20 ), .CP(
        ClockA), .CDN(n2216), .Q(n3012) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[16]  ( .D(\SerDes_U2/Des_U1/N19 ), .CP(
        ClockA), .CDN(n2215), .Q(n3013) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[15]  ( .D(\SerDes_U2/Des_U1/N18 ), .CP(
        ClockA), .CDN(n2216), .Q(n3014) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[14]  ( .D(\SerDes_U2/Des_U1/N17 ), .CP(
        ClockA), .CDN(n2219), .Q(n3015) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[13]  ( .D(\SerDes_U2/Des_U1/N16 ), .CP(
        ClockA), .CDN(n2230), .Q(n3016) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[12]  ( .D(\SerDes_U2/Des_U1/N15 ), .CP(
        ClockA), .CDN(n2216), .Q(n3017) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[11]  ( .D(\SerDes_U2/Des_U1/N14 ), .CP(
        ClockA), .CDN(n2233), .Q(n3018) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[10]  ( .D(\SerDes_U2/Des_U1/N13 ), .CP(
        ClockA), .CDN(n2217), .Q(n3019) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[9]  ( .D(\SerDes_U2/Des_U1/N12 ), .CP(
        ClockA), .CDN(n2218), .Q(n3020) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[8]  ( .D(\SerDes_U2/Des_U1/N11 ), .CP(
        ClockA), .CDN(n2216), .Q(n3021) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[7]  ( .D(\SerDes_U2/Des_U1/N10 ), .CP(
        ClockA), .CDN(n2218), .Q(n3022) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[6]  ( .D(\SerDes_U2/Des_U1/N9 ), .CP(
        ClockA), .CDN(n2216), .Q(n3023) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[5]  ( .D(\SerDes_U2/Des_U1/N8 ), .CP(
        ClockA), .CDN(n2226), .Q(n3024) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[4]  ( .D(\SerDes_U2/Des_U1/N7 ), .CP(
        ClockA), .CDN(n2217), .Q(n3025) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[3]  ( .D(\SerDes_U2/Des_U1/N6 ), .CP(
        ClockA), .CDN(n2216), .Q(n3026) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[2]  ( .D(\SerDes_U2/Des_U1/N5 ), .CP(
        ClockA), .CDN(n2217), .Q(n3027) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[1]  ( .D(\SerDes_U2/Des_U1/N4 ), .CP(
        ClockA), .CDN(n2216), .Q(n3028) );
  DFCNQD1 \SerDes_U2/Des_U1/ParBuf_reg[0]  ( .D(\SerDes_U2/Des_U1/N3 ), .CP(
        ClockA), .CDN(n2217), .Q(n3029) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[31]  ( .D(\SerDes_U1/Des_U1/N34 ), .CP(
        ClockB), .CDN(n2233), .Q(n3030) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[30]  ( .D(\SerDes_U1/Des_U1/N33 ), .CP(
        ClockB), .CDN(n2233), .Q(n3031) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[29]  ( .D(\SerDes_U1/Des_U1/N32 ), .CP(
        ClockB), .CDN(n2233), .Q(n3032) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[28]  ( .D(\SerDes_U1/Des_U1/N31 ), .CP(
        ClockB), .CDN(n2233), .Q(n3033) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[27]  ( .D(\SerDes_U1/Des_U1/N30 ), .CP(
        ClockB), .CDN(n2232), .Q(n3034) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[26]  ( .D(\SerDes_U1/Des_U1/N29 ), .CP(
        ClockB), .CDN(n2232), .Q(n3035) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[25]  ( .D(\SerDes_U1/Des_U1/N28 ), .CP(
        ClockB), .CDN(n2232), .Q(n3036) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[24]  ( .D(\SerDes_U1/Des_U1/N27 ), .CP(
        ClockB), .CDN(n2232), .Q(n3037) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[23]  ( .D(\SerDes_U1/Des_U1/N26 ), .CP(
        ClockB), .CDN(n2232), .Q(n3038) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[22]  ( .D(\SerDes_U1/Des_U1/N25 ), .CP(
        ClockB), .CDN(n2232), .Q(n3039) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[21]  ( .D(\SerDes_U1/Des_U1/N24 ), .CP(
        ClockB), .CDN(n2232), .Q(n3040) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[20]  ( .D(\SerDes_U1/Des_U1/N23 ), .CP(
        ClockB), .CDN(n2232), .Q(n3041) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[19]  ( .D(\SerDes_U1/Des_U1/N22 ), .CP(
        ClockB), .CDN(n2232), .Q(n3042) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[18]  ( .D(\SerDes_U1/Des_U1/N21 ), .CP(
        ClockB), .CDN(n2231), .Q(n3043) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[17]  ( .D(\SerDes_U1/Des_U1/N20 ), .CP(
        ClockB), .CDN(n2231), .Q(n3044) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[16]  ( .D(\SerDes_U1/Des_U1/N19 ), .CP(
        ClockB), .CDN(n2231), .Q(n3045) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[15]  ( .D(\SerDes_U1/Des_U1/N18 ), .CP(
        ClockB), .CDN(n2231), .Q(n3046) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[14]  ( .D(\SerDes_U1/Des_U1/N17 ), .CP(
        ClockB), .CDN(n2231), .Q(n3047) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[13]  ( .D(\SerDes_U1/Des_U1/N16 ), .CP(
        ClockB), .CDN(n2231), .Q(n3048) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[12]  ( .D(\SerDes_U1/Des_U1/N15 ), .CP(
        ClockB), .CDN(n2231), .Q(n3049) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[11]  ( .D(\SerDes_U1/Des_U1/N14 ), .CP(
        ClockB), .CDN(n2231), .Q(n3050) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[10]  ( .D(\SerDes_U1/Des_U1/N13 ), .CP(
        ClockB), .CDN(n2231), .Q(n3051) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[9]  ( .D(\SerDes_U1/Des_U1/N12 ), .CP(
        ClockB), .CDN(n2231), .Q(n3052) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[8]  ( .D(\SerDes_U1/Des_U1/N11 ), .CP(
        ClockB), .CDN(n2230), .Q(n3053) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[7]  ( .D(\SerDes_U1/Des_U1/N10 ), .CP(
        ClockB), .CDN(n2230), .Q(n3054) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[6]  ( .D(\SerDes_U1/Des_U1/N9 ), .CP(
        ClockB), .CDN(n2230), .Q(n3055) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[5]  ( .D(\SerDes_U1/Des_U1/N8 ), .CP(
        ClockB), .CDN(n2230), .Q(n3056) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[4]  ( .D(\SerDes_U1/Des_U1/N7 ), .CP(
        ClockB), .CDN(n2230), .Q(n3057) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[3]  ( .D(\SerDes_U1/Des_U1/N6 ), .CP(
        ClockB), .CDN(n2230), .Q(n3058) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[2]  ( .D(\SerDes_U1/Des_U1/N5 ), .CP(
        ClockB), .CDN(n2230), .Q(n3059) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[1]  ( .D(\SerDes_U1/Des_U1/N4 ), .CP(
        ClockB), .CDN(n2230), .Q(n3060) );
  DFCNQD1 \SerDes_U1/Des_U1/ParBuf_reg[0]  ( .D(\SerDes_U1/Des_U1/N3 ), .CP(
        ClockB), .CDN(n2230), .Q(n3061) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[63]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ), .CPN(n2291), .CDN(n2208), 
        .QN(n1004) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[63]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ), .CPN(n2274), .CDN(n2195), 
        .QN(n856) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2228), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2227), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2232), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2268), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2202), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2221), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2223), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2224), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2226), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2215), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2217), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2310), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2219), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2220), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2260), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2216), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2269), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2230), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2229), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2220), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2223), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2226), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2304), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2184), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2201), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(n2305), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2237), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .CP(\SerDes_U2/Rx_ParClk ), 
        .CDN(n2201), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] )
         );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2213), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2215), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2260), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2232), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2233), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2226), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2228), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2229), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2221), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2214), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2224), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2318), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2224), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2201), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2319), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2203), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2202), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N55 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[26]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[29]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N82 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[30]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[30]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N83 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[29]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[26]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N79 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[25]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[22]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N75 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[21]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[18]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N71 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[17]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N54 ), .CP(n2351), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N58 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[6]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[9]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N62 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[10]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[13]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N66 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[14]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[14]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N67 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[13]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[10]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N63 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[9]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[6]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N59 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[17]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N70 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[18]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[21]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N74 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[22]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[25]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N78 ), .CP(n2351), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2186), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2187), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2264), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2214), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2210), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2200), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2215), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2266), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2258), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2200), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2316), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2206), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2242), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2202), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2248), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2247), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2246), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2210), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2190), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2187), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2183), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2201), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2202), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2203), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2217), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2248), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2247), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2246), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2266), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2314), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2203), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2241), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N57 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N53 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[27]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N80 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[28]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[31]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N84 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[31]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[28]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N81 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[27]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[24]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N77 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[23]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ), .CP(n2349), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[20]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N73 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[19]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[16]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N69 ), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[15]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N56 ), .CP(n2351), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[7]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N60 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[8]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[11]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N64 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[12]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ), .CP(n2351), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[15]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N68 ), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[16]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n1239), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .QN(n1385) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n1238), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .QN(n1386) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1235), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .QN(n1387) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1234), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .QN(n1388) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[12]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N65 ), .CP(n2349), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[11]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[8]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N61 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf_reg[7]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ), .CP(n2349), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[19]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N72 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[20]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[23]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N76 ), .CP(n2351), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf_reg[24]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ), .CP(n2351), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n1132), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .QN(n1392) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n1131), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .QN(n1393) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1127), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2195), 
        .QN(n1316) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1126), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2195), 
        .QN(n1317) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n1224), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .QN(n1389) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1220), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .QN(n1390) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1219), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2205), 
        .QN(n1391) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2199), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2245), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2248), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2199), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2211), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2206), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2214), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2213), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2210), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2183), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2184), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2193), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2312), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2211), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2228), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2189), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2236), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2189), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2213), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2307), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2220), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2223), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2224), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2308), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2226), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2228), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n1042), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1394) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[0]  ( .D(n1041), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1395) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n1040), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1396) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1039), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1318) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[0]  ( .D(n1038), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1319) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1037), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .QN(n1320) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[8]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ), .CPN(n2296), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ), .QN(n910) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[9]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[8] ), .CPN(n2292), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ), .QN(n912) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[10]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[9] ), .CPN(n2297), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ), .QN(n914) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[11]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[10] ), .CPN(n2289), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ), .QN(n916) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[12]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[11] ), .CPN(n2292), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ), .QN(n918) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[13]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[12] ), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2214), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ), .QN(n920) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[14]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[13] ), .CPN(n2290), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ), .QN(n922) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[15]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[14] ), .CPN(n2290), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ), .QN(n924) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[18]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2212), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ), .QN(n997) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[19]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[18] ), .CPN(n2295), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ), .QN(n1003) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[22]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ), .CPN(n2297), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ), .QN(n2992) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[24]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ), .CPN(n2296), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ), .QN(n926) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[25]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[24] ), .CPN(n2295), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ), .QN(n928) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[26]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[25] ), .CPN(n2297), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ), .QN(n930) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[27]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[26] ), .CPN(n2289), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ), .QN(n932) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[28]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[27] ), .CPN(n2290), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ), .QN(n934) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[29]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[28] ), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2211), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ), .QN(n936) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[30]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[29] ), .CPN(n2298), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ), .QN(n938) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[31]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[30] ), .CPN(n2291), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ), .QN(n940) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[32]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[31] ), .CPN(n2295), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ), .QN(n2991) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[34]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ), .CPN(n2294), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ), .QN(n989) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[35]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[34] ), .CPN(n2294), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ), .QN(n990) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[38]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ), .CPN(n2294), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ), .QN(n2993) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[40]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ), .CPN(n2294), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ), .QN(n942) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[41]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[40] ), .CPN(n2294), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ), .QN(n944) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[42]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[41] ), .CPN(n2293), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ), .QN(n946) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[43]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[42] ), .CPN(n2293), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ), .QN(n948) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[44]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[43] ), .CPN(n2293), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ), .QN(n950) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[45]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[44] ), .CPN(n2293), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ), .QN(n952) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[46]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[45] ), .CPN(n2293), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ), .QN(n954) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[47]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[46] ), .CPN(n2293), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ), .QN(n956) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[48]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[47] ), .CPN(n2293), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ), .QN(n985) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[53]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ), .QN(n2995) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[55]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ), .QN(n2994) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[56]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[55] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ), .QN(n958) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[57]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[56] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ), .QN(n960) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[58]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[57] ), .CPN(n2292), .CDN(n2208), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ), .QN(n962) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[59]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[58] ), .CPN(n2292), .CDN(n2208), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ), .QN(n964) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[60]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[59] ), .CPN(n2291), .CDN(n2208), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ), .QN(n966) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[61]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[60] ), .CPN(n2291), .CDN(n2208), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ), .QN(n968) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[62]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[61] ), .CPN(n2291), .CDN(n2208), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[62] ), .QN(n970) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[31]  ( .D(n1209), .CPN(
        n2291), .CDN(n2208), .QN(n1352) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[30]  ( .D(n1208), .CPN(
        n2291), .CDN(n2183), .QN(n1351) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[29]  ( .D(n1207), .CPN(
        n2291), .CDN(n2183), .QN(n1350) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[28]  ( .D(n1206), .CPN(
        n2291), .CDN(n2183), .QN(n1349) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[27]  ( .D(n1205), .CPN(
        n2291), .CDN(n2183), .QN(n1348) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[26]  ( .D(n1204), .CPN(
        n2290), .CDN(n2183), .QN(n1347) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[25]  ( .D(n1203), .CPN(
        n2290), .CDN(n2183), .QN(n1346) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[24]  ( .D(n1202), .CPN(
        n2290), .CDN(n2183), .QN(n1345) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[23]  ( .D(n1201), .CPN(
        n2290), .CDN(n2183), .QN(n1344) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[22]  ( .D(n1200), .CPN(
        n2290), .CDN(n2183), .QN(n1343) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[21]  ( .D(n1199), .CPN(
        n2290), .CDN(n2184), .QN(n1342) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[20]  ( .D(n1198), .CPN(
        n2290), .CDN(n2184), .QN(n1341) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[19]  ( .D(n1197), .CPN(
        n2290), .CDN(n2184), .QN(n1340) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[18]  ( .D(n1196), .CPN(
        n2290), .CDN(n2184), .QN(n1339) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[17]  ( .D(n1195), .CPN(
        n2289), .CDN(n2184), .QN(n1338) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[16]  ( .D(n1194), .CPN(
        n2289), .CDN(n2184), .QN(n1337) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[15]  ( .D(n1193), .CPN(
        n2289), .CDN(n2184), .QN(n1336) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[14]  ( .D(n1192), .CPN(
        n2289), .CDN(n2184), .QN(n1335) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[13]  ( .D(n1191), .CPN(
        n2289), .CDN(n2184), .QN(n1334) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[12]  ( .D(n1190), .CPN(
        n2289), .CDN(n2184), .QN(n1333) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[11]  ( .D(n1189), .CPN(
        n2289), .CDN(n2185), .QN(n1332) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[10]  ( .D(n1188), .CPN(
        n2289), .CDN(n2185), .QN(n1331) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[9]  ( .D(n1187), .CPN(n2289), .CDN(n2185), .QN(n1330) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[8]  ( .D(n1186), .CPN(n2296), .CDN(n2185), .QN(n1329) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[7]  ( .D(n1185), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2185), .QN(n1328) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[6]  ( .D(n1184), .CPN(n2296), .CDN(n2185), .QN(n1327) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[5]  ( .D(n1183), .CPN(n2298), .CDN(n2185), .QN(n1326) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[4]  ( .D(n1182), .CPN(n2295), .CDN(n2185), .QN(n1325) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[3]  ( .D(n1181), .CPN(n2297), .CDN(n2185), .QN(n1324) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[2]  ( .D(n1180), .CPN(n2296), .CDN(n2185), .QN(n1323) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[1]  ( .D(n1179), .CPN(n2295), .CDN(n2186), .QN(n1322) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/Decoder_reg[0]  ( .D(n1178), .CPN(n2296), .CDN(n2186), .QN(n1321) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[8]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ), .QN(n762) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[9]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[8] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ), .QN(n764) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[10]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[9] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ), .QN(n766) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[11]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[10] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ), .QN(n768) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[12]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[11] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ), .QN(n770) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[13]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[12] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ), .QN(n772) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[14]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[13] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ), .QN(n774) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[15]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[14] ), .CPN(n2279), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ), .QN(n776) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[18]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ), .QN(n849) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[19]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[18] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ), .QN(n855) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[22]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ), .QN(n2979) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[24]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ), .CPN(n2278), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ), .QN(n778) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[25]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[24] ), .CPN(n2278), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ), .QN(n780) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[26]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[25] ), .CPN(n2278), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ), .QN(n782) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[27]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[26] ), .CPN(n2278), .CDN(n2201), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ), .QN(n784) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[28]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[27] ), .CPN(n2278), .CDN(n2201), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ), .QN(n786) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[29]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[28] ), .CPN(n2278), .CDN(n2201), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ), .QN(n788) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[30]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[29] ), .CPN(n2278), .CDN(n2201), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ), .QN(n790) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[31]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[30] ), .CPN(n2278), .CDN(n2183), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ), .QN(n792) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[32]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[31] ), .CPN(n2278), .CDN(n2192), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ), .QN(n2978) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[34]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ), .CPN(n2277), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ), .QN(n841) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[35]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[34] ), .CPN(n2277), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ), .QN(n842) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[38]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ), .QN(n2980) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[40]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ), .QN(n794) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[41]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[40] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ), .QN(n796) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[42]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[41] ), .CPN(n2276), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ), .QN(n798) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[43]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[42] ), .CPN(n2276), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ), .QN(n800) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[44]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[43] ), .CPN(n2276), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ), .QN(n802) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[45]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[44] ), .CPN(n2276), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ), .QN(n804) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[46]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[45] ), .CPN(n2276), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ), .QN(n806) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[47]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[46] ), .CPN(n2276), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ), .QN(n808) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[48]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[47] ), .CPN(n2276), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ), .QN(n837) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[53]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ), .CPN(n2275), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ), .QN(n2982) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[55]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ), .CPN(n2275), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ), .QN(n2981) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[56]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[55] ), .CPN(n2275), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ), .QN(n810) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[57]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[56] ), .CPN(n2275), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ), .QN(n812) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[58]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[57] ), .CPN(n2275), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ), .QN(n814) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[59]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[58] ), .CPN(n2275), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ), .QN(n816) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[60]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[59] ), .CPN(n2274), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ), .QN(n818) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[61]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[60] ), .CPN(n2274), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ), .QN(n820) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[62]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[61] ), .CPN(n2274), .CDN(n2195), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[62] ), .QN(n822) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[31]  ( .D(n1118), .CPN(
        n2274), .CDN(n2194), .QN(n1384) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[30]  ( .D(n1117), .CPN(
        n2274), .CDN(n2193), .QN(n1383) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[29]  ( .D(n1116), .CPN(
        n2274), .CDN(n2193), .QN(n1382) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[28]  ( .D(n1115), .CPN(
        n2274), .CDN(n2193), .QN(n1381) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[27]  ( .D(n1114), .CPN(
        n2274), .CDN(n2193), .QN(n1380) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[26]  ( .D(n1113), .CPN(
        n2273), .CDN(n2193), .QN(n1379) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[25]  ( .D(n1112), .CPN(
        n2273), .CDN(n2193), .QN(n1378) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[24]  ( .D(n1111), .CPN(
        n2273), .CDN(n2193), .QN(n1377) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[23]  ( .D(n1110), .CPN(
        n2273), .CDN(n2193), .QN(n1376) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[22]  ( .D(n1109), .CPN(
        n2273), .CDN(n2193), .QN(n1375) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[21]  ( .D(n1108), .CPN(
        n2273), .CDN(n2192), .QN(n1374) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[20]  ( .D(n1107), .CPN(
        n2273), .CDN(n2192), .QN(n1373) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[19]  ( .D(n1106), .CPN(
        n2273), .CDN(n2192), .QN(n1372) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[18]  ( .D(n1105), .CPN(
        n2273), .CDN(n2192), .QN(n1371) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[17]  ( .D(n1104), .CPN(
        n2272), .CDN(n2192), .QN(n1370) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[16]  ( .D(n1103), .CPN(
        n2272), .CDN(n2192), .QN(n1369) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[15]  ( .D(n1102), .CPN(
        n2272), .CDN(n2192), .QN(n1368) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[14]  ( .D(n1101), .CPN(
        n2272), .CDN(n2192), .QN(n1367) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[13]  ( .D(n1100), .CPN(
        n2272), .CDN(n2192), .QN(n1366) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[12]  ( .D(n1099), .CPN(
        n2272), .CDN(n2191), .QN(n1365) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[11]  ( .D(n1098), .CPN(
        n2272), .CDN(n2191), .QN(n1364) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[10]  ( .D(n1097), .CPN(
        n2272), .CDN(n2191), .QN(n1363) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[9]  ( .D(n1096), .CPN(n2272), .CDN(n2191), .QN(n1362) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[8]  ( .D(n1095), .CPN(n2271), .CDN(n2191), .QN(n1361) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[7]  ( .D(n1094), .CPN(n2271), .CDN(n2191), .QN(n1360) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[6]  ( .D(n1093), .CPN(n2271), .CDN(n2191), .QN(n1359) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[5]  ( .D(n1092), .CPN(n2271), .CDN(n2191), .QN(n1358) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[4]  ( .D(n1091), .CPN(n2271), .CDN(n2191), .QN(n1357) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[3]  ( .D(n1090), .CPN(n2271), .CDN(n2191), .QN(n1356) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[2]  ( .D(n1089), .CPN(n2271), .CDN(n2190), .QN(n1355) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[1]  ( .D(n1088), .CPN(n2271), .CDN(n2190), .QN(n1354) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/Decoder_reg[0]  ( .D(n1087), .CPN(n2271), .CDN(n2190), .QN(n1353) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[1]  ( .D(n1245), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .QN(n1030) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[0]  ( .D(n1243), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .QN(n1024) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[2]  ( .D(n1241), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .Q(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .QN(n1018) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[1]  ( .D(n1138), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2190), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .QN(n871) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[0]  ( .D(n1136), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2193), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .QN(n864) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[2]  ( .D(n1134), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .QN(n858) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[1]  ( .D(n1229), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .QN(n1016) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[0]  ( .D(n1227), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .QN(n1011) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState_reg[2]  ( .D(n1222), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .QN(n1006) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[1]  ( .D(n1047), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2205), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .QN(n723) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[0]  ( .D(n1045), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .QN(n717) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [31]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2187), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2261), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2251), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [23]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2250), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [21]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [19]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [17]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [15]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [13]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [9]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [7]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2246), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [5]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [3]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [1]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [0]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [2]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2213), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [4]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [6]), .E(n2321), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [10]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [12]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [14]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [16]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [20]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [22]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [26]), .E(n2322), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2262), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        \SerDes_U2/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .CP(\SerDes_U2/Rx_ParClk ), .CDN(n2215), .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2200), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2206), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2253), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2421), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2257), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[14][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2201), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2199), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2212), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2203), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2199), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2223), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2419), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[13][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2215), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2413), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[10][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2229), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2206), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2206), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2248), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2246), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2266), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2411), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[9][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2184), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2184), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2193), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2213), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2203), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2187), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2193), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2211), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2405), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2224), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2201), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2183), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2184), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2187), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2403), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2214), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2226), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2218), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2232), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2230), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2228), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2226), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2224), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2223), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2221), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2220), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2218), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2215), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2397), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2206), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2228), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2226), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2232), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2233), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2224), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2223), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2220), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2184), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2266), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2245), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2265), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2202), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2395), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2201), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2222), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2265), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2248), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2187), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2193), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2218), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2266), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2226), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2221), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2423), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[15][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2226), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2182), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2217), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2257), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2193), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2227), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2266), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2417), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[12][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2243), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2183), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2221), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2253), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2249), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2246), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2216), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2415), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2244), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[11][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2200), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2237), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2221), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2213), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2244), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2263), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2252), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2259), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2256), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2200), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2215), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2270), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2217), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2192), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2260), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2267), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2268), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2231), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n1247), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2200), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2217), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2214), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2212), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2409), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2206), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[8][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2183), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2238), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2239), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2407), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2213), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2183), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2265), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2248), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2269), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2184), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2185), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2187), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2200), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2217), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2203), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2264), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2248), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2401), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2247), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2246), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2249), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2253), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2254), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2255), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2240), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2183), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2191), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2205), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2208), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2207), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2245), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2251), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2234), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2242), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2241), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2261), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2219), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2220), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2222), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2399), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2223), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2224), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2225), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [31]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2194), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [29]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2246), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [27]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2191), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2195), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2196), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [21]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2198), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [19]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2197), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [17]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2212), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [15]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2214), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2209), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [11]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2210), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [9]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2204), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [7]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [5]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [3]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [1]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [0]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [4]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [6]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [8]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [10]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [12]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2235), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [14]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [20]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [22]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [24]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .E(n2393), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [28]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        \SerDes_U1/Des_U1/DecodeToFIFO [30]), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .CP(\SerDes_U1/Rx_ParClk ), .CDN(n2236), .Q(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2262), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [0]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2193), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [1]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ), .E(n2348), .CP(ClockA), 
        .CDN(n2232), .Q(\SerDes_U1/Ser_U1/FIFO_Out [2]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ), .E(n2348), .CP(ClockA), 
        .CDN(n2235), .Q(\SerDes_U1/Ser_U1/FIFO_Out [3]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ), .E(n2348), .CP(ClockA), 
        .CDN(n2208), .Q(\SerDes_U1/Ser_U1/FIFO_Out [4]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ), .E(n2348), .CP(ClockA), 
        .CDN(n2259), .Q(\SerDes_U1/Ser_U1/FIFO_Out [5]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ), .E(n2348), .CP(ClockA), 
        .CDN(n2195), .Q(\SerDes_U1/Ser_U1/FIFO_Out [6]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ), .E(n2348), .CP(ClockA), 
        .CDN(n2215), .Q(\SerDes_U1/Ser_U1/FIFO_Out [7]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ), .E(n2348), .CP(ClockA), 
        .CDN(n2227), .Q(\SerDes_U1/Ser_U1/FIFO_Out [8]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ), .E(n2348), .CP(ClockA), 
        .CDN(n2192), .Q(\SerDes_U1/Ser_U1/FIFO_Out [9]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ), .E(n2348), .CP(ClockA), 
        .CDN(n2258), .Q(\SerDes_U1/Ser_U1/FIFO_Out [10]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ), .E(n2348), .CP(ClockA), 
        .CDN(n2257), .Q(\SerDes_U1/Ser_U1/FIFO_Out [11]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ), .E(n2348), .CP(ClockA), 
        .CDN(n2267), .Q(\SerDes_U1/Ser_U1/FIFO_Out [12]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2224), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [13]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2210), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [14]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2214), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [15]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2270), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [16]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2256), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [17]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2259), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [18]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2242), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [19]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2182), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [20]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2261), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [21]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ), .E(n2348), .CP(ClockA), 
        .CDN(n2265), .Q(\SerDes_U1/Ser_U1/FIFO_Out [22]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2265), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [23]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ), .E(n2348), .CP(ClockA), 
        .CDN(n2254), .Q(\SerDes_U1/Ser_U1/FIFO_Out [24]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2253), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [25]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ), .E(n2348), .CP(ClockA), 
        .CDN(n2191), .Q(\SerDes_U1/Ser_U1/FIFO_Out [26]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2261), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [27]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ), .E(n2348), .CP(ClockA), 
        .CDN(n2254), .Q(\SerDes_U1/Ser_U1/FIFO_Out [28]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2255), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [29]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ), .E(n2348), .CP(ClockA), 
        .CDN(n2182), .Q(\SerDes_U1/Ser_U1/FIFO_Out [30]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2250), 
        .Q(\SerDes_U1/Ser_U1/FIFO_Out [31]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        InParDataA[0]), .E(n2328), .CP(ClockA), .CDN(n2199), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2212), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2188), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2184), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        InParDataA[4]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2267), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        InParDataA[5]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2206), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        InParDataA[6]), .E(n2328), .CP(ClockA), .CDN(n2206), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        InParDataA[7]), .E(n2327), .CP(ClockA), .CDN(n2242), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        InParDataA[8]), .E(n2328), .CP(ClockA), .CDN(n2184), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        InParDataA[9]), .E(n2327), .CP(ClockA), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        InParDataA[10]), .E(n2327), .CP(ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        InParDataA[11]), .E(n2327), .CP(ClockA), .CDN(n2253), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        InParDataA[12]), .E(n2327), .CP(ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        InParDataA[13]), .E(n2327), .CP(ClockA), .CDN(n2261), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        InParDataA[14]), .E(n2327), .CP(ClockA), .CDN(n2255), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        InParDataA[15]), .E(n2327), .CP(ClockA), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        InParDataA[16]), .E(n2327), .CP(ClockA), .CDN(n2251), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        InParDataA[17]), .E(n2327), .CP(ClockA), .CDN(n2211), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        InParDataA[18]), .E(n2327), .CP(ClockA), .CDN(n2259), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        InParDataA[19]), .E(n2327), .CP(ClockA), .CDN(n2215), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        InParDataA[20]), .E(n2328), .CP(ClockA), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        InParDataA[21]), .E(n2328), .CP(ClockA), .CDN(n2198), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        InParDataA[22]), .E(n2328), .CP(ClockA), .CDN(n2236), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        InParDataA[23]), .E(n2328), .CP(ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        InParDataA[24]), .E(n2328), .CP(ClockA), .CDN(n2251), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        InParDataA[25]), .E(n2328), .CP(ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        InParDataA[26]), .E(n2328), .CP(ClockA), .CDN(n2270), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        InParDataA[27]), .E(n2328), .CP(ClockA), .CDN(n2184), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        InParDataA[28]), .E(n2328), .CP(ClockA), .CDN(n2234), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        InParDataA[29]), .E(n2328), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2245), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .CP(
        ClockA), .CDN(n2202), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        InParDataA[0]), .E(n2333), .CP(ClockA), .CDN(n2244), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2270), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        InParDataA[4]), .E(n2333), .CP(ClockA), .CDN(n2256), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        InParDataA[5]), .E(n2333), .CP(ClockA), .CDN(n2257), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        InParDataA[6]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2265), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        InParDataA[7]), .E(n2333), .CP(ClockA), .CDN(n2248), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        InParDataA[8]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        InParDataA[9]), .E(n2333), .CP(ClockA), .CDN(n2246), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        InParDataA[10]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2251), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        InParDataA[11]), .E(n2333), .CP(ClockA), .CDN(n2228), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        InParDataA[12]), .E(n2333), .CP(ClockA), .CDN(n2245), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        InParDataA[13]), .E(n2333), .CP(ClockA), .CDN(n2243), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        InParDataA[14]), .E(n2333), .CP(ClockA), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        InParDataA[15]), .E(n2333), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        InParDataA[16]), .E(n2333), .CP(ClockA), .CDN(n2253), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        InParDataA[17]), .E(n2333), .CP(ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        InParDataA[18]), .E(n2333), .CP(ClockA), .CDN(n2264), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        InParDataA[19]), .E(n2333), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        InParDataA[20]), .E(n2333), .CP(ClockA), .CDN(n2201), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        InParDataA[21]), .E(n2333), .CP(ClockA), .CDN(n2194), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        InParDataA[22]), .E(n2333), .CP(ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        InParDataA[23]), .E(n2333), .CP(ClockA), .CDN(n2255), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        InParDataA[24]), .E(n2333), .CP(ClockA), .CDN(n2209), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        InParDataA[25]), .E(n2333), .CP(ClockA), .CDN(n2238), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        InParDataA[26]), .E(n2333), .CP(ClockA), .CDN(n2220), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        InParDataA[27]), .E(n2333), .CP(ClockA), .CDN(n2229), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        InParDataA[28]), .E(n2333), .CP(ClockA), .CDN(n2248), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        InParDataA[29]), .E(n2333), .CP(ClockA), .CDN(n2204), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .CP(
        ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        InParDataA[0]), .E(n2342), .CP(ClockA), .CDN(n2200), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2213), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2221), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2194), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        InParDataA[4]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        InParDataA[5]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2192), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        InParDataA[6]), .E(n2342), .CP(ClockA), .CDN(n2207), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        InParDataA[7]), .E(n2341), .CP(ClockA), .CDN(n2195), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        InParDataA[8]), .E(n2342), .CP(ClockA), .CDN(n2261), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        InParDataA[9]), .E(n2341), .CP(ClockA), .CDN(n2261), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        InParDataA[10]), .E(n2341), .CP(ClockA), .CDN(n2264), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        InParDataA[11]), .E(n2341), .CP(ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        InParDataA[12]), .E(n2341), .CP(ClockA), .CDN(n2265), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        InParDataA[13]), .E(n2341), .CP(ClockA), .CDN(n2248), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        InParDataA[14]), .E(n2341), .CP(ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        InParDataA[15]), .E(n2341), .CP(ClockA), .CDN(n2246), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        InParDataA[16]), .E(n2341), .CP(ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        InParDataA[17]), .E(n2341), .CP(ClockA), .CDN(n2244), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        InParDataA[18]), .E(n2341), .CP(ClockA), .CDN(n2245), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        InParDataA[19]), .E(n2341), .CP(ClockA), .CDN(n2243), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        InParDataA[20]), .E(n2342), .CP(ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        InParDataA[21]), .E(n2342), .CP(ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        InParDataA[22]), .E(n2342), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        InParDataA[23]), .E(n2342), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        InParDataA[24]), .E(n2342), .CP(ClockA), .CDN(n2251), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        InParDataA[25]), .E(n2342), .CP(ClockA), .CDN(n2240), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        InParDataA[26]), .E(n2342), .CP(ClockA), .CDN(n2231), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        InParDataA[27]), .E(n2342), .CP(ClockA), .CDN(n2256), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        InParDataA[28]), .E(n2342), .CP(ClockA), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        InParDataA[29]), .E(n2342), .CP(ClockA), .CDN(n2217), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2255), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .CP(
        ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        InParDataA[0]), .E(n2337), .CP(ClockA), .CDN(n2240), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2237), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2190), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2242), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        InParDataA[4]), .E(n2337), .CP(ClockA), .CDN(n2246), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        InParDataA[5]), .E(n2337), .CP(ClockA), .CDN(n2241), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        InParDataA[6]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2219), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        InParDataA[7]), .E(n2337), .CP(ClockA), .CDN(n2211), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        InParDataA[8]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2233), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        InParDataA[9]), .E(n2337), .CP(ClockA), .CDN(n2251), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        InParDataA[10]), .E(n2337), .CP(ClockA), .CDN(n2239), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        InParDataA[11]), .E(n2337), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        InParDataA[12]), .E(n2337), .CP(ClockA), .CDN(n2220), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        InParDataA[13]), .E(n2337), .CP(ClockA), .CDN(n2239), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        InParDataA[14]), .E(n2337), .CP(ClockA), .CDN(n2219), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        InParDataA[15]), .E(n2337), .CP(ClockA), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        InParDataA[16]), .E(n2337), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        InParDataA[17]), .E(n2337), .CP(ClockA), .CDN(n2208), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        InParDataA[18]), .E(n2337), .CP(ClockA), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        InParDataA[19]), .E(n2337), .CP(ClockA), .CDN(n2214), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        InParDataA[20]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2267), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        InParDataA[21]), .E(n2337), .CP(ClockA), .CDN(n2241), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        InParDataA[22]), .E(n2337), .CP(ClockA), .CDN(n2264), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        InParDataA[23]), .E(n2337), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        InParDataA[24]), .E(n2337), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        InParDataA[25]), .E(n2337), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        InParDataA[26]), .E(n2337), .CP(ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        InParDataA[27]), .E(n2337), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        InParDataA[28]), .E(n2337), .CP(ClockA), .CDN(n2229), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        InParDataA[29]), .E(n2337), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2211), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .CP(
        ClockA), .CDN(n2216), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        InParDataA[0]), .E(n2339), .CP(ClockA), .CDN(n2233), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2270), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2205), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2188), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        InParDataA[4]), .E(n2339), .CP(ClockA), .CDN(n2242), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        InParDataA[5]), .E(n2339), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        InParDataA[6]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2241), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        InParDataA[7]), .E(n2339), .CP(ClockA), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        InParDataA[8]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        InParDataA[9]), .E(n2339), .CP(ClockA), .CDN(n2239), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        InParDataA[10]), .E(n2339), .CP(ClockA), .CDN(n2270), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        InParDataA[11]), .E(n2339), .CP(ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        InParDataA[12]), .E(n2339), .CP(ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        InParDataA[13]), .E(n2339), .CP(ClockA), .CDN(n2257), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        InParDataA[14]), .E(n2339), .CP(ClockA), .CDN(n2256), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        InParDataA[15]), .E(n2339), .CP(ClockA), .CDN(n2188), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        InParDataA[16]), .E(n2339), .CP(ClockA), .CDN(n2253), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        InParDataA[17]), .E(n2339), .CP(ClockA), .CDN(n2209), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        InParDataA[18]), .E(n2339), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        InParDataA[19]), .E(n2339), .CP(ClockA), .CDN(n2267), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        InParDataA[20]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2201), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        InParDataA[21]), .E(n2339), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        InParDataA[22]), .E(n2339), .CP(ClockA), .CDN(n2269), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        InParDataA[23]), .E(n2339), .CP(ClockA), .CDN(n2211), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        InParDataA[24]), .E(n2339), .CP(ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        InParDataA[25]), .E(n2339), .CP(ClockA), .CDN(n2228), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        InParDataA[26]), .E(n2339), .CP(ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        InParDataA[27]), .E(n2339), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        InParDataA[28]), .E(n2339), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        InParDataA[29]), .E(n2339), .CP(ClockA), .CDN(n1247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2203), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .CP(
        ClockA), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ) );
  DFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SDN(n2257), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]) );
  DFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SDN(n2229), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]) );
  DFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .SDN(n2256), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]) );
  DFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .SDN(n2189), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        InParDataA[0]), .E(n2331), .CP(ClockA), .CDN(n2200), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2256), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        InParDataA[4]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2185), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        InParDataA[5]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2210), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        InParDataA[6]), .E(n2331), .CP(ClockA), .CDN(n2199), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        InParDataA[7]), .E(n2330), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        InParDataA[8]), .E(n2331), .CP(ClockA), .CDN(n2242), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        InParDataA[9]), .E(n2330), .CP(ClockA), .CDN(n2218), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        InParDataA[10]), .E(n2330), .CP(ClockA), .CDN(n2217), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        InParDataA[11]), .E(n2330), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        InParDataA[12]), .E(n2330), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        InParDataA[13]), .E(n2330), .CP(ClockA), .CDN(n2241), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        InParDataA[14]), .E(n2330), .CP(ClockA), .CDN(n2218), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        InParDataA[15]), .E(n2330), .CP(ClockA), .CDN(n2202), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        InParDataA[16]), .E(n2330), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        InParDataA[17]), .E(n2330), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        InParDataA[18]), .E(n2330), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        InParDataA[19]), .E(n2330), .CP(ClockA), .CDN(n2199), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        InParDataA[20]), .E(n2331), .CP(ClockA), .CDN(n2211), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        InParDataA[21]), .E(n2331), .CP(ClockA), .CDN(n2187), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        InParDataA[22]), .E(n2331), .CP(ClockA), .CDN(n2197), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        InParDataA[23]), .E(n2331), .CP(ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        InParDataA[24]), .E(n2331), .CP(ClockA), .CDN(n2269), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        InParDataA[25]), .E(n2331), .CP(ClockA), .CDN(n2231), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        InParDataA[26]), .E(n2331), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        InParDataA[27]), .E(n2331), .CP(ClockA), .CDN(n2199), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        InParDataA[28]), .E(n2331), .CP(ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        InParDataA[29]), .E(n2331), .CP(ClockA), .CDN(n2197), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2235), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .CP(
        ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        InParDataA[0]), .E(n2335), .CP(ClockA), .CDN(n2217), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2267), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2269), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2235), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        InParDataA[4]), .E(n2335), .CP(ClockA), .CDN(n2257), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        InParDataA[5]), .E(n2335), .CP(ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        InParDataA[6]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        InParDataA[7]), .E(n2335), .CP(ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        InParDataA[8]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        InParDataA[9]), .E(n2335), .CP(ClockA), .CDN(n2229), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        InParDataA[10]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2243), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        InParDataA[11]), .E(n2335), .CP(ClockA), .CDN(n1247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        InParDataA[12]), .E(n2335), .CP(ClockA), .CDN(n2248), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        InParDataA[13]), .E(n2335), .CP(ClockA), .CDN(n2231), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        InParDataA[14]), .E(n2335), .CP(ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        InParDataA[15]), .E(n2335), .CP(ClockA), .CDN(n2262), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        InParDataA[16]), .E(n2335), .CP(ClockA), .CDN(n2257), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        InParDataA[17]), .E(n2335), .CP(ClockA), .CDN(n2256), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        InParDataA[18]), .E(n2335), .CP(ClockA), .CDN(n2189), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        InParDataA[19]), .E(n2335), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        InParDataA[20]), .E(n2335), .CP(ClockA), .CDN(n2245), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        InParDataA[21]), .E(n2335), .CP(ClockA), .CDN(n2265), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        InParDataA[22]), .E(n2335), .CP(ClockA), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        InParDataA[23]), .E(n2335), .CP(ClockA), .CDN(n2258), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        InParDataA[24]), .E(n2335), .CP(ClockA), .CDN(n2210), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        InParDataA[25]), .E(n2335), .CP(ClockA), .CDN(n2234), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        InParDataA[26]), .E(n2335), .CP(ClockA), .CDN(n2250), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        InParDataA[27]), .E(n2335), .CP(ClockA), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        InParDataA[28]), .E(n2335), .CP(ClockA), .CDN(n2224), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        InParDataA[29]), .E(n2335), .CP(ClockA), .CDN(n2269), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .CP(
        ClockA), .CDN(n2244), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        InParDataA[0]), .E(n2345), .CP(ClockA), .CDN(n2259), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        InParDataA[1]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2213), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        InParDataA[2]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2268), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        InParDataA[3]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2189), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        InParDataA[4]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2217), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        InParDataA[5]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        InParDataA[6]), .E(n2345), .CP(ClockA), .CDN(n2243), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        InParDataA[7]), .E(n2344), .CP(ClockA), .CDN(n2238), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        InParDataA[8]), .E(n2345), .CP(ClockA), .CDN(n2196), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        InParDataA[9]), .E(n2344), .CP(ClockA), .CDN(n2230), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        InParDataA[10]), .E(n2344), .CP(ClockA), .CDN(n2253), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        InParDataA[11]), .E(n2344), .CP(ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        InParDataA[12]), .E(n2344), .CP(ClockA), .CDN(n2244), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        InParDataA[13]), .E(n2344), .CP(ClockA), .CDN(n2245), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        InParDataA[14]), .E(n2344), .CP(ClockA), .CDN(n2243), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        InParDataA[15]), .E(n2344), .CP(ClockA), .CDN(n2265), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        InParDataA[16]), .E(n2344), .CP(ClockA), .CDN(n2248), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        InParDataA[17]), .E(n2344), .CP(ClockA), .CDN(n2247), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        InParDataA[18]), .E(n2344), .CP(ClockA), .CDN(n2246), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        InParDataA[19]), .E(n2344), .CP(ClockA), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        InParDataA[20]), .E(n2345), .CP(ClockA), .CDN(n2254), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        InParDataA[21]), .E(n2345), .CP(ClockA), .CDN(n2223), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        InParDataA[22]), .E(n2345), .CP(ClockA), .CDN(n2260), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        InParDataA[23]), .E(n2345), .CP(ClockA), .CDN(n2252), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        InParDataA[24]), .E(n2345), .CP(ClockA), .CDN(n2246), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        InParDataA[25]), .E(n2345), .CP(ClockA), .CDN(n2192), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        InParDataA[26]), .E(n2345), .CP(ClockA), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        InParDataA[27]), .E(n2345), .CP(ClockA), .CDN(n2182), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        InParDataA[28]), .E(n2345), .CP(ClockA), .CDN(n2208), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        InParDataA[29]), .E(n2345), .CP(ClockA), .CDN(n2257), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        InParDataA[30]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2266), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        InParDataA[31]), .E(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .CP(
        ClockA), .CDN(n2195), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[4]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N42 ), .E(\SerDes_U1/SerLineValid ), .CP(
        n2293), .CDN(n2261), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[4]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N42 ), .E(\SerDes_U2/SerLineValid ), .CP(
        n2285), .CDN(n2250), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ) );
  DFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1221), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(n2961) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[2]  ( .D(n1143), 
        .CPN(n2289), .CDN(n2189), .Q(n2955) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[2]  ( .D(n1052), 
        .CPN(n2283), .CDN(n2205), .Q(n2946) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n1121), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .CP(
        \SerDes_U2/Rx_ParClk ), .CDN(n1121), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[36]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[35] ), .CPN(n2294), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[51]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[36]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[35] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[51]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ), .CPN(n2275), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .E(n1298), .CP(ClockB), 
        .CDN(n2250), .Q(\SerDes_U2/Ser_U1/FIFO_Out [31]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ), .E(n1298), .CP(ClockB), 
        .CDN(n2266), .Q(\SerDes_U2/Ser_U1/FIFO_Out [30]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ), .E(n2425), .CP(ClockB), 
        .CDN(n2236), .Q(\SerDes_U2/Ser_U1/FIFO_Out [29]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ), .E(n1298), .CP(ClockB), 
        .CDN(n2235), .Q(\SerDes_U2/Ser_U1/FIFO_Out [28]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ), .E(n1298), .CP(ClockB), 
        .CDN(n2187), .Q(\SerDes_U2/Ser_U1/FIFO_Out [27]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ), .E(n1298), .CP(ClockB), 
        .CDN(n2193), .Q(\SerDes_U2/Ser_U1/FIFO_Out [26]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ), .E(n1298), .CP(ClockB), 
        .CDN(n2199), .Q(\SerDes_U2/Ser_U1/FIFO_Out [25]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ), .E(n1298), .CP(ClockB), 
        .CDN(n2228), .Q(\SerDes_U2/Ser_U1/FIFO_Out [24]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ), .E(n1298), .CP(ClockB), 
        .CDN(n2215), .Q(\SerDes_U2/Ser_U1/FIFO_Out [23]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ), .E(n1298), .CP(ClockB), 
        .CDN(n2266), .Q(\SerDes_U2/Ser_U1/FIFO_Out [22]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ), .E(n1298), .CP(ClockB), 
        .CDN(n2188), .Q(\SerDes_U2/Ser_U1/FIFO_Out [21]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ), .E(n2425), .CP(ClockB), 
        .CDN(n2263), .Q(\SerDes_U2/Ser_U1/FIFO_Out [20]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ), .E(n1298), .CP(ClockB), 
        .CDN(n2233), .Q(\SerDes_U2/Ser_U1/FIFO_Out [19]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ), .E(n1298), .CP(ClockB), 
        .CDN(n2267), .Q(\SerDes_U2/Ser_U1/FIFO_Out [18]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ), .E(n2425), .CP(ClockB), 
        .CDN(n2249), .Q(\SerDes_U2/Ser_U1/FIFO_Out [17]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ), .E(n1298), .CP(ClockB), 
        .CDN(n2200), .Q(\SerDes_U2/Ser_U1/FIFO_Out [16]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ), .E(n2425), .CP(ClockB), 
        .CDN(n2202), .Q(\SerDes_U2/Ser_U1/FIFO_Out [15]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ), .E(n1298), .CP(ClockB), 
        .CDN(n2215), .Q(\SerDes_U2/Ser_U1/FIFO_Out [14]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ), .E(n2425), .CP(ClockB), 
        .CDN(n2245), .Q(\SerDes_U2/Ser_U1/FIFO_Out [13]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ), .E(n1298), .CP(ClockB), 
        .CDN(n2192), .Q(\SerDes_U2/Ser_U1/FIFO_Out [12]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ), .E(n2425), .CP(ClockB), 
        .CDN(n2246), .Q(\SerDes_U2/Ser_U1/FIFO_Out [11]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ), .E(n1298), .CP(ClockB), 
        .CDN(n2267), .Q(\SerDes_U2/Ser_U1/FIFO_Out [10]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ), .E(n2425), .CP(ClockB), 
        .CDN(n2237), .Q(\SerDes_U2/Ser_U1/FIFO_Out [9]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ), .E(n2425), .CP(ClockB), 
        .CDN(n2197), .Q(\SerDes_U2/Ser_U1/FIFO_Out [8]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ), .E(n2425), .CP(ClockB), 
        .CDN(n2263), .Q(\SerDes_U2/Ser_U1/FIFO_Out [7]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ), .E(n2425), .CP(ClockB), 
        .CDN(n2187), .Q(\SerDes_U2/Ser_U1/FIFO_Out [6]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ), .E(n2425), .CP(ClockB), 
        .CDN(n2228), .Q(\SerDes_U2/Ser_U1/FIFO_Out [5]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ), .E(n2425), .CP(ClockB), 
        .CDN(n2230), .Q(\SerDes_U2/Ser_U1/FIFO_Out [4]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ), .E(n2425), .CP(ClockB), 
        .CDN(n2236), .Q(\SerDes_U2/Ser_U1/FIFO_Out [3]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ), .E(n2425), .CP(ClockB), 
        .CDN(n2227), .Q(\SerDes_U2/Ser_U1/FIFO_Out [2]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ), .E(n2425), .CP(ClockB), 
        .CDN(n2228), .Q(\SerDes_U2/Ser_U1/FIFO_Out [1]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ), .E(n2425), .CP(ClockB), 
        .CDN(n2226), .Q(\SerDes_U2/Ser_U1/FIFO_Out [0]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2234), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2233), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2234), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N2 ), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [1]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N3 ), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [2]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N4 ), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [3]) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[3]  ( .D(n1142), 
        .CPN(n2294), .CDN(n2189), .Q(n2958), .QN(n1312) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[3]  ( .D(n1051), 
        .CPN(n2286), .CDN(n2205), .Q(n2949), .QN(n1313) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n2228), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N2 ), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n2217), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [1]) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N3 ), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [2]) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N4 ), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n2217), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [3]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1212), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[52]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[52]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ), .CPN(n2275), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState_reg[2]  ( .D(n1044), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .Q(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .CP(
        \SerDes_U1/Rx_ParClk ), .CDN(n1212), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRxToDecode ), .CPN(n2289), .CDN(n2215), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[1]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ), .CPN(n2297), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[2]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ), .CPN(n2289), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[4]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ), .CPN(n2293), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[5]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ), .CPN(n2295), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRxToDecode ), .CPN(n2281), .CDN(n2198), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[1]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ), .CPN(n2281), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[2]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ), .CPN(n2281), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[4]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ), .CPN(n2281), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[5]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ), .CPN(n2281), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[6]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ), .CPN(n2295), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[16]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[15] ), .CPN(n2295), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[17]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ), .CPN(n2298), .CDN(n2214), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[20]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[19] ), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2214), .Q(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[21]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ), .CPN(n2296), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[23]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[22] ), .CPN(n2298), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[33]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[32] ), .CPN(n2294), .CDN(n2211), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[37]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ), .CPN(n2294), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[39]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[38] ), .CPN(n2294), .CDN(n2210), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[49]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[48] ), .CPN(n2293), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[50]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ), .CPN(n2293), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[54]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[53] ), .CPN(n2292), .CDN(n2209), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[6]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ), .CPN(n2280), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[16]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[15] ), .CPN(n2279), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[17]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[20]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[19] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[21]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[23]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[22] ), .CPN(n2279), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[33]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[32] ), .CPN(n2277), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[37]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[39]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[38] ), .CPN(n2277), .CDN(n2197), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[49]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[48] ), .CPN(n2276), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[50]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ), .CPN(n2276), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[54]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[53] ), .CPN(n2275), .CDN(n2196), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ) );
  DFCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), .Q(
        n2976), .QN(n1309) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[3]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ), .CPN(n2292), .CDN(n2213), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[3]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ), .CPN(n2281), .CDN(n2198), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR_reg[7]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ), .CPN(n2291), .CDN(n2212), 
        .Q(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR_reg[7]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ), .CPN(n2280), .CDN(n2199), 
        .Q(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[3]  ( .D(n1240), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .Q(n2963) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n1237), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .Q(n2964) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[3]  ( .D(n1236), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .Q(n2966) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/OldReadAr_reg[2]  ( .D(n1233), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), 
        .Q(n2965) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[3]  ( .D(n1133), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(n2951) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n1130), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(n2950) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[2]  ( .D(n1225), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(n2959) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/OldWriteAr_reg[1]  ( .D(n1223), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(n2960) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][31]  ( .D(
        InParDataB[31]), .E(n2385), .CP(ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2224), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2225), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][23]  ( .D(
        InParDataB[23]), .E(n2385), .CP(ClockB), .CDN(n2231), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][21]  ( .D(
        InParDataB[21]), .E(n2385), .CP(ClockB), .CDN(n2230), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][17]  ( .D(
        InParDataB[17]), .E(n2385), .CP(ClockB), .CDN(n2226), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][13]  ( .D(
        InParDataB[13]), .E(n2385), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][11]  ( .D(
        InParDataB[11]), .E(n2385), .CP(ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][9]  ( .D(
        InParDataB[9]), .E(n2385), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][7]  ( .D(
        InParDataB[7]), .E(n2385), .CP(ClockB), .CDN(n2199), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][5]  ( .D(
        InParDataB[5]), .E(n2385), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][3]  ( .D(
        InParDataB[3]), .E(n2385), .CP(ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][1]  ( .D(
        InParDataB[1]), .E(n2385), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][0]  ( .D(
        InParDataB[0]), .E(n2385), .CP(ClockB), .CDN(n2184), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][2]  ( .D(
        InParDataB[2]), .E(n2385), .CP(ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][4]  ( .D(
        InParDataB[4]), .E(n2385), .CP(ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][6]  ( .D(
        InParDataB[6]), .E(n2385), .CP(ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][10]  ( .D(
        InParDataB[10]), .E(n2385), .CP(ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][12]  ( .D(
        InParDataB[12]), .E(n2385), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][14]  ( .D(
        InParDataB[14]), .E(n2385), .CP(ClockB), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][16]  ( .D(
        InParDataB[16]), .E(n2385), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][18]  ( .D(
        InParDataB[18]), .E(n2385), .CP(ClockB), .CDN(n2231), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][20]  ( .D(
        InParDataB[20]), .E(n2385), .CP(ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][22]  ( .D(
        InParDataB[22]), .E(n2385), .CP(ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][24]  ( .D(
        InParDataB[24]), .E(n2385), .CP(ClockB), .CDN(n2199), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][26]  ( .D(
        InParDataB[26]), .E(n2385), .CP(ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[14][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .CP(
        ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][31]  ( .D(
        InParDataB[31]), .E(n2383), .CP(ClockB), .CDN(n2206), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][23]  ( .D(
        InParDataB[23]), .E(n2383), .CP(ClockB), .CDN(n2254), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][21]  ( .D(
        InParDataB[21]), .E(n2383), .CP(ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][17]  ( .D(
        InParDataB[17]), .E(n2383), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2206), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][13]  ( .D(
        InParDataB[13]), .E(n2383), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][11]  ( .D(
        InParDataB[11]), .E(n2383), .CP(ClockB), .CDN(n2192), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][9]  ( .D(
        InParDataB[9]), .E(n2383), .CP(ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][7]  ( .D(
        InParDataB[7]), .E(n2383), .CP(ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][5]  ( .D(
        InParDataB[5]), .E(n2383), .CP(ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][3]  ( .D(
        InParDataB[3]), .E(n2383), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][1]  ( .D(
        InParDataB[1]), .E(n2383), .CP(ClockB), .CDN(n2215), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][0]  ( .D(
        InParDataB[0]), .E(n2383), .CP(ClockB), .CDN(n2233), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][2]  ( .D(
        InParDataB[2]), .E(n2383), .CP(ClockB), .CDN(n2200), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][4]  ( .D(
        InParDataB[4]), .E(n2383), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][6]  ( .D(
        InParDataB[6]), .E(n2383), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][10]  ( .D(
        InParDataB[10]), .E(n2383), .CP(ClockB), .CDN(n2223), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][12]  ( .D(
        InParDataB[12]), .E(n2383), .CP(ClockB), .CDN(n2207), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][14]  ( .D(
        InParDataB[14]), .E(n2383), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][16]  ( .D(
        InParDataB[16]), .E(n2383), .CP(ClockB), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][18]  ( .D(
        InParDataB[18]), .E(n2383), .CP(ClockB), .CDN(n2233), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][20]  ( .D(
        InParDataB[20]), .E(n2383), .CP(ClockB), .CDN(n2198), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][22]  ( .D(
        InParDataB[22]), .E(n2383), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][24]  ( .D(
        InParDataB[24]), .E(n2383), .CP(ClockB), .CDN(n2189), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][26]  ( .D(
        InParDataB[26]), .E(n2383), .CP(ClockB), .CDN(n2234), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[13][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .CP(
        ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][31]  ( .D(
        InParDataB[31]), .E(n2377), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2230), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][23]  ( .D(
        InParDataB[23]), .E(n2377), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][21]  ( .D(
        InParDataB[21]), .E(n2377), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][17]  ( .D(
        InParDataB[17]), .E(n2377), .CP(ClockB), .CDN(n2249), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][13]  ( .D(
        InParDataB[13]), .E(n2377), .CP(ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][11]  ( .D(
        InParDataB[11]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][9]  ( .D(
        InParDataB[9]), .E(n2377), .CP(ClockB), .CDN(n2223), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][7]  ( .D(
        InParDataB[7]), .E(n2377), .CP(ClockB), .CDN(n2260), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][5]  ( .D(
        InParDataB[5]), .E(n2377), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][3]  ( .D(
        InParDataB[3]), .E(n2377), .CP(ClockB), .CDN(n2239), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][1]  ( .D(
        InParDataB[1]), .E(n2377), .CP(ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][0]  ( .D(
        InParDataB[0]), .E(n2377), .CP(ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][2]  ( .D(
        InParDataB[2]), .E(n2377), .CP(ClockB), .CDN(n2263), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][4]  ( .D(
        InParDataB[4]), .E(n2377), .CP(ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][6]  ( .D(
        InParDataB[6]), .E(n2377), .CP(ClockB), .CDN(n2257), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][8]  ( .D(
        InParDataB[8]), .E(n2377), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][10]  ( .D(
        InParDataB[10]), .E(n2377), .CP(ClockB), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][12]  ( .D(
        InParDataB[12]), .E(n2377), .CP(ClockB), .CDN(n2234), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][14]  ( .D(
        InParDataB[14]), .E(n2377), .CP(ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][16]  ( .D(
        InParDataB[16]), .E(n2377), .CP(ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][18]  ( .D(
        InParDataB[18]), .E(n2377), .CP(ClockB), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][20]  ( .D(
        InParDataB[20]), .E(n2377), .CP(ClockB), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][22]  ( .D(
        InParDataB[22]), .E(n2377), .CP(ClockB), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][24]  ( .D(
        InParDataB[24]), .E(n2377), .CP(ClockB), .CDN(n2223), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][26]  ( .D(
        InParDataB[26]), .E(n2377), .CP(ClockB), .CDN(n2224), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2225), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[10][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .CP(
        ClockB), .CDN(n2232), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][31]  ( .D(
        InParDataB[31]), .E(n2375), .CP(ClockB), .CDN(n2198), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2211), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][23]  ( .D(
        InParDataB[23]), .E(n2375), .CP(ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][21]  ( .D(
        InParDataB[21]), .E(n2375), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][19]  ( .D(
        InParDataB[19]), .E(n2375), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2234), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][15]  ( .D(
        InParDataB[15]), .E(n2375), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][11]  ( .D(
        InParDataB[11]), .E(n2375), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][9]  ( .D(
        InParDataB[9]), .E(n2375), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][7]  ( .D(
        InParDataB[7]), .E(n2375), .CP(ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][5]  ( .D(
        InParDataB[5]), .E(n2375), .CP(ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][3]  ( .D(
        InParDataB[3]), .E(n2375), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][1]  ( .D(
        InParDataB[1]), .E(n2375), .CP(ClockB), .CDN(n2211), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][0]  ( .D(
        InParDataB[0]), .E(n2375), .CP(ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][2]  ( .D(
        InParDataB[2]), .E(n2375), .CP(ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][4]  ( .D(
        InParDataB[4]), .E(n2375), .CP(ClockB), .CDN(n2232), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][6]  ( .D(
        InParDataB[6]), .E(n2375), .CP(ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2192), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][10]  ( .D(
        InParDataB[10]), .E(n2375), .CP(ClockB), .CDN(n2231), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][12]  ( .D(
        InParDataB[12]), .E(n2375), .CP(ClockB), .CDN(n2210), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][14]  ( .D(
        InParDataB[14]), .E(n2375), .CP(ClockB), .CDN(n2209), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][16]  ( .D(
        InParDataB[16]), .E(n2375), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][18]  ( .D(
        InParDataB[18]), .E(n2375), .CP(ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][20]  ( .D(
        InParDataB[20]), .E(n2375), .CP(ClockB), .CDN(n2206), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][22]  ( .D(
        InParDataB[22]), .E(n2375), .CP(ClockB), .CDN(n2207), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][24]  ( .D(
        InParDataB[24]), .E(n2375), .CP(ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][26]  ( .D(
        InParDataB[26]), .E(n2375), .CP(ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2204), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[9][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .CP(
        ClockB), .CDN(n2200), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][31]  ( .D(
        InParDataB[31]), .E(n2369), .CP(ClockB), .CDN(n2184), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n1247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][23]  ( .D(
        InParDataB[23]), .E(n2369), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][21]  ( .D(
        InParDataB[21]), .E(n2369), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][17]  ( .D(
        InParDataB[17]), .E(n2369), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2223), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][13]  ( .D(
        InParDataB[13]), .E(n2369), .CP(ClockB), .CDN(n2263), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][11]  ( .D(
        InParDataB[11]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][9]  ( .D(
        InParDataB[9]), .E(n2369), .CP(ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][7]  ( .D(
        InParDataB[7]), .E(n2369), .CP(ClockB), .CDN(n2257), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][5]  ( .D(
        InParDataB[5]), .E(n2369), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][3]  ( .D(
        InParDataB[3]), .E(n2369), .CP(ClockB), .CDN(n1247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][1]  ( .D(
        InParDataB[1]), .E(n2369), .CP(ClockB), .CDN(n2182), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][0]  ( .D(
        InParDataB[0]), .E(n2369), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][2]  ( .D(
        InParDataB[2]), .E(n2369), .CP(ClockB), .CDN(n2268), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][4]  ( .D(
        InParDataB[4]), .E(n2369), .CP(ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][6]  ( .D(
        InParDataB[6]), .E(n2369), .CP(ClockB), .CDN(n2249), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][8]  ( .D(
        InParDataB[8]), .E(n2369), .CP(ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][10]  ( .D(
        InParDataB[10]), .E(n2369), .CP(ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][12]  ( .D(
        InParDataB[12]), .E(n2369), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][14]  ( .D(
        InParDataB[14]), .E(n2369), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][16]  ( .D(
        InParDataB[16]), .E(n2369), .CP(ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][18]  ( .D(
        InParDataB[18]), .E(n2369), .CP(ClockB), .CDN(n2199), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][20]  ( .D(
        InParDataB[20]), .E(n2369), .CP(ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][22]  ( .D(
        InParDataB[22]), .E(n2369), .CP(ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][24]  ( .D(
        InParDataB[24]), .E(n2369), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][26]  ( .D(
        InParDataB[26]), .E(n2369), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[6][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .CP(
        ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][31]  ( .D(
        InParDataB[31]), .E(n2367), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][23]  ( .D(
        InParDataB[23]), .E(n2367), .CP(ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][21]  ( .D(
        InParDataB[21]), .E(n2367), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][19]  ( .D(
        InParDataB[19]), .E(n2367), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][15]  ( .D(
        InParDataB[15]), .E(n2367), .CP(ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2204), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][11]  ( .D(
        InParDataB[11]), .E(n2367), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][9]  ( .D(
        InParDataB[9]), .E(n2367), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][7]  ( .D(
        InParDataB[7]), .E(n2367), .CP(ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][5]  ( .D(
        InParDataB[5]), .E(n2367), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][3]  ( .D(
        InParDataB[3]), .E(n2367), .CP(ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][1]  ( .D(
        InParDataB[1]), .E(n2367), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][0]  ( .D(
        InParDataB[0]), .E(n2367), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][2]  ( .D(
        InParDataB[2]), .E(n2367), .CP(ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][4]  ( .D(
        InParDataB[4]), .E(n2367), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][6]  ( .D(
        InParDataB[6]), .E(n2367), .CP(ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2254), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][10]  ( .D(
        InParDataB[10]), .E(n2367), .CP(ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][12]  ( .D(
        InParDataB[12]), .E(n2367), .CP(ClockB), .CDN(n2250), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][14]  ( .D(
        InParDataB[14]), .E(n2367), .CP(ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][16]  ( .D(
        InParDataB[16]), .E(n2367), .CP(ClockB), .CDN(n2230), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][18]  ( .D(
        InParDataB[18]), .E(n2367), .CP(ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][20]  ( .D(
        InParDataB[20]), .E(n2367), .CP(ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][22]  ( .D(
        InParDataB[22]), .E(n2367), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][24]  ( .D(
        InParDataB[24]), .E(n2367), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][26]  ( .D(
        InParDataB[26]), .E(n2367), .CP(ClockB), .CDN(n2197), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[5][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .CP(
        ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][31]  ( .D(
        InParDataB[31]), .E(n2361), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2195), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][23]  ( .D(
        InParDataB[23]), .E(n2361), .CP(ClockB), .CDN(n2198), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][21]  ( .D(
        InParDataB[21]), .E(n2361), .CP(ClockB), .CDN(n2199), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][19]  ( .D(
        InParDataB[19]), .E(n2361), .CP(ClockB), .CDN(n2197), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][15]  ( .D(
        InParDataB[15]), .E(n2361), .CP(ClockB), .CDN(n2197), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2229), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][11]  ( .D(
        InParDataB[11]), .E(n2361), .CP(ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][9]  ( .D(
        InParDataB[9]), .E(n2361), .CP(ClockB), .CDN(n2226), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][7]  ( .D(
        InParDataB[7]), .E(n2361), .CP(ClockB), .CDN(n2260), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][5]  ( .D(
        InParDataB[5]), .E(n2361), .CP(ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][3]  ( .D(
        InParDataB[3]), .E(n2361), .CP(ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][1]  ( .D(
        InParDataB[1]), .E(n2361), .CP(ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][0]  ( .D(
        InParDataB[0]), .E(n2361), .CP(ClockB), .CDN(n2268), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][2]  ( .D(
        InParDataB[2]), .E(n2361), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][4]  ( .D(
        InParDataB[4]), .E(n2361), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][6]  ( .D(
        InParDataB[6]), .E(n2361), .CP(ClockB), .CDN(n2268), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][10]  ( .D(
        InParDataB[10]), .E(n2361), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][12]  ( .D(
        InParDataB[12]), .E(n2361), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][14]  ( .D(
        InParDataB[14]), .E(n2361), .CP(ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][16]  ( .D(
        InParDataB[16]), .E(n2361), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][18]  ( .D(
        InParDataB[18]), .E(n2361), .CP(ClockB), .CDN(n2260), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][20]  ( .D(
        InParDataB[20]), .E(n2361), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][22]  ( .D(
        InParDataB[22]), .E(n2361), .CP(ClockB), .CDN(n1247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][24]  ( .D(
        InParDataB[24]), .E(n2361), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][26]  ( .D(
        InParDataB[26]), .E(n2361), .CP(ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[2][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .CP(
        ClockB), .CDN(n2206), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][31]  ( .D(
        InParDataB[31]), .E(n2359), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2230), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][23]  ( .D(
        InParDataB[23]), .E(n2359), .CP(ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][21]  ( .D(
        InParDataB[21]), .E(n2359), .CP(ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][17]  ( .D(
        InParDataB[17]), .E(n2359), .CP(ClockB), .CDN(n2190), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2182), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][13]  ( .D(
        InParDataB[13]), .E(n2359), .CP(ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][11]  ( .D(
        InParDataB[11]), .E(n2359), .CP(ClockB), .CDN(n2189), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][9]  ( .D(
        InParDataB[9]), .E(n2359), .CP(ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][7]  ( .D(
        InParDataB[7]), .E(n2359), .CP(ClockB), .CDN(n2240), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][5]  ( .D(
        InParDataB[5]), .E(n2359), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][3]  ( .D(
        InParDataB[3]), .E(n2359), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][1]  ( .D(
        InParDataB[1]), .E(n2359), .CP(ClockB), .CDN(n2225), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][0]  ( .D(
        InParDataB[0]), .E(n2359), .CP(ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][2]  ( .D(
        InParDataB[2]), .E(n2359), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][4]  ( .D(
        InParDataB[4]), .E(n2359), .CP(ClockB), .CDN(n2207), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][6]  ( .D(
        InParDataB[6]), .E(n2359), .CP(ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][10]  ( .D(
        InParDataB[10]), .E(n2359), .CP(ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][12]  ( .D(
        InParDataB[12]), .E(n2359), .CP(ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][14]  ( .D(
        InParDataB[14]), .E(n2359), .CP(ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][16]  ( .D(
        InParDataB[16]), .E(n2359), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][18]  ( .D(
        InParDataB[18]), .E(n2359), .CP(ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][20]  ( .D(
        InParDataB[20]), .E(n2359), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][22]  ( .D(
        InParDataB[22]), .E(n2359), .CP(ClockB), .CDN(n2209), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][24]  ( .D(
        InParDataB[24]), .E(n2359), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][26]  ( .D(
        InParDataB[26]), .E(n2359), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2257), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[1][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .CP(
        ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[3]  ( .D(n1129), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(n2952) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/OldReadAr_reg[1]  ( .D(n1128), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(n2953) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][31]  ( .D(
        InParDataB[31]), .E(n2387), .CP(ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n1247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][23]  ( .D(
        InParDataB[23]), .E(n2387), .CP(ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][21]  ( .D(
        InParDataB[21]), .E(n2387), .CP(ClockB), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][19]  ( .D(
        InParDataB[19]), .E(n2387), .CP(ClockB), .CDN(n2240), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2185), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][15]  ( .D(
        InParDataB[15]), .E(n2387), .CP(ClockB), .CDN(n2238), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][11]  ( .D(
        InParDataB[11]), .E(n2387), .CP(ClockB), .CDN(n2210), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][9]  ( .D(
        InParDataB[9]), .E(n2387), .CP(ClockB), .CDN(n2182), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][7]  ( .D(
        InParDataB[7]), .E(n2387), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][5]  ( .D(
        InParDataB[5]), .E(n2387), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][3]  ( .D(
        InParDataB[3]), .E(n2387), .CP(ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][1]  ( .D(
        InParDataB[1]), .E(n2387), .CP(ClockB), .CDN(n2226), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][0]  ( .D(
        InParDataB[0]), .E(n2387), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][2]  ( .D(
        InParDataB[2]), .E(n2387), .CP(ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][4]  ( .D(
        InParDataB[4]), .E(n2387), .CP(ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][6]  ( .D(
        InParDataB[6]), .E(n2387), .CP(ClockB), .CDN(n2257), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2223), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][10]  ( .D(
        InParDataB[10]), .E(n2387), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][12]  ( .D(
        InParDataB[12]), .E(n2387), .CP(ClockB), .CDN(n2192), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][14]  ( .D(
        InParDataB[14]), .E(n2387), .CP(ClockB), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][16]  ( .D(
        InParDataB[16]), .E(n2387), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][18]  ( .D(
        InParDataB[18]), .E(n2387), .CP(ClockB), .CDN(n2215), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][20]  ( .D(
        InParDataB[20]), .E(n2387), .CP(ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][22]  ( .D(
        InParDataB[22]), .E(n2387), .CP(ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][24]  ( .D(
        InParDataB[24]), .E(n2387), .CP(ClockB), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][26]  ( .D(
        InParDataB[26]), .E(n2387), .CP(ClockB), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[15][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .CP(
        ClockB), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][31]  ( .D(
        InParDataB[31]), .E(n2381), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2185), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][23]  ( .D(
        InParDataB[23]), .E(n2381), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][21]  ( .D(
        InParDataB[21]), .E(n2381), .CP(ClockB), .CDN(n2232), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][19]  ( .D(
        InParDataB[19]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][17]  ( .D(
        InParDataB[17]), .E(n2381), .CP(ClockB), .CDN(n2196), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][15]  ( .D(
        InParDataB[15]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][13]  ( .D(
        InParDataB[13]), .E(n2381), .CP(ClockB), .CDN(n2195), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][11]  ( .D(
        InParDataB[11]), .E(n2381), .CP(ClockB), .CDN(n2250), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][9]  ( .D(
        InParDataB[9]), .E(n2381), .CP(ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][7]  ( .D(
        InParDataB[7]), .E(n2381), .CP(ClockB), .CDN(n2187), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][5]  ( .D(
        InParDataB[5]), .E(n2381), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][3]  ( .D(
        InParDataB[3]), .E(n2381), .CP(ClockB), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][1]  ( .D(
        InParDataB[1]), .E(n2381), .CP(ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][0]  ( .D(
        InParDataB[0]), .E(n2381), .CP(ClockB), .CDN(n2230), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][2]  ( .D(
        InParDataB[2]), .E(n2381), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][4]  ( .D(
        InParDataB[4]), .E(n2381), .CP(ClockB), .CDN(n2232), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][6]  ( .D(
        InParDataB[6]), .E(n2381), .CP(ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][10]  ( .D(
        InParDataB[10]), .E(n2381), .CP(ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][12]  ( .D(
        InParDataB[12]), .E(n2381), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][14]  ( .D(
        InParDataB[14]), .E(n2381), .CP(ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][16]  ( .D(
        InParDataB[16]), .E(n2381), .CP(ClockB), .CDN(n2192), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][18]  ( .D(
        InParDataB[18]), .E(n2381), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][20]  ( .D(
        InParDataB[20]), .E(n2381), .CP(ClockB), .CDN(n2219), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][22]  ( .D(
        InParDataB[22]), .E(n2381), .CP(ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][24]  ( .D(
        InParDataB[24]), .E(n2381), .CP(ClockB), .CDN(n2192), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][26]  ( .D(
        InParDataB[26]), .E(n2381), .CP(ClockB), .CDN(n2190), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2242), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[12][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .CP(
        ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][31]  ( .D(
        InParDataB[31]), .E(n2379), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2260), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2211), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2235), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][23]  ( .D(
        InParDataB[23]), .E(n2379), .CP(ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][21]  ( .D(
        InParDataB[21]), .E(n2379), .CP(ClockB), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][19]  ( .D(
        InParDataB[19]), .E(n2379), .CP(ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][15]  ( .D(
        InParDataB[15]), .E(n2379), .CP(ClockB), .CDN(n2238), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2239), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][11]  ( .D(
        InParDataB[11]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][9]  ( .D(
        InParDataB[9]), .E(n2379), .CP(ClockB), .CDN(n2197), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][7]  ( .D(
        InParDataB[7]), .E(n2379), .CP(ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][5]  ( .D(
        InParDataB[5]), .E(n2379), .CP(ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][3]  ( .D(
        InParDataB[3]), .E(n2379), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][1]  ( .D(
        InParDataB[1]), .E(n2379), .CP(ClockB), .CDN(n2250), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][0]  ( .D(
        InParDataB[0]), .E(n2379), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][2]  ( .D(
        InParDataB[2]), .E(n2379), .CP(ClockB), .CDN(n2264), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][4]  ( .D(
        InParDataB[4]), .E(n2379), .CP(ClockB), .CDN(n2254), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][6]  ( .D(
        InParDataB[6]), .E(n2379), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][8]  ( .D(
        InParDataB[8]), .E(n2379), .CP(ClockB), .CDN(n2259), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][10]  ( .D(
        InParDataB[10]), .E(n2379), .CP(ClockB), .CDN(n2190), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][12]  ( .D(
        InParDataB[12]), .E(n2379), .CP(ClockB), .CDN(n2234), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][14]  ( .D(
        InParDataB[14]), .E(n2379), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][16]  ( .D(
        InParDataB[16]), .E(n2379), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][18]  ( .D(
        InParDataB[18]), .E(n2379), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][20]  ( .D(
        InParDataB[20]), .E(n2379), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][22]  ( .D(
        InParDataB[22]), .E(n2379), .CP(ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][24]  ( .D(
        InParDataB[24]), .E(n2379), .CP(ClockB), .CDN(n2184), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][26]  ( .D(
        InParDataB[26]), .E(n2379), .CP(ClockB), .CDN(n2185), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[11][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .CP(
        ClockB), .CDN(n2187), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][31]  ( .D(
        InParDataB[31]), .E(n2373), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2220), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][23]  ( .D(
        InParDataB[23]), .E(n2373), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][21]  ( .D(
        InParDataB[21]), .E(n2373), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][19]  ( .D(
        InParDataB[19]), .E(n2373), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][15]  ( .D(
        InParDataB[15]), .E(n2373), .CP(ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][11]  ( .D(
        InParDataB[11]), .E(n2373), .CP(ClockB), .CDN(n2218), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][9]  ( .D(
        InParDataB[9]), .E(n2373), .CP(ClockB), .CDN(n2216), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][7]  ( .D(
        InParDataB[7]), .E(n2373), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][5]  ( .D(
        InParDataB[5]), .E(n2373), .CP(ClockB), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][3]  ( .D(
        InParDataB[3]), .E(n2373), .CP(ClockB), .CDN(n2240), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][1]  ( .D(
        InParDataB[1]), .E(n2373), .CP(ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][0]  ( .D(
        InParDataB[0]), .E(n2373), .CP(ClockB), .CDN(n2239), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][2]  ( .D(
        InParDataB[2]), .E(n2373), .CP(ClockB), .CDN(n2238), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][4]  ( .D(
        InParDataB[4]), .E(n2373), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][6]  ( .D(
        InParDataB[6]), .E(n2373), .CP(ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][10]  ( .D(
        InParDataB[10]), .E(n2373), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][12]  ( .D(
        InParDataB[12]), .E(n2373), .CP(ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][14]  ( .D(
        InParDataB[14]), .E(n2373), .CP(ClockB), .CDN(n2240), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][16]  ( .D(
        InParDataB[16]), .E(n2373), .CP(ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][18]  ( .D(
        InParDataB[18]), .E(n2373), .CP(ClockB), .CDN(n2233), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][20]  ( .D(
        InParDataB[20]), .E(n2373), .CP(ClockB), .CDN(n2195), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][22]  ( .D(
        InParDataB[22]), .E(n2373), .CP(ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][24]  ( .D(
        InParDataB[24]), .E(n2373), .CP(ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][26]  ( .D(
        InParDataB[26]), .E(n2373), .CP(ClockB), .CDN(n2222), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[8][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .CP(
        ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][31]  ( .D(
        InParDataB[31]), .E(n2371), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2258), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][23]  ( .D(
        InParDataB[23]), .E(n2371), .CP(ClockB), .CDN(n2195), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][21]  ( .D(
        InParDataB[21]), .E(n2371), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][19]  ( .D(
        InParDataB[19]), .E(n2371), .CP(ClockB), .CDN(n2187), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2254), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][15]  ( .D(
        InParDataB[15]), .E(n2371), .CP(ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][11]  ( .D(
        InParDataB[11]), .E(n2371), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][9]  ( .D(
        InParDataB[9]), .E(n2371), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][7]  ( .D(
        InParDataB[7]), .E(n2371), .CP(ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][5]  ( .D(
        InParDataB[5]), .E(n2371), .CP(ClockB), .CDN(n2246), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][3]  ( .D(
        InParDataB[3]), .E(n2371), .CP(ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][1]  ( .D(
        InParDataB[1]), .E(n2371), .CP(ClockB), .CDN(n2224), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][0]  ( .D(
        InParDataB[0]), .E(n2371), .CP(ClockB), .CDN(n2249), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][2]  ( .D(
        InParDataB[2]), .E(n2371), .CP(ClockB), .CDN(n2225), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][4]  ( .D(
        InParDataB[4]), .E(n2371), .CP(ClockB), .CDN(n2263), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][6]  ( .D(
        InParDataB[6]), .E(n2371), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][10]  ( .D(
        InParDataB[10]), .E(n2371), .CP(ClockB), .CDN(n2239), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][12]  ( .D(
        InParDataB[12]), .E(n2371), .CP(ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][14]  ( .D(
        InParDataB[14]), .E(n2371), .CP(ClockB), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][16]  ( .D(
        InParDataB[16]), .E(n2371), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][18]  ( .D(
        InParDataB[18]), .E(n2371), .CP(ClockB), .CDN(n2232), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][20]  ( .D(
        InParDataB[20]), .E(n2371), .CP(ClockB), .CDN(n2238), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][22]  ( .D(
        InParDataB[22]), .E(n2371), .CP(ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][24]  ( .D(
        InParDataB[24]), .E(n2371), .CP(ClockB), .CDN(n2250), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][26]  ( .D(
        InParDataB[26]), .E(n2371), .CP(ClockB), .CDN(n2249), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[7][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .CP(
        ClockB), .CDN(n2263), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][31]  ( .D(
        InParDataB[31]), .E(n2365), .CP(ClockB), .CDN(n2249), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2250), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2234), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][23]  ( .D(
        InParDataB[23]), .E(n2365), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][21]  ( .D(
        InParDataB[21]), .E(n2365), .CP(ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][19]  ( .D(
        InParDataB[19]), .E(n2365), .CP(ClockB), .CDN(n2262), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][15]  ( .D(
        InParDataB[15]), .E(n2365), .CP(ClockB), .CDN(n2224), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][11]  ( .D(
        InParDataB[11]), .E(n2365), .CP(ClockB), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][9]  ( .D(
        InParDataB[9]), .E(n2365), .CP(ClockB), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][7]  ( .D(
        InParDataB[7]), .E(n2365), .CP(ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][5]  ( .D(
        InParDataB[5]), .E(n2365), .CP(ClockB), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][3]  ( .D(
        InParDataB[3]), .E(n2365), .CP(ClockB), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][1]  ( .D(
        InParDataB[1]), .E(n2365), .CP(ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][0]  ( .D(
        InParDataB[0]), .E(n2365), .CP(ClockB), .CDN(n2244), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][2]  ( .D(
        InParDataB[2]), .E(n2365), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][4]  ( .D(
        InParDataB[4]), .E(n2365), .CP(ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][6]  ( .D(
        InParDataB[6]), .E(n2365), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][10]  ( .D(
        InParDataB[10]), .E(n2365), .CP(ClockB), .CDN(n2217), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][12]  ( .D(
        InParDataB[12]), .E(n2365), .CP(ClockB), .CDN(n2253), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][14]  ( .D(
        InParDataB[14]), .E(n2365), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][16]  ( .D(
        InParDataB[16]), .E(n2365), .CP(ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][18]  ( .D(
        InParDataB[18]), .E(n2365), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][20]  ( .D(
        InParDataB[20]), .E(n2365), .CP(ClockB), .CDN(n2182), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][22]  ( .D(
        InParDataB[22]), .E(n2365), .CP(ClockB), .CDN(n2199), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][24]  ( .D(
        InParDataB[24]), .E(n2365), .CP(ClockB), .CDN(n2211), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][26]  ( .D(
        InParDataB[26]), .E(n2365), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[4][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .CP(
        ClockB), .CDN(n2198), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][31]  ( .D(
        InParDataB[31]), .E(n2363), .CP(ClockB), .CDN(n2226), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2241), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2215), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][23]  ( .D(
        InParDataB[23]), .E(n2363), .CP(ClockB), .CDN(n2200), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][21]  ( .D(
        InParDataB[21]), .E(n2363), .CP(ClockB), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][19]  ( .D(
        InParDataB[19]), .E(n2363), .CP(ClockB), .CDN(n2209), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2266), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][15]  ( .D(
        InParDataB[15]), .E(n2363), .CP(ClockB), .CDN(n2204), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2205), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][11]  ( .D(
        InParDataB[11]), .E(n2363), .CP(ClockB), .CDN(n2208), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][9]  ( .D(
        InParDataB[9]), .E(n2363), .CP(ClockB), .CDN(n2207), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][7]  ( .D(
        InParDataB[7]), .E(n2363), .CP(ClockB), .CDN(n2206), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][5]  ( .D(
        InParDataB[5]), .E(n2363), .CP(ClockB), .CDN(n2212), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][3]  ( .D(
        InParDataB[3]), .E(n2363), .CP(ClockB), .CDN(n2214), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][1]  ( .D(
        InParDataB[1]), .E(n2363), .CP(ClockB), .CDN(n2213), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][0]  ( .D(
        InParDataB[0]), .E(n2363), .CP(ClockB), .CDN(n2211), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][2]  ( .D(
        InParDataB[2]), .E(n2363), .CP(ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][4]  ( .D(
        InParDataB[4]), .E(n2363), .CP(ClockB), .CDN(n2216), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][6]  ( .D(
        InParDataB[6]), .E(n2363), .CP(ClockB), .CDN(n2183), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2184), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][10]  ( .D(
        InParDataB[10]), .E(n2363), .CP(ClockB), .CDN(n2185), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][12]  ( .D(
        InParDataB[12]), .E(n2363), .CP(ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][14]  ( .D(
        InParDataB[14]), .E(n2363), .CP(ClockB), .CDN(n2187), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][16]  ( .D(
        InParDataB[16]), .E(n2363), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][18]  ( .D(
        InParDataB[18]), .E(n2363), .CP(ClockB), .CDN(n2189), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][20]  ( .D(
        InParDataB[20]), .E(n2363), .CP(ClockB), .CDN(n2190), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][22]  ( .D(
        InParDataB[22]), .E(n2363), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][24]  ( .D(
        InParDataB[24]), .E(n2363), .CP(ClockB), .CDN(n2215), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][26]  ( .D(
        InParDataB[26]), .E(n2363), .CP(ClockB), .CDN(n2268), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2265), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[3][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .CP(
        ClockB), .CDN(n2248), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][31]  ( .D(
        InParDataB[31]), .E(n2357), .CP(ClockB), .CDN(n2252), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][29]  ( .D(
        InParDataB[29]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2268), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][27]  ( .D(
        InParDataB[27]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][25]  ( .D(
        InParDataB[25]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2191), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][23]  ( .D(
        InParDataB[23]), .E(n2357), .CP(ClockB), .CDN(n2243), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][21]  ( .D(
        InParDataB[21]), .E(n2357), .CP(ClockB), .CDN(n2270), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][19]  ( .D(
        InParDataB[19]), .E(n2357), .CP(ClockB), .CDN(n2256), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][17]  ( .D(
        InParDataB[17]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2255), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][15]  ( .D(
        InParDataB[15]), .E(n2357), .CP(ClockB), .CDN(n2251), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][13]  ( .D(
        InParDataB[13]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n1247), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][11]  ( .D(
        InParDataB[11]), .E(n2357), .CP(ClockB), .CDN(n2257), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][9]  ( .D(
        InParDataB[9]), .E(n2357), .CP(ClockB), .CDN(n2200), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][7]  ( .D(
        InParDataB[7]), .E(n2357), .CP(ClockB), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][5]  ( .D(
        InParDataB[5]), .E(n2357), .CP(ClockB), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][3]  ( .D(
        InParDataB[3]), .E(n2357), .CP(ClockB), .CDN(n2210), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][1]  ( .D(
        InParDataB[1]), .E(n2357), .CP(ClockB), .CDN(n2197), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][0]  ( .D(
        InParDataB[0]), .E(n2357), .CP(ClockB), .CDN(n2215), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][2]  ( .D(
        InParDataB[2]), .E(n2357), .CP(ClockB), .CDN(n2260), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][4]  ( .D(
        InParDataB[4]), .E(n2357), .CP(ClockB), .CDN(n2207), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][6]  ( .D(
        InParDataB[6]), .E(n2357), .CP(ClockB), .CDN(n2203), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][8]  ( .D(
        InParDataB[8]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2261), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][10]  ( .D(
        InParDataB[10]), .E(n2357), .CP(ClockB), .CDN(n2263), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][12]  ( .D(
        InParDataB[12]), .E(n2357), .CP(ClockB), .CDN(n2254), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][14]  ( .D(
        InParDataB[14]), .E(n2357), .CP(ClockB), .CDN(n2186), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][16]  ( .D(
        InParDataB[16]), .E(n2357), .CP(ClockB), .CDN(n2188), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][18]  ( .D(
        InParDataB[18]), .E(n2357), .CP(ClockB), .CDN(n2193), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][20]  ( .D(
        InParDataB[20]), .E(n2357), .CP(ClockB), .CDN(n2245), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][22]  ( .D(
        InParDataB[22]), .E(n2357), .CP(ClockB), .CDN(n2201), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][24]  ( .D(
        InParDataB[24]), .E(n2357), .CP(ClockB), .CDN(n2194), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][26]  ( .D(
        InParDataB[26]), .E(n2357), .CP(ClockB), .CDN(n2202), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][28]  ( .D(
        InParDataB[28]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2189), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage_reg[0][30]  ( .D(
        InParDataB[30]), .E(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .CP(
        ClockB), .CDN(n2190), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ), .CP(ClockA), .CDN(
        n1218), .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .CP(ClockA), .CDN(
        n1218), .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ) );
  DFCND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n1218), .Q(n2984), .QN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ) );
  DFCND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n1212), .Q(n2987), .QN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ) );
  DFCND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n1217), .Q(n2968), .QN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N7 ) );
  DFCND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[0]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n1121), .Q(n2974), .QN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N7 ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2233), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N1 ), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2227), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr [0]) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N1 ), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr [0]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ), .CP(ClockB), .CDN(
        n1217), .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .CP(ClockB), .CDN(
        n1217), .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2217), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2234), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2183), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidr_reg  ( .D(n1139), .CPN(n2292), 
        .CDN(n2190), .Q(n2954) );
  EDFCNQD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[1]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N39 ), .E(\SerDes_U1/SerLineValid ), .CP(
        n2296), .CDN(n2193), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[1]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N39 ), .E(\SerDes_U2/SerLineValid ), .CP(
        n2284), .CDN(n2191), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ) );
  DFCND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n1218), .Q(n2985), .QN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ) );
  DFCND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n1212), .Q(n2988), .QN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ) );
  DFCND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n1217), .Q(n2969), .QN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N19 ) );
  DFCND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/CounterClockN_reg[1]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n1121), .Q(n2975), .QN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N19 ) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteCmdr_reg  ( .D(n1226), 
        .CPN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), 
        .Q(n2986), .QN(n1311) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2234), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2218), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[2]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N40 ), .E(\SerDes_U1/SerLineValid ), .CP(
        n2292), .CDN(n2244), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[3]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N41 ), .E(\SerDes_U1/SerLineValid ), .CP(
        n2294), .CDN(n2268), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[2]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N40 ), .E(\SerDes_U2/SerLineValid ), .CP(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[3]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N41 ), .E(\SerDes_U2/SerLineValid ), .CP(
        n2282), .CDN(n2270), .Q(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutReg_reg  ( .D(
        n1213), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), 
        .CDN(n2226), .Q(\SerDes_U1/Tx_SerClk ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/ClockOutReg_reg  ( .D(
        n1122), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), 
        .CDN(n2228), .Q(\SerDes_U2/Tx_SerClk ) );
  DFCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), .Q(
        n2970), .QN(n1300) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[0]  ( .D(n1145), 
        .CPN(n2293), .CDN(n2189), .Q(n2957) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[0]  ( .D(n1054), 
        .CPN(\SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2205), .Q(n2948)
         );
  DFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[1]  ( .D(
        n1141), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2221), .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] )
         );
  DFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[1]  ( .D(
        n1050), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2231), .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] )
         );
  DFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[1]  ( .D(
        n1214), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2263), .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] )
         );
  DFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[1]  ( .D(
        n1123), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2244), .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] )
         );
  DFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[4]  ( .D(
        n1211), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2270), .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] )
         );
  DFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[4]  ( .D(
        n1120), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2270), .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] )
         );
  DFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[4]  ( .D(
        n1216), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2193), .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] )
         );
  DFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[4]  ( .D(
        n1125), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2213), .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] )
         );
  EDFCNQD1 \SerDes_U1/Des_U1/DesDec_Rx1/Count32_reg[0]  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N38 ), .E(\SerDes_U1/SerLineValid ), .CP(
        n2291), .CDN(n2255), .Q(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/DesDec_Rx1/Count32_reg[0]  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N38 ), .E(\SerDes_U2/SerLineValid ), .CP(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2226), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2218), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2249), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2263), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[5]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[0]  ( .D(n1177), .CPN(n2291), .CDN(n2186), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [0]), .QN(n908) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[1]  ( .D(n1176), .CPN(n2298), .CDN(n2186), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [1]), .QN(n907) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[2]  ( .D(n1175), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2186), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [2]), .QN(n906) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[3]  ( .D(n1174), .CPN(n2295), .CDN(n2186), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [3]), .QN(n905) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[4]  ( .D(n1173), .CPN(n2298), .CDN(n2186), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [4]), .QN(n904) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[5]  ( .D(n1172), .CPN(n2297), .CDN(n2186), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [5]), .QN(n903) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[6]  ( .D(n1171), .CPN(n2296), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [6]), .QN(n902) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[7]  ( .D(n1170), .CPN(n2297), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [7]), .QN(n901) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[8]  ( .D(n1169), .CPN(n2295), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [8]), .QN(n900) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[9]  ( .D(n1168), .CPN(n2296), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [9]), .QN(n899) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[10]  ( .D(n1167), .CPN(
        n2297), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [10]), .QN(n898) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[11]  ( .D(n1166), .CPN(
        n2295), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [11]), .QN(n897) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[12]  ( .D(n1165), .CPN(
        n2297), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [12]), .QN(n896) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[13]  ( .D(n1164), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2187), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [13]), .QN(n895) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[14]  ( .D(n1163), .CPN(
        n2296), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [14]), .QN(n894) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[15]  ( .D(n1162), .CPN(
        n2296), .CDN(n2187), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [15]), .QN(n893) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[16]  ( .D(n1161), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [16]), .QN(n892) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[17]  ( .D(n1160), .CPN(
        n2297), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [17]), .QN(n891) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[18]  ( .D(n1159), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [18]), .QN(n890) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[19]  ( .D(n1158), .CPN(
        n2295), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [19]), .QN(n889) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[20]  ( .D(n1157), .CPN(
        n2293), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [20]), .QN(n888) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[21]  ( .D(n1156), .CPN(
        n2297), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [21]), .QN(n887) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[22]  ( .D(n1155), .CPN(
        n2290), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [22]), .QN(n886) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[23]  ( .D(n1154), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [23]), .QN(n885) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[24]  ( .D(n1153), .CPN(
        n2298), .CDN(n2188), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [24]), .QN(n884) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[25]  ( .D(n1152), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2188), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [25]), .QN(n883) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[26]  ( .D(n1151), .CPN(
        \SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2189), .Q(
        \SerDes_U1/Des_U1/DecodeToFIFO [26]), .QN(n882) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[27]  ( .D(n1150), .CPN(
        n2297), .CDN(n2189), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [27]), .QN(n881) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[28]  ( .D(n1149), .CPN(
        n2291), .CDN(n2189), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [28]), .QN(n880) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[29]  ( .D(n1148), .CPN(
        n2295), .CDN(n2189), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [29]), .QN(n879) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[30]  ( .D(n1147), .CPN(
        n2294), .CDN(n2189), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [30]), .QN(n878) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParOutr_reg[31]  ( .D(n1146), .CPN(
        n2298), .CDN(n2189), .Q(\SerDes_U1/Des_U1/DecodeToFIFO [31]), .QN(n877) );
  DFSNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[0]  ( .D(
        n1140), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2264), .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] )
         );
  DFSNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[0]  ( .D(
        n1049), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .SDN(
        n2252), .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] )
         );
  DFSNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[0]  ( .D(
        n1215), .CP(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2260), .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] )
         );
  DFSNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[0]  ( .D(
        n1124), .CP(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .SDN(
        n2259), .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] )
         );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/ParValidTimer_reg[1]  ( .D(n1144), 
        .CPN(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2189), .Q(n2956)
         );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidTimer_reg[1]  ( .D(n1053), 
        .CPN(n2272), .CDN(n2205), .Q(n2947) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ), .CDN(n2222), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParValidr_reg  ( .D(n1048), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2205), .Q(n2945) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteCmdr_reg  ( .D(n1043), 
        .CPN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2203), 
        .Q(n2977) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2246), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2234), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2233), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2217), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2218), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2216), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/UnLoad_reg  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N79 ), .CPN(n2298), .CDN(n2186), .QN(
        n1307) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/UnLoad_reg  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N79 ), .CPN(n2286), .CDN(n2190), .QN(
        n1308) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2234), 
        .Q(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2229), 
        .Q(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ), .CDN(n2227), 
        .Q(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), .CDN(n2217), 
        .Q(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ) );
  DFCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), .Q(
        n2989), .QN(n1315) );
  DFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2218), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2266), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ), .CP(
        \SerDes_U1/Des_U1/SerialClk ), .CDN(n2233), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/MCntr1/N5 ), .CP(
        \SerDes_U2/Des_U1/SerialClk ), .CDN(n2226), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/CtrCarry ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2225), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/MCntr1/N5 ), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2228), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/CtrCarry ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2186), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[5]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N13 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[5]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N13 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ) );
  DFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2239), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]) );
  DFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [1]), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2221), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteCmdr_reg  ( .D(n1242), 
        .CPN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), 
        .Q(n2973) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteCmdr_reg  ( .D(n1135), 
        .CPN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2194), 
        .Q(n2990) );
  DFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [0]), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2229), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2204), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2259), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2255), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[2]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2236), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ) );
  DFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutReg_reg  ( .D(
        n1210), .CP(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), 
        .CDN(n2233), .Q(\SerDes_U1/Des_U1/SerialClk ) );
  DFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/ClockOutReg_reg  ( .D(
        n1119), .CP(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ), 
        .CDN(n2226), .Q(\SerDes_U2/Des_U1/SerialClk ) );
  DFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2222), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ) );
  DFNCND1 \SerDes_U1/Des_U1/DesDec_Rx1/doParSync_reg  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N47 ), .CPN(n2298), .CDN(n2186), .Q(n2996) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/doParSync_reg  ( .D(
        \SerDes_U2/Des_U1/DesDec_Rx1/N47 ), .CPN(n2285), .CDN(n2190), .Q(n2983) );
  DFCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [2]), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2202), .Q(
        n2972), .QN(n1310) );
  EDFCNQD1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ), .E(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ) );
  EDFCNQD1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ), .E(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/SampleWire ), .CDN(n2258), .Q(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ), .E(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2263), .Q(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor_reg[3]  ( 
        .D(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ), .E(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CP(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/SampleWire ), .CDN(n2237), .Q(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2185), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]) );
  DFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [1]), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2232), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ) );
  DFCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/NextState [0]), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), .Q(
        n2971), .QN(n1301) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2184), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2244), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[0]  ( .D(n1086), .CPN(n2271), .CDN(n2190), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [0]), .QN(n760) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[1]  ( .D(n1085), .CPN(n2273), .CDN(n2190), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [1]), .QN(n759) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[2]  ( .D(n1084), .CPN(n2282), .CDN(n2213), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [2]), .QN(n758) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[3]  ( .D(n1083), .CPN(n2283), .CDN(n2215), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [3]), .QN(n757) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[4]  ( .D(n1082), .CPN(n2284), .CDN(n2213), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [4]), .QN(n756) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[5]  ( .D(n1081), .CPN(n2285), .CDN(n2215), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [5]), .QN(n755) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[6]  ( .D(n1080), .CPN(n2285), .CDN(n2214), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [6]), .QN(n754) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[7]  ( .D(n1079), .CPN(n2286), .CDN(n2208), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [7]), .QN(n753) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[8]  ( .D(n1078), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2208), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [8]), .QN(n752) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[9]  ( .D(n1077), .CPN(n2284), .CDN(n2208), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [9]), .QN(n751) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[10]  ( .D(n1076), .CPN(
        n2286), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [10]), .QN(n750) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[11]  ( .D(n1075), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2207), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [11]), .QN(n749) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[12]  ( .D(n1074), .CPN(
        n2286), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [12]), .QN(n748) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[13]  ( .D(n1073), .CPN(
        n2285), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [13]), .QN(n747) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[14]  ( .D(n1072), .CPN(
        n2284), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [14]), .QN(n746) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[15]  ( .D(n1071), .CPN(
        n2283), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [15]), .QN(n745) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[16]  ( .D(n1070), .CPN(
        n2282), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [16]), .QN(n744) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[17]  ( .D(n1069), .CPN(
        n2283), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [17]), .QN(n743) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[18]  ( .D(n1068), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2207), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [18]), .QN(n742) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[19]  ( .D(n1067), .CPN(
        n2282), .CDN(n2207), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [19]), .QN(n741) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[20]  ( .D(n1066), .CPN(
        n2286), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [20]), .QN(n740) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[21]  ( .D(n1065), .CPN(
        n2284), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [21]), .QN(n739) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[22]  ( .D(n1064), .CPN(
        n2281), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [22]), .QN(n738) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[23]  ( .D(n1063), .CPN(
        n2274), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [23]), .QN(n737) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[24]  ( .D(n1062), .CPN(
        \SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .CDN(n2206), .Q(
        \SerDes_U2/Des_U1/DecodeToFIFO [24]), .QN(n736) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[25]  ( .D(n1061), .CPN(
        n2286), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [25]), .QN(n735) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[26]  ( .D(n1060), .CPN(
        n2283), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [26]), .QN(n734) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[27]  ( .D(n1059), .CPN(
        n2284), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [27]), .QN(n733) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[28]  ( .D(n1058), .CPN(
        n2285), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [28]), .QN(n732) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[29]  ( .D(n1057), .CPN(
        n2281), .CDN(n2206), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [29]), .QN(n731) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[30]  ( .D(n1056), .CPN(
        n2282), .CDN(n2205), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [30]), .QN(n730) );
  DFNCND1 \SerDes_U2/Des_U1/DesDec_Rx1/ParOutr_reg[31]  ( .D(n1055), .CPN(
        n2283), .CDN(n2205), .Q(\SerDes_U2/Des_U1/DecodeToFIFO [31]), .QN(n729) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/SerValidr_reg  ( .D(n1036), .CP(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2218), .Q(
        \SerDes_U2/SerLineValid ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/SerValidr_reg  ( .D(n1035), .CP(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .CDN(n2222), .Q(
        \SerDes_U1/SerLineValid ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2187), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[4]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N12 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[4]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N12 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2184), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2240), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[3]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N11 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N11 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/WriteAr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2245), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N10 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N10 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2231), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2182), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2269), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[3]  ( .D(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ), .E(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2267), .Q(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2186), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2185), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ), .E(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2198), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2250), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2264), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2262), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ), .CP(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2243), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2183), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2209), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadAr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ), .CP(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2210), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ) );
  DFNCND1 \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadCmdr_reg  ( .D(n1244), .CPN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2201), .Q(
        n1298), .QN(n1314) );
  DFNCND1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/ReadCmdr_reg  ( .D(n1137), .CPN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2190), .Q(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .QN(n869) );
  DFNCND1 \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/ReadCmdr_reg  ( .D(n1228), .CPN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClock ), .CDN(n2204), .Q(
        \SerDes_U1/Ser_U1/FIFO_Tx1/SM_MemReadCmd ), .QN(n1015) );
  DFNCND1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/ReadCmdr_reg  ( .D(n1046), .CPN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClock ), .CDN(n2205), .Q(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .QN(n721) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr_reg  ( .D(n2352), .CP(
        ClockA), .CDN(n2217), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr_reg  ( .D(n2350), .CP(
        ClockB), .CDN(n2230), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[1]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N9 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[1]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N9 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ) );
  DFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N_reg[0]  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N8 ), .CP(\SerDes_U1/Tx_SerClk ), .CDN(
        n2226), .Q(\SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ) );
  DFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N_reg[0]  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N8 ), .CP(\SerDes_U2/Tx_SerClk ), .CDN(
        n2228), .Q(\SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ) );
  EDFCNQD1 \SerDes_U1/Ser_U1/SerEnc_Tx1/SerOutr_reg  ( .D(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 ), .E(n2997), .CP(
        \SerDes_U1/Tx_SerClk ), .CDN(n2254), .Q(
        \SerDes_U1/Des_U1/SerRxToDecode ) );
  EDFCNQD1 \SerDes_U2/Ser_U1/SerEnc_Tx1/SerOutr_reg  ( .D(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ), .E(n2997), .CP(
        \SerDes_U2/Tx_SerClk ), .CDN(n2237), .Q(
        \SerDes_U2/Des_U1/SerRxToDecode ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2261), 
        .Q(\SerDes_U2/Des_U1/N34 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2207), 
        .Q(\SerDes_U2/Des_U1/N33 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ), .E(n2347), .CP(ClockA), 
        .CDN(n2206), .Q(\SerDes_U2/Des_U1/N32 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2252), 
        .Q(\SerDes_U2/Des_U1/N31 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2247), 
        .Q(\SerDes_U2/Des_U1/N30 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2200), 
        .Q(\SerDes_U2/Des_U1/N29 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2248), 
        .Q(\SerDes_U2/Des_U1/N28 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2218), 
        .Q(\SerDes_U2/Des_U1/N27 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2202), 
        .Q(\SerDes_U2/Des_U1/N26 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2251), 
        .Q(\SerDes_U2/Des_U1/N25 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2254), 
        .Q(\SerDes_U2/Des_U1/N24 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2253), 
        .Q(\SerDes_U2/Des_U1/N23 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ), .E(n2347), .CP(ClockA), 
        .CDN(n2201), .Q(\SerDes_U2/Des_U1/N22 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2242), 
        .Q(\SerDes_U2/Des_U1/N21 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ), .E(n2347), .CP(ClockA), 
        .CDN(n2256), .Q(\SerDes_U2/Des_U1/N20 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2241), 
        .Q(\SerDes_U2/Des_U1/N19 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ), .E(n2347), .CP(ClockA), 
        .CDN(n2231), .Q(\SerDes_U2/Des_U1/N18 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2266), 
        .Q(\SerDes_U2/Des_U1/N17 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ), .E(n2347), .CP(ClockA), 
        .CDN(n2221), .Q(\SerDes_U2/Des_U1/N16 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2211), 
        .Q(\SerDes_U2/Des_U1/N15 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ), .E(n2347), .CP(ClockA), 
        .CDN(n2219), .Q(\SerDes_U2/Des_U1/N14 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ), .E(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockA), .CDN(n2220), 
        .Q(\SerDes_U2/Des_U1/N13 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ), .E(n2347), .CP(ClockA), 
        .CDN(n2222), .Q(\SerDes_U2/Des_U1/N12 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ), .E(n2347), .CP(ClockA), 
        .CDN(n2223), .Q(\SerDes_U2/Des_U1/N11 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ), .E(n2347), .CP(ClockA), 
        .CDN(n2224), .Q(\SerDes_U2/Des_U1/N10 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ), .E(n2347), .CP(ClockA), 
        .CDN(n2225), .Q(\SerDes_U2/Des_U1/N9 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ), .E(n2347), .CP(ClockA), 
        .CDN(n2230), .Q(\SerDes_U2/Des_U1/N8 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ), .E(n2347), .CP(ClockA), 
        .CDN(n2229), .Q(\SerDes_U2/Des_U1/N7 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ), .E(n2347), .CP(ClockA), 
        .CDN(n2226), .Q(\SerDes_U2/Des_U1/N6 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ), .E(n2347), .CP(ClockA), 
        .CDN(n2214), .Q(\SerDes_U2/Des_U1/N5 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ), .E(n2347), .CP(ClockA), 
        .CDN(n2212), .Q(\SerDes_U2/Des_U1/N4 ) );
  EDFCNQD1 \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ), .E(n2347), .CP(ClockA), 
        .CDN(n2206), .Q(\SerDes_U2/Des_U1/N3 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[31]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2259), 
        .Q(\SerDes_U1/Des_U1/N34 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[30]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2246), 
        .Q(\SerDes_U1/Des_U1/N33 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[29]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ), .E(n2426), .CP(ClockB), 
        .CDN(n2250), .Q(\SerDes_U1/Des_U1/N32 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[28]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ), .E(n2426), .CP(ClockB), 
        .CDN(n2244), .Q(\SerDes_U1/Des_U1/N31 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[27]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ), .E(n2426), .CP(ClockB), 
        .CDN(n2270), .Q(\SerDes_U1/Des_U1/N30 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[26]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ), .E(n2426), .CP(ClockB), 
        .CDN(n2204), .Q(\SerDes_U1/Des_U1/N29 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[25]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ), .E(n2426), .CP(ClockB), 
        .CDN(n2187), .Q(\SerDes_U1/Des_U1/N28 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[24]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ), .E(n2426), .CP(ClockB), 
        .CDN(n2242), .Q(\SerDes_U1/Des_U1/N27 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[23]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ), .E(n2426), .CP(ClockB), 
        .CDN(n2248), .Q(\SerDes_U1/Des_U1/N26 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[22]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ), .E(n2426), .CP(ClockB), 
        .CDN(n2241), .Q(\SerDes_U1/Des_U1/N25 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[21]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ), .E(n2426), .CP(ClockB), 
        .CDN(n2220), .Q(\SerDes_U1/Des_U1/N24 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[20]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ), .E(n2426), .CP(ClockB), 
        .CDN(n2238), .Q(\SerDes_U1/Des_U1/N23 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[19]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ), .E(n2426), .CP(ClockB), 
        .CDN(n2227), .Q(\SerDes_U1/Des_U1/N22 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[18]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2218), 
        .Q(\SerDes_U1/Des_U1/N21 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[17]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2255), 
        .Q(\SerDes_U1/Des_U1/N20 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[16]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2183), 
        .Q(\SerDes_U1/Des_U1/N19 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[15]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2264), 
        .Q(\SerDes_U1/Des_U1/N18 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[14]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2253), 
        .Q(\SerDes_U1/Des_U1/N17 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[13]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2231), 
        .Q(\SerDes_U1/Des_U1/N16 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[12]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2262), 
        .Q(\SerDes_U1/Des_U1/N15 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[11]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2196), 
        .Q(\SerDes_U1/Des_U1/N14 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[10]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2238), 
        .Q(\SerDes_U1/Des_U1/N13 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[9]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ), .E(n2426), .CP(ClockB), 
        .CDN(n2258), .Q(\SerDes_U1/Des_U1/N12 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[8]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2223), 
        .Q(\SerDes_U1/Des_U1/N11 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[7]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ), .E(n2426), .CP(ClockB), 
        .CDN(n2182), .Q(\SerDes_U1/Des_U1/N10 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[6]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2234), 
        .Q(\SerDes_U1/Des_U1/N9 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[5]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ), .E(n2426), .CP(ClockB), 
        .CDN(n2263), .Q(\SerDes_U1/Des_U1/N8 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[4]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2254), 
        .Q(\SerDes_U1/Des_U1/N7 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[3]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ), .E(n2426), .CP(ClockB), 
        .CDN(n2253), .Q(\SerDes_U1/Des_U1/N6 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[2]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2252), 
        .Q(\SerDes_U1/Des_U1/N5 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[1]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ), .E(n2426), .CP(ClockB), 
        .CDN(n2264), .Q(\SerDes_U1/Des_U1/N4 ) );
  EDFCNQD1 \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/DataOr_reg[0]  ( .D(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ), .E(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_MemReadCmd ), .CP(ClockB), .CDN(n2249), 
        .Q(\SerDes_U1/Des_U1/N3 ) );
  DFSND1 \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .CP(ClockA), .SDN(
        n2237), .QN(n1218) );
  DFSND1 \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .CP(ClockB), .SDN(
        n2200), .QN(n1217) );
  DFSND1 \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .CP(
        \SerDes_U1/Rx_ParClk ), .SDN(n2239), .QN(n1212) );
  DFSND1 \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .CP(
        \SerDes_U2/Rx_ParClk ), .SDN(n2238), .QN(n1121) );
  EDFCNQD4 \SerDes_U1/Des_U1/DesDec_Rx1/ParClkr_reg  ( .D(
        \SerDes_U1/Des_U1/DesDec_Rx1/N37 ), .E(
        \SerDes_U1/Des_U1/DesDec_Rx1/N43 ), .CP(n2298), .CDN(n2182), .Q(
        \SerDes_U1/Rx_ParClk ) );
  NR2D1 U1027 ( .A1(n2582), .A2(n2892), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ) );
  NR2D1 U1028 ( .A1(n2809), .A2(n2818), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ) );
  NR2D1 U1029 ( .A1(n2814), .A2(n2817), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ) );
  NR2D1 U1030 ( .A1(n2809), .A2(n2817), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ) );
  NR2D1 U1031 ( .A1(n2815), .A2(n2809), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ) );
  NR2D1 U1032 ( .A1(n2815), .A2(n2816), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ) );
  NR2D1 U1033 ( .A1(n2815), .A2(n2808), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ) );
  NR2D1 U1034 ( .A1(n2808), .A2(n2818), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ) );
  NR2D1 U1035 ( .A1(n2808), .A2(n2819), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ) );
  NR2D1 U1036 ( .A1(n2925), .A2(n2928), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ) );
  INR2D1 U1037 ( .A1(n2990), .B1(n2916), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ) );
  NR2D1 U1038 ( .A1(n2925), .A2(n2926), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ) );
  NR2D1 U1039 ( .A1(n2917), .A2(n2929), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ) );
  NR2D1 U1040 ( .A1(n2917), .A2(n2930), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ) );
  NR2D1 U1041 ( .A1(n2567), .A2(n2892), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ) );
  NR2D1 U1042 ( .A1(n2567), .A2(n2891), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ) );
  NR2D1 U1043 ( .A1(n2582), .A2(n2891), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ) );
  NR2D2 U1044 ( .A1(n1299), .A2(Reset), .ZN(n1296) );
  INVD1 U1045 ( .I(Reset), .ZN(n1247) );
  INVD0 U1046 ( .I(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), .ZN(n2300) );
  INR2D1 U1047 ( .A1(n2931), .B1(n2932), .ZN(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ) );
  INVD0 U1048 ( .I(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), .ZN(n2288) );
  INR2D1 U1049 ( .A1(n2843), .B1(n2844), .ZN(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ) );
  NR2D1 U1050 ( .A1(n2816), .A2(n2819), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ) );
  NR2D1 U1051 ( .A1(n2814), .A2(n2819), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ) );
  NR2D1 U1052 ( .A1(n2816), .A2(n2818), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ) );
  INR2D1 U1053 ( .A1(n2973), .B1(n2807), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ) );
  NR2D1 U1054 ( .A1(n2816), .A2(n2817), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ) );
  NR2D1 U1055 ( .A1(n2814), .A2(n2815), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ) );
  NR2D1 U1056 ( .A1(n2809), .A2(n2819), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ) );
  NR2D1 U1057 ( .A1(n2808), .A2(n2817), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ) );
  NR2D1 U1058 ( .A1(n2927), .A2(n2930), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ) );
  NR2D1 U1059 ( .A1(n2925), .A2(n2930), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ) );
  NR2D1 U1060 ( .A1(n2927), .A2(n2929), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ) );
  NR2D1 U1061 ( .A1(n2927), .A2(n2928), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ) );
  NR2D1 U1062 ( .A1(n2926), .A2(n2927), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ) );
  NR2D1 U1063 ( .A1(n2918), .A2(n2930), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ) );
  NR2D1 U1064 ( .A1(n2918), .A2(n2929), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ) );
  NR2D1 U1065 ( .A1(n2917), .A2(n2928), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ) );
  NR2D1 U1066 ( .A1(n2918), .A2(n2928), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ) );
  NR2D1 U1067 ( .A1(n2926), .A2(n2917), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ) );
  NR2D1 U1068 ( .A1(n2926), .A2(n2918), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ) );
  NR2D1 U1069 ( .A1(n2763), .A2(n2842), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ) );
  NR2D1 U1070 ( .A1(n2762), .A2(n2839), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ) );
  NR2D1 U1071 ( .A1(n2762), .A2(n2842), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ) );
  NR2D1 U1072 ( .A1(n2763), .A2(n2839), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ) );
  OR2D1 U1073 ( .A1(n1302), .A2(Reset), .Z(n1297) );
  MUX2ND0 U1074 ( .I0(n1542), .I1(n1543), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1303) );
  MUX2ND0 U1075 ( .I0(n1546), .I1(n1547), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1304) );
  MUX2ND0 U1076 ( .I0(n1534), .I1(n1535), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1305) );
  MUX2ND0 U1077 ( .I0(n1538), .I1(n1539), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1306) );
  MUX2ND0 U1078 ( .I0(n1544), .I1(n1545), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1397) );
  MUX2ND0 U1079 ( .I0(n1548), .I1(n1549), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1398) );
  MUX2ND0 U1080 ( .I0(n1536), .I1(n1537), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1399) );
  MUX2ND0 U1081 ( .I0(n1540), .I1(n1541), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(n1400) );
  CKBD0 U1082 ( .CLK(n2144), .C(n1402) );
  CKNXD16 U1083 ( .I(n1402), .ZN(OutParDataB[29]) );
  CKBD0 U1084 ( .CLK(n2143), .C(n1404) );
  CKNXD16 U1085 ( .I(n1404), .ZN(OutParDataB[28]) );
  CKBD0 U1086 ( .CLK(n2145), .C(n1406) );
  CKNXD16 U1087 ( .I(n1406), .ZN(OutParDataB[30]) );
  CKBD0 U1088 ( .CLK(n2142), .C(n1408) );
  CKNXD16 U1089 ( .I(n1408), .ZN(OutParDataB[27]) );
  CKBD0 U1090 ( .CLK(n2140), .C(n1410) );
  CKNXD16 U1091 ( .I(n1410), .ZN(OutParDataB[25]) );
  CKBD0 U1092 ( .CLK(n2141), .C(n1412) );
  CKNXD16 U1093 ( .I(n1412), .ZN(OutParDataB[26]) );
  CKBD0 U1094 ( .CLK(n2139), .C(n1414) );
  CKNXD16 U1095 ( .I(n1414), .ZN(OutParDataB[24]) );
  CKBD0 U1096 ( .CLK(n2146), .C(n1416) );
  CKNXD16 U1097 ( .I(n1416), .ZN(OutParDataB[31]) );
  CKBD0 U1098 ( .CLK(n2118), .C(n1418) );
  CKNXD16 U1099 ( .I(n1418), .ZN(OutParDataB[3]) );
  CKBD0 U1100 ( .CLK(n2116), .C(n1420) );
  CKNXD16 U1101 ( .I(n1420), .ZN(OutParDataB[1]) );
  CKBD0 U1102 ( .CLK(n2117), .C(n1422) );
  CKNXD16 U1103 ( .I(n1422), .ZN(OutParDataB[2]) );
  CKBD0 U1104 ( .CLK(n2138), .C(n1424) );
  CKNXD16 U1105 ( .I(n1424), .ZN(OutParDataB[23]) );
  CKBD0 U1106 ( .CLK(n2136), .C(n1426) );
  CKNXD16 U1107 ( .I(n1426), .ZN(OutParDataB[21]) );
  CKBD0 U1108 ( .CLK(n2137), .C(n1428) );
  CKNXD16 U1109 ( .I(n1428), .ZN(OutParDataB[22]) );
  CKBD0 U1110 ( .CLK(n2135), .C(n1430) );
  CKNXD16 U1111 ( .I(n1430), .ZN(OutParDataB[20]) );
  CKBD0 U1112 ( .CLK(n2119), .C(n1432) );
  CKNXD16 U1113 ( .I(n1432), .ZN(OutParDataB[4]) );
  CKBD0 U1114 ( .CLK(n2120), .C(n1434) );
  CKNXD16 U1115 ( .I(n1434), .ZN(OutParDataB[5]) );
  CKBD0 U1116 ( .CLK(n2115), .C(n1436) );
  CKNXD16 U1117 ( .I(n1436), .ZN(OutParDataB[0]) );
  CKBD0 U1118 ( .CLK(n2122), .C(n1438) );
  CKNXD16 U1119 ( .I(n1438), .ZN(OutParDataB[7]) );
  CKBD0 U1120 ( .CLK(n2134), .C(n1440) );
  CKNXD16 U1121 ( .I(n1440), .ZN(OutParDataB[19]) );
  CKBD0 U1122 ( .CLK(n2132), .C(n1442) );
  CKNXD16 U1123 ( .I(n1442), .ZN(OutParDataB[17]) );
  CKBD0 U1124 ( .CLK(n2133), .C(n1444) );
  CKNXD16 U1125 ( .I(n1444), .ZN(OutParDataB[18]) );
  CKBD0 U1126 ( .CLK(n2131), .C(n1446) );
  CKNXD16 U1127 ( .I(n1446), .ZN(OutParDataB[16]) );
  CKBD0 U1128 ( .CLK(n2121), .C(n1448) );
  CKNXD16 U1129 ( .I(n1448), .ZN(OutParDataB[6]) );
  CKBD0 U1130 ( .CLK(n2125), .C(n1450) );
  CKNXD16 U1131 ( .I(n1450), .ZN(OutParDataB[10]) );
  CKBD0 U1132 ( .CLK(n2123), .C(n1452) );
  CKNXD16 U1133 ( .I(n1452), .ZN(OutParDataB[8]) );
  CKBD0 U1134 ( .CLK(n2124), .C(n1454) );
  CKNXD16 U1135 ( .I(n1454), .ZN(OutParDataB[9]) );
  CKBD0 U1136 ( .CLK(n2130), .C(n1456) );
  CKNXD16 U1137 ( .I(n1456), .ZN(OutParDataB[15]) );
  CKBD0 U1138 ( .CLK(n2128), .C(n1458) );
  CKNXD16 U1139 ( .I(n1458), .ZN(OutParDataB[13]) );
  CKBD0 U1140 ( .CLK(n2129), .C(n1460) );
  CKNXD16 U1141 ( .I(n1460), .ZN(OutParDataB[14]) );
  CKBD0 U1142 ( .CLK(n2127), .C(n1462) );
  CKNXD16 U1143 ( .I(n1462), .ZN(OutParDataB[12]) );
  CKBD0 U1144 ( .CLK(n2126), .C(n1464) );
  CKNXD16 U1145 ( .I(n1464), .ZN(OutParDataB[11]) );
  CKBD0 U1146 ( .CLK(n2164), .C(n1466) );
  CKNXD16 U1147 ( .I(n1466), .ZN(OutParDataA[17]) );
  CKBD0 U1148 ( .CLK(n2163), .C(n1468) );
  CKNXD16 U1149 ( .I(n1468), .ZN(OutParDataA[16]) );
  CKBD0 U1150 ( .CLK(n2165), .C(n1470) );
  CKNXD16 U1151 ( .I(n1470), .ZN(OutParDataA[18]) );
  CKBD0 U1152 ( .CLK(n2162), .C(n1472) );
  CKNXD16 U1153 ( .I(n1472), .ZN(OutParDataA[15]) );
  CKBD0 U1154 ( .CLK(n2160), .C(n1474) );
  CKNXD16 U1155 ( .I(n1474), .ZN(OutParDataA[13]) );
  CKBD0 U1156 ( .CLK(n2161), .C(n1476) );
  CKNXD16 U1157 ( .I(n1476), .ZN(OutParDataA[14]) );
  CKBD0 U1158 ( .CLK(n2159), .C(n1478) );
  CKNXD16 U1159 ( .I(n1478), .ZN(OutParDataA[12]) );
  CKBD0 U1160 ( .CLK(n2166), .C(n1480) );
  CKNXD16 U1161 ( .I(n1480), .ZN(OutParDataA[19]) );
  CKBD0 U1162 ( .CLK(n2168), .C(n1482) );
  CKNXD16 U1163 ( .I(n1482), .ZN(OutParDataA[21]) );
  CKBD0 U1164 ( .CLK(n2167), .C(n1484) );
  CKNXD16 U1165 ( .I(n1484), .ZN(OutParDataA[20]) );
  CKBD0 U1166 ( .CLK(n2169), .C(n1486) );
  CKNXD16 U1167 ( .I(n1486), .ZN(OutParDataA[22]) );
  CKBD0 U1168 ( .CLK(n2158), .C(n1488) );
  CKNXD16 U1169 ( .I(n1488), .ZN(OutParDataA[11]) );
  CKBD0 U1170 ( .CLK(n2156), .C(n1490) );
  CKNXD16 U1171 ( .I(n1490), .ZN(OutParDataA[9]) );
  CKBD0 U1172 ( .CLK(n2157), .C(n1492) );
  CKNXD16 U1173 ( .I(n1492), .ZN(OutParDataA[10]) );
  CKBD0 U1174 ( .CLK(n2155), .C(n1494) );
  CKNXD16 U1175 ( .I(n1494), .ZN(OutParDataA[8]) );
  CKBD0 U1176 ( .CLK(n2170), .C(n1496) );
  CKNXD16 U1177 ( .I(n1496), .ZN(OutParDataA[23]) );
  CKBD0 U1178 ( .CLK(n2172), .C(n1498) );
  CKNXD16 U1179 ( .I(n1498), .ZN(OutParDataA[25]) );
  CKBD0 U1180 ( .CLK(n2171), .C(n1500) );
  CKNXD16 U1181 ( .I(n1500), .ZN(OutParDataA[24]) );
  CKBD0 U1182 ( .CLK(n2173), .C(n1502) );
  CKNXD16 U1183 ( .I(n1502), .ZN(OutParDataA[26]) );
  CKBD0 U1184 ( .CLK(n2154), .C(n1504) );
  CKNXD16 U1185 ( .I(n1504), .ZN(OutParDataA[7]) );
  CKBD0 U1186 ( .CLK(n2152), .C(n1506) );
  CKNXD16 U1187 ( .I(n1506), .ZN(OutParDataA[5]) );
  CKBD0 U1188 ( .CLK(n2153), .C(n1508) );
  CKNXD16 U1189 ( .I(n1508), .ZN(OutParDataA[6]) );
  CKBD0 U1190 ( .CLK(n2151), .C(n1510) );
  CKNXD16 U1191 ( .I(n1510), .ZN(OutParDataA[4]) );
  CKBD0 U1192 ( .CLK(n2174), .C(n1512) );
  CKNXD16 U1193 ( .I(n1512), .ZN(OutParDataA[27]) );
  CKBD0 U1194 ( .CLK(n2176), .C(n1514) );
  CKNXD16 U1195 ( .I(n1514), .ZN(OutParDataA[29]) );
  CKBD0 U1196 ( .CLK(n2175), .C(n1516) );
  CKNXD16 U1197 ( .I(n1516), .ZN(OutParDataA[28]) );
  CKBD0 U1198 ( .CLK(n2177), .C(n1518) );
  CKNXD16 U1199 ( .I(n1518), .ZN(OutParDataA[30]) );
  CKBD0 U1200 ( .CLK(n2150), .C(n1520) );
  CKNXD16 U1201 ( .I(n1520), .ZN(OutParDataA[3]) );
  CKBD0 U1202 ( .CLK(n2148), .C(n1522) );
  CKNXD16 U1203 ( .I(n1522), .ZN(OutParDataA[1]) );
  CKBD0 U1204 ( .CLK(n2149), .C(n1524) );
  CKNXD16 U1205 ( .I(n1524), .ZN(OutParDataA[2]) );
  CKBD0 U1206 ( .CLK(n2147), .C(n1526) );
  CKNXD16 U1207 ( .I(n1526), .ZN(OutParDataA[0]) );
  CKBD0 U1208 ( .CLK(n2178), .C(n1528) );
  CKNXD16 U1209 ( .I(n1528), .ZN(OutParDataA[31]) );
  BUFFD1 U1210 ( .I(n2245), .Z(n2227) );
  BUFFD1 U1211 ( .I(n2245), .Z(n2228) );
  BUFFD1 U1212 ( .I(n2244), .Z(n2229) );
  BUFFD1 U1213 ( .I(n2245), .Z(n2226) );
  BUFFD1 U1214 ( .I(n2246), .Z(n2225) );
  BUFFD1 U1215 ( .I(n2246), .Z(n2224) );
  BUFFD1 U1216 ( .I(n2246), .Z(n2223) );
  BUFFD1 U1217 ( .I(n2247), .Z(n2222) );
  BUFFD1 U1218 ( .I(n2247), .Z(n2221) );
  BUFFD1 U1219 ( .I(n2247), .Z(n2220) );
  BUFFD1 U1220 ( .I(n2248), .Z(n2219) );
  BUFFD1 U1221 ( .I(n2243), .Z(n2234) );
  BUFFD1 U1222 ( .I(n2242), .Z(n2236) );
  BUFFD1 U1223 ( .I(n2242), .Z(n2235) );
  BUFFD1 U1224 ( .I(n2241), .Z(n2240) );
  BUFFD1 U1225 ( .I(n2241), .Z(n2239) );
  BUFFD1 U1226 ( .I(n2241), .Z(n2238) );
  BUFFD1 U1227 ( .I(n2242), .Z(n2237) );
  BUFFD1 U1228 ( .I(n2248), .Z(n2218) );
  BUFFD1 U1229 ( .I(n2260), .Z(n2184) );
  BUFFD1 U1230 ( .I(n2260), .Z(n2183) );
  BUFFD1 U1231 ( .I(n2253), .Z(n2203) );
  BUFFD1 U1232 ( .I(n2252), .Z(n2206) );
  BUFFD1 U1233 ( .I(n2252), .Z(n2207) );
  BUFFD1 U1234 ( .I(n2257), .Z(n2191) );
  BUFFD1 U1235 ( .I(n2256), .Z(n2196) );
  BUFFD1 U1236 ( .I(n2255), .Z(n2197) );
  BUFFD1 U1237 ( .I(n2257), .Z(n2192) );
  BUFFD1 U1238 ( .I(n2254), .Z(n2200) );
  BUFFD1 U1239 ( .I(n2255), .Z(n2199) );
  BUFFD1 U1240 ( .I(n2255), .Z(n2198) );
  BUFFD1 U1241 ( .I(n2256), .Z(n2195) );
  BUFFD1 U1242 ( .I(n2256), .Z(n2194) );
  BUFFD1 U1243 ( .I(n2257), .Z(n2193) );
  BUFFD1 U1244 ( .I(n2258), .Z(n2190) );
  BUFFD1 U1245 ( .I(n2258), .Z(n2189) );
  BUFFD1 U1246 ( .I(n2258), .Z(n2188) );
  BUFFD1 U1247 ( .I(n2259), .Z(n2187) );
  BUFFD1 U1248 ( .I(n2259), .Z(n2186) );
  BUFFD1 U1249 ( .I(n2259), .Z(n2185) );
  BUFFD1 U1250 ( .I(n2252), .Z(n2208) );
  BUFFD1 U1251 ( .I(n2251), .Z(n2209) );
  BUFFD1 U1252 ( .I(n2251), .Z(n2210) );
  BUFFD1 U1253 ( .I(n2251), .Z(n2211) );
  BUFFD1 U1254 ( .I(n2250), .Z(n2213) );
  BUFFD1 U1255 ( .I(n2250), .Z(n2214) );
  BUFFD1 U1256 ( .I(n2250), .Z(n2212) );
  BUFFD1 U1257 ( .I(n2253), .Z(n2205) );
  BUFFD1 U1258 ( .I(n2253), .Z(n2204) );
  BUFFD1 U1259 ( .I(n2254), .Z(n2202) );
  BUFFD1 U1260 ( .I(n2254), .Z(n2201) );
  BUFFD1 U1261 ( .I(n2243), .Z(n2233) );
  BUFFD1 U1262 ( .I(n2248), .Z(n2217) );
  BUFFD1 U1263 ( .I(n2243), .Z(n2232) );
  BUFFD1 U1264 ( .I(n2244), .Z(n2230) );
  BUFFD1 U1265 ( .I(n2249), .Z(n2216) );
  BUFFD1 U1266 ( .I(n2244), .Z(n2231) );
  BUFFD1 U1267 ( .I(n2249), .Z(n2215) );
  BUFFD1 U1268 ( .I(n2191), .Z(n2241) );
  BUFFD1 U1269 ( .I(n2262), .Z(n2255) );
  BUFFD1 U1270 ( .I(n2262), .Z(n2256) );
  BUFFD1 U1271 ( .I(n2262), .Z(n2257) );
  BUFFD1 U1272 ( .I(n2261), .Z(n2258) );
  BUFFD1 U1273 ( .I(n2261), .Z(n2259) );
  BUFFD1 U1274 ( .I(n2263), .Z(n2252) );
  BUFFD1 U1275 ( .I(n2264), .Z(n2251) );
  BUFFD1 U1276 ( .I(n2264), .Z(n2250) );
  BUFFD1 U1277 ( .I(n2264), .Z(n2249) );
  BUFFD1 U1278 ( .I(n2266), .Z(n2243) );
  BUFFD1 U1279 ( .I(n2266), .Z(n2245) );
  BUFFD1 U1280 ( .I(n2192), .Z(n2242) );
  BUFFD1 U1281 ( .I(n2265), .Z(n2246) );
  BUFFD1 U1282 ( .I(n2263), .Z(n2253) );
  BUFFD1 U1283 ( .I(n2265), .Z(n2247) );
  BUFFD1 U1284 ( .I(n2263), .Z(n2254) );
  BUFFD1 U1285 ( .I(n2266), .Z(n2244) );
  BUFFD1 U1286 ( .I(n2265), .Z(n2248) );
  BUFFD1 U1287 ( .I(n2261), .Z(n2260) );
  BUFFD1 U1288 ( .I(n2269), .Z(n2262) );
  BUFFD1 U1289 ( .I(n2269), .Z(n2261) );
  BUFFD1 U1290 ( .I(n2268), .Z(n2264) );
  BUFFD1 U1291 ( .I(n2268), .Z(n2263) );
  BUFFD1 U1292 ( .I(n2267), .Z(n2266) );
  BUFFD1 U1293 ( .I(n2267), .Z(n2265) );
  BUFFD1 U1294 ( .I(n2270), .Z(n2269) );
  BUFFD1 U1295 ( .I(n2270), .Z(n2268) );
  BUFFD1 U1296 ( .I(n2270), .Z(n2267) );
  BUFFD1 U1297 ( .I(n2114), .Z(n2113) );
  BUFFD1 U1298 ( .I(n2114), .Z(n2112) );
  BUFFD1 U1299 ( .I(n2011), .Z(n2010) );
  BUFFD1 U1300 ( .I(n2011), .Z(n2009) );
  BUFFD1 U1301 ( .I(n1755), .Z(n1757) );
  BUFFD1 U1302 ( .I(n1755), .Z(n1758) );
  BUFFD1 U1303 ( .I(n1755), .Z(n1759) );
  BUFFD1 U1304 ( .I(n1896), .Z(n1898) );
  BUFFD1 U1305 ( .I(n1758), .Z(n1760) );
  BUFFD1 U1306 ( .I(n1895), .Z(n1899) );
  BUFFD1 U1307 ( .I(n1895), .Z(n1900) );
  BUFFD1 U1308 ( .I(n2114), .Z(n2111) );
  BUFFD1 U1309 ( .I(n2011), .Z(n2008) );
  BUFFD1 U1310 ( .I(n2110), .Z(n2109) );
  BUFFD1 U1311 ( .I(n2007), .Z(n2006) );
  BUFFD1 U1312 ( .I(n1899), .Z(n1897) );
  BUFFD1 U1313 ( .I(n1891), .Z(n1892) );
  BUFFD1 U1314 ( .I(n1751), .Z(n1753) );
  BUFFD1 U1315 ( .I(n1751), .Z(n1754) );
  BUFFD1 U1316 ( .I(n1892), .Z(n1893) );
  BUFFD1 U1317 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1894) );
  BUFFD1 U1318 ( .I(n1753), .Z(n1752) );
  BUFFD1 U1319 ( .I(n2285), .Z(n2271) );
  BUFFD1 U1320 ( .I(n2285), .Z(n2272) );
  BUFFD1 U1321 ( .I(n2285), .Z(n2273) );
  BUFFD1 U1322 ( .I(n2284), .Z(n2274) );
  BUFFD1 U1323 ( .I(n2284), .Z(n2275) );
  BUFFD1 U1324 ( .I(n2283), .Z(n2276) );
  BUFFD1 U1325 ( .I(n2283), .Z(n2277) );
  BUFFD1 U1326 ( .I(n2282), .Z(n2278) );
  BUFFD1 U1327 ( .I(n2282), .Z(n2279) );
  BUFFD1 U1328 ( .I(n2283), .Z(n2280) );
  BUFFD1 U1329 ( .I(n2290), .Z(n2289) );
  BUFFD1 U1330 ( .I(n2294), .Z(n2290) );
  BUFFD1 U1331 ( .I(n2297), .Z(n2291) );
  BUFFD1 U1332 ( .I(n2297), .Z(n2292) );
  BUFFD1 U1333 ( .I(n2296), .Z(n2293) );
  BUFFD1 U1334 ( .I(n2296), .Z(n2294) );
  BUFFD1 U1335 ( .I(n2182), .Z(n2270) );
  INVD1 U1336 ( .I(n2303), .ZN(n2108) );
  INVD1 U1337 ( .I(n2355), .ZN(n1890) );
  INVD1 U1338 ( .I(n2391), .ZN(n1750) );
  INVD1 U1339 ( .I(n2392), .ZN(n1749) );
  INVD1 U1340 ( .I(n2356), .ZN(n1889) );
  BUFFD1 U1341 ( .I(n2282), .Z(n2281) );
  INVD1 U1342 ( .I(n2288), .ZN(n2287) );
  INVD1 U1343 ( .I(n2300), .ZN(n2299) );
  INVD1 U1344 ( .I(n2311), .ZN(n2310) );
  INVD1 U1345 ( .I(n2313), .ZN(n2312) );
  INVD1 U1346 ( .I(n2394), .ZN(n2393) );
  INVD1 U1347 ( .I(n2402), .ZN(n2401) );
  INVD1 U1348 ( .I(n2410), .ZN(n2409) );
  INVD1 U1349 ( .I(n2418), .ZN(n2417) );
  INVD1 U1350 ( .I(n2420), .ZN(n2419) );
  INVD1 U1351 ( .I(n2422), .ZN(n2421) );
  INVD1 U1352 ( .I(n2336), .ZN(n2335) );
  INVD1 U1353 ( .I(n2334), .ZN(n2333) );
  INVD1 U1354 ( .I(n2358), .ZN(n2357) );
  INVD1 U1355 ( .I(n2366), .ZN(n2365) );
  INVD1 U1356 ( .I(n2374), .ZN(n2373) );
  INVD1 U1357 ( .I(n2382), .ZN(n2381) );
  INVD1 U1358 ( .I(n2384), .ZN(n2383) );
  INVD1 U1359 ( .I(n2386), .ZN(n2385) );
  INVD1 U1360 ( .I(n2317), .ZN(n2316) );
  INVD1 U1361 ( .I(n2396), .ZN(n2395) );
  INVD1 U1362 ( .I(n2398), .ZN(n2397) );
  INVD1 U1363 ( .I(n2404), .ZN(n2403) );
  INVD1 U1364 ( .I(n2406), .ZN(n2405) );
  INVD1 U1365 ( .I(n2424), .ZN(n2423) );
  INVD1 U1366 ( .I(n2360), .ZN(n2359) );
  INVD1 U1367 ( .I(n2362), .ZN(n2361) );
  INVD1 U1368 ( .I(n2368), .ZN(n2367) );
  INVD1 U1369 ( .I(n2370), .ZN(n2369) );
  INVD1 U1370 ( .I(n2315), .ZN(n2314) );
  INVD1 U1371 ( .I(n2400), .ZN(n2399) );
  INVD1 U1372 ( .I(n2412), .ZN(n2411) );
  INVD1 U1373 ( .I(n2414), .ZN(n2413) );
  INVD1 U1374 ( .I(n2416), .ZN(n2415) );
  INVD1 U1375 ( .I(n2340), .ZN(n2339) );
  INVD1 U1376 ( .I(n2338), .ZN(n2337) );
  INVD1 U1377 ( .I(n2364), .ZN(n2363) );
  INVD1 U1378 ( .I(n2376), .ZN(n2375) );
  INVD1 U1379 ( .I(n2378), .ZN(n2377) );
  INVD1 U1380 ( .I(n2380), .ZN(n2379) );
  INVD1 U1381 ( .I(n2388), .ZN(n2387) );
  INVD1 U1382 ( .I(n2320), .ZN(n2319) );
  INVD1 U1383 ( .I(n2320), .ZN(n2318) );
  INVD1 U1384 ( .I(n2323), .ZN(n2322) );
  INVD1 U1385 ( .I(n2323), .ZN(n2321) );
  INVD1 U1386 ( .I(n2346), .ZN(n2345) );
  INVD1 U1387 ( .I(n2346), .ZN(n2344) );
  INVD1 U1388 ( .I(n2343), .ZN(n2342) );
  INVD1 U1389 ( .I(n2343), .ZN(n2341) );
  INVD1 U1390 ( .I(n1297), .ZN(n2181) );
  INVD1 U1391 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N193 ), .ZN(n2311) );
  INVD1 U1392 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N226 ), .ZN(n2313) );
  INVD1 U1393 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N132 ), .ZN(n2394) );
  INVD1 U1394 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N264 ), .ZN(n2402) );
  INVD1 U1395 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N396 ), .ZN(n2410) );
  INVD1 U1396 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N528 ), .ZN(n2418) );
  INVD1 U1397 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N561 ), .ZN(n2420) );
  INVD1 U1398 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N594 ), .ZN(n2422) );
  INVD1 U1399 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N226 ), .ZN(n2336) );
  INVD1 U1400 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N193 ), .ZN(n2334) );
  INVD1 U1401 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N132 ), .ZN(n2358) );
  INVD1 U1402 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N264 ), .ZN(n2366) );
  INVD1 U1403 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N396 ), .ZN(n2374) );
  INVD1 U1404 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N528 ), .ZN(n2382) );
  INVD1 U1405 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N561 ), .ZN(n2384) );
  INVD1 U1406 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N594 ), .ZN(n2386) );
  INVD1 U1407 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N165 ), .ZN(n2396) );
  INVD1 U1408 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N198 ), .ZN(n2398) );
  INVD1 U1409 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N297 ), .ZN(n2404) );
  INVD1 U1410 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N330 ), .ZN(n2406) );
  INVD1 U1411 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N429 ), .ZN(n2412) );
  INVD1 U1412 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N462 ), .ZN(n2414) );
  INVD1 U1413 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N165 ), .ZN(n2360) );
  INVD1 U1414 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N198 ), .ZN(n2362) );
  INVD1 U1415 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N297 ), .ZN(n2368) );
  INVD1 U1416 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N330 ), .ZN(n2370) );
  INVD1 U1417 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N429 ), .ZN(n2376) );
  INVD1 U1418 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N462 ), .ZN(n2378) );
  INVD1 U1419 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N292 ), .ZN(n2317) );
  INVD1 U1420 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N231 ), .ZN(n2400) );
  INVD1 U1421 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N495 ), .ZN(n2416) );
  INVD1 U1422 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N627 ), .ZN(n2424) );
  INVD1 U1423 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N231 ), .ZN(n2364) );
  INVD1 U1424 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N495 ), .ZN(n2380) );
  INVD1 U1425 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N627 ), .ZN(n2388) );
  INVD1 U1426 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N259 ), .ZN(n2315) );
  INVD1 U1427 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N292 ), .ZN(n2340) );
  INVD1 U1428 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N259 ), .ZN(n2338) );
  INVD1 U1429 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ), .ZN(n2320) );
  INVD1 U1430 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ), .ZN(n2323) );
  INVD1 U1431 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ), .ZN(n2346) );
  INVD1 U1432 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ), .ZN(n2343) );
  BUFFD1 U1433 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .Z(n1755) );
  BUFFD1 U1434 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .Z(n1896) );
  BUFFD1 U1435 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1891) );
  BUFFD1 U1436 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .Z(n2114) );
  BUFFD1 U1437 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .Z(n2011) );
  BUFFD1 U1438 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .Z(n2110) );
  BUFFD1 U1439 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .Z(n2007) );
  BUFFD1 U1440 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .Z(n1756) );
  BUFFD1 U1441 ( .I(n1247), .Z(n2182) );
  BUFFD1 U1442 ( .I(n2286), .Z(n2285) );
  BUFFD1 U1443 ( .I(n2286), .Z(n2284) );
  BUFFD1 U1444 ( .I(n2286), .Z(n2283) );
  BUFFD1 U1445 ( .I(n2295), .Z(n2297) );
  BUFFD1 U1446 ( .I(n2298), .Z(n2296) );
  BUFFD1 U1447 ( .I(n2275), .Z(n2282) );
  BUFFD1 U1448 ( .I(n2298), .Z(n2295) );
  BUFFD1 U1449 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1751) );
  BUFFD1 U1450 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .Z(n1895) );
  INVD1 U1451 ( .I(n2326), .ZN(n2005) );
  INVD1 U1452 ( .I(n2408), .ZN(n2407) );
  INVD1 U1453 ( .I(n2372), .ZN(n2371) );
  INVD1 U1454 ( .I(n2306), .ZN(n2305) );
  INVD1 U1455 ( .I(n2306), .ZN(n2304) );
  INVD1 U1456 ( .I(n2309), .ZN(n2308) );
  INVD1 U1457 ( .I(n2309), .ZN(n2307) );
  INVD1 U1458 ( .I(n2332), .ZN(n2331) );
  INVD1 U1459 ( .I(n2332), .ZN(n2330) );
  INVD1 U1460 ( .I(n2329), .ZN(n2328) );
  INVD1 U1461 ( .I(n2329), .ZN(n2327) );
  INVD1 U1462 ( .I(n721), .ZN(n2347) );
  INVD1 U1463 ( .I(n869), .ZN(n2426) );
  INVD1 U1464 ( .I(n1015), .ZN(n2348) );
  INVD1 U1465 ( .I(n1314), .ZN(n2425) );
  INVD1 U1466 ( .I(n2350), .ZN(n2349) );
  INVD1 U1467 ( .I(n2352), .ZN(n2351) );
  BUFFD1 U1468 ( .I(\SerDes_U2/Des_U1/DesDec_Rx1/SerClock ), .Z(n2286) );
  BUFFD1 U1469 ( .I(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock ), .Z(n2298) );
  INVD1 U1470 ( .I(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), .ZN(n2350) );
  INVD1 U1471 ( .I(\SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .ZN(n2352) );
  INVD1 U1472 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N363 ), .ZN(n2372) );
  INVD1 U1473 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N363 ), .ZN(n2408) );
  INVD1 U1474 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ), .ZN(n2306) );
  INVD1 U1475 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ), .ZN(n2309) );
  INVD1 U1476 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ), .ZN(n2332) );
  INVD1 U1477 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ), .ZN(n2329) );
  INVD1 U1478 ( .I(n2434), .ZN(n2431) );
  INVD1 U1479 ( .I(n2430), .ZN(n2427) );
  MUX4ND0 U1480 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2110), .ZN(n2032) );
  MUX4ND0 U1481 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2035) );
  MUX4ND0 U1482 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .S0(n2114), .S1(
        n2110), .ZN(n2038) );
  MUX4ND0 U1483 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .S0(n2114), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2041) );
  MUX4ND0 U1484 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2044) );
  MUX4ND0 U1485 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .S0(n2114), 
        .S1(n2110), .ZN(n2047) );
  MUX4ND0 U1486 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2110), .ZN(n2050) );
  MUX4ND0 U1487 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .S0(n2114), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2053) );
  MUX4ND0 U1488 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .S0(n2114), 
        .S1(n2110), .ZN(n2056) );
  MUX4ND0 U1489 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .S0(n2114), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2059) );
  MUX4ND0 U1490 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2062) );
  MUX4ND0 U1491 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .S0(n2111), 
        .S1(n2110), .ZN(n2065) );
  MUX4ND0 U1492 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .S0(n2114), 
        .S1(n2110), .ZN(n2068) );
  MUX4ND0 U1493 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2110), .ZN(n2071) );
  MUX4ND0 U1494 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .S0(n2114), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2074) );
  MUX4ND0 U1495 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .S0(n2114), 
        .S1(n2110), .ZN(n2089) );
  MUX4ND0 U1496 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2092) );
  MUX4ND0 U1497 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2109), .ZN(n2095) );
  MUX4ND0 U1498 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .S0(n2111), 
        .S1(n2110), .ZN(n2098) );
  MUX4ND0 U1499 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2007), .ZN(n1995) );
  MUX4ND0 U1500 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .S0(n2011), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1992) );
  MUX4ND0 U1501 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .S0(n2011), 
        .S1(n2007), .ZN(n1989) );
  MUX4ND0 U1502 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2007), .ZN(n1986) );
  MUX4ND0 U1503 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1971) );
  MUX4ND0 U1504 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .S0(n2011), 
        .S1(n2007), .ZN(n1968) );
  MUX4ND0 U1505 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .S0(n2011), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1965) );
  MUX4ND0 U1506 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1962) );
  MUX4ND0 U1507 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2007), .ZN(n1959) );
  MUX4ND0 U1508 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .S0(n2011), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1956) );
  MUX4ND0 U1509 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .S0(n2008), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1953) );
  MUX4ND0 U1510 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .S0(n2011), 
        .S1(n2007), .ZN(n1950) );
  MUX4ND0 U1511 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1947) );
  MUX4ND0 U1512 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .S0(n2011), 
        .S1(n2007), .ZN(n1944) );
  MUX4ND0 U1513 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2007), .ZN(n1941) );
  MUX4ND0 U1514 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .S0(n2011), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1938) );
  MUX4ND0 U1515 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .S0(n2011), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1935) );
  MUX4ND0 U1516 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1932) );
  MUX4ND0 U1517 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .S0(n2008), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1929) );
  MUX4ND0 U1518 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .S0(n2114), .S1(
        n2110), .ZN(n2014) );
  MUX4ND0 U1519 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2109), .ZN(n2017) );
  MUX4ND0 U1520 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .S0(n2114), .S1(
        n2110), .ZN(n2020) );
  MUX4ND0 U1521 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .S0(n2111), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2023) );
  MUX4ND0 U1522 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .S0(n2112), .S1(
        n2109), .ZN(n2026) );
  MUX4ND0 U1523 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .S0(n2114), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2029) );
  MUX4ND0 U1524 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .S0(n2114), 
        .S1(n2110), .ZN(n2077) );
  MUX4ND0 U1525 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .S0(n2113), 
        .S1(n2110), .ZN(n2080) );
  MUX4ND0 U1526 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2083) );
  MUX4ND0 U1527 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .S0(n2114), 
        .S1(n2110), .ZN(n2086) );
  MUX4ND0 U1528 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(n2110), .ZN(n2101) );
  MUX4ND0 U1529 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .S0(n2114), 
        .S1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2104) );
  MUX4ND0 U1530 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2107) );
  MUX4ND0 U1531 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n2004) );
  MUX4ND0 U1532 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .S0(n2008), 
        .S1(n2007), .ZN(n2001) );
  MUX4ND0 U1533 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .S0(n2011), 
        .S1(n2007), .ZN(n1998) );
  MUX4ND0 U1534 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .S0(n2011), 
        .S1(n2007), .ZN(n1983) );
  MUX4ND0 U1535 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .S0(n2011), 
        .S1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1980) );
  MUX4ND0 U1536 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .S0(n2011), 
        .S1(n2007), .ZN(n1977) );
  MUX4ND0 U1537 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .S0(n2010), 
        .S1(n2007), .ZN(n1974) );
  MUX4ND0 U1538 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .S0(n2011), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1926) );
  MUX4ND0 U1539 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2006), .ZN(n1923) );
  MUX4ND0 U1540 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2007), .ZN(n1920) );
  MUX4ND0 U1541 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .S0(n2009), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n1917) );
  MUX4ND0 U1542 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .S1(n2006), .ZN(n1914) );
  MUX4ND0 U1543 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .S0(n2011), .S1(
        n2006), .ZN(n1911) );
  AN2D1 U1544 ( .A1(n2431), .A2(n2432), .Z(\SerDes_U2/Ser_U1/SerEnc_Tx1/N24 )
         );
  AN2D1 U1545 ( .A1(n2427), .A2(n2428), .Z(\SerDes_U1/Ser_U1/SerEnc_Tx1/N24 )
         );
  ND2D1 U1546 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .ZN(n2434) );
  ND2D1 U1547 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .ZN(n2430) );
  INVD1 U1548 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .ZN(n2734) );
  INVD1 U1549 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .ZN(n2391) );
  MUX4D0 U1550 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][2] ), .S0(n1757), 
        .S1(n1753), .Z(n1629) );
  MUX4D0 U1551 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][3] ), .S0(n1759), 
        .S1(n1753), .Z(n1633) );
  MUX4D0 U1552 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][4] ), .S0(n1760), 
        .S1(n1753), .Z(n1637) );
  MUX4D0 U1553 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][5] ), .S0(n1755), 
        .S1(n1754), .Z(n1641) );
  MUX4D0 U1554 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][6] ), .S0(n1757), 
        .S1(n1754), .Z(n1645) );
  MUX4D0 U1555 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][7] ), .S0(n1759), 
        .S1(n1754), .Z(n1649) );
  MUX4D0 U1556 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][8] ), .S0(n1755), 
        .S1(n1752), .Z(n1653) );
  MUX4D0 U1557 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][9] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1751), .Z(n1657) );
  MUX4D0 U1558 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][10] ), .S0(n1755), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1661) );
  MUX4D0 U1559 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][11] ), .S0(n1755), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1665) );
  MUX4D0 U1560 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][12] ), .S0(n1756), 
        .S1(n1751), .Z(n1669) );
  MUX4D0 U1561 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][13] ), .S0(n1756), 
        .S1(n1753), .Z(n1673) );
  MUX4D0 U1562 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][14] ), .S0(n1756), 
        .S1(n1754), .Z(n1677) );
  MUX4D0 U1563 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][15] ), .S0(n1756), 
        .S1(n1752), .Z(n1681) );
  MUX4D0 U1564 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][16] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1753), .Z(n1685) );
  MUX4D0 U1565 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][17] ), .S0(n1757), 
        .S1(n1751), .Z(n1689) );
  MUX4D0 U1566 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][18] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1693) );
  MUX4D0 U1567 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][19] ), .S0(n1757), 
        .S1(n1752), .Z(n1697) );
  MUX4D0 U1568 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][20] ), .S0(n1758), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1701) );
  MUX4D0 U1569 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][21] ), .S0(n1758), 
        .S1(n1752), .Z(n1705) );
  MUX4D0 U1570 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][22] ), .S0(n1758), 
        .S1(n1752), .Z(n1709) );
  MUX4D0 U1571 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][23] ), .S0(n1759), 
        .S1(n1753), .Z(n1713) );
  MUX4D0 U1572 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][24] ), .S0(n1759), 
        .S1(n1751), .Z(n1717) );
  MUX4D0 U1573 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][25] ), .S0(n1759), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1721) );
  MUX4D0 U1574 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][26] ), .S0(n1755), 
        .S1(n1753), .Z(n1725) );
  MUX4D0 U1575 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][27] ), .S0(n1756), 
        .S1(n1752), .Z(n1729) );
  MUX4D0 U1576 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][28] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1754), .Z(n1733) );
  MUX4D0 U1577 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][29] ), .S0(n1760), 
        .S1(n1751), .Z(n1737) );
  MUX4D0 U1578 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][30] ), .S0(n1760), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1741) );
  MUX4D0 U1579 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][31] ), .S0(n1760), 
        .S1(n1752), .Z(n1745) );
  MUX4D0 U1580 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][2] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1893), .Z(n1769) );
  MUX4D0 U1581 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][3] ), .S0(n1896), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1773) );
  MUX4D0 U1582 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][4] ), .S0(n1895), 
        .S1(n1891), .Z(n1777) );
  MUX4D0 U1583 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][5] ), .S0(n1898), 
        .S1(n1891), .Z(n1781) );
  MUX4D0 U1584 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][6] ), .S0(n1898), 
        .S1(n1892), .Z(n1785) );
  MUX4D0 U1585 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][7] ), .S0(n1898), 
        .S1(n1891), .Z(n1789) );
  MUX4D0 U1586 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][8] ), .S0(n1897), 
        .S1(n1891), .Z(n1793) );
  MUX4D0 U1587 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][9] ), .S0(n1896), 
        .S1(n1891), .Z(n1797) );
  MUX4D0 U1588 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][10] ), .S0(n1899), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1801) );
  MUX4D0 U1589 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][11] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1805) );
  MUX4D0 U1590 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][12] ), .S0(n1900), 
        .S1(n1893), .Z(n1809) );
  MUX4D0 U1591 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][13] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1813) );
  MUX4D0 U1592 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][14] ), .S0(n1898), 
        .S1(n1893), .Z(n1817) );
  MUX4D0 U1593 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][15] ), .S0(n1895), 
        .S1(n1891), .Z(n1821) );
  MUX4D0 U1594 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][16] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1892), .Z(n1825) );
  MUX4D0 U1595 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][17] ), .S0(n1900), 
        .S1(n1892), .Z(n1829) );
  MUX4D0 U1596 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][18] ), .S0(n1900), 
        .S1(n1892), .Z(n1833) );
  MUX4D0 U1597 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][19] ), .S0(n1896), 
        .S1(n1892), .Z(n1837) );
  MUX4D0 U1598 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][20] ), .S0(n1896), 
        .S1(n1894), .Z(n1841) );
  MUX4D0 U1599 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][21] ), .S0(n1898), 
        .S1(n1893), .Z(n1845) );
  MUX4D0 U1600 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][22] ), .S0(n1895), 
        .S1(n1892), .Z(n1849) );
  MUX4D0 U1601 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][23] ), .S0(n1895), 
        .S1(n1891), .Z(n1853) );
  MUX4D0 U1602 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][24] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1857) );
  MUX4D0 U1603 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][25] ), .S0(n1897), 
        .S1(n1894), .Z(n1861) );
  MUX4D0 U1604 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][26] ), .S0(n1899), 
        .S1(n1893), .Z(n1865) );
  MUX4D0 U1605 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][27] ), .S0(n1899), 
        .S1(n1893), .Z(n1869) );
  MUX4D0 U1606 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][28] ), .S0(n1899), 
        .S1(n1893), .Z(n1873) );
  MUX4D0 U1607 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][29] ), .S0(n1900), 
        .S1(n1894), .Z(n1877) );
  MUX4D0 U1608 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][30] ), .S0(n1900), 
        .S1(n1894), .Z(n1881) );
  MUX4D0 U1609 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][31] ), .S0(n1900), 
        .S1(n1894), .Z(n1885) );
  MUX4D0 U1610 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][0] ), .S0(n1897), 
        .S1(n1892), .Z(n1761) );
  MUX4D0 U1611 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[12][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[13][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[14][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[15][1] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1765) );
  MUX4D0 U1612 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][0] ), .S0(n1758), 
        .S1(n1752), .Z(n1621) );
  MUX4D0 U1613 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[12][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[13][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[14][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[15][1] ), .S0(n1755), 
        .S1(n1752), .Z(n1625) );
  INVD1 U1614 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(n2303) );
  MUX4ND0 U1615 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[0] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[1] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[2] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[3] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1534) );
  MUX4ND0 U1616 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[4] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[5] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[6] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[7] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1535) );
  MUX4ND0 U1617 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[24] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[25] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[26] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[27] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1536) );
  MUX4ND0 U1618 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[28] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[29] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[30] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[31] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1537) );
  MUX4ND0 U1619 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[16] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[17] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[18] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[19] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1538) );
  MUX4ND0 U1620 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[20] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[21] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[22] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[23] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1539) );
  MUX4ND0 U1621 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[8] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[9] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[10] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[11] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1540) );
  MUX4ND0 U1622 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[12] ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[13] ), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[14] ), .I3(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/InBuf[15] ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1541) );
  MUX4ND0 U1623 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[0] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[1] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[2] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[3] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1542) );
  MUX4ND0 U1624 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[4] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[5] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[6] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[7] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1543) );
  MUX4ND0 U1625 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[24] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[25] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[26] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[27] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1544) );
  MUX4ND0 U1626 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[28] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[29] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[30] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[31] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1545) );
  MUX4ND0 U1627 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[16] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[17] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[18] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[19] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1546) );
  MUX4ND0 U1628 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[20] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[21] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[22] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[23] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1547) );
  MUX4ND0 U1629 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[8] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[9] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[10] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[11] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1548) );
  MUX4ND0 U1630 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[12] ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[13] ), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[14] ), .I3(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/InBuf[15] ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .S1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .ZN(n1549) );
  INVD1 U1631 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .ZN(n2392) );
  INVD1 U1632 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .ZN(n2354) );
  INVD1 U1633 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .ZN(n2302) );
  INVD1 U1634 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .ZN(n2356) );
  INVD1 U1635 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .ZN(n2353) );
  INVD1 U1636 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .ZN(n2630) );
  MUX4D0 U1637 ( .I0(n1624), .I1(n1622), .I2(n1623), .I3(n1621), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ) );
  MUX4D0 U1638 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][0] ), .S0(n1760), .S1(
        n1752), .Z(n1623) );
  MUX4D0 U1639 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][0] ), .S0(n1757), 
        .S1(n1752), .Z(n1622) );
  MUX4D0 U1640 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .S0(n1759), .S1(
        n1752), .Z(n1624) );
  MUX4D0 U1641 ( .I0(n1628), .I1(n1626), .I2(n1627), .I3(n1625), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ) );
  MUX4D0 U1642 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][1] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1752), .Z(n1627) );
  MUX4D0 U1643 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][1] ), .S0(n1758), 
        .S1(n1752), .Z(n1626) );
  MUX4D0 U1644 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1752), .Z(n1628) );
  MUX4D0 U1645 ( .I0(n1632), .I1(n1630), .I2(n1631), .I3(n1629), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ) );
  MUX4D0 U1646 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][2] ), .S0(n1758), .S1(
        n1753), .Z(n1631) );
  MUX4D0 U1647 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][2] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1753), .Z(n1630) );
  MUX4D0 U1648 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .S0(n1756), .S1(
        n1753), .Z(n1632) );
  MUX4D0 U1649 ( .I0(n1636), .I1(n1634), .I2(n1635), .I3(n1633), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ) );
  MUX4D0 U1650 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][3] ), .S0(n1759), .S1(
        n1753), .Z(n1635) );
  MUX4D0 U1651 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][3] ), .S0(n1757), 
        .S1(n1753), .Z(n1634) );
  MUX4D0 U1652 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .S0(n1755), .S1(
        n1753), .Z(n1636) );
  MUX4D0 U1653 ( .I0(n1640), .I1(n1638), .I2(n1639), .I3(n1637), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ) );
  MUX4D0 U1654 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][4] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1753), .Z(n1639) );
  MUX4D0 U1655 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][4] ), .S0(n1756), 
        .S1(n1753), .Z(n1638) );
  MUX4D0 U1656 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .S0(n1760), .S1(
        n1753), .Z(n1640) );
  MUX4D0 U1657 ( .I0(n1644), .I1(n1642), .I2(n1643), .I3(n1641), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ) );
  MUX4D0 U1658 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][5] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1754), .Z(n1643) );
  MUX4D0 U1659 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][5] ), .S0(n1756), 
        .S1(n1754), .Z(n1642) );
  MUX4D0 U1660 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .S0(n1760), .S1(
        n1754), .Z(n1644) );
  MUX4D0 U1661 ( .I0(n1648), .I1(n1646), .I2(n1647), .I3(n1645), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ) );
  MUX4D0 U1662 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][6] ), .S0(n1755), .S1(
        n1754), .Z(n1647) );
  MUX4D0 U1663 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][6] ), .S0(n1756), 
        .S1(n1754), .Z(n1646) );
  MUX4D0 U1664 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .S0(n1758), .S1(
        n1754), .Z(n1648) );
  MUX4D0 U1665 ( .I0(n1652), .I1(n1650), .I2(n1651), .I3(n1649), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ) );
  MUX4D0 U1666 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][7] ), .S0(n1760), .S1(
        n1754), .Z(n1651) );
  MUX4D0 U1667 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][7] ), .S0(n1759), 
        .S1(n1754), .Z(n1650) );
  MUX4D0 U1668 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .S0(n1757), .S1(
        n1754), .Z(n1652) );
  MUX4D0 U1669 ( .I0(n1656), .I1(n1654), .I2(n1655), .I3(n1653), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ) );
  MUX4D0 U1670 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][8] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1753), .Z(n1655) );
  MUX4D0 U1671 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][8] ), .S0(n1757), 
        .S1(n1751), .Z(n1654) );
  MUX4D0 U1672 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .S0(n1756), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1656) );
  MUX4D0 U1673 ( .I0(n1660), .I1(n1658), .I2(n1659), .I3(n1657), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ) );
  MUX4D0 U1674 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][9] ), .S0(n1756), .S1(
        n1753), .Z(n1659) );
  MUX4D0 U1675 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][9] ), .S0(n1755), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1658) );
  MUX4D0 U1676 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .S0(n1756), .S1(
        n1754), .Z(n1660) );
  MUX4D0 U1677 ( .I0(n1664), .I1(n1662), .I2(n1663), .I3(n1661), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ) );
  MUX4D0 U1678 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][10] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1663) );
  MUX4D0 U1679 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][10] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1752), .Z(n1662) );
  MUX4D0 U1680 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1752), .Z(n1664) );
  MUX4D0 U1681 ( .I0(n1668), .I1(n1666), .I2(n1667), .I3(n1665), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ) );
  MUX4D0 U1682 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][11] ), .S0(n1755), 
        .S1(n1751), .Z(n1667) );
  MUX4D0 U1683 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][11] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1666) );
  MUX4D0 U1684 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .S0(n1758), 
        .S1(n1752), .Z(n1668) );
  MUX4D0 U1685 ( .I0(n1672), .I1(n1670), .I2(n1671), .I3(n1669), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ) );
  MUX4D0 U1686 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][12] ), .S0(n1758), 
        .S1(n1751), .Z(n1671) );
  MUX4D0 U1687 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][12] ), .S0(n1755), 
        .S1(n1752), .Z(n1670) );
  MUX4D0 U1688 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .S0(n1756), 
        .S1(n1754), .Z(n1672) );
  MUX4D0 U1689 ( .I0(n1676), .I1(n1674), .I2(n1675), .I3(n1673), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ) );
  MUX4D0 U1690 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][13] ), .S0(n1755), 
        .S1(n1753), .Z(n1675) );
  MUX4D0 U1691 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][13] ), .S0(n1756), 
        .S1(n1751), .Z(n1674) );
  MUX4D0 U1692 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1676) );
  MUX4D0 U1693 ( .I0(n1680), .I1(n1678), .I2(n1679), .I3(n1677), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ) );
  MUX4D0 U1694 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][14] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1753), .Z(n1679) );
  MUX4D0 U1695 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][14] ), .S0(n1756), 
        .S1(n1752), .Z(n1678) );
  MUX4D0 U1696 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .S0(n1755), 
        .S1(n1754), .Z(n1680) );
  MUX4D0 U1697 ( .I0(n1684), .I1(n1682), .I2(n1683), .I3(n1681), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ) );
  MUX4D0 U1698 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][15] ), .S0(n1756), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1683) );
  MUX4D0 U1699 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][15] ), .S0(n1755), 
        .S1(n1751), .Z(n1682) );
  MUX4D0 U1700 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .S0(n1759), 
        .S1(n1754), .Z(n1684) );
  MUX4D0 U1701 ( .I0(n1688), .I1(n1686), .I2(n1687), .I3(n1685), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ) );
  MUX4D0 U1702 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][16] ), .S0(n1755), 
        .S1(n1752), .Z(n1687) );
  MUX4D0 U1703 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][16] ), .S0(n1758), 
        .S1(n1754), .Z(n1686) );
  MUX4D0 U1704 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .S0(n1756), 
        .S1(n1752), .Z(n1688) );
  MUX4D0 U1705 ( .I0(n1692), .I1(n1690), .I2(n1691), .I3(n1689), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ) );
  MUX4D0 U1706 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][17] ), .S0(n1757), 
        .S1(n1751), .Z(n1691) );
  MUX4D0 U1707 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][17] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1690) );
  MUX4D0 U1708 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1692) );
  MUX4D0 U1709 ( .I0(n1696), .I1(n1694), .I2(n1695), .I3(n1693), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ) );
  MUX4D0 U1710 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][18] ), .S0(n1757), 
        .S1(n1751), .Z(n1695) );
  MUX4D0 U1711 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][18] ), .S0(n1757), 
        .S1(n1752), .Z(n1694) );
  MUX4D0 U1712 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1696) );
  MUX4D0 U1713 ( .I0(n1700), .I1(n1698), .I2(n1699), .I3(n1697), .S0(n1749), 
        .S1(n1750), .Z(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ) );
  MUX4D0 U1714 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][19] ), .S0(n1757), 
        .S1(n1753), .Z(n1699) );
  MUX4D0 U1715 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][19] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1698) );
  MUX4D0 U1716 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .S0(n1757), 
        .S1(n1751), .Z(n1700) );
  MUX4D0 U1717 ( .I0(n1704), .I1(n1702), .I2(n1703), .I3(n1701), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ) );
  MUX4D0 U1718 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][20] ), .S0(n1758), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1703) );
  MUX4D0 U1719 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][20] ), .S0(n1758), 
        .S1(n1751), .Z(n1702) );
  MUX4D0 U1720 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .S0(n1758), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1704) );
  MUX4D0 U1721 ( .I0(n1708), .I1(n1706), .I2(n1707), .I3(n1705), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ) );
  MUX4D0 U1722 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][21] ), .S0(n1758), 
        .S1(n1751), .Z(n1707) );
  MUX4D0 U1723 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][21] ), .S0(n1758), 
        .S1(n1753), .Z(n1706) );
  MUX4D0 U1724 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .S0(n1758), 
        .S1(n1751), .Z(n1708) );
  MUX4D0 U1725 ( .I0(n1712), .I1(n1710), .I2(n1711), .I3(n1709), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ) );
  MUX4D0 U1726 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][22] ), .S0(n1758), 
        .S1(n1751), .Z(n1711) );
  MUX4D0 U1727 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][22] ), .S0(n1758), 
        .S1(n1753), .Z(n1710) );
  MUX4D0 U1728 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .S0(n1758), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1712) );
  MUX4D0 U1729 ( .I0(n1716), .I1(n1714), .I2(n1715), .I3(n1713), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ) );
  MUX4D0 U1730 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][23] ), .S0(n1759), 
        .S1(n1751), .Z(n1715) );
  MUX4D0 U1731 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][23] ), .S0(n1759), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1714) );
  MUX4D0 U1732 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .S0(n1759), 
        .S1(n1754), .Z(n1716) );
  MUX4D0 U1733 ( .I0(n1720), .I1(n1718), .I2(n1719), .I3(n1717), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ) );
  MUX4D0 U1734 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][24] ), .S0(n1759), 
        .S1(n1751), .Z(n1719) );
  MUX4D0 U1735 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][24] ), .S0(n1759), 
        .S1(n1754), .Z(n1718) );
  MUX4D0 U1736 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .S0(n1759), 
        .S1(n1751), .Z(n1720) );
  MUX4D0 U1737 ( .I0(n1724), .I1(n1722), .I2(n1723), .I3(n1721), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ) );
  MUX4D0 U1738 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][25] ), .S0(n1759), 
        .S1(n1751), .Z(n1723) );
  MUX4D0 U1739 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][25] ), .S0(n1759), 
        .S1(n1752), .Z(n1722) );
  MUX4D0 U1740 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .S0(n1759), 
        .S1(n1754), .Z(n1724) );
  MUX4D0 U1741 ( .I0(n1728), .I1(n1726), .I2(n1727), .I3(n1725), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ) );
  MUX4D0 U1742 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][26] ), .S0(n1755), 
        .S1(n1753), .Z(n1727) );
  MUX4D0 U1743 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][26] ), .S0(n1759), 
        .S1(n1751), .Z(n1726) );
  MUX4D0 U1744 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .S0(n1755), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1728) );
  MUX4D0 U1745 ( .I0(n1732), .I1(n1730), .I2(n1731), .I3(n1729), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ) );
  MUX4D0 U1746 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][27] ), .S0(n1757), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1731) );
  MUX4D0 U1747 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][27] ), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .S1(n1752), .Z(n1730) );
  MUX4D0 U1748 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .S0(n1756), 
        .S1(n1754), .Z(n1732) );
  MUX4D0 U1749 ( .I0(n1736), .I1(n1734), .I2(n1735), .I3(n1733), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(n1750), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ) );
  MUX4D0 U1750 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][28] ), .S0(n1760), 
        .S1(n1752), .Z(n1735) );
  MUX4D0 U1751 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][28] ), .S0(n1756), 
        .S1(n1753), .Z(n1734) );
  MUX4D0 U1752 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .S0(n1760), 
        .S1(n1751), .Z(n1736) );
  MUX4D0 U1753 ( .I0(n1740), .I1(n1738), .I2(n1739), .I3(n1737), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N52 ) );
  MUX4D0 U1754 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][29] ), .S0(n1760), 
        .S1(n1753), .Z(n1739) );
  MUX4D0 U1755 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][29] ), .S0(n1760), 
        .S1(n1752), .Z(n1738) );
  MUX4D0 U1756 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .S0(n1760), 
        .S1(n1754), .Z(n1740) );
  MUX4D0 U1757 ( .I0(n1744), .I1(n1742), .I2(n1743), .I3(n1741), .S0(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N51 ) );
  MUX4D0 U1758 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][30] ), .S0(n1760), 
        .S1(n1754), .Z(n1743) );
  MUX4D0 U1759 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][30] ), .S0(n1760), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .Z(n1742) );
  MUX4D0 U1760 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .S0(n1760), 
        .S1(n1751), .Z(n1744) );
  MUX4D0 U1761 ( .I0(n1748), .I1(n1746), .I2(n1747), .I3(n1745), .S0(n1749), 
        .S1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ) );
  MUX4D0 U1762 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[7][31] ), .S0(n1760), 
        .S1(n1754), .Z(n1747) );
  MUX4D0 U1763 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[8][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[9][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[10][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[11][31] ), .S0(n1760), 
        .S1(n1751), .Z(n1746) );
  MUX4D0 U1764 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .I2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), .I3(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .S0(n1760), 
        .S1(n1754), .Z(n1748) );
  MUX4D0 U1765 ( .I0(n1764), .I1(n1762), .I2(n1763), .I3(n1761), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ) );
  MUX4D0 U1766 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][0] ), .S0(n1897), .S1(
        n1894), .Z(n1763) );
  MUX4D0 U1767 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][0] ), .S0(n1897), 
        .S1(n1893), .Z(n1762) );
  MUX4D0 U1768 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .S0(n1897), .S1(
        n1891), .Z(n1764) );
  MUX4D0 U1769 ( .I0(n1768), .I1(n1766), .I2(n1767), .I3(n1765), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ) );
  MUX4D0 U1770 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][1] ), .S0(n1897), .S1(
        n1893), .Z(n1767) );
  MUX4D0 U1771 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][1] ), .S0(n1897), 
        .S1(n1892), .Z(n1766) );
  MUX4D0 U1772 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .S0(n1897), .S1(
        n1894), .Z(n1768) );
  MUX4D0 U1773 ( .I0(n1772), .I1(n1770), .I2(n1771), .I3(n1769), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ) );
  MUX4D0 U1774 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][2] ), .S0(n1895), .S1(
        n1894), .Z(n1771) );
  MUX4D0 U1775 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][2] ), .S0(n1896), 
        .S1(n1893), .Z(n1770) );
  MUX4D0 U1776 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .S0(n1896), .S1(
        n1891), .Z(n1772) );
  MUX4D0 U1777 ( .I0(n1776), .I1(n1774), .I2(n1775), .I3(n1773), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ) );
  MUX4D0 U1778 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][3] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1893), .Z(n1775) );
  MUX4D0 U1779 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][3] ), .S0(n1896), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1774) );
  MUX4D0 U1780 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .S0(n1895), .S1(
        n1892), .Z(n1776) );
  MUX4D0 U1781 ( .I0(n1780), .I1(n1778), .I2(n1779), .I3(n1777), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ) );
  MUX4D0 U1782 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][4] ), .S0(n1895), .S1(
        n1891), .Z(n1779) );
  MUX4D0 U1783 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][4] ), .S0(n1895), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1778) );
  MUX4D0 U1784 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1780) );
  MUX4D0 U1785 ( .I0(n1784), .I1(n1782), .I2(n1783), .I3(n1781), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ) );
  MUX4D0 U1786 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][5] ), .S0(n1898), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1783) );
  MUX4D0 U1787 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][5] ), .S0(n1898), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1782) );
  MUX4D0 U1788 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .S0(n1898), .S1(
        n1893), .Z(n1784) );
  MUX4D0 U1789 ( .I0(n1788), .I1(n1786), .I2(n1787), .I3(n1785), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ) );
  MUX4D0 U1790 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][6] ), .S0(n1898), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1787) );
  MUX4D0 U1791 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][6] ), .S0(n1898), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1786) );
  MUX4D0 U1792 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .S0(n1898), .S1(
        n1891), .Z(n1788) );
  MUX4D0 U1793 ( .I0(n1792), .I1(n1790), .I2(n1791), .I3(n1789), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ) );
  MUX4D0 U1794 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][7] ), .S0(n1898), .S1(
        n1894), .Z(n1791) );
  MUX4D0 U1795 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][7] ), .S0(n1898), 
        .S1(n1892), .Z(n1790) );
  MUX4D0 U1796 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .S0(n1898), .S1(
        n1893), .Z(n1792) );
  MUX4D0 U1797 ( .I0(n1796), .I1(n1794), .I2(n1795), .I3(n1793), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ) );
  MUX4D0 U1798 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][8] ), .S0(n1898), .S1(
        n1891), .Z(n1795) );
  MUX4D0 U1799 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][8] ), .S0(n1895), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1794) );
  MUX4D0 U1800 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1796) );
  MUX4D0 U1801 ( .I0(n1800), .I1(n1798), .I2(n1799), .I3(n1797), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ) );
  MUX4D0 U1802 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][9] ), .S0(n1896), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1799) );
  MUX4D0 U1803 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][9] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1798) );
  MUX4D0 U1804 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .S0(n1900), .S1(
        n1891), .Z(n1800) );
  MUX4D0 U1805 ( .I0(n1804), .I1(n1802), .I2(n1803), .I3(n1801), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ) );
  MUX4D0 U1806 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][10] ), .S0(n1895), 
        .S1(n1893), .Z(n1803) );
  MUX4D0 U1807 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][10] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1802) );
  MUX4D0 U1808 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .S0(n1899), 
        .S1(n1891), .Z(n1804) );
  MUX4D0 U1809 ( .I0(n1808), .I1(n1806), .I2(n1807), .I3(n1805), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ) );
  MUX4D0 U1810 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][11] ), .S0(n1895), 
        .S1(n1891), .Z(n1807) );
  MUX4D0 U1811 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][11] ), .S0(n1898), 
        .S1(n1894), .Z(n1806) );
  MUX4D0 U1812 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .S0(n1896), 
        .S1(n1891), .Z(n1808) );
  MUX4D0 U1813 ( .I0(n1812), .I1(n1810), .I2(n1811), .I3(n1809), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ) );
  MUX4D0 U1814 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][12] ), .S0(n1899), 
        .S1(n1893), .Z(n1811) );
  MUX4D0 U1815 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][12] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1810) );
  MUX4D0 U1816 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .S0(n1896), 
        .S1(n1891), .Z(n1812) );
  MUX4D0 U1817 ( .I0(n1816), .I1(n1814), .I2(n1815), .I3(n1813), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ) );
  MUX4D0 U1818 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][13] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1815) );
  MUX4D0 U1819 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][13] ), .S0(n1897), 
        .S1(n1894), .Z(n1814) );
  MUX4D0 U1820 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .S0(n1900), 
        .S1(n1891), .Z(n1816) );
  MUX4D0 U1821 ( .I0(n1820), .I1(n1818), .I2(n1819), .I3(n1817), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ) );
  MUX4D0 U1822 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][14] ), .S0(n1900), 
        .S1(n1893), .Z(n1819) );
  MUX4D0 U1823 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][14] ), .S0(n1899), 
        .S1(n1894), .Z(n1818) );
  MUX4D0 U1824 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .S0(n1896), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1820) );
  MUX4D0 U1825 ( .I0(n1824), .I1(n1822), .I2(n1823), .I3(n1821), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ) );
  MUX4D0 U1826 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][15] ), .S0(n1898), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1823) );
  MUX4D0 U1827 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][15] ), .S0(n1898), 
        .S1(n1892), .Z(n1822) );
  MUX4D0 U1828 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .S0(n1895), 
        .S1(n1891), .Z(n1824) );
  MUX4D0 U1829 ( .I0(n1828), .I1(n1826), .I2(n1827), .I3(n1825), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ) );
  MUX4D0 U1830 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][16] ), .S0(n1896), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1827) );
  MUX4D0 U1831 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][16] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1893), .Z(n1826) );
  MUX4D0 U1832 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .S0(n1895), 
        .S1(n1894), .Z(n1828) );
  MUX4D0 U1833 ( .I0(n1832), .I1(n1830), .I2(n1831), .I3(n1829), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ) );
  MUX4D0 U1834 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][17] ), .S0(n1897), 
        .S1(n1892), .Z(n1831) );
  MUX4D0 U1835 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][17] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1892), .Z(n1830) );
  MUX4D0 U1836 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .S0(n1895), 
        .S1(n1892), .Z(n1832) );
  MUX4D0 U1837 ( .I0(n1836), .I1(n1834), .I2(n1835), .I3(n1833), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ) );
  MUX4D0 U1838 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][18] ), .S0(n1895), 
        .S1(n1892), .Z(n1835) );
  MUX4D0 U1839 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][18] ), .S0(n1896), 
        .S1(n1892), .Z(n1834) );
  MUX4D0 U1840 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1892), .Z(n1836) );
  MUX4D0 U1841 ( .I0(n1840), .I1(n1838), .I2(n1839), .I3(n1837), .S0(n1889), 
        .S1(n1890), .Z(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ) );
  MUX4D0 U1842 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][19] ), .S0(n1899), 
        .S1(n1892), .Z(n1839) );
  MUX4D0 U1843 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][19] ), .S0(n1898), 
        .S1(n1892), .Z(n1838) );
  MUX4D0 U1844 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1892), .Z(n1840) );
  MUX4D0 U1845 ( .I0(n1844), .I1(n1842), .I2(n1843), .I3(n1841), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ) );
  MUX4D0 U1846 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][20] ), .S0(n1896), 
        .S1(n1894), .Z(n1843) );
  MUX4D0 U1847 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][20] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1842) );
  MUX4D0 U1848 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1844) );
  MUX4D0 U1849 ( .I0(n1848), .I1(n1846), .I2(n1847), .I3(n1845), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ) );
  MUX4D0 U1850 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][21] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1847) );
  MUX4D0 U1851 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][21] ), .S0(n1895), 
        .S1(n1892), .Z(n1846) );
  MUX4D0 U1852 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .S0(n1900), 
        .S1(n1893), .Z(n1848) );
  MUX4D0 U1853 ( .I0(n1852), .I1(n1850), .I2(n1851), .I3(n1849), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ) );
  MUX4D0 U1854 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][22] ), .S0(n1897), 
        .S1(n1894), .Z(n1851) );
  MUX4D0 U1855 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][22] ), .S0(n1899), 
        .S1(n1892), .Z(n1850) );
  MUX4D0 U1856 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .S0(n1897), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1852) );
  MUX4D0 U1857 ( .I0(n1856), .I1(n1854), .I2(n1855), .I3(n1853), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ) );
  MUX4D0 U1858 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][23] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1894), .Z(n1855) );
  MUX4D0 U1859 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][23] ), .S0(n1895), 
        .S1(n1892), .Z(n1854) );
  MUX4D0 U1860 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .S0(n1896), 
        .S1(n1892), .Z(n1856) );
  MUX4D0 U1861 ( .I0(n1860), .I1(n1858), .I2(n1859), .I3(n1857), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ) );
  MUX4D0 U1862 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][24] ), .S0(n1895), 
        .S1(n1894), .Z(n1859) );
  MUX4D0 U1863 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][24] ), .S0(n1896), 
        .S1(n1892), .Z(n1858) );
  MUX4D0 U1864 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .S0(n1896), 
        .S1(n1891), .Z(n1860) );
  MUX4D0 U1865 ( .I0(n1864), .I1(n1862), .I2(n1863), .I3(n1861), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ) );
  MUX4D0 U1866 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][25] ), .S0(n1896), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .Z(n1863) );
  MUX4D0 U1867 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][25] ), .S0(n1897), 
        .S1(n1892), .Z(n1862) );
  MUX4D0 U1868 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), .S1(n1891), .Z(n1864) );
  MUX4D0 U1869 ( .I0(n1868), .I1(n1866), .I2(n1867), .I3(n1865), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ) );
  MUX4D0 U1870 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][26] ), .S0(n1899), 
        .S1(n1893), .Z(n1867) );
  MUX4D0 U1871 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][26] ), .S0(n1899), 
        .S1(n1893), .Z(n1866) );
  MUX4D0 U1872 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .S0(n1899), 
        .S1(n1893), .Z(n1868) );
  MUX4D0 U1873 ( .I0(n1872), .I1(n1870), .I2(n1871), .I3(n1869), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ) );
  MUX4D0 U1874 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][27] ), .S0(n1899), 
        .S1(n1893), .Z(n1871) );
  MUX4D0 U1875 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][27] ), .S0(n1899), 
        .S1(n1893), .Z(n1870) );
  MUX4D0 U1876 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .S0(n1899), 
        .S1(n1893), .Z(n1872) );
  MUX4D0 U1877 ( .I0(n1876), .I1(n1874), .I2(n1875), .I3(n1873), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ) );
  MUX4D0 U1878 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][28] ), .S0(n1899), 
        .S1(n1893), .Z(n1875) );
  MUX4D0 U1879 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][28] ), .S0(n1899), 
        .S1(n1893), .Z(n1874) );
  MUX4D0 U1880 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .S0(n1899), 
        .S1(n1893), .Z(n1876) );
  MUX4D0 U1881 ( .I0(n1880), .I1(n1878), .I2(n1879), .I3(n1877), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N52 ) );
  MUX4D0 U1882 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][29] ), .S0(n1900), 
        .S1(n1894), .Z(n1879) );
  MUX4D0 U1883 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][29] ), .S0(n1900), 
        .S1(n1894), .Z(n1878) );
  MUX4D0 U1884 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .S0(n1900), 
        .S1(n1894), .Z(n1880) );
  MUX4D0 U1885 ( .I0(n1884), .I1(n1882), .I2(n1883), .I3(n1881), .S0(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .S1(n1890), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N51 ) );
  MUX4D0 U1886 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][30] ), .S0(n1900), 
        .S1(n1894), .Z(n1883) );
  MUX4D0 U1887 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][30] ), .S0(n1900), 
        .S1(n1894), .Z(n1882) );
  MUX4D0 U1888 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .S0(n1900), 
        .S1(n1894), .Z(n1884) );
  MUX4D0 U1889 ( .I0(n1888), .I1(n1886), .I2(n1887), .I3(n1885), .S0(n1889), 
        .S1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .Z(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ) );
  MUX4D0 U1890 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[4][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[5][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[6][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[7][31] ), .S0(n1900), 
        .S1(n1894), .Z(n1887) );
  MUX4D0 U1891 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[8][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[9][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[10][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[11][31] ), .S0(n1900), 
        .S1(n1894), .Z(n1886) );
  MUX4D0 U1892 ( .I0(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .I2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), .I3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .S0(n1900), 
        .S1(n1894), .Z(n1888) );
  INVD1 U1893 ( .I(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .ZN(n2355) );
  INVD1 U1894 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .ZN(n2390) );
  INVD1 U1895 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .ZN(n2325) );
  INVD1 U1896 ( .I(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), .ZN(n2389) );
  INVD1 U1897 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .ZN(n2542) );
  INVD2 U1898 ( .I(n1308), .ZN(n2179) );
  INVD2 U1899 ( .I(n1307), .ZN(n2180) );
  INVD1 U1900 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n2324) );
  INVD1 U1901 ( .I(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n2301) );
  INVD1 U1902 ( .I(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), .ZN(n2432) );
  INVD1 U1903 ( .I(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), .ZN(n2428) );
  INVD1 U1904 ( .I(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(n2326) );
  INR2D1 U1905 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), .B1(n2433), .ZN(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ) );
  INR2D1 U1906 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), .B1(n2429), .ZN(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N26 ) );
  TIEH U1907 ( .Z(n2997) );
  MUX2ND0 U1908 ( .I0(n1901), .I1(n1902), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ) );
  MUX2ND0 U1909 ( .I0(n1903), .I1(n1904), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ) );
  MUX2ND0 U1910 ( .I0(n1902), .I1(n1901), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ) );
  MUX2ND0 U1911 ( .I0(n1904), .I1(n1903), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ) );
  MUX2ND0 U1912 ( .I0(n1304), .I1(n1397), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1902) );
  MUX2ND0 U1913 ( .I0(n1303), .I1(n1398), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1901) );
  MUX2ND0 U1914 ( .I0(n1397), .I1(n1303), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1904) );
  MUX2ND0 U1915 ( .I0(n1398), .I1(n1304), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1903) );
  MUX2ND0 U1916 ( .I0(n1905), .I1(n1906), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N29 ) );
  MUX2ND0 U1917 ( .I0(n1907), .I1(n1908), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N27 ) );
  MUX2ND0 U1918 ( .I0(n1906), .I1(n1905), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N25 ) );
  MUX2ND0 U1919 ( .I0(n1908), .I1(n1907), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N23 ) );
  MUX2ND0 U1920 ( .I0(n1306), .I1(n1399), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1906) );
  MUX2ND0 U1921 ( .I0(n1305), .I1(n1400), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1905) );
  MUX2ND0 U1922 ( .I0(n1399), .I1(n1305), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1908) );
  MUX2ND0 U1923 ( .I0(n1400), .I1(n1306), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), 
        .ZN(n1907) );
  MUX3ND0 U1924 ( .I0(n1909), .I1(n1910), .I2(n1911), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N84 ) );
  MUX3ND0 U1925 ( .I0(n1912), .I1(n1913), .I2(n1914), .S0(n2007), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N83 ) );
  MUX3ND0 U1926 ( .I0(n1915), .I1(n1916), .I2(n1917), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N82 ) );
  MUX3ND0 U1927 ( .I0(n1918), .I1(n1919), .I2(n1920), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N81 ) );
  MUX3ND0 U1928 ( .I0(n1921), .I1(n1922), .I2(n1923), .S0(n2007), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N80 ) );
  MUX3ND0 U1929 ( .I0(n1924), .I1(n1925), .I2(n1926), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N79 ) );
  MUX3ND0 U1930 ( .I0(n1927), .I1(n1928), .I2(n1929), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n2005), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N78 ) );
  MUX3ND0 U1931 ( .I0(n1930), .I1(n1931), .I2(n1932), .S0(n2007), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N77 ) );
  MUX3ND0 U1932 ( .I0(n1933), .I1(n1934), .I2(n1935), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N76 ) );
  MUX3ND0 U1933 ( .I0(n1936), .I1(n1937), .I2(n1938), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n2005), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N75 ) );
  MUX3ND0 U1934 ( .I0(n1939), .I1(n1940), .I2(n1941), .S0(n2007), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N74 ) );
  MUX3ND0 U1935 ( .I0(n1942), .I1(n1943), .I2(n1944), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N73 ) );
  MUX3ND0 U1936 ( .I0(n1945), .I1(n1946), .I2(n1947), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n2005), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N72 ) );
  MUX3ND0 U1937 ( .I0(n1948), .I1(n1949), .I2(n1950), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N71 ) );
  MUX3ND0 U1938 ( .I0(n1951), .I1(n1952), .I2(n1953), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N70 ) );
  MUX3ND0 U1939 ( .I0(n1954), .I1(n1955), .I2(n1956), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N69 ) );
  MUX3ND0 U1940 ( .I0(n1957), .I1(n1958), .I2(n1959), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N68 ) );
  MUX3ND0 U1941 ( .I0(n1960), .I1(n1961), .I2(n1962), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N67 ) );
  MUX3ND0 U1942 ( .I0(n1963), .I1(n1964), .I2(n1965), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N66 ) );
  MUX3ND0 U1943 ( .I0(n1966), .I1(n1967), .I2(n1968), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N65 ) );
  MUX3ND0 U1944 ( .I0(n1969), .I1(n1970), .I2(n1971), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N64 ) );
  MUX3ND0 U1945 ( .I0(n1972), .I1(n1973), .I2(n1974), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N63 ) );
  MUX3ND0 U1946 ( .I0(n1975), .I1(n1976), .I2(n1977), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N62 ) );
  MUX3ND0 U1947 ( .I0(n1978), .I1(n1979), .I2(n1980), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N61 ) );
  MUX3ND0 U1948 ( .I0(n1981), .I1(n1982), .I2(n1983), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N60 ) );
  MUX3ND0 U1949 ( .I0(n1984), .I1(n1985), .I2(n1986), .S0(n2006), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N59 ) );
  MUX3ND0 U1950 ( .I0(n1987), .I1(n1988), .I2(n1989), .S0(n2007), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N58 ) );
  MUX3ND0 U1951 ( .I0(n1990), .I1(n1991), .I2(n1992), .S0(n2006), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N57 ) );
  MUX3ND0 U1952 ( .I0(n1993), .I1(n1994), .I2(n1995), .S0(n2007), .S1(n2005), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N56 ) );
  MUX3ND0 U1953 ( .I0(n1996), .I1(n1997), .I2(n1998), .S0(n2007), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N55 ) );
  MUX3ND0 U1954 ( .I0(n1999), .I1(n2000), .I2(n2001), .S0(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .S1(n2005), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N54 ) );
  MUX3ND0 U1955 ( .I0(n2002), .I1(n2003), .I2(n2004), .S0(n2007), .S1(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N53 ) );
  MUX2ND0 U1956 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][0] ), .S(n2008), 
        .ZN(n1910) );
  MUX2ND0 U1957 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][0] ), .S(n2008), 
        .ZN(n1909) );
  MUX2ND0 U1958 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][1] ), .S(n2008), 
        .ZN(n1913) );
  MUX2ND0 U1959 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][1] ), .S(n2008), 
        .ZN(n1912) );
  MUX2ND0 U1960 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][2] ), .S(n2008), 
        .ZN(n1916) );
  MUX2ND0 U1961 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][2] ), .S(n2008), 
        .ZN(n1915) );
  MUX2ND0 U1962 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][3] ), .S(n2008), 
        .ZN(n1919) );
  MUX2ND0 U1963 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][3] ), .S(n2008), 
        .ZN(n1918) );
  MUX2ND0 U1964 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][4] ), .S(n2008), 
        .ZN(n1922) );
  MUX2ND0 U1965 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][4] ), .S(n2008), 
        .ZN(n1921) );
  MUX2ND0 U1966 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][5] ), .S(n2008), 
        .ZN(n1925) );
  MUX2ND0 U1967 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][5] ), .S(n2008), 
        .ZN(n1924) );
  MUX2ND0 U1968 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][6] ), .S(n2009), 
        .ZN(n1928) );
  MUX2ND0 U1969 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][6] ), .S(n2009), 
        .ZN(n1927) );
  MUX2ND0 U1970 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][7] ), .S(n2009), 
        .ZN(n1931) );
  MUX2ND0 U1971 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][7] ), .S(n2009), 
        .ZN(n1930) );
  MUX2ND0 U1972 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][8] ), .S(n2009), 
        .ZN(n1934) );
  MUX2ND0 U1973 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][8] ), .S(n2009), 
        .ZN(n1933) );
  MUX2ND0 U1974 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][9] ), .S(n2009), 
        .ZN(n1937) );
  MUX2ND0 U1975 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][9] ), .S(n2009), 
        .ZN(n1936) );
  MUX2ND0 U1976 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][10] ), .S(n2009), 
        .ZN(n1940) );
  MUX2ND0 U1977 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][10] ), .S(n2009), 
        .ZN(n1939) );
  MUX2ND0 U1978 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][11] ), .S(n2009), 
        .ZN(n1943) );
  MUX2ND0 U1979 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][11] ), .S(n2009), 
        .ZN(n1942) );
  MUX2ND0 U1980 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][12] ), .S(n2009), 
        .ZN(n1946) );
  MUX2ND0 U1981 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][12] ), .S(n2009), 
        .ZN(n1945) );
  MUX2ND0 U1982 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][13] ), .S(n2010), 
        .ZN(n1949) );
  MUX2ND0 U1983 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][13] ), .S(n2010), 
        .ZN(n1948) );
  MUX2ND0 U1984 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][14] ), .S(n2010), 
        .ZN(n1952) );
  MUX2ND0 U1985 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][14] ), .S(n2010), 
        .ZN(n1951) );
  MUX2ND0 U1986 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][15] ), .S(n2010), 
        .ZN(n1955) );
  MUX2ND0 U1987 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][15] ), .S(n2010), 
        .ZN(n1954) );
  MUX2ND0 U1988 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][16] ), .S(n2010), 
        .ZN(n1958) );
  MUX2ND0 U1989 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][16] ), .S(n2010), 
        .ZN(n1957) );
  MUX2ND0 U1990 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][17] ), .S(n2010), 
        .ZN(n1961) );
  MUX2ND0 U1991 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][17] ), .S(n2010), 
        .ZN(n1960) );
  MUX2ND0 U1992 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][18] ), .S(n2010), 
        .ZN(n1964) );
  MUX2ND0 U1993 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][18] ), .S(n2009), 
        .ZN(n1963) );
  MUX2ND0 U1994 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][19] ), .S(n2010), 
        .ZN(n1967) );
  MUX2ND0 U1995 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][19] ), .S(n2010), 
        .ZN(n1966) );
  MUX2ND0 U1996 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][20] ), .S(n2011), 
        .ZN(n1970) );
  MUX2ND0 U1997 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][20] ), .S(n2010), 
        .ZN(n1969) );
  MUX2ND0 U1998 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][21] ), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n1973) );
  MUX2ND0 U1999 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][21] ), .S(n2010), 
        .ZN(n1972) );
  MUX2ND0 U2000 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][22] ), .S(n2009), 
        .ZN(n1976) );
  MUX2ND0 U2001 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][22] ), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n1975) );
  MUX2ND0 U2002 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][23] ), .S(n2010), 
        .ZN(n1979) );
  MUX2ND0 U2003 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][23] ), .S(n2008), 
        .ZN(n1978) );
  MUX2ND0 U2004 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][24] ), .S(n2010), 
        .ZN(n1982) );
  MUX2ND0 U2005 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][24] ), .S(n2011), 
        .ZN(n1981) );
  MUX2ND0 U2006 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][25] ), .S(n2010), 
        .ZN(n1985) );
  MUX2ND0 U2007 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][25] ), .S(n2010), 
        .ZN(n1984) );
  MUX2ND0 U2008 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][26] ), .S(n2009), 
        .ZN(n1988) );
  MUX2ND0 U2009 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][26] ), .S(n2010), 
        .ZN(n1987) );
  MUX2ND0 U2010 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][27] ), .S(n2010), 
        .ZN(n1991) );
  MUX2ND0 U2011 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][27] ), .S(n2009), 
        .ZN(n1990) );
  MUX2ND0 U2012 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][28] ), .S(n2009), 
        .ZN(n1994) );
  MUX2ND0 U2013 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][28] ), .S(n2009), 
        .ZN(n1993) );
  MUX2ND0 U2014 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][29] ), .S(n2009), 
        .ZN(n1997) );
  MUX2ND0 U2015 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][29] ), .S(n2008), 
        .ZN(n1996) );
  MUX2ND0 U2016 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][30] ), .S(n2008), 
        .ZN(n2000) );
  MUX2ND0 U2017 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][30] ), .S(n2008), 
        .ZN(n1999) );
  MUX2ND0 U2018 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[2][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[3][31] ), .S(n2008), 
        .ZN(n2003) );
  MUX2ND0 U2019 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/Storage[1][31] ), .S(n2008), 
        .ZN(n2002) );
  MUX3ND0 U2020 ( .I0(n2012), .I1(n2013), .I2(n2014), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N84 ) );
  MUX3ND0 U2021 ( .I0(n2015), .I1(n2016), .I2(n2017), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N83 ) );
  MUX3ND0 U2022 ( .I0(n2018), .I1(n2019), .I2(n2020), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N82 ) );
  MUX3ND0 U2023 ( .I0(n2021), .I1(n2022), .I2(n2023), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N81 ) );
  MUX3ND0 U2024 ( .I0(n2024), .I1(n2025), .I2(n2026), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N80 ) );
  MUX3ND0 U2025 ( .I0(n2027), .I1(n2028), .I2(n2029), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N79 ) );
  MUX3ND0 U2026 ( .I0(n2030), .I1(n2031), .I2(n2032), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N78 ) );
  MUX3ND0 U2027 ( .I0(n2033), .I1(n2034), .I2(n2035), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N77 ) );
  MUX3ND0 U2028 ( .I0(n2036), .I1(n2037), .I2(n2038), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N76 ) );
  MUX3ND0 U2029 ( .I0(n2039), .I1(n2040), .I2(n2041), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N75 ) );
  MUX3ND0 U2030 ( .I0(n2042), .I1(n2043), .I2(n2044), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N74 ) );
  MUX3ND0 U2031 ( .I0(n2045), .I1(n2046), .I2(n2047), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N73 ) );
  MUX3ND0 U2032 ( .I0(n2048), .I1(n2049), .I2(n2050), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N72 ) );
  MUX3ND0 U2033 ( .I0(n2051), .I1(n2052), .I2(n2053), .S0(n2110), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N71 ) );
  MUX3ND0 U2034 ( .I0(n2054), .I1(n2055), .I2(n2056), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n2108), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N70 ) );
  MUX3ND0 U2035 ( .I0(n2057), .I1(n2058), .I2(n2059), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n2108), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N69 ) );
  MUX3ND0 U2036 ( .I0(n2060), .I1(n2061), .I2(n2062), .S0(n2110), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N68 ) );
  MUX3ND0 U2037 ( .I0(n2063), .I1(n2064), .I2(n2065), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N67 ) );
  MUX3ND0 U2038 ( .I0(n2066), .I1(n2067), .I2(n2068), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n2108), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N66 ) );
  MUX3ND0 U2039 ( .I0(n2069), .I1(n2070), .I2(n2071), .S0(n2110), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N65 ) );
  MUX3ND0 U2040 ( .I0(n2072), .I1(n2073), .I2(n2074), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N64 ) );
  MUX3ND0 U2041 ( .I0(n2075), .I1(n2076), .I2(n2077), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(n2108), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N63 ) );
  MUX3ND0 U2042 ( .I0(n2078), .I1(n2079), .I2(n2080), .S0(n2110), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N62 ) );
  MUX3ND0 U2043 ( .I0(n2081), .I1(n2082), .I2(n2083), .S0(n2109), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N61 ) );
  MUX3ND0 U2044 ( .I0(n2084), .I1(n2085), .I2(n2086), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N60 ) );
  MUX3ND0 U2045 ( .I0(n2087), .I1(n2088), .I2(n2089), .S0(n2110), .S1(n2108), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N59 ) );
  MUX3ND0 U2046 ( .I0(n2090), .I1(n2091), .I2(n2092), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N58 ) );
  MUX3ND0 U2047 ( .I0(n2093), .I1(n2094), .I2(n2095), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N57 ) );
  MUX3ND0 U2048 ( .I0(n2096), .I1(n2097), .I2(n2098), .S0(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N56 ) );
  MUX3ND0 U2049 ( .I0(n2099), .I1(n2100), .I2(n2101), .S0(n2110), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N55 ) );
  MUX3ND0 U2050 ( .I0(n2102), .I1(n2103), .I2(n2104), .S0(n2110), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N54 ) );
  MUX3ND0 U2051 ( .I0(n2105), .I1(n2106), .I2(n2107), .S0(n2109), .S1(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N53 ) );
  MUX2ND0 U2052 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][0] ), .S(n2111), 
        .ZN(n2013) );
  MUX2ND0 U2053 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][0] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][0] ), .S(n2111), 
        .ZN(n2012) );
  MUX2ND0 U2054 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][1] ), .S(n2111), 
        .ZN(n2016) );
  MUX2ND0 U2055 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][1] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][1] ), .S(n2111), 
        .ZN(n2015) );
  MUX2ND0 U2056 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][2] ), .S(n2111), 
        .ZN(n2019) );
  MUX2ND0 U2057 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][2] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][2] ), .S(n2111), 
        .ZN(n2018) );
  MUX2ND0 U2058 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][3] ), .S(n2111), 
        .ZN(n2022) );
  MUX2ND0 U2059 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][3] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][3] ), .S(n2111), 
        .ZN(n2021) );
  MUX2ND0 U2060 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][4] ), .S(n2111), 
        .ZN(n2025) );
  MUX2ND0 U2061 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][4] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][4] ), .S(n2111), 
        .ZN(n2024) );
  MUX2ND0 U2062 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][5] ), .S(n2111), 
        .ZN(n2028) );
  MUX2ND0 U2063 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][5] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][5] ), .S(n2111), 
        .ZN(n2027) );
  MUX2ND0 U2064 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][6] ), .S(n2112), 
        .ZN(n2031) );
  MUX2ND0 U2065 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][6] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][6] ), .S(n2112), 
        .ZN(n2030) );
  MUX2ND0 U2066 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][7] ), .S(n2112), 
        .ZN(n2034) );
  MUX2ND0 U2067 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][7] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][7] ), .S(n2112), 
        .ZN(n2033) );
  MUX2ND0 U2068 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][8] ), .S(n2112), 
        .ZN(n2037) );
  MUX2ND0 U2069 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][8] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][8] ), .S(n2112), 
        .ZN(n2036) );
  MUX2ND0 U2070 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][9] ), .S(n2112), 
        .ZN(n2040) );
  MUX2ND0 U2071 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][9] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][9] ), .S(n2112), 
        .ZN(n2039) );
  MUX2ND0 U2072 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][10] ), .S(n2112), 
        .ZN(n2043) );
  MUX2ND0 U2073 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][10] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][10] ), .S(n2112), 
        .ZN(n2042) );
  MUX2ND0 U2074 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][11] ), .S(n2112), 
        .ZN(n2046) );
  MUX2ND0 U2075 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][11] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][11] ), .S(n2112), 
        .ZN(n2045) );
  MUX2ND0 U2076 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][12] ), .S(n2112), 
        .ZN(n2049) );
  MUX2ND0 U2077 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][12] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][12] ), .S(n2112), 
        .ZN(n2048) );
  MUX2ND0 U2078 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][13] ), .S(n2113), 
        .ZN(n2052) );
  MUX2ND0 U2079 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][13] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][13] ), .S(n2113), 
        .ZN(n2051) );
  MUX2ND0 U2080 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][14] ), .S(n2113), 
        .ZN(n2055) );
  MUX2ND0 U2081 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][14] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][14] ), .S(n2113), 
        .ZN(n2054) );
  MUX2ND0 U2082 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][15] ), .S(n2113), 
        .ZN(n2058) );
  MUX2ND0 U2083 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][15] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][15] ), .S(n2113), 
        .ZN(n2057) );
  MUX2ND0 U2084 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][16] ), .S(n2113), 
        .ZN(n2061) );
  MUX2ND0 U2085 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][16] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][16] ), .S(n2113), 
        .ZN(n2060) );
  MUX2ND0 U2086 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][17] ), .S(n2113), 
        .ZN(n2064) );
  MUX2ND0 U2087 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][17] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][17] ), .S(n2113), 
        .ZN(n2063) );
  MUX2ND0 U2088 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][18] ), .S(n2113), 
        .ZN(n2067) );
  MUX2ND0 U2089 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][18] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][18] ), .S(n2112), 
        .ZN(n2066) );
  MUX2ND0 U2090 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][19] ), .S(n2113), 
        .ZN(n2070) );
  MUX2ND0 U2091 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][19] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][19] ), .S(n2113), 
        .ZN(n2069) );
  MUX2ND0 U2092 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][20] ), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n2073) );
  MUX2ND0 U2093 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][20] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][20] ), .S(n2113), 
        .ZN(n2072) );
  MUX2ND0 U2094 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][21] ), .S(n2114), 
        .ZN(n2076) );
  MUX2ND0 U2095 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][21] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][21] ), .S(n2113), 
        .ZN(n2075) );
  MUX2ND0 U2096 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][22] ), .S(n2112), 
        .ZN(n2079) );
  MUX2ND0 U2097 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][22] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][22] ), .S(n2114), 
        .ZN(n2078) );
  MUX2ND0 U2098 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][23] ), .S(n2113), 
        .ZN(n2082) );
  MUX2ND0 U2099 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][23] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][23] ), .S(n2111), 
        .ZN(n2081) );
  MUX2ND0 U2100 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][24] ), .S(n2113), 
        .ZN(n2085) );
  MUX2ND0 U2101 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][24] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][24] ), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n2084) );
  MUX2ND0 U2102 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][25] ), .S(n2113), 
        .ZN(n2088) );
  MUX2ND0 U2103 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][25] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][25] ), .S(n2113), 
        .ZN(n2087) );
  MUX2ND0 U2104 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][26] ), .S(n2112), 
        .ZN(n2091) );
  MUX2ND0 U2105 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][26] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][26] ), .S(n2113), 
        .ZN(n2090) );
  MUX2ND0 U2106 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][27] ), .S(n2113), 
        .ZN(n2094) );
  MUX2ND0 U2107 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][27] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][27] ), .S(n2112), 
        .ZN(n2093) );
  MUX2ND0 U2108 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][28] ), .S(n2112), 
        .ZN(n2097) );
  MUX2ND0 U2109 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][28] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][28] ), .S(n2112), 
        .ZN(n2096) );
  MUX2ND0 U2110 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][29] ), .S(n2112), 
        .ZN(n2100) );
  MUX2ND0 U2111 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][29] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][29] ), .S(n2111), 
        .ZN(n2099) );
  MUX2ND0 U2112 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][30] ), .S(n2111), 
        .ZN(n2103) );
  MUX2ND0 U2113 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][30] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][30] ), .S(n2111), 
        .ZN(n2102) );
  MUX2ND0 U2114 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[2][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[3][31] ), .S(n2111), 
        .ZN(n2106) );
  MUX2ND0 U2115 ( .I0(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[0][31] ), 
        .I1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/Storage[1][31] ), .S(n2111), 
        .ZN(n2105) );
  CKND0 U2116 ( .CLK(n3061), .CN(n2115) );
  CKND0 U2117 ( .CLK(n3060), .CN(n2116) );
  CKND0 U2118 ( .CLK(n3059), .CN(n2117) );
  CKND0 U2119 ( .CLK(n3058), .CN(n2118) );
  CKND0 U2120 ( .CLK(n3057), .CN(n2119) );
  CKND0 U2121 ( .CLK(n3056), .CN(n2120) );
  CKND0 U2122 ( .CLK(n3055), .CN(n2121) );
  CKND0 U2123 ( .CLK(n3054), .CN(n2122) );
  CKND0 U2124 ( .CLK(n3053), .CN(n2123) );
  CKND0 U2125 ( .CLK(n3052), .CN(n2124) );
  CKND0 U2126 ( .CLK(n3051), .CN(n2125) );
  CKND0 U2127 ( .CLK(n3050), .CN(n2126) );
  CKND0 U2128 ( .CLK(n3049), .CN(n2127) );
  CKND0 U2129 ( .CLK(n3048), .CN(n2128) );
  CKND0 U2130 ( .CLK(n3047), .CN(n2129) );
  CKND0 U2131 ( .CLK(n3046), .CN(n2130) );
  CKND0 U2132 ( .CLK(n3045), .CN(n2131) );
  CKND0 U2133 ( .CLK(n3044), .CN(n2132) );
  CKND0 U2134 ( .CLK(n3043), .CN(n2133) );
  CKND0 U2135 ( .CLK(n3042), .CN(n2134) );
  CKND0 U2136 ( .CLK(n3041), .CN(n2135) );
  CKND0 U2137 ( .CLK(n3040), .CN(n2136) );
  CKND0 U2138 ( .CLK(n3039), .CN(n2137) );
  CKND0 U2139 ( .CLK(n3038), .CN(n2138) );
  CKND0 U2140 ( .CLK(n3037), .CN(n2139) );
  CKND0 U2141 ( .CLK(n3036), .CN(n2140) );
  CKND0 U2142 ( .CLK(n3035), .CN(n2141) );
  CKND0 U2143 ( .CLK(n3034), .CN(n2142) );
  CKND0 U2144 ( .CLK(n3033), .CN(n2143) );
  CKND0 U2145 ( .CLK(n3032), .CN(n2144) );
  CKND0 U2146 ( .CLK(n3031), .CN(n2145) );
  CKND0 U2147 ( .CLK(n3030), .CN(n2146) );
  CKND0 U2148 ( .CLK(n3029), .CN(n2147) );
  CKND0 U2149 ( .CLK(n3028), .CN(n2148) );
  CKND0 U2150 ( .CLK(n3027), .CN(n2149) );
  CKND0 U2151 ( .CLK(n3026), .CN(n2150) );
  CKND0 U2152 ( .CLK(n3025), .CN(n2151) );
  CKND0 U2153 ( .CLK(n3024), .CN(n2152) );
  CKND0 U2154 ( .CLK(n3023), .CN(n2153) );
  CKND0 U2155 ( .CLK(n3022), .CN(n2154) );
  CKND0 U2156 ( .CLK(n3021), .CN(n2155) );
  CKND0 U2157 ( .CLK(n3020), .CN(n2156) );
  CKND0 U2158 ( .CLK(n3019), .CN(n2157) );
  CKND0 U2159 ( .CLK(n3018), .CN(n2158) );
  CKND0 U2160 ( .CLK(n3017), .CN(n2159) );
  CKND0 U2161 ( .CLK(n3016), .CN(n2160) );
  CKND0 U2162 ( .CLK(n3015), .CN(n2161) );
  CKND0 U2163 ( .CLK(n3014), .CN(n2162) );
  CKND0 U2164 ( .CLK(n3013), .CN(n2163) );
  CKND0 U2165 ( .CLK(n3012), .CN(n2164) );
  CKND0 U2166 ( .CLK(n3011), .CN(n2165) );
  CKND0 U2167 ( .CLK(n3010), .CN(n2166) );
  CKND0 U2168 ( .CLK(n3009), .CN(n2167) );
  CKND0 U2169 ( .CLK(n3008), .CN(n2168) );
  CKND0 U2170 ( .CLK(n3007), .CN(n2169) );
  CKND0 U2171 ( .CLK(n3006), .CN(n2170) );
  CKND0 U2172 ( .CLK(n3005), .CN(n2171) );
  CKND0 U2173 ( .CLK(n3004), .CN(n2172) );
  CKND0 U2174 ( .CLK(n3003), .CN(n2173) );
  CKND0 U2175 ( .CLK(n3002), .CN(n2174) );
  CKND0 U2176 ( .CLK(n3001), .CN(n2175) );
  CKND0 U2177 ( .CLK(n3000), .CN(n2176) );
  CKND0 U2178 ( .CLK(n2999), .CN(n2177) );
  CKND0 U2179 ( .CLK(n2998), .CN(n2178) );
  OR2D1 U2180 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N2 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N3 ), .Z(n2429) );
  MUX2ND0 U2181 ( .I0(n2430), .I1(n2429), .S(\SerDes_U1/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(\SerDes_U1/Ser_U1/SerEnc_Tx1/N28 ) );
  OR2D1 U2182 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N2 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N3 ), .Z(n2433) );
  MUX2ND0 U2183 ( .I0(n2434), .I1(n2433), .S(\SerDes_U2/Ser_U1/SerEnc_Tx1/N4 ), 
        .ZN(\SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ) );
  OAI31D0 U2184 ( .A1(n2435), .A2(Reset), .A3(n2436), .B(n2437), .ZN(n1246) );
  OAI21D0 U2185 ( .A1(n2438), .A2(Reset), .B(n2967), .ZN(n2437) );
  AOI21D0 U2186 ( .A1(n2971), .A2(n2972), .B(n2439), .ZN(n2438) );
  NR3D0 U2187 ( .A1(n1302), .A2(n2350), .A3(n2440), .ZN(n2436) );
  MUX2ND0 U2188 ( .I0(n2441), .I1(n1030), .S(n2442), .ZN(n1245) );
  AOI211D0 U2189 ( .A1(n2443), .A2(n2444), .B(n2445), .C(n2439), .ZN(n2441) );
  OAI22D0 U2190 ( .A1(n2446), .A2(n2447), .B1(n2448), .B2(n2446), .ZN(n2445)
         );
  MUX2D0 U2191 ( .I0(n2448), .I1(n2449), .S(n2971), .Z(n2443) );
  ND4D0 U2192 ( .A1(n2450), .A2(n2451), .A3(n2452), .A4(n2453), .ZN(n2448) );
  NR3D0 U2193 ( .A1(n2454), .A2(n2455), .A3(n2456), .ZN(n2453) );
  XNR2D0 U2194 ( .A1(n2457), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .ZN(n2456) );
  XNR2D0 U2195 ( .A1(n2458), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), 
        .ZN(n2454) );
  OAI33D0 U2196 ( .A1(n2459), .A2(n2460), .A3(n2461), .B1(n2462), .B2(n2463), 
        .B3(n2464), .ZN(n1244) );
  XNR2D0 U2197 ( .A1(n2966), .A2(n2356), .ZN(n2461) );
  XNR2D0 U2198 ( .A1(n2965), .A2(n2355), .ZN(n2460) );
  ND3D0 U2199 ( .A1(n2465), .A2(n2466), .A3(n2467), .ZN(n2459) );
  XNR2D0 U2200 ( .A1(n2353), .A2(n1388), .ZN(n2467) );
  XNR2D0 U2201 ( .A1(n2354), .A2(n1387), .ZN(n2465) );
  MUX2ND0 U2202 ( .I0(n2468), .I1(n1024), .S(n2442), .ZN(n1243) );
  AOI32D0 U2203 ( .A1(n2444), .A2(n2469), .A3(n2470), .B1(n2971), .B2(n2471), 
        .ZN(n2468) );
  OAI21D0 U2204 ( .A1(n2472), .A2(n1300), .B(n1310), .ZN(n2471) );
  NR4D0 U2205 ( .A1(n2470), .A2(n2473), .A3(n2474), .A4(n2475), .ZN(n2472) );
  XNR2D0 U2206 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n2476), 
        .ZN(n2475) );
  XNR2D0 U2207 ( .A1(n2477), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), 
        .ZN(n2474) );
  XNR2D0 U2208 ( .A1(n2478), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n2473) );
  OAI31D0 U2209 ( .A1(n2479), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), 
        .A3(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .B(n2480), .ZN(n2469) );
  MUX2ND0 U2210 ( .I0(n2481), .I1(n2482), .S(n2355), .ZN(n2480) );
  OAI32D0 U2211 ( .A1(n2483), .A2(n2356), .A3(n2450), .B1(n2451), .B2(n2484), 
        .ZN(n2482) );
  OAI32D0 U2212 ( .A1(n2483), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .A3(n2451), .B1(n2450), .B2(n2484), .ZN(n2481) );
  CKND2D0 U2213 ( .A1(n2485), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .ZN(n2484) );
  XNR2D0 U2214 ( .A1(n2457), .A2(n2356), .ZN(n2485) );
  MUX2ND0 U2215 ( .I0(n2486), .I1(n2487), .S(n2355), .ZN(n2479) );
  NR2D0 U2216 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), .A2(n2450), 
        .ZN(n2487) );
  NR2D0 U2217 ( .A1(n2356), .A2(n2451), .ZN(n2486) );
  OAI33D0 U2218 ( .A1(n2488), .A2(n2489), .A3(n2490), .B1(n2491), .B2(n2439), 
        .B3(n2464), .ZN(n1242) );
  XNR2D0 U2219 ( .A1(n2963), .A2(n2457), .ZN(n2490) );
  XNR2D0 U2220 ( .A1(n2964), .A2(n2458), .ZN(n2489) );
  ND3D0 U2221 ( .A1(n2492), .A2(n2493), .A3(n2494), .ZN(n2488) );
  XNR2D0 U2222 ( .A1(n2495), .A2(n1386), .ZN(n2494) );
  XNR2D0 U2223 ( .A1(n2496), .A2(n1385), .ZN(n2492) );
  MUX2ND0 U2224 ( .I0(n2497), .I1(n1018), .S(n2442), .ZN(n1241) );
  OA211D0 U2225 ( .A1(n2970), .A2(n1301), .B(n2498), .C(n2499), .Z(n2442) );
  AOI22D0 U2226 ( .A1(n2972), .A2(n2500), .B1(n2439), .B2(n2501), .ZN(n2499)
         );
  AO31D0 U2227 ( .A1(n2181), .A2(\SerDes_U2/Ser_U1/SerEnc_Tx1/HalfParClkr ), 
        .A3(InParValidB), .B(n1301), .Z(n2500) );
  AOI21D0 U2228 ( .A1(n2971), .A2(n2502), .B(n2463), .ZN(n2497) );
  IOA22D0 U2229 ( .B1(n1300), .B2(n2449), .A1(n2447), .A2(n2972), .ZN(n2502)
         );
  ND4D0 U2230 ( .A1(n2503), .A2(n2470), .A3(n2504), .A4(n2478), .ZN(n2447) );
  CKND2D0 U2231 ( .A1(n2451), .A2(n2450), .ZN(n2478) );
  CKND2D0 U2232 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n2354), 
        .ZN(n2450) );
  CKND2D0 U2233 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N45 ), .A2(n2496), 
        .ZN(n2451) );
  XNR2D0 U2234 ( .A1(n2505), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .ZN(n2504) );
  CKND2D0 U2235 ( .A1(n2506), .A2(n2483), .ZN(n2505) );
  MUX2ND0 U2236 ( .I0(n2496), .I1(n2507), .S(n2457), .ZN(n2506) );
  NR2D0 U2237 ( .A1(n2496), .A2(n2458), .ZN(n2507) );
  XNR3D0 U2238 ( .A1(n2458), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), 
        .A3(n2355), .ZN(n2503) );
  IND4D0 U2239 ( .A1(n2470), .B1(n2508), .B2(n2509), .B3(n2510), .ZN(n2449) );
  XNR2D0 U2240 ( .A1(n2511), .A2(n2354), .ZN(n2510) );
  XNR2D0 U2241 ( .A1(n2356), .A2(n2512), .ZN(n2509) );
  XNR2D0 U2242 ( .A1(n2513), .A2(n2355), .ZN(n2508) );
  INR2D0 U2243 ( .A1(n2452), .B1(n2455), .ZN(n2470) );
  NR2D0 U2244 ( .A1(n2353), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n2455) );
  CKND2D0 U2245 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .A2(n2353), 
        .ZN(n2452) );
  MUX2D0 U2246 ( .I0(n2963), .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), 
        .S(n2493), .Z(n1240) );
  MUX2ND0 U2247 ( .I0(n1385), .I1(n2496), .S(n2493), .ZN(n1239) );
  MUX2ND0 U2248 ( .I0(n1386), .I1(n2495), .S(n2493), .ZN(n1238) );
  MUX2D0 U2249 ( .I0(n2964), .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .S(n2493), .Z(n1237) );
  OA21D0 U2250 ( .A1(n2439), .A2(n2464), .B(n2501), .Z(n2493) );
  CKND0 U2251 ( .CLK(n2498), .CN(n2464) );
  MUX2D0 U2252 ( .I0(n2966), .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N47 ), 
        .S(n2466), .Z(n1236) );
  MUX2ND0 U2253 ( .I0(n1387), .I1(n2354), .S(n2466), .ZN(n1235) );
  MUX2ND0 U2254 ( .I0(n1388), .I1(n2353), .S(n2466), .ZN(n1234) );
  MUX2D0 U2255 ( .I0(n2965), .I1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), 
        .S(n2466), .Z(n1233) );
  AN3D0 U2256 ( .A1(n2181), .A2(InParValidB), .A3(n2514), .Z(n2466) );
  AOI21D0 U2257 ( .A1(n2498), .A2(n2435), .B(n2350), .ZN(n2514) );
  INR2D0 U2258 ( .A1(n2446), .B1(n2444), .ZN(n2498) );
  ND3D0 U2259 ( .A1(n2972), .A2(n1300), .A3(n2971), .ZN(n2446) );
  OAI31D0 U2260 ( .A1(n2515), .A2(Reset), .A3(n2501), .B(n2516), .ZN(n1232) );
  OAI21D0 U2261 ( .A1(n2517), .A2(Reset), .B(n1302), .ZN(n2516) );
  AOI21D0 U2262 ( .A1(n2444), .A2(n1301), .B(n2439), .ZN(n2517) );
  NR2D0 U2263 ( .A1(n1300), .A2(n2972), .ZN(n2444) );
  NR2D0 U2264 ( .A1(n2440), .A2(n2967), .ZN(n2501) );
  CKND0 U2265 ( .CLK(InParValidB), .CN(n2440) );
  OAI31D0 U2266 ( .A1(n2518), .A2(Reset), .A3(n2519), .B(n2520), .ZN(n1231) );
  OAI21D0 U2267 ( .A1(Reset), .A2(n2521), .B(n1299), .ZN(n2520) );
  OAI22D0 U2268 ( .A1(n2522), .A2(n1401), .B1(n2523), .B2(n2524), .ZN(n1230)
         );
  OAI31D0 U2269 ( .A1(n1299), .A2(n2352), .A3(n2525), .B(n2199), .ZN(n2524) );
  AOI21D0 U2270 ( .A1(n2518), .A2(n2526), .B(Reset), .ZN(n2522) );
  MUX2ND0 U2271 ( .I0(n2527), .I1(n1016), .S(n2528), .ZN(n1229) );
  NR2D0 U2272 ( .A1(n2529), .A2(n2530), .ZN(n2527) );
  MUX2ND0 U2273 ( .I0(n2531), .I1(n2532), .S(n2533), .ZN(n2530) );
  OAI21D0 U2274 ( .A1(n2534), .A2(n2535), .B(n2536), .ZN(n2532) );
  CKND0 U2275 ( .CLK(n2537), .CN(n2534) );
  OAI21D0 U2276 ( .A1(n2538), .A2(n2539), .B(n2540), .ZN(n2531) );
  MUX2ND0 U2277 ( .I0(n2535), .I1(n2541), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n2539) );
  OA211D0 U2278 ( .A1(n2005), .A2(n2542), .B(n2543), .C(n2544), .Z(n2535) );
  NR2D0 U2279 ( .A1(n2545), .A2(n2546), .ZN(n2544) );
  NR2D0 U2280 ( .A1(n2547), .A2(n2543), .ZN(n2538) );
  MUX2ND0 U2281 ( .I0(n2548), .I1(n2549), .S(n2550), .ZN(n1228) );
  IND4D0 U2282 ( .A1(n2551), .B1(n2552), .B2(n2553), .B3(n2554), .ZN(n2549) );
  XNR2D0 U2283 ( .A1(n2324), .A2(n1390), .ZN(n2554) );
  XNR2D0 U2284 ( .A1(n2325), .A2(n1391), .ZN(n2553) );
  XNR2D0 U2285 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n2961), 
        .ZN(n2552) );
  MUX2ND0 U2286 ( .I0(n2555), .I1(n1011), .S(n2528), .ZN(n1227) );
  AOI21D0 U2287 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A2(
        n2556), .B(n2536), .ZN(n2555) );
  OAI31D0 U2288 ( .A1(n2557), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A3(n2546), .B(
        n2558), .ZN(n2556) );
  OAI31D0 U2289 ( .A1(n2559), .A2(n2560), .A3(n2561), .B(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n2558) );
  XNR2D0 U2290 ( .A1(n2562), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .ZN(n2559) );
  MUX2ND0 U2291 ( .I0(n2563), .I1(n2564), .S(n2325), .ZN(n2557) );
  NR2D0 U2292 ( .A1(n2565), .A2(n2566), .ZN(n2564) );
  XNR2D0 U2293 ( .A1(n2542), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), 
        .ZN(n2566) );
  OAI22D0 U2294 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n2567), 
        .B1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .B2(n2543), .ZN(
        n2563) );
  OAI33D0 U2295 ( .A1(n2568), .A2(n2569), .A3(n2570), .B1(n1311), .B2(n2529), 
        .B3(n2550), .ZN(n1226) );
  XNR2D0 U2296 ( .A1(n2959), .A2(n2542), .ZN(n2570) );
  XNR2D0 U2297 ( .A1(n2960), .A2(n2565), .ZN(n2569) );
  OAI211D0 U2298 ( .A1(n2529), .A2(n2571), .B(n2519), .C(n2572), .ZN(n2568) );
  XNR2D0 U2299 ( .A1(n2573), .A2(n1389), .ZN(n2572) );
  MUX2D0 U2300 ( .I0(n2959), .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .S(n2574), .Z(n1225) );
  MUX2ND0 U2301 ( .I0(n1389), .I1(n2573), .S(n2574), .ZN(n1224) );
  MUX2D0 U2302 ( .I0(n2960), .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), 
        .S(n2574), .Z(n1223) );
  OA21D0 U2303 ( .A1(n2529), .A2(n2571), .B(n2519), .Z(n2574) );
  MUX2ND0 U2304 ( .I0(n2575), .I1(n1006), .S(n2528), .ZN(n1222) );
  AOI211D0 U2305 ( .A1(n2533), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .B(n2571), .C(n2576), .ZN(n2528) );
  AO22D0 U2306 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        n2577), .B1(n2519), .B2(n2529), .Z(n2576) );
  NR2D0 U2307 ( .A1(n2525), .A2(n2962), .ZN(n2519) );
  CKND0 U2308 ( .CLK(InParValidA), .CN(n2525) );
  CKND2D0 U2309 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .A2(
        n2551), .ZN(n2577) );
  OAI221D0 U2310 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        n2578), .B1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .B2(
        n2537), .C(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(
        n2575) );
  OAI211D0 U2311 ( .A1(n2579), .A2(n2580), .B(n2545), .C(n2560), .ZN(n2537) );
  CKND0 U2312 ( .CLK(n2546), .CN(n2560) );
  MUX2ND0 U2313 ( .I0(n2581), .I1(n2567), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(n2580) );
  CKND2D0 U2314 ( .A1(n2582), .A2(n2567), .ZN(n2581) );
  NR2D0 U2315 ( .A1(n2565), .A2(n2543), .ZN(n2579) );
  OA211D0 U2316 ( .A1(n2543), .A2(n2547), .B(n2541), .C(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .Z(n2578) );
  AN3D0 U2317 ( .A1(n2561), .A2(n2546), .A3(n2583), .Z(n2541) );
  MUX2ND0 U2318 ( .I0(n2584), .I1(n2585), .S(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .ZN(n2583) );
  NR2D0 U2319 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .A2(n2547), 
        .ZN(n2585) );
  OAI21D0 U2320 ( .A1(n2542), .A2(n2324), .B(n2586), .ZN(n2584) );
  XNR2D0 U2321 ( .A1(n2573), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(n2546) );
  XNR2D0 U2322 ( .A1(n2545), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n2561) );
  XNR2D0 U2323 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n2325), 
        .ZN(n2545) );
  CKND2D0 U2324 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n2542), 
        .ZN(n2543) );
  MUX2D0 U2325 ( .I0(n2961), .I1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), 
        .S(n2587), .Z(n1221) );
  MUX2ND0 U2326 ( .I0(n1390), .I1(n2324), .S(n2587), .ZN(n1220) );
  MUX2ND0 U2327 ( .I0(n1391), .I1(n2325), .S(n2587), .ZN(n1219) );
  INR2D0 U2328 ( .A1(n2550), .B1(n2551), .ZN(n2587) );
  ND3D0 U2329 ( .A1(InParValidA), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/HalfParClkr ), .A3(n1296), .ZN(n2551) );
  IND2D0 U2330 ( .A1(n2571), .B1(n2523), .ZN(n2550) );
  MUX2ND0 U2331 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .I1(
        n2526), .S(n2533), .ZN(n2571) );
  CKND0 U2332 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .CN(
        n2533) );
  AO222D0 U2333 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ), .A2(
        n2588), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ), .B2(n2589), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .C2(n2590), 
        .Z(n1216) );
  AO222D0 U2334 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ), .A2(
        n2588), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ), .B2(n2589), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .C2(n2590), 
        .Z(n1215) );
  AO222D0 U2335 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ), .A2(
        n2588), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ), .B2(n2589), .C1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .C2(n2590), 
        .Z(n1214) );
  CKND0 U2336 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CN(
        n2590) );
  AN2D0 U2337 ( .A1(n2591), .A2(n2592), .Z(n2589) );
  AN3D0 U2338 ( .A1(n2593), .A2(n2594), .A3(n2595), .Z(n2588) );
  CKXOR2D0 U2339 ( .A1(\SerDes_U1/Tx_SerClk ), .A2(n2596), .Z(n1213) );
  AO222D0 U2340 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ), .A2(
        n2597), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ), .B2(n2598), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .C2(n2599), 
        .Z(n1211) );
  XNR2D0 U2341 ( .A1(n2600), .A2(\SerDes_U1/Des_U1/SerialClk ), .ZN(n1210) );
  MUX2ND0 U2342 ( .I0(n1352), .I1(n1004), .S(n2299), .ZN(n1209) );
  MUX2ND0 U2343 ( .I0(n1351), .I1(n970), .S(n2299), .ZN(n1208) );
  MUX2ND0 U2344 ( .I0(n1350), .I1(n968), .S(n2299), .ZN(n1207) );
  MUX2ND0 U2345 ( .I0(n1349), .I1(n966), .S(n2299), .ZN(n1206) );
  MUX2ND0 U2346 ( .I0(n1348), .I1(n964), .S(n2299), .ZN(n1205) );
  MUX2ND0 U2347 ( .I0(n1347), .I1(n962), .S(n2299), .ZN(n1204) );
  MUX2ND0 U2348 ( .I0(n1346), .I1(n960), .S(n2299), .ZN(n1203) );
  MUX2ND0 U2349 ( .I0(n1345), .I1(n958), .S(n2299), .ZN(n1202) );
  MUX2ND0 U2350 ( .I0(n1344), .I1(n956), .S(n2299), .ZN(n1201) );
  MUX2ND0 U2351 ( .I0(n1343), .I1(n954), .S(n2299), .ZN(n1200) );
  MUX2ND0 U2352 ( .I0(n1342), .I1(n952), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1199) );
  MUX2ND0 U2353 ( .I0(n1341), .I1(n950), .S(n2299), .ZN(n1198) );
  MUX2ND0 U2354 ( .I0(n1340), .I1(n948), .S(n2299), .ZN(n1197) );
  MUX2ND0 U2355 ( .I0(n1339), .I1(n946), .S(n2299), .ZN(n1196) );
  MUX2ND0 U2356 ( .I0(n1338), .I1(n944), .S(n2299), .ZN(n1195) );
  MUX2ND0 U2357 ( .I0(n1337), .I1(n942), .S(n2299), .ZN(n1194) );
  MUX2ND0 U2358 ( .I0(n1336), .I1(n940), .S(n2299), .ZN(n1193) );
  MUX2ND0 U2359 ( .I0(n1335), .I1(n938), .S(n2299), .ZN(n1192) );
  MUX2ND0 U2360 ( .I0(n1334), .I1(n936), .S(n2299), .ZN(n1191) );
  MUX2ND0 U2361 ( .I0(n1333), .I1(n934), .S(n2299), .ZN(n1190) );
  MUX2ND0 U2362 ( .I0(n1332), .I1(n932), .S(n2299), .ZN(n1189) );
  MUX2ND0 U2363 ( .I0(n1331), .I1(n930), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1188) );
  MUX2ND0 U2364 ( .I0(n1330), .I1(n928), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1187) );
  MUX2ND0 U2365 ( .I0(n1329), .I1(n926), .S(n2299), .ZN(n1186) );
  MUX2ND0 U2366 ( .I0(n1328), .I1(n924), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1185) );
  MUX2ND0 U2367 ( .I0(n1327), .I1(n922), .S(n2299), .ZN(n1184) );
  MUX2ND0 U2368 ( .I0(n1326), .I1(n920), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1183) );
  MUX2ND0 U2369 ( .I0(n1325), .I1(n918), .S(n2299), .ZN(n1182) );
  MUX2ND0 U2370 ( .I0(n1324), .I1(n916), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1181) );
  MUX2ND0 U2371 ( .I0(n1323), .I1(n914), .S(n2299), .ZN(n1180) );
  MUX2ND0 U2372 ( .I0(n1322), .I1(n912), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1179) );
  MUX2ND0 U2373 ( .I0(n1321), .I1(n910), .S(\SerDes_U1/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1178) );
  MUX2ND0 U2374 ( .I0(n908), .I1(n1321), .S(n2180), .ZN(n1177) );
  MUX2ND0 U2375 ( .I0(n907), .I1(n1322), .S(n2180), .ZN(n1176) );
  MUX2ND0 U2376 ( .I0(n906), .I1(n1323), .S(n2180), .ZN(n1175) );
  MUX2ND0 U2377 ( .I0(n905), .I1(n1324), .S(n2180), .ZN(n1174) );
  MUX2ND0 U2378 ( .I0(n904), .I1(n1325), .S(n2180), .ZN(n1173) );
  MUX2ND0 U2379 ( .I0(n903), .I1(n1326), .S(n2180), .ZN(n1172) );
  MUX2ND0 U2380 ( .I0(n902), .I1(n1327), .S(n2180), .ZN(n1171) );
  MUX2ND0 U2381 ( .I0(n901), .I1(n1328), .S(n2180), .ZN(n1170) );
  MUX2ND0 U2382 ( .I0(n900), .I1(n1329), .S(n2180), .ZN(n1169) );
  MUX2ND0 U2383 ( .I0(n899), .I1(n1330), .S(n2180), .ZN(n1168) );
  MUX2ND0 U2384 ( .I0(n898), .I1(n1331), .S(n2180), .ZN(n1167) );
  MUX2ND0 U2385 ( .I0(n897), .I1(n1332), .S(n2180), .ZN(n1166) );
  MUX2ND0 U2386 ( .I0(n896), .I1(n1333), .S(n2180), .ZN(n1165) );
  MUX2ND0 U2387 ( .I0(n895), .I1(n1334), .S(n2180), .ZN(n1164) );
  MUX2ND0 U2388 ( .I0(n894), .I1(n1335), .S(n2180), .ZN(n1163) );
  MUX2ND0 U2389 ( .I0(n893), .I1(n1336), .S(n2180), .ZN(n1162) );
  MUX2ND0 U2390 ( .I0(n892), .I1(n1337), .S(n2180), .ZN(n1161) );
  MUX2ND0 U2391 ( .I0(n891), .I1(n1338), .S(n2180), .ZN(n1160) );
  MUX2ND0 U2392 ( .I0(n890), .I1(n1339), .S(n2180), .ZN(n1159) );
  MUX2ND0 U2393 ( .I0(n889), .I1(n1340), .S(n2180), .ZN(n1158) );
  MUX2ND0 U2394 ( .I0(n888), .I1(n1341), .S(n2180), .ZN(n1157) );
  MUX2ND0 U2395 ( .I0(n887), .I1(n1342), .S(n2180), .ZN(n1156) );
  MUX2ND0 U2396 ( .I0(n886), .I1(n1343), .S(n2180), .ZN(n1155) );
  MUX2ND0 U2397 ( .I0(n885), .I1(n1344), .S(n2180), .ZN(n1154) );
  MUX2ND0 U2398 ( .I0(n884), .I1(n1345), .S(n2180), .ZN(n1153) );
  MUX2ND0 U2399 ( .I0(n883), .I1(n1346), .S(n2180), .ZN(n1152) );
  MUX2ND0 U2400 ( .I0(n882), .I1(n1347), .S(n2180), .ZN(n1151) );
  MUX2ND0 U2401 ( .I0(n881), .I1(n1348), .S(n2180), .ZN(n1150) );
  MUX2ND0 U2402 ( .I0(n880), .I1(n1349), .S(n2180), .ZN(n1149) );
  MUX2ND0 U2403 ( .I0(n879), .I1(n1350), .S(n2180), .ZN(n1148) );
  MUX2ND0 U2404 ( .I0(n878), .I1(n1351), .S(n2180), .ZN(n1147) );
  MUX2ND0 U2405 ( .I0(n877), .I1(n1352), .S(n2180), .ZN(n1146) );
  NR2D0 U2406 ( .A1(n2180), .A2(n2601), .ZN(n1145) );
  XNR2D0 U2407 ( .A1(n2957), .A2(n1312), .ZN(n2601) );
  NR2D0 U2408 ( .A1(n2180), .A2(n2602), .ZN(n1144) );
  CKXOR2D0 U2409 ( .A1(n2956), .A2(n2603), .Z(n2602) );
  NR2D0 U2410 ( .A1(n2180), .A2(n2604), .ZN(n1143) );
  XNR2D0 U2411 ( .A1(n2605), .A2(n2955), .ZN(n2604) );
  INR2D0 U2412 ( .A1(n2956), .B1(n2603), .ZN(n2605) );
  CKND2D0 U2413 ( .A1(n2957), .A2(n1312), .ZN(n2603) );
  NR2D0 U2414 ( .A1(n2180), .A2(n2606), .ZN(n1142) );
  AOI31D0 U2415 ( .A1(n2956), .A2(n2957), .A3(n2955), .B(n2958), .ZN(n2606) );
  AO222D0 U2416 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ), .A2(
        n2597), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ), .B2(n2598), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .C2(n2599), 
        .Z(n1141) );
  AO222D0 U2417 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ), .A2(
        n2597), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ), .B2(n2598), .C1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .C2(n2599), 
        .Z(n1140) );
  CKND0 U2418 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CN(
        n2599) );
  AN2D0 U2419 ( .A1(n2607), .A2(n2608), .Z(n2598) );
  AN3D0 U2420 ( .A1(n2609), .A2(n2610), .A3(n2611), .Z(n2597) );
  IND2D0 U2421 ( .A1(n2180), .B1(n2612), .ZN(n1139) );
  OAI21D0 U2422 ( .A1(\SerDes_U1/Rx_ParClk ), .A2(n1312), .B(n2954), .ZN(n2612) );
  MUX2ND0 U2423 ( .I0(n871), .I1(n2613), .S(n2614), .ZN(n1138) );
  AOI211D0 U2424 ( .A1(n2615), .A2(n1315), .B(n2616), .C(n2617), .ZN(n2613) );
  AOI211D0 U2425 ( .A1(n2618), .A2(n2619), .B(n2620), .C(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .ZN(n2616) );
  ND4D0 U2426 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(n2619) );
  MUX2ND0 U2427 ( .I0(n2625), .I1(n2626), .S(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(n2615) );
  CKND2D0 U2428 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2627), .ZN(n2626) );
  AN4D0 U2429 ( .A1(n2624), .A2(n2623), .A3(n2622), .A4(n2621), .Z(n2625) );
  OA211D0 U2430 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n2391), 
        .B(n2628), .C(n2629), .Z(n2621) );
  AOI21D0 U2431 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .A2(n2630), 
        .B(n2631), .ZN(n2629) );
  AOI22D0 U2432 ( .A1(n2392), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), 
        .B1(n2391), .B2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .ZN(
        n2622) );
  OAI33D0 U2433 ( .A1(n2632), .A2(n869), .A3(n2633), .B1(n2634), .B2(n2635), 
        .B3(n2636), .ZN(n1137) );
  XNR2D0 U2434 ( .A1(n2952), .A2(n2392), .ZN(n2636) );
  XNR2D0 U2435 ( .A1(n2953), .A2(n2390), .ZN(n2635) );
  IND3D0 U2436 ( .A1(n2637), .B1(n2638), .B2(n2639), .ZN(n2634) );
  XNR2D0 U2437 ( .A1(n2391), .A2(n1317), .ZN(n2639) );
  XNR2D0 U2438 ( .A1(n2389), .A2(n1316), .ZN(n2638) );
  OAI211D0 U2439 ( .A1(n864), .A2(n2614), .B(n2640), .C(n2641), .ZN(n1136) );
  AOI31D0 U2440 ( .A1(n2642), .A2(n2643), .A3(n2644), .B(n2645), .ZN(n2641) );
  OAI31D0 U2441 ( .A1(n2646), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), 
        .A3(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .B(n2647), .ZN(n2643) );
  MUX2ND0 U2442 ( .I0(n2648), .I1(n2649), .S(n2391), .ZN(n2647) );
  OAI32D0 U2443 ( .A1(n2650), .A2(n2392), .A3(n2624), .B1(n2628), .B2(n2651), 
        .ZN(n2649) );
  OAI32D0 U2444 ( .A1(n2650), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), 
        .A3(n2628), .B1(n2624), .B2(n2651), .ZN(n2648) );
  CKND2D0 U2445 ( .A1(n2652), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n2651) );
  XNR2D0 U2446 ( .A1(n2630), .A2(n2392), .ZN(n2652) );
  MUX2ND0 U2447 ( .I0(n2653), .I1(n2654), .S(n2391), .ZN(n2646) );
  NR2D0 U2448 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .A2(n2624), 
        .ZN(n2654) );
  NR2D0 U2449 ( .A1(n2392), .A2(n2628), .ZN(n2653) );
  ND3D0 U2450 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2655), .A3(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(
        n2640) );
  ND4D0 U2451 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(n2655) );
  XNR2D0 U2452 ( .A1(n2660), .A2(n2661), .ZN(n2658) );
  XNR2D0 U2453 ( .A1(n2630), .A2(n2662), .ZN(n2657) );
  XNR2D0 U2454 ( .A1(n2663), .A2(n2664), .ZN(n2656) );
  OAI32D0 U2455 ( .A1(n2665), .A2(n2666), .A3(n2667), .B1(n2632), .B2(n2668), 
        .ZN(n1135) );
  XNR2D0 U2456 ( .A1(n2951), .A2(n2630), .ZN(n2667) );
  XNR2D0 U2457 ( .A1(n2950), .A2(n2664), .ZN(n2666) );
  ND3D0 U2458 ( .A1(n2669), .A2(n2670), .A3(n2671), .ZN(n2665) );
  XNR2D0 U2459 ( .A1(n2660), .A2(n1393), .ZN(n2671) );
  XNR2D0 U2460 ( .A1(n2672), .A2(n1392), .ZN(n2669) );
  OAI221D0 U2461 ( .A1(n2673), .A2(n2620), .B1(n858), .B2(n2614), .C(n2674), 
        .ZN(n1134) );
  AOI31D0 U2462 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A3(n2675), .B(
        n2633), .ZN(n2674) );
  CKND0 U2463 ( .CLK(n2676), .CN(n2633) );
  CKND0 U2464 ( .CLK(n2627), .CN(n2675) );
  ND4D0 U2465 ( .A1(n2677), .A2(n2678), .A3(n2679), .A4(n2659), .ZN(n2627) );
  XNR2D0 U2466 ( .A1(n2392), .A2(n2680), .ZN(n2679) );
  XNR2D0 U2467 ( .A1(n2681), .A2(n2390), .ZN(n2678) );
  XNR2D0 U2468 ( .A1(n2682), .A2(n2391), .ZN(n2677) );
  OR2D0 U2469 ( .A1(n2954), .A2(n2683), .Z(n2614) );
  CKND0 U2470 ( .CLK(n2618), .CN(n2673) );
  ND4D0 U2471 ( .A1(n2684), .A2(n2642), .A3(n2685), .A4(n2661), .ZN(n2618) );
  CKND2D0 U2472 ( .A1(n2628), .A2(n2624), .ZN(n2661) );
  CKND2D0 U2473 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n2390), 
        .ZN(n2624) );
  CKND2D0 U2474 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .A2(n2672), 
        .ZN(n2628) );
  XNR2D0 U2475 ( .A1(n2686), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), 
        .ZN(n2685) );
  CKND2D0 U2476 ( .A1(n2687), .A2(n2650), .ZN(n2686) );
  MUX2ND0 U2477 ( .I0(n2672), .I1(n2688), .S(n2630), .ZN(n2687) );
  NR2D0 U2478 ( .A1(n2672), .A2(n2664), .ZN(n2688) );
  CKND0 U2479 ( .CLK(n2659), .CN(n2642) );
  IND2D0 U2480 ( .A1(n2631), .B1(n2623), .ZN(n2659) );
  CKND2D0 U2481 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .A2(n2389), 
        .ZN(n2623) );
  NR2D0 U2482 ( .A1(n2389), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), 
        .ZN(n2631) );
  XNR3D0 U2483 ( .A1(n2664), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), 
        .A3(n2391), .ZN(n2684) );
  MUX2D0 U2484 ( .I0(n2951), .I1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), 
        .S(n2670), .Z(n1133) );
  MUX2ND0 U2485 ( .I0(n1392), .I1(n2672), .S(n2670), .ZN(n1132) );
  MUX2ND0 U2486 ( .I0(n1393), .I1(n2660), .S(n2670), .ZN(n1131) );
  MUX2D0 U2487 ( .I0(n2950), .I1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .S(n2670), .Z(n1130) );
  AN2D0 U2488 ( .A1(n2954), .A2(n2632), .Z(n2670) );
  OAI221D0 U2489 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2620), .B1(n2989), .B2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .C(n2689), .ZN(
        n2632) );
  MUX2D0 U2490 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N47 ), .I1(n2952), 
        .S(n2637), .Z(n1129) );
  MUX2D0 U2491 ( .I0(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N45 ), .I1(n2953), 
        .S(n2637), .Z(n1128) );
  MUX2ND0 U2492 ( .I0(n2389), .I1(n1316), .S(n2637), .ZN(n1127) );
  MUX2ND0 U2493 ( .I0(n2391), .I1(n1317), .S(n2637), .ZN(n1126) );
  NR2D0 U2494 ( .A1(n2645), .A2(n2644), .ZN(n2637) );
  CKND0 U2495 ( .CLK(n2689), .CN(n2644) );
  CKND2D0 U2496 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n1315), .ZN(n2689) );
  AO222D0 U2497 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N31 ), .A2(
        n2690), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N39 ), .B2(n2691), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .C2(n2692), 
        .Z(n1125) );
  AO222D0 U2498 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N27 ), .A2(
        n2690), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N35 ), .B2(n2691), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .C2(n2692), 
        .Z(n1124) );
  AO222D0 U2499 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N28 ), .A2(
        n2690), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N36 ), .B2(n2691), .C1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .C2(n2692), 
        .Z(n1123) );
  CKND0 U2500 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ), .CN(
        n2692) );
  AN2D0 U2501 ( .A1(n2693), .A2(n2694), .Z(n2691) );
  AN3D0 U2502 ( .A1(n2695), .A2(n2696), .A3(n2697), .Z(n2690) );
  CKXOR2D0 U2503 ( .A1(\SerDes_U2/Tx_SerClk ), .A2(n2698), .Z(n1122) );
  AO222D0 U2504 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N31 ), .A2(
        n2699), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N39 ), .B2(n2700), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .C2(n2701), 
        .Z(n1120) );
  XNR2D0 U2505 ( .A1(n2702), .A2(\SerDes_U2/Des_U1/SerialClk ), .ZN(n1119) );
  MUX2ND0 U2506 ( .I0(n1384), .I1(n856), .S(n2287), .ZN(n1118) );
  MUX2ND0 U2507 ( .I0(n1383), .I1(n822), .S(n2287), .ZN(n1117) );
  MUX2ND0 U2508 ( .I0(n1382), .I1(n820), .S(n2287), .ZN(n1116) );
  MUX2ND0 U2509 ( .I0(n1381), .I1(n818), .S(n2287), .ZN(n1115) );
  MUX2ND0 U2510 ( .I0(n1380), .I1(n816), .S(n2287), .ZN(n1114) );
  MUX2ND0 U2511 ( .I0(n1379), .I1(n814), .S(n2287), .ZN(n1113) );
  MUX2ND0 U2512 ( .I0(n1378), .I1(n812), .S(n2287), .ZN(n1112) );
  MUX2ND0 U2513 ( .I0(n1377), .I1(n810), .S(n2287), .ZN(n1111) );
  MUX2ND0 U2514 ( .I0(n1376), .I1(n808), .S(n2287), .ZN(n1110) );
  MUX2ND0 U2515 ( .I0(n1375), .I1(n806), .S(n2287), .ZN(n1109) );
  MUX2ND0 U2516 ( .I0(n1374), .I1(n804), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1108) );
  MUX2ND0 U2517 ( .I0(n1373), .I1(n802), .S(n2287), .ZN(n1107) );
  MUX2ND0 U2518 ( .I0(n1372), .I1(n800), .S(n2287), .ZN(n1106) );
  MUX2ND0 U2519 ( .I0(n1371), .I1(n798), .S(n2287), .ZN(n1105) );
  MUX2ND0 U2520 ( .I0(n1370), .I1(n796), .S(n2287), .ZN(n1104) );
  MUX2ND0 U2521 ( .I0(n1369), .I1(n794), .S(n2287), .ZN(n1103) );
  MUX2ND0 U2522 ( .I0(n1368), .I1(n792), .S(n2287), .ZN(n1102) );
  MUX2ND0 U2523 ( .I0(n1367), .I1(n790), .S(n2287), .ZN(n1101) );
  MUX2ND0 U2524 ( .I0(n1366), .I1(n788), .S(n2287), .ZN(n1100) );
  MUX2ND0 U2525 ( .I0(n1365), .I1(n786), .S(n2287), .ZN(n1099) );
  MUX2ND0 U2526 ( .I0(n1364), .I1(n784), .S(n2287), .ZN(n1098) );
  MUX2ND0 U2527 ( .I0(n1363), .I1(n782), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1097) );
  MUX2ND0 U2528 ( .I0(n1362), .I1(n780), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1096) );
  MUX2ND0 U2529 ( .I0(n1361), .I1(n778), .S(n2287), .ZN(n1095) );
  MUX2ND0 U2530 ( .I0(n1360), .I1(n776), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1094) );
  MUX2ND0 U2531 ( .I0(n1359), .I1(n774), .S(n2287), .ZN(n1093) );
  MUX2ND0 U2532 ( .I0(n1358), .I1(n772), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1092) );
  MUX2ND0 U2533 ( .I0(n1357), .I1(n770), .S(n2287), .ZN(n1091) );
  MUX2ND0 U2534 ( .I0(n1356), .I1(n768), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1090) );
  MUX2ND0 U2535 ( .I0(n1355), .I1(n766), .S(n2287), .ZN(n1089) );
  MUX2ND0 U2536 ( .I0(n1354), .I1(n764), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1088) );
  MUX2ND0 U2537 ( .I0(n1353), .I1(n762), .S(\SerDes_U2/Des_U1/DesDec_Rx1/N79 ), 
        .ZN(n1087) );
  MUX2ND0 U2538 ( .I0(n760), .I1(n1353), .S(n2179), .ZN(n1086) );
  MUX2ND0 U2539 ( .I0(n759), .I1(n1354), .S(n2179), .ZN(n1085) );
  MUX2ND0 U2540 ( .I0(n758), .I1(n1355), .S(n2179), .ZN(n1084) );
  MUX2ND0 U2541 ( .I0(n757), .I1(n1356), .S(n2179), .ZN(n1083) );
  MUX2ND0 U2542 ( .I0(n756), .I1(n1357), .S(n2179), .ZN(n1082) );
  MUX2ND0 U2543 ( .I0(n755), .I1(n1358), .S(n2179), .ZN(n1081) );
  MUX2ND0 U2544 ( .I0(n754), .I1(n1359), .S(n2179), .ZN(n1080) );
  MUX2ND0 U2545 ( .I0(n753), .I1(n1360), .S(n2179), .ZN(n1079) );
  MUX2ND0 U2546 ( .I0(n752), .I1(n1361), .S(n2179), .ZN(n1078) );
  MUX2ND0 U2547 ( .I0(n751), .I1(n1362), .S(n2179), .ZN(n1077) );
  MUX2ND0 U2548 ( .I0(n750), .I1(n1363), .S(n2179), .ZN(n1076) );
  MUX2ND0 U2549 ( .I0(n749), .I1(n1364), .S(n2179), .ZN(n1075) );
  MUX2ND0 U2550 ( .I0(n748), .I1(n1365), .S(n2179), .ZN(n1074) );
  MUX2ND0 U2551 ( .I0(n747), .I1(n1366), .S(n2179), .ZN(n1073) );
  MUX2ND0 U2552 ( .I0(n746), .I1(n1367), .S(n2179), .ZN(n1072) );
  MUX2ND0 U2553 ( .I0(n745), .I1(n1368), .S(n2179), .ZN(n1071) );
  MUX2ND0 U2554 ( .I0(n744), .I1(n1369), .S(n2179), .ZN(n1070) );
  MUX2ND0 U2555 ( .I0(n743), .I1(n1370), .S(n2179), .ZN(n1069) );
  MUX2ND0 U2556 ( .I0(n742), .I1(n1371), .S(n2179), .ZN(n1068) );
  MUX2ND0 U2557 ( .I0(n741), .I1(n1372), .S(n2179), .ZN(n1067) );
  MUX2ND0 U2558 ( .I0(n740), .I1(n1373), .S(n2179), .ZN(n1066) );
  MUX2ND0 U2559 ( .I0(n739), .I1(n1374), .S(n2179), .ZN(n1065) );
  MUX2ND0 U2560 ( .I0(n738), .I1(n1375), .S(n2179), .ZN(n1064) );
  MUX2ND0 U2561 ( .I0(n737), .I1(n1376), .S(n2179), .ZN(n1063) );
  MUX2ND0 U2562 ( .I0(n736), .I1(n1377), .S(n2179), .ZN(n1062) );
  MUX2ND0 U2563 ( .I0(n735), .I1(n1378), .S(n2179), .ZN(n1061) );
  MUX2ND0 U2564 ( .I0(n734), .I1(n1379), .S(n2179), .ZN(n1060) );
  MUX2ND0 U2565 ( .I0(n733), .I1(n1380), .S(n2179), .ZN(n1059) );
  MUX2ND0 U2566 ( .I0(n732), .I1(n1381), .S(n2179), .ZN(n1058) );
  MUX2ND0 U2567 ( .I0(n731), .I1(n1382), .S(n2179), .ZN(n1057) );
  MUX2ND0 U2568 ( .I0(n730), .I1(n1383), .S(n2179), .ZN(n1056) );
  MUX2ND0 U2569 ( .I0(n729), .I1(n1384), .S(n2179), .ZN(n1055) );
  NR2D0 U2570 ( .A1(n2179), .A2(n2703), .ZN(n1054) );
  XNR2D0 U2571 ( .A1(n2948), .A2(n1313), .ZN(n2703) );
  NR2D0 U2572 ( .A1(n2179), .A2(n2704), .ZN(n1053) );
  CKXOR2D0 U2573 ( .A1(n2947), .A2(n2705), .Z(n2704) );
  NR2D0 U2574 ( .A1(n2179), .A2(n2706), .ZN(n1052) );
  XNR2D0 U2575 ( .A1(n2707), .A2(n2946), .ZN(n2706) );
  INR2D0 U2576 ( .A1(n2947), .B1(n2705), .ZN(n2707) );
  CKND2D0 U2577 ( .A1(n2948), .A2(n1313), .ZN(n2705) );
  NR2D0 U2578 ( .A1(n2179), .A2(n2708), .ZN(n1051) );
  AOI31D0 U2579 ( .A1(n2947), .A2(n2948), .A3(n2946), .B(n2949), .ZN(n2708) );
  AO222D0 U2580 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N28 ), .A2(
        n2699), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N36 ), .B2(n2700), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .C2(n2701), 
        .Z(n1050) );
  AO222D0 U2581 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N27 ), .A2(
        n2699), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N35 ), .B2(n2700), .C1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .C2(n2701), 
        .Z(n1049) );
  CKND0 U2582 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ), .CN(
        n2701) );
  AN2D0 U2583 ( .A1(n2709), .A2(n2710), .Z(n2700) );
  AN3D0 U2584 ( .A1(n2711), .A2(n2712), .A3(n2713), .Z(n2699) );
  IND2D0 U2585 ( .A1(n2179), .B1(n2714), .ZN(n1048) );
  OAI21D0 U2586 ( .A1(\SerDes_U2/Rx_ParClk ), .A2(n1313), .B(n2945), .ZN(n2714) );
  MUX2ND0 U2587 ( .I0(n723), .I1(n2715), .S(n2716), .ZN(n1047) );
  AOI32D0 U2588 ( .A1(n2717), .A2(n2718), .A3(n2719), .B1(n2720), .B2(n1309), 
        .ZN(n2715) );
  IOA22D0 U2589 ( .B1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .B2(
        n2721), .A1(n2722), .A2(n2723), .ZN(n2720) );
  NR4D0 U2590 ( .A1(n2724), .A2(n2725), .A3(n2726), .A4(n2718), .ZN(n2721) );
  OAI32D0 U2591 ( .A1(n2726), .A2(n2724), .A3(n2725), .B1(n2727), .B2(n2728), 
        .ZN(n2717) );
  CKND0 U2592 ( .CLK(n2729), .CN(n2728) );
  OA22D0 U2593 ( .A1(n2730), .A2(n2731), .B1(n2732), .B2(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .Z(n2727) );
  OAI221D0 U2594 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .A2(n2733), 
        .B1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), .B2(n2734), .C(n2730), 
        .ZN(n2725) );
  OAI22D0 U2595 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n2302), 
        .B1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .B2(n2301), .ZN(
        n2726) );
  OAI31D0 U2596 ( .A1(n2735), .A2(n721), .A3(n2736), .B(n2737), .ZN(n1046) );
  IND4D0 U2597 ( .A1(n2738), .B1(n2739), .B2(n2740), .B3(n2741), .ZN(n2737) );
  XNR2D0 U2598 ( .A1(n2301), .A2(n1319), .ZN(n2741) );
  XNR2D0 U2599 ( .A1(n2302), .A2(n1320), .ZN(n2740) );
  XNR2D0 U2600 ( .A1(n2303), .A2(n1318), .ZN(n2739) );
  OAI211D0 U2601 ( .A1(n717), .A2(n2716), .B(n2742), .C(n2743), .ZN(n1045) );
  AOI31D0 U2602 ( .A1(n2744), .A2(n1309), .A3(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .B(n2719), .ZN(
        n2743) );
  OAI32D0 U2603 ( .A1(n2745), .A2(n2730), .A3(n2731), .B1(n2746), .B2(n2732), 
        .ZN(n2744) );
  CKND2D0 U2604 ( .A1(n2747), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), 
        .ZN(n2732) );
  AOI22D0 U2605 ( .A1(n2724), .A2(n2748), .B1(n2749), .B2(n2303), .ZN(n2746)
         );
  NR2D0 U2606 ( .A1(n2303), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n2724) );
  CKND2D0 U2607 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n2302), 
        .ZN(n2730) );
  XNR2D0 U2608 ( .A1(n2734), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N50 ), 
        .ZN(n2745) );
  OAI31D0 U2609 ( .A1(n2750), .A2(n2747), .A3(n2751), .B(n2723), .ZN(n2742) );
  XNR2D0 U2610 ( .A1(n2748), .A2(n2752), .ZN(n2751) );
  XNR2D0 U2611 ( .A1(n2753), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .ZN(n2750) );
  CKND0 U2612 ( .CLK(n2754), .CN(n2716) );
  OAI211D0 U2613 ( .A1(n2755), .A2(n2722), .B(n2756), .C(n2757), .ZN(n1044) );
  AOI21D0 U2614 ( .A1(n2754), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/NextState [2]), .B(n2758), .ZN(
        n2757) );
  AOI31D0 U2615 ( .A1(n2759), .A2(n2729), .A3(n2747), .B(n2760), .ZN(n2758) );
  CKND0 U2616 ( .CLK(n2731), .CN(n2747) );
  CKXOR2D0 U2617 ( .A1(n2303), .A2(n2761), .Z(n2729) );
  CKND2D0 U2618 ( .A1(n2762), .A2(n2763), .ZN(n2761) );
  XNR2D0 U2619 ( .A1(n2748), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), 
        .ZN(n2759) );
  NR2D0 U2620 ( .A1(n2764), .A2(n2945), .ZN(n2754) );
  ND3D0 U2621 ( .A1(n2765), .A2(n2731), .A3(n2766), .ZN(n2722) );
  XNR2D0 U2622 ( .A1(n2767), .A2(n2302), .ZN(n2766) );
  XNR2D0 U2623 ( .A1(n2733), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), 
        .ZN(n2731) );
  XNR2D0 U2624 ( .A1(n2303), .A2(n2768), .ZN(n2765) );
  CKND0 U2625 ( .CLK(n2723), .CN(n2755) );
  NR2D0 U2626 ( .A1(n2718), .A2(n2769), .ZN(n2723) );
  MUX2ND0 U2627 ( .I0(n2770), .I1(n2771), .S(n2735), .ZN(n1043) );
  ND4D0 U2628 ( .A1(n2772), .A2(n2945), .A3(n2773), .A4(n2774), .ZN(n2771) );
  XNR2D0 U2629 ( .A1(n2733), .A2(n1395), .ZN(n2774) );
  XNR2D0 U2630 ( .A1(n2748), .A2(n1396), .ZN(n2773) );
  XNR2D0 U2631 ( .A1(n2734), .A2(n1394), .ZN(n2772) );
  MUX2ND0 U2632 ( .I0(n1394), .I1(n2734), .S(n2775), .ZN(n1042) );
  MUX2ND0 U2633 ( .I0(n1395), .I1(n2733), .S(n2775), .ZN(n1041) );
  MUX2ND0 U2634 ( .I0(n1396), .I1(n2748), .S(n2775), .ZN(n1040) );
  AN2D0 U2635 ( .A1(n2945), .A2(n2735), .Z(n2775) );
  OAI22D0 U2636 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2760), .B1(n2976), .B2(n2776), .ZN(n2735) );
  NR2D0 U2637 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2769), .ZN(n2776) );
  MUX2ND0 U2638 ( .I0(n2303), .I1(n1318), .S(n2738), .ZN(n1039) );
  MUX2ND0 U2639 ( .I0(n2301), .I1(n1319), .S(n2738), .ZN(n1038) );
  MUX2ND0 U2640 ( .I0(n2302), .I1(n1320), .S(n2738), .ZN(n1037) );
  AOI21D0 U2641 ( .A1(n1309), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .B(n2719), .ZN(
        n2738) );
  AO22D0 U2642 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ), .A2(
        n2697), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ), .B2(n2693), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ) );
  MUX2ND0 U2643 ( .I0(n2777), .I1(n2778), .S(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .ZN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ) );
  CKND2D0 U2644 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        n2694), .ZN(n2778) );
  ND3D0 U2645 ( .A1(n2779), .A2(n2696), .A3(n2780), .ZN(n2694) );
  ND4D0 U2646 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .ZN(n2780) );
  IND3D0 U2647 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .B1(
        n2696), .B2(n2695), .ZN(n2777) );
  CKND2D0 U2648 ( .A1(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .ZN(n2695) );
  AO22D0 U2649 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ), .A2(
        n2697), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ), .B2(n2693), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ) );
  AO22D0 U2650 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ), .A2(
        n2697), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ), .B2(n2693), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ) );
  AN2D0 U2651 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .Z(n2693) );
  NR2D0 U2652 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .ZN(n2697) );
  INR2D0 U2653 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ), .B1(
        n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ) );
  INR2D0 U2654 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ), .B1(
        n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ) );
  INR2D0 U2655 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ), .B1(
        n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ) );
  INR2D0 U2656 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ), .B1(
        n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ) );
  INR2D0 U2657 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ), .B1(
        n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ) );
  INR2D0 U2658 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ), .B1(n2698), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ) );
  OA21D0 U2659 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), 
        .A2(n2696), .B(n2781), .Z(n2698) );
  IOA22D0 U2660 ( .B1(n2782), .B2(n2783), .A1(n2696), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .ZN(n2781)
         );
  AOI221D0 U2661 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .A2(n2779), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .B2(n2784), .C(n2785), .ZN(n2783) );
  AOI221D0 U2662 ( .A1(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(n2786), .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B2(n2787), 
        .C(n2788), .ZN(n2785) );
  IAO21D0 U2663 ( .A1(n2787), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .ZN(n2788)
         );
  OAI32D0 U2664 ( .A1(n2789), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .A3(n2790), 
        .B1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .B2(
        n2791), .ZN(n2787) );
  AN2D0 U2665 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), 
        .A2(n2791), .Z(n2790) );
  CKND0 U2666 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .CN(n2791) );
  CKND0 U2667 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .CN(n2789) );
  CKND0 U2668 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .CN(n2786) );
  CKND0 U2669 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .CN(n2784) );
  NR2D0 U2670 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), 
        .A2(n2779), .ZN(n2782) );
  CKND0 U2671 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .CN(n2779) );
  CKND0 U2672 ( .CLK(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .CN(n2696) );
  AN2D0 U2673 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]), .A2(
        n1247), .Z(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ) );
  CKXOR2D0 U2674 ( .A1(n2968), .A2(n2969), .Z(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ) );
  XNR2D0 U2675 ( .A1(n2792), .A2(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ) );
  OAI221D0 U2676 ( .A1(n2968), .A2(n2793), .B1(n2969), .B2(n2792), .C(n2794), 
        .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ) );
  CKND0 U2677 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .CN(
        n2794) );
  NR2D0 U2678 ( .A1(n2792), .A2(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .ZN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ) );
  CKND0 U2679 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .CN(n2792) );
  IAO21D0 U2680 ( .A1(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .A2(
        n2969), .B(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .ZN(n2793) );
  CKND0 U2681 ( .CLK(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U2/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ) );
  AN2D0 U2682 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [31]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N84 ) );
  AN2D0 U2683 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [30]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N83 ) );
  AN2D0 U2684 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [29]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N82 ) );
  AN2D0 U2685 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [28]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N81 ) );
  AN2D0 U2686 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [27]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N80 ) );
  AN2D0 U2687 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [26]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N79 ) );
  AN2D0 U2688 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [25]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N78 ) );
  AN2D0 U2689 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [24]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N77 ) );
  AN2D0 U2690 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [23]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N76 ) );
  AN2D0 U2691 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [22]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N75 ) );
  AN2D0 U2692 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [21]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N74 ) );
  AN2D0 U2693 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [20]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N73 ) );
  AN2D0 U2694 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [19]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N72 ) );
  AN2D0 U2695 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [18]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N71 ) );
  AN2D0 U2696 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [17]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N70 ) );
  AN2D0 U2697 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [16]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N69 ) );
  AN2D0 U2698 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [15]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N68 ) );
  AN2D0 U2699 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [14]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N67 ) );
  AN2D0 U2700 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [13]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N66 ) );
  AN2D0 U2701 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [12]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N65 ) );
  AN2D0 U2702 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [11]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N64 ) );
  AN2D0 U2703 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [10]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N63 ) );
  AN2D0 U2704 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [9]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N62 ) );
  AN2D0 U2705 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [8]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N61 ) );
  AN2D0 U2706 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [7]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N60 ) );
  AN2D0 U2707 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [6]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N59 ) );
  AN2D0 U2708 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [5]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N58 ) );
  AN2D0 U2709 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [4]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N57 ) );
  AN2D0 U2710 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [3]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N56 ) );
  AN2D0 U2711 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [2]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N55 ) );
  AN2D0 U2712 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [1]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N54 ) );
  AN2D0 U2713 ( .A1(\SerDes_U2/Ser_U1/FIFO_Out [0]), .A2(n2181), .Z(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N53 ) );
  OAI31D0 U2714 ( .A1(n2795), .A2(n2796), .A3(n2797), .B(n2798), .ZN(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N31 ) );
  OAI21D0 U2715 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N23 ), .A2(n2799), .B(n2800), .ZN(n2798) );
  MUX2ND0 U2716 ( .I0(n2801), .I1(n2802), .S(n2799), .ZN(n2800) );
  MUX3ND0 U2717 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/N25 ), .I1(n2803), .I2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N24 ), .S0(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .S1(n2804), .ZN(n2802) );
  NR2D0 U2718 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .ZN(n2804) );
  MUX2D0 U2719 ( .I0(n2805), .I1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N26 ), .S(n2796), 
        .Z(n2803) );
  AN2D0 U2720 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N27 ), .A2(n2797), .Z(n2805)
         );
  IND2D0 U2721 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .B1(n2797), .ZN(
        n2799) );
  CKND0 U2722 ( .CLK(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), .CN(n2797) );
  OAI21D0 U2723 ( .A1(\SerDes_U2/Ser_U1/SerEnc_Tx1/N6 ), .A2(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .B(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .ZN(n2796) );
  MUX2ND0 U2724 ( .I0(\SerDes_U2/Ser_U1/SerEnc_Tx1/N29 ), .I1(
        \SerDes_U2/Ser_U1/SerEnc_Tx1/N28 ), .S(n2801), .ZN(n2795) );
  CKND0 U2725 ( .CLK(\SerDes_U2/Ser_U1/SerEnc_Tx1/N5 ), .CN(n2801) );
  CKND0 U2726 ( .CLK(ClockB), .CN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U2727 ( .A1(n2515), .A2(n2435), .A3(n2491), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N71 ) );
  OAI22D0 U2728 ( .A1(n2435), .A2(n2356), .B1(n2512), .B2(n2491), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N70 ) );
  OA211D0 U2729 ( .A1(n2806), .A2(n2457), .B(n2807), .C(n2483), .Z(n2512) );
  OAI22D0 U2730 ( .A1(n2435), .A2(n2355), .B1(n2513), .B2(n2491), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N69 ) );
  XNR2D0 U2731 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n2806), 
        .ZN(n2513) );
  OAI22D0 U2732 ( .A1(n2435), .A2(n2354), .B1(n2511), .B2(n2491), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N68 ) );
  AN2D0 U2733 ( .A1(n2808), .A2(n2809), .Z(n2511) );
  OAI22D0 U2734 ( .A1(n2435), .A2(n2353), .B1(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .B2(n2491), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N67 ) );
  CKND2D0 U2735 ( .A1(n2973), .A2(n2435), .ZN(n2491) );
  CKND0 U2736 ( .CLK(n2463), .CN(n2435) );
  NR3D0 U2737 ( .A1(n1301), .A2(n1310), .A3(n1300), .ZN(n2463) );
  NR2D0 U2738 ( .A1(n2477), .A2(n2462), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N51 ) );
  XNR2D0 U2739 ( .A1(n2810), .A2(n2356), .ZN(n2477) );
  CKND2D0 U2740 ( .A1(n2515), .A2(n2462), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N50 ) );
  NR2D0 U2741 ( .A1(n2462), .A2(n2476), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ) );
  OAI21D0 U2742 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), .A2(n2811), 
        .B(n2810), .ZN(n2476) );
  CKND2D0 U2743 ( .A1(n2811), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N46 ), 
        .ZN(n2810) );
  NR2D0 U2744 ( .A1(n2354), .A2(n2353), .ZN(n2811) );
  MUX2ND0 U2745 ( .I0(n2812), .I1(n2813), .S(n2354), .ZN(
        \SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ) );
  OR2D0 U2746 ( .A1(n2462), .A2(n2353), .Z(n2813) );
  CKND0 U2747 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ), .CN(n2812) );
  NR2D0 U2748 ( .A1(n2462), .A2(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_Mem1/N44 ), 
        .ZN(\SerDes_U2/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ) );
  CKND2D0 U2749 ( .A1(n1298), .A2(n2515), .ZN(n2462) );
  CKND0 U2750 ( .CLK(n2439), .CN(n2515) );
  NR3D0 U2751 ( .A1(n2971), .A2(n2970), .A3(n2972), .ZN(n2439) );
  ND3D0 U2752 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .A3(n2973), .ZN(n2815)
         );
  IND2D0 U2753 ( .A1(n2483), .B1(n2973), .ZN(n2817) );
  CKND2D0 U2754 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .A2(n2458), 
        .ZN(n2483) );
  ND3D0 U2755 ( .A1(n2806), .A2(n2457), .A3(
        \SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .ZN(n2807) );
  ND3D0 U2756 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n2457), 
        .A3(n2973), .ZN(n2818) );
  CKND0 U2757 ( .CLK(n2806), .CN(n2814) );
  NR2D0 U2758 ( .A1(n2496), .A2(n2495), .ZN(n2806) );
  CKND2D0 U2759 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n2495), 
        .ZN(n2809) );
  CKND2D0 U2760 ( .A1(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .A2(n2496), 
        .ZN(n2808) );
  ND3D0 U2761 ( .A1(n2458), .A2(n2457), .A3(n2973), .ZN(n2819) );
  CKND0 U2762 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [3]), .CN(n2457)
         );
  CKND0 U2763 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .CN(n2458)
         );
  CKND2D0 U2764 ( .A1(n2495), .A2(n2496), .ZN(n2816) );
  CKND0 U2765 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .CN(n2496)
         );
  CKND0 U2766 ( .CLK(\SerDes_U2/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .CN(n2495)
         );
  AO22D0 U2767 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ), .A2(
        n2713), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ), .B2(n2709), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ) );
  MUX2ND0 U2768 ( .I0(n2820), .I1(n2821), .S(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .ZN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ) );
  CKND2D0 U2769 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        n2710), .ZN(n2821) );
  ND3D0 U2770 ( .A1(n2822), .A2(n2712), .A3(n2823), .ZN(n2710) );
  ND4D0 U2771 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .ZN(n2823) );
  IND3D0 U2772 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .B1(
        n2712), .B2(n2711), .ZN(n2820) );
  CKND2D0 U2773 ( .A1(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n2711) );
  AO22D0 U2774 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ), .A2(
        n2713), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ), .B2(n2709), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ) );
  AO22D0 U2775 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ), .A2(
        n2713), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ), .B2(n2709), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ) );
  AN2D0 U2776 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .Z(n2709) );
  NR2D0 U2777 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .ZN(n2713) );
  AN2D0 U2778 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ), .A2(n2702), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ) );
  AN2D0 U2779 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ), .A2(n2702), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ) );
  AN2D0 U2780 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ), .A2(n2702), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ) );
  AN2D0 U2781 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ), .A2(n2702), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ) );
  AN2D0 U2782 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ), .A2(n2702), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ) );
  AN2D0 U2783 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ), .A2(n2702), 
        .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ) );
  OAI21D0 U2784 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), 
        .A2(n2712), .B(n2824), .ZN(n2702) );
  IOA22D0 U2785 ( .B1(n2825), .B2(n2826), .A1(n2712), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .ZN(n2824)
         );
  AOI221D0 U2786 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .A2(n2822), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .B2(n2827), .C(n2828), .ZN(n2826) );
  AOI221D0 U2787 ( .A1(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(n2829), .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B2(n2830), 
        .C(n2831), .ZN(n2828) );
  IAO21D0 U2788 ( .A1(n2830), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .ZN(n2831)
         );
  OAI32D0 U2789 ( .A1(n2832), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .A3(n2833), 
        .B1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .B2(
        n2834), .ZN(n2830) );
  AN2D0 U2790 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), 
        .A2(n2834), .Z(n2833) );
  CKND0 U2791 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .CN(n2834) );
  CKND0 U2792 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .CN(n2832) );
  CKND0 U2793 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .CN(n2829) );
  CKND0 U2794 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .CN(n2827) );
  NR2D0 U2795 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), 
        .A2(n2822), .ZN(n2825) );
  CKND0 U2796 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .CN(n2822) );
  CKND0 U2797 ( .CLK(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .CN(n2712) );
  AN2D0 U2798 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]), .A2(
        n2211), .Z(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ) );
  CKXOR2D0 U2799 ( .A1(n2974), .A2(n2975), .Z(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ) );
  XNR2D0 U2800 ( .A1(n2835), .A2(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ) );
  OAI221D0 U2801 ( .A1(n2974), .A2(n2836), .B1(n2975), .B2(n2835), .C(n2837), 
        .ZN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ) );
  CKND0 U2802 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .CN(
        n2837) );
  NR2D0 U2803 ( .A1(n2835), .A2(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .ZN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ) );
  CKND0 U2804 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .CN(n2835) );
  IAO21D0 U2805 ( .A1(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .A2(
        n2975), .B(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .ZN(n2836) );
  CKND0 U2806 ( .CLK(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U2/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ) );
  CKND2D0 U2807 ( .A1(\SerDes_U2/Rx_ParClk ), .A2(ClockA), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ) );
  IND3D0 U2808 ( .A1(n2977), .B1(n2756), .B2(n2764), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N66 ) );
  OAI22D0 U2809 ( .A1(n2303), .A2(n2756), .B1(n2768), .B2(n2770), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N65 ) );
  AN2D0 U2810 ( .A1(n2838), .A2(n2762), .Z(n2768) );
  MUX2D0 U2811 ( .I0(n2734), .I1(n2763), .S(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .Z(n2838) );
  OAI22D0 U2812 ( .A1(n2302), .A2(n2756), .B1(n2767), .B2(n2770), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N64 ) );
  CKND2D0 U2813 ( .A1(n2977), .A2(n2756), .ZN(n2770) );
  XNR2D0 U2814 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .ZN(n2767) );
  MUX2ND0 U2815 ( .I0(n2301), .I1(n2839), .S(n2756), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N63 ) );
  CKND0 U2816 ( .CLK(n2736), .CN(n2756) );
  NR2D0 U2817 ( .A1(n2718), .A2(n2760), .ZN(n2736) );
  CKND0 U2818 ( .CLK(n2719), .CN(n2760) );
  NR2D0 U2819 ( .A1(n1309), .A2(n2769), .ZN(n2719) );
  NR2D0 U2820 ( .A1(n2753), .A2(n2840), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ) );
  XNR2D0 U2821 ( .A1(n2303), .A2(n2841), .ZN(n2753) );
  CKND2D0 U2822 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N49 ), .A2(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .ZN(n2841) );
  CKND2D0 U2823 ( .A1(n721), .A2(n2764), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ) );
  INR2D0 U2824 ( .A1(n2752), .B1(n2840), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ) );
  XNR2D0 U2825 ( .A1(n2302), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), 
        .ZN(n2752) );
  NR2D0 U2826 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N48 ), .A2(n2840), 
        .ZN(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/N46 ) );
  IND2D0 U2827 ( .A1(n721), .B1(n2764), .ZN(n2840) );
  ND3D0 U2828 ( .A1(n2718), .A2(n1309), .A3(n2769), .ZN(n2764) );
  CKND0 U2829 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .CN(
        n2769) );
  CKND0 U2830 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .CN(
        n2718) );
  NR3D0 U2831 ( .A1(n2839), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N99 ) );
  NR3D0 U2832 ( .A1(n2842), .A2(n2748), .A3(n2734), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N358 ) );
  NR3D0 U2833 ( .A1(n2839), .A2(n2748), .A3(n2734), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N325 ) );
  CKND0 U2834 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .CN(n2748)
         );
  CKND0 U2835 ( .CLK(n2749), .CN(n2762) );
  NR2D0 U2836 ( .A1(n2734), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), 
        .ZN(n2749) );
  CKND2D0 U2837 ( .A1(n2977), .A2(n2733), .ZN(n2839) );
  CKND0 U2838 ( .CLK(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .CN(n2733)
         );
  CKND2D0 U2839 ( .A1(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n2734), 
        .ZN(n2763) );
  NR3D0 U2840 ( .A1(n2842), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U2/Des_U1/FIFO_Rx1/FIFO_Mem1/N160 ) );
  CKND2D0 U2841 ( .A1(n2977), .A2(\SerDes_U2/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), 
        .ZN(n2842) );
  AN2D0 U2842 ( .A1(\SerDes_U2/Des_U1/SerialClk ), .A2(
        \SerDes_U2/SerLineValid ), .Z(\SerDes_U2/Des_U1/DesDec_Rx1/SerClock )
         );
  NR2D0 U2843 ( .A1(n2843), .A2(n2844), .ZN(\SerDes_U2/Des_U1/DesDec_Rx1/N47 )
         );
  CKND2D0 U2844 ( .A1(n2845), .A2(n2846), .ZN(n2844) );
  NR4D0 U2845 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[7] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[6] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[5] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[4] ), .ZN(n2846) );
  NR4D0 U2846 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[3] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[2] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[1] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[0] ), .ZN(n2845) );
  AN4D0 U2847 ( .A1(n2847), .A2(n2848), .A3(n2849), .A4(n2850), .Z(n2843) );
  NR4D0 U2848 ( .A1(n2851), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[50] ), 
        .A3(n855), .A4(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[49] ), .ZN(n2850)
         );
  ND3D0 U2849 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[52] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[51] ), .A3(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[36] ), .ZN(n2851) );
  NR4D0 U2850 ( .A1(n2852), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[21] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[33] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[20] ), .ZN(n2849) );
  ND3D0 U2851 ( .A1(n841), .A2(n837), .A3(n842), .ZN(n2852) );
  NR4D0 U2852 ( .A1(n2853), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[39] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[54] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[37] ), .ZN(n2848) );
  ND3D0 U2853 ( .A1(n2982), .A2(n849), .A3(n2981), .ZN(n2853) );
  NR4D0 U2854 ( .A1(n2854), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[17] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[23] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/FrameSR[16] ), .ZN(n2847) );
  ND3D0 U2855 ( .A1(n2979), .A2(n2980), .A3(n2978), .ZN(n2854) );
  OA21D0 U2856 ( .A1(n2855), .A2(n2983), .B(\SerDes_U2/SerLineValid ), .Z(
        \SerDes_U2/Des_U1/DesDec_Rx1/N43 ) );
  NR4D0 U2857 ( .A1(n2856), .A2(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[2] ), 
        .A3(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[4] ), .A4(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[3] ), .ZN(n2855) );
  OR2D0 U2858 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/Count32[1] ), .A2(
        \SerDes_U2/Des_U1/DesDec_Rx1/Count32[0] ), .Z(n2856) );
  INR2D0 U2859 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N34 ), .B1(n2983), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N42 ) );
  INR2D0 U2860 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N33 ), .B1(n2983), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N41 ) );
  INR2D0 U2861 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N32 ), .B1(n2983), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N40 ) );
  INR2D0 U2862 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N31 ), .B1(n2983), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N39 ) );
  INR2D0 U2863 ( .A1(\SerDes_U2/Des_U1/DesDec_Rx1/N30 ), .B1(n2983), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N38 ) );
  NR2D0 U2864 ( .A1(n2983), .A2(\SerDes_U2/Rx_ParClk ), .ZN(
        \SerDes_U2/Des_U1/DesDec_Rx1/N37 ) );
  AO22D0 U2865 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N32 ), .A2(
        n2595), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N40 ), .B2(n2591), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N55 ) );
  MUX2ND0 U2866 ( .I0(n2857), .I1(n2858), .S(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .ZN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N54 ) );
  CKND2D0 U2867 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        n2592), .ZN(n2858) );
  ND3D0 U2868 ( .A1(n2859), .A2(n2594), .A3(n2860), .ZN(n2592) );
  ND4D0 U2869 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .ZN(n2860) );
  IND3D0 U2870 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .B1(
        n2594), .B2(n2593), .ZN(n2857) );
  CKND2D0 U2871 ( .A1(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .ZN(n2593) );
  AO22D0 U2872 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N30 ), .A2(
        n2595), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N38 ), .B2(n2591), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N51 ) );
  AO22D0 U2873 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N29 ), .A2(
        n2595), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N37 ), .B2(n2591), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N49 ) );
  AN2D0 U2874 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .Z(n2591) );
  NR2D0 U2875 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [0]), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/AdjFreq [1]), .ZN(n2595) );
  INR2D0 U2876 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N14 ), .B1(
        n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N21 ) );
  INR2D0 U2877 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N13 ), .B1(
        n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N20 ) );
  INR2D0 U2878 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N12 ), .B1(
        n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N19 ) );
  INR2D0 U2879 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N11 ), .B1(
        n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N18 ) );
  INR2D0 U2880 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N10 ), .B1(
        n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N17 ) );
  INR2D0 U2881 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N9 ), .B1(n2596), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/N16 ) );
  OA21D0 U2882 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), 
        .A2(n2594), .B(n2861), .Z(n2596) );
  IOA22D0 U2883 ( .B1(n2862), .B2(n2863), .A1(n2594), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[5] ), .ZN(n2861)
         );
  AOI221D0 U2884 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), .A2(n2859), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .B2(n2864), .C(n2865), .ZN(n2863) );
  AOI221D0 U2885 ( .A1(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .A2(n2866), .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B2(n2867), 
        .C(n2868), .ZN(n2865) );
  IAO21D0 U2886 ( .A1(n2867), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[2] ), .ZN(n2868)
         );
  OAI32D0 U2887 ( .A1(n2869), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[0] ), .A3(n2870), 
        .B1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), .B2(
        n2871), .ZN(n2867) );
  AN2D0 U2888 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[1] ), 
        .A2(n2871), .Z(n2870) );
  CKND0 U2889 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[1] ), .CN(n2871) );
  CKND0 U2890 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[0] ), .CN(n2869) );
  CKND0 U2891 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[3] ), 
        .CN(n2866) );
  CKND0 U2892 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[3] ), .CN(n2864) );
  NR2D0 U2893 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastDivvy[4] ), 
        .A2(n2859), .ZN(n2862) );
  CKND0 U2894 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[4] ), .CN(n2859) );
  CKND0 U2895 ( .CLK(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/DivideFactor[5] ), .CN(n2594) );
  AN2D0 U2896 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/WireD [5]), .A2(
        n2264), .Z(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/VFO1/FastClock ) );
  CKXOR2D0 U2897 ( .A1(n2984), .A2(n2985), .Z(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N8 ) );
  XNR2D0 U2898 ( .A1(n2872), .A2(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N6 ) );
  OAI221D0 U2899 ( .A1(n2984), .A2(n2873), .B1(n2985), .B2(n2872), .C(n2874), 
        .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N20 ) );
  CKND0 U2900 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ), .CN(
        n2874) );
  NR2D0 U2901 ( .A1(n2872), .A2(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .ZN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N9 ) );
  CKND0 U2902 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .CN(n2872) );
  IAO21D0 U2903 ( .A1(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ), .A2(
        n2985), .B(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[1] ), 
        .ZN(n2873) );
  CKND0 U2904 ( .CLK(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U1/Ser_U1/SerTx_Tx1/PLL_TxU1/Comp1/N5 ) );
  AN2D0 U2905 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [31]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N84 ) );
  AN2D0 U2906 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [30]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N83 ) );
  AN2D0 U2907 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [29]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N82 ) );
  AN2D0 U2908 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [28]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N81 ) );
  AN2D0 U2909 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [27]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N80 ) );
  AN2D0 U2910 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [26]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N79 ) );
  AN2D0 U2911 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [25]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N78 ) );
  AN2D0 U2912 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [24]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N77 ) );
  AN2D0 U2913 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [23]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N76 ) );
  AN2D0 U2914 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [22]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N75 ) );
  AN2D0 U2915 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [21]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N74 ) );
  AN2D0 U2916 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [20]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N73 ) );
  AN2D0 U2917 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [19]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N72 ) );
  AN2D0 U2918 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [18]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N71 ) );
  AN2D0 U2919 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [17]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N70 ) );
  AN2D0 U2920 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [16]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N69 ) );
  AN2D0 U2921 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [15]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N68 ) );
  AN2D0 U2922 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [14]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N67 ) );
  AN2D0 U2923 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [13]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N66 ) );
  AN2D0 U2924 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [12]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N65 ) );
  AN2D0 U2925 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [11]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N64 ) );
  AN2D0 U2926 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [10]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N63 ) );
  AN2D0 U2927 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [9]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N62 ) );
  AN2D0 U2928 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [8]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N61 ) );
  AN2D0 U2929 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [7]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N60 ) );
  AN2D0 U2930 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [6]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N59 ) );
  AN2D0 U2931 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [5]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N58 ) );
  AN2D0 U2932 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [4]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N57 ) );
  AN2D0 U2933 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [3]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N56 ) );
  AN2D0 U2934 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [2]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N55 ) );
  AN2D0 U2935 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [1]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N54 ) );
  AN2D0 U2936 ( .A1(\SerDes_U1/Ser_U1/FIFO_Out [0]), .A2(n1296), .Z(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N53 ) );
  OAI31D0 U2937 ( .A1(n2875), .A2(n2876), .A3(n2877), .B(n2878), .ZN(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N31 ) );
  OAI21D0 U2938 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N23 ), .A2(n2879), .B(n2880), .ZN(n2878) );
  MUX2ND0 U2939 ( .I0(n2881), .I1(n2882), .S(n2879), .ZN(n2880) );
  MUX3ND0 U2940 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/N25 ), .I1(n2883), .I2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N24 ), .S0(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .S1(n2884), .ZN(n2882) );
  NR2D0 U2941 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .ZN(n2884) );
  MUX2D0 U2942 ( .I0(n2885), .I1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N26 ), .S(n2876), 
        .Z(n2883) );
  AN2D0 U2943 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N27 ), .A2(n2877), .Z(n2885)
         );
  IND2D0 U2944 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .B1(n2877), .ZN(
        n2879) );
  CKND0 U2945 ( .CLK(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), .CN(n2877) );
  OAI21D0 U2946 ( .A1(\SerDes_U1/Ser_U1/SerEnc_Tx1/N6 ), .A2(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .B(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/Sh_N[5] ), .ZN(n2876) );
  MUX2ND0 U2947 ( .I0(\SerDes_U1/Ser_U1/SerEnc_Tx1/N29 ), .I1(
        \SerDes_U1/Ser_U1/SerEnc_Tx1/N28 ), .S(n2881), .ZN(n2875) );
  CKND0 U2948 ( .CLK(\SerDes_U1/Ser_U1/SerEnc_Tx1/N5 ), .CN(n2881) );
  CKND0 U2949 ( .CLK(ClockA), .CN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U2950 ( .A1(n2523), .A2(n1311), .A3(n2518), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N66 ) );
  OAI21D0 U2951 ( .A1(n2542), .A2(n2886), .B(n2887), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N65 ) );
  MUX2ND0 U2952 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .I1(n2888), 
        .S(n2523), .ZN(n2887) );
  NR2D0 U2953 ( .A1(n2586), .A2(n1311), .ZN(n2888) );
  CKND0 U2954 ( .CLK(n2547), .CN(n2586) );
  OAI21D0 U2955 ( .A1(n2582), .A2(n2573), .B(n2567), .ZN(n2547) );
  OAI21D0 U2956 ( .A1(n2565), .A2(n2886), .B(n2889), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N64 ) );
  MUX2ND0 U2957 ( .I0(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .I1(n2890), 
        .S(n2523), .ZN(n2889) );
  NR2D0 U2958 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n2891), 
        .ZN(n2890) );
  OAI21D0 U2959 ( .A1(n2523), .A2(n2324), .B(n2886), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N63 ) );
  IND2D0 U2960 ( .A1(n2892), .B1(n2523), .ZN(n2886) );
  CKND2D0 U2961 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .A2(
        n2536), .ZN(n2523) );
  CKND0 U2962 ( .CLK(n2526), .CN(n2536) );
  CKND2D0 U2963 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .ZN(n2526) );
  NR2D0 U2964 ( .A1(n2562), .A2(n2548), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N49 ) );
  CKXOR2D0 U2965 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N50 ), .A2(n2893), 
        .Z(n2562) );
  CKND2D0 U2966 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N49 ), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), .ZN(n2893) );
  CKND2D0 U2967 ( .A1(n1015), .A2(n2518), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N48 ) );
  CKND0 U2968 ( .CLK(n2529), .CN(n2518) );
  MUX2ND0 U2969 ( .I0(n2894), .I1(n2895), .S(n2325), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N47 ) );
  CKND2D0 U2970 ( .A1(n2896), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(n2895) );
  CKND0 U2971 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ), .CN(n2894) );
  NR2D0 U2972 ( .A1(n2548), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N48 ), 
        .ZN(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/N46 ) );
  CKND0 U2973 ( .CLK(n2896), .CN(n2548) );
  NR2D0 U2974 ( .A1(n2529), .A2(n1015), .ZN(n2896) );
  NR2D0 U2975 ( .A1(n2521), .A2(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[1] ), .ZN(n2529) );
  IND2D0 U2976 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[0] ), .B1(
        n2540), .ZN(n2521) );
  CKND0 U2977 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_SM1/CurState[2] ), .CN(
        n2540) );
  NR3D0 U2978 ( .A1(n2892), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N99 ) );
  NR3D0 U2979 ( .A1(n2891), .A2(n2542), .A3(n2565), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N358 ) );
  NR3D0 U2980 ( .A1(n2892), .A2(n2542), .A3(n2565), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N325 ) );
  CKND2D0 U2981 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), .A2(n2565), 
        .ZN(n2567) );
  CKND0 U2982 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .CN(n2565)
         );
  CKND2D0 U2983 ( .A1(n2986), .A2(n2573), .ZN(n2892) );
  CKND0 U2984 ( .CLK(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), .CN(n2573)
         );
  CKND2D0 U2985 ( .A1(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .A2(n2542), 
        .ZN(n2582) );
  NR3D0 U2986 ( .A1(n2891), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [2]), 
        .A3(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [1]), .ZN(
        \SerDes_U1/Ser_U1/FIFO_Tx1/FIFO_Mem1/N160 ) );
  CKND2D0 U2987 ( .A1(n2986), .A2(\SerDes_U1/Ser_U1/FIFO_Tx1/SM_WriteAddr [0]), 
        .ZN(n2891) );
  AO22D0 U2988 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N32 ), .A2(
        n2611), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N40 ), .B2(n2607), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N55 ) );
  MUX2ND0 U2989 ( .I0(n2897), .I1(n2898), .S(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .ZN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N54 ) );
  CKND2D0 U2990 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        n2608), .ZN(n2898) );
  ND3D0 U2991 ( .A1(n2899), .A2(n2610), .A3(n2900), .ZN(n2608) );
  ND4D0 U2992 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .A3(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .A4(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .ZN(n2900) );
  IND3D0 U2993 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .B1(
        n2610), .B2(n2609), .ZN(n2897) );
  CKND2D0 U2994 ( .A1(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n2609) );
  AO22D0 U2995 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N30 ), .A2(
        n2611), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N38 ), .B2(n2607), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N51 ) );
  AO22D0 U2996 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N29 ), .A2(
        n2611), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N37 ), .B2(n2607), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N49 ) );
  AN2D0 U2997 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .Z(n2607) );
  NR2D0 U2998 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [0]), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/AdjFreq [1]), .ZN(n2611) );
  AN2D0 U2999 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N14 ), .A2(n2600), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N21 ) );
  AN2D0 U3000 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N13 ), .A2(n2600), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N20 ) );
  AN2D0 U3001 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N12 ), .A2(n2600), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N19 ) );
  AN2D0 U3002 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N11 ), .A2(n2600), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N18 ) );
  AN2D0 U3003 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N10 ), .A2(n2600), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N17 ) );
  AN2D0 U3004 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N9 ), .A2(n2600), 
        .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/N16 ) );
  OAI21D0 U3005 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), 
        .A2(n2610), .B(n2901), .ZN(n2600) );
  IOA22D0 U3006 ( .B1(n2902), .B2(n2903), .A1(n2610), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[5] ), .ZN(n2901)
         );
  AOI221D0 U3007 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), .A2(n2899), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .B2(n2904), .C(n2905), .ZN(n2903) );
  AOI221D0 U3008 ( .A1(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(n2906), .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B2(n2907), 
        .C(n2908), .ZN(n2905) );
  IAO21D0 U3009 ( .A1(n2907), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[2] ), .B(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[2] ), .ZN(n2908)
         );
  OAI32D0 U3010 ( .A1(n2909), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[0] ), .A3(n2910), 
        .B1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), .B2(
        n2911), .ZN(n2907) );
  AN2D0 U3011 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[1] ), 
        .A2(n2911), .Z(n2910) );
  CKND0 U3012 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[1] ), .CN(n2911) );
  CKND0 U3013 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[0] ), .CN(n2909) );
  CKND0 U3014 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[3] ), 
        .CN(n2906) );
  CKND0 U3015 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[3] ), .CN(n2904) );
  NR2D0 U3016 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastDivvy[4] ), 
        .A2(n2899), .ZN(n2902) );
  CKND0 U3017 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[4] ), .CN(n2899) );
  CKND0 U3018 ( .CLK(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/DivideFactor[5] ), .CN(n2610) );
  AN2D0 U3019 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/WireD [5]), .A2(
        n2257), .Z(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/VFO1/FastClock ) );
  CKXOR2D0 U3020 ( .A1(n2987), .A2(n2988), .Z(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N8 ) );
  XNR2D0 U3021 ( .A1(n2912), .A2(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), .ZN(
        \SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N6 ) );
  OAI221D0 U3022 ( .A1(n2987), .A2(n2913), .B1(n2988), .B2(n2912), .C(n2914), 
        .ZN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N20 ) );
  CKND0 U3023 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ), .CN(
        n2914) );
  NR2D0 U3024 ( .A1(n2912), .A2(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .ZN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N9 ) );
  CKND0 U3025 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .CN(n2912) );
  IAO21D0 U3026 ( .A1(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ), .A2(
        n2988), .B(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .ZN(n2913) );
  CKND0 U3027 ( .CLK(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/ClockInN[0] ), 
        .CN(\SerDes_U1/Des_U1/SerRx_Rx1/PLL_RxU1/Comp1/N5 ) );
  CKND2D0 U3028 ( .A1(\SerDes_U1/Rx_ParClk ), .A2(ClockB), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/StateClockRaw ) );
  ND3D0 U3029 ( .A1(n2683), .A2(n2676), .A3(n2668), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N71 ) );
  OAI22D0 U3030 ( .A1(n2392), .A2(n2676), .B1(n2680), .B2(n2668), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N70 ) );
  OA211D0 U3031 ( .A1(n2915), .A2(n2630), .B(n2916), .C(n2650), .Z(n2680) );
  OAI22D0 U3032 ( .A1(n2391), .A2(n2676), .B1(n2682), .B2(n2668), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N69 ) );
  XNR2D0 U3033 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n2915), 
        .ZN(n2682) );
  OAI22D0 U3034 ( .A1(n2390), .A2(n2676), .B1(n2681), .B2(n2668), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N68 ) );
  AN2D0 U3035 ( .A1(n2917), .A2(n2918), .Z(n2681) );
  OAI22D0 U3036 ( .A1(n2389), .A2(n2676), .B1(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .B2(n2668), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N67 ) );
  CKND2D0 U3037 ( .A1(n2990), .A2(n2676), .ZN(n2668) );
  CKND2D0 U3038 ( .A1(n2645), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .ZN(n2676) );
  CKND0 U3039 ( .CLK(n2620), .CN(n2645) );
  CKND2D0 U3040 ( .A1(n2989), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(n2620) );
  NR2D0 U3041 ( .A1(n2662), .A2(n2919), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N51 ) );
  XNR2D0 U3042 ( .A1(n2920), .A2(n2392), .ZN(n2662) );
  CKND2D0 U3043 ( .A1(n2683), .A2(n2919), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N50 ) );
  CKND0 U3044 ( .CLK(n2617), .CN(n2683) );
  NR2D0 U3045 ( .A1(n2663), .A2(n2919), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N49 ) );
  OAI21D0 U3046 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), .A2(n2921), 
        .B(n2920), .ZN(n2663) );
  CKND2D0 U3047 ( .A1(n2921), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N46 ), 
        .ZN(n2920) );
  NR2D0 U3048 ( .A1(n2389), .A2(n2390), .ZN(n2921) );
  MUX2ND0 U3049 ( .I0(n2922), .I1(n2923), .S(n2390), .ZN(
        \SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N48 ) );
  CKND2D0 U3050 ( .A1(n2924), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), 
        .ZN(n2923) );
  CKND0 U3051 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ), .CN(n2922) );
  NR2D0 U3052 ( .A1(n2919), .A2(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_Mem1/N44 ), 
        .ZN(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/N47 ) );
  CKND0 U3053 ( .CLK(n2924), .CN(n2919) );
  NR2D0 U3054 ( .A1(n869), .A2(n2617), .ZN(n2924) );
  NR3D0 U3055 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[1] ), .A2(
        n2989), .A3(\SerDes_U1/Des_U1/FIFO_Rx1/FIFO_SM1/CurState[0] ), .ZN(
        n2617) );
  ND3D0 U3056 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .A2(
        \SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A3(n2990), .ZN(n2926)
         );
  IND2D0 U3057 ( .A1(n2650), .B1(n2990), .ZN(n2928) );
  CKND2D0 U3058 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [3]), .A2(n2664), 
        .ZN(n2650) );
  ND3D0 U3059 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n2630), 
        .A3(n2915), .ZN(n2916) );
  ND3D0 U3060 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .A2(n2630), 
        .A3(n2990), .ZN(n2929) );
  CKND0 U3061 ( .CLK(n2915), .CN(n2925) );
  NR2D0 U3062 ( .A1(n2660), .A2(n2672), .ZN(n2915) );
  CKND2D0 U3063 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .A2(n2660), 
        .ZN(n2918) );
  CKND2D0 U3064 ( .A1(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .A2(n2672), 
        .ZN(n2917) );
  ND3D0 U3065 ( .A1(n2664), .A2(n2630), .A3(n2990), .ZN(n2930) );
  CKND0 U3066 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [2]), .CN(n2664)
         );
  CKND2D0 U3067 ( .A1(n2660), .A2(n2672), .ZN(n2927) );
  CKND0 U3068 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [1]), .CN(n2672)
         );
  CKND0 U3069 ( .CLK(\SerDes_U1/Des_U1/FIFO_Rx1/SM_WriteAddr [0]), .CN(n2660)
         );
  AN2D0 U3070 ( .A1(\SerDes_U1/Des_U1/SerialClk ), .A2(
        \SerDes_U1/SerLineValid ), .Z(\SerDes_U1/Des_U1/DesDec_Rx1/SerClock )
         );
  NR2D0 U3071 ( .A1(n2931), .A2(n2932), .ZN(\SerDes_U1/Des_U1/DesDec_Rx1/N47 )
         );
  CKND2D0 U3072 ( .A1(n2933), .A2(n2934), .ZN(n2932) );
  NR4D0 U3073 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[7] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[6] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[5] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[4] ), .ZN(n2934) );
  NR4D0 U3074 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[3] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[2] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[1] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[0] ), .ZN(n2933) );
  AN4D0 U3075 ( .A1(n2935), .A2(n2936), .A3(n2937), .A4(n2938), .Z(n2931) );
  NR4D0 U3076 ( .A1(n2939), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[50] ), 
        .A3(n1003), .A4(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[49] ), .ZN(n2938)
         );
  ND3D0 U3077 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[52] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[51] ), .A3(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[36] ), .ZN(n2939) );
  NR4D0 U3078 ( .A1(n2940), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[21] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[33] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[20] ), .ZN(n2937) );
  ND3D0 U3079 ( .A1(n989), .A2(n985), .A3(n990), .ZN(n2940) );
  NR4D0 U3080 ( .A1(n2941), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[39] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[54] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[37] ), .ZN(n2936) );
  ND3D0 U3081 ( .A1(n2995), .A2(n997), .A3(n2994), .ZN(n2941) );
  NR4D0 U3082 ( .A1(n2942), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[17] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[23] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/FrameSR[16] ), .ZN(n2935) );
  ND3D0 U3083 ( .A1(n2992), .A2(n2993), .A3(n2991), .ZN(n2942) );
  OA21D0 U3084 ( .A1(n2943), .A2(n2996), .B(\SerDes_U1/SerLineValid ), .Z(
        \SerDes_U1/Des_U1/DesDec_Rx1/N43 ) );
  NR4D0 U3085 ( .A1(n2944), .A2(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[2] ), 
        .A3(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[4] ), .A4(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[3] ), .ZN(n2943) );
  OR2D0 U3086 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/Count32[1] ), .A2(
        \SerDes_U1/Des_U1/DesDec_Rx1/Count32[0] ), .Z(n2944) );
  INR2D0 U3087 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N34 ), .B1(n2996), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N42 ) );
  INR2D0 U3088 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N33 ), .B1(n2996), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N41 ) );
  INR2D0 U3089 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N32 ), .B1(n2996), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N40 ) );
  INR2D0 U3090 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N31 ), .B1(n2996), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N39 ) );
  INR2D0 U3091 ( .A1(\SerDes_U1/Des_U1/DesDec_Rx1/N30 ), .B1(n2996), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N38 ) );
  NR2D0 U3092 ( .A1(n2996), .A2(\SerDes_U1/Rx_ParClk ), .ZN(
        \SerDes_U1/Des_U1/DesDec_Rx1/N37 ) );
endmodule


module FullDup_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_2 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_4 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_5 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_6 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_7 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_8 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_9 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_3 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_10 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_11 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_12 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_inc_13 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_4 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FullDup_DW01_dec_5 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

