
module fifo_cntrl ( clk, rstN, wrN, rdN, empty, full, mem_empty_even, 
    mem_empty_odd, mem_full_even, mem_full_odd, ldN_even, ldN_odd, 
    out_sel_odd_evenN, rdN_even, wrN_even, rdN_odd, wrN_odd );
input  clk, rstN, wrN, rdN, mem_empty_even, mem_empty_odd, mem_full_even, 
    mem_full_odd;
output empty, full, ldN_even, ldN_odd, out_sel_odd_evenN, rdN_even, wrN_even, 
    rdN_odd, wrN_odd;
    wire N5, N9, in_sel_odd_evenN, N17, mem_empty_even_dly, mem_empty_odd_dly, 
        dout_avail_even, N49, dout_avail_odd, N66, wrN_even_dly_by_rdN, 
        wrN_odd_dly_by_rdN, ldN_even_dly, ldN_odd_dly, N75, N77, N78, N108, 
        N110, n7, n8, n10, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
        n22, n24;
    xor2a2 U4 ( .A(N17), .B(wrN), .Y(n8) );
    and2b2 U5 ( .A(n14), .B(n13), .Y(rdN_odd) );
    and2b2 U6 ( .A(n7), .B(n12), .Y(rdN_even) );
    xor2a2 U7 ( .A(N5), .B(rdN), .Y(n10) );
    inv1a1 U8 ( .A(rstN), .Y(N9) );
    mx2d3 U9 ( .D0(n18), .D1(n21), .S(mem_empty_odd), .Y(N110) );
    mx2d3 U10 ( .D0(n19), .D1(n22), .S(mem_empty_even), .Y(N108) );
    inv1a1 U11 ( .A(mem_empty_odd), .Y(N66) );
    inv1a1 U12 ( .A(mem_empty_even), .Y(N49) );
    clk1a15 U13 ( .A(n16), .Y(wrN_odd) );
    clk1a15 U14 ( .A(n15), .Y(wrN_even) );
    oa1a3 U15 ( .A(ldN_odd_dly), .B(n14), .C(wrN_odd_dly_by_rdN), .Y(n16) );
    inv1a3 U16 ( .A(n20), .Y(n14) );
    oa1a3 U17 ( .A(ldN_even_dly), .B(n7), .C(wrN_even_dly_by_rdN), .Y(n15) );
    or2b2 U18 ( .A(N17), .B(wrN), .Y(ldN_even) );
    and2a3 U19 ( .A(mem_full_even), .B(mem_full_odd), .Y(full) );
    inv1a3 U20 ( .A(out_sel_odd_evenN), .Y(N5) );
    fdmf1a3 ldN_odd_dly_reg ( .D0(N9), .D1(1'b1), .S(ldN_odd), .CLK(clk), .Q(
        ldN_odd_dly) );
    fdf1a3 ldN_even_dly_reg ( .D(N75), .CLK(clk), .Q(ldN_even_dly) );
    fdf1a3 wrN_odd_dly_by_rdN_reg ( .D(N78), .CLK(clk), .Q(wrN_odd_dly_by_rdN)
         );
    fdf1a3 wrN_even_dly_by_rdN_reg ( .D(N77), .CLK(clk), .Q(
        wrN_even_dly_by_rdN) );
    fdef2a3 dout_avail_odd_reg ( .D(N66), .E(N110), .CLK(clk), .CLR(rstN), .Q(
        dout_avail_odd) );
    inv1a1 U21 ( .A(dout_avail_odd), .Y(n17) );
    fdef2a3 dout_avail_even_reg ( .D(N49), .E(N108), .CLK(clk), .CLR(rstN), 
        .Q(dout_avail_even) );
    inv1a1 U22 ( .A(dout_avail_even), .Y(n24) );
    fdf2a3 mem_empty_odd_dly_reg ( .D(mem_empty_odd), .CLK(clk), .CLR(rstN), 
        .Q(mem_empty_odd_dly) );
    inv1a1 U23 ( .A(mem_empty_odd_dly), .Y(n18) );
    fdf2a3 mem_empty_even_dly_reg ( .D(mem_empty_even), .CLK(clk), .CLR(rstN), 
        .Q(mem_empty_even_dly) );
    inv1a1 U24 ( .A(mem_empty_even_dly), .Y(n19) );
    and3d2 U25 ( .A(rdN), .B(out_sel_odd_evenN), .C(mem_empty_even), .Y(n7) );
    inv1a3 U26 ( .A(in_sel_odd_evenN), .Y(N17) );
    or2b2 U27 ( .A(in_sel_odd_evenN), .B(wrN), .Y(ldN_odd) );
    fdf2a3 in_sel_odd_evenN_reg ( .D(n8), .CLK(clk), .CLR(rstN), .Q(
        in_sel_odd_evenN) );
    fdf2a9 out_sel_odd_evenN_reg ( .D(n10), .CLK(clk), .CLR(rstN), .Q(
        out_sel_odd_evenN) );
    and2b2 U29 ( .A(dout_avail_even), .B(n17), .Y(empty) );
    or2b2 U30 ( .A(rstN), .B(ldN_even), .Y(N75) );
    or3c2 U31 ( .A(rstN), .B(n7), .C(ldN_even_dly), .Y(N77) );
    or3c2 U32 ( .A(rstN), .B(n14), .C(ldN_odd_dly), .Y(N78) );
    or3c2 U33 ( .A(out_sel_odd_evenN), .B(N66), .C(rdN), .Y(n20) );
    or3c2 U34 ( .A(n17), .B(mem_empty_odd_dly), .C(mem_empty_odd), .Y(n13) );
    or3c2 U35 ( .A(n24), .B(mem_empty_even_dly), .C(mem_empty_even), .Y(n12)
         );
    or2b2 U36 ( .A(out_sel_odd_evenN), .B(rdN), .Y(n21) );
    or2b2 U37 ( .A(N5), .B(rdN), .Y(n22) );
endmodule


module ram16X8_0 ( data, addr, oe, wrN, clk );
inout  [7:0] data;
input  [3:0] addr;
input  oe, wrN, clk;
    wire \ram0[7] , \ram0[6] , \ram0[5] , \ram0[4] , \ram0[3] , \ram0[2] , 
        \ram0[1] , \ram0[0] , \ram1[7] , \ram1[6] , \ram1[5] , \ram1[4] , 
        \ram1[3] , \ram1[2] , \ram1[1] , \ram1[0] , \ram2[7] , \ram2[6] , 
        \ram2[5] , \ram2[4] , \ram2[3] , \ram2[2] , \ram2[1] , \ram2[0] , 
        \ram3[7] , \ram3[6] , \ram3[5] , \ram3[4] , \ram3[3] , \ram3[2] , 
        \ram3[1] , \ram3[0] , \ram4[7] , \ram4[6] , \ram4[5] , \ram4[4] , 
        \ram4[3] , \ram4[2] , \ram4[1] , \ram4[0] , \ram5[7] , \ram5[6] , 
        \ram5[5] , \ram5[4] , \ram5[3] , \ram5[2] , \ram5[1] , \ram5[0] , 
        \ram6[7] , \ram6[6] , \ram6[5] , \ram6[4] , \ram6[3] , \ram6[2] , 
        \ram6[1] , \ram6[0] , \ram7[7] , \ram7[6] , \ram7[5] , \ram7[4] , 
        \ram7[3] , \ram7[2] , \ram7[1] , \ram7[0] , \ram8[7] , \ram8[6] , 
        \ram8[5] , \ram8[4] , \ram8[3] , \ram8[2] , \ram8[1] , \ram8[0] , 
        \ram9[7] , \ram9[6] , \ram9[5] , \ram9[4] , \ram9[3] , \ram9[2] , 
        \ram9[1] , \ram9[0] , \ram10[7] , \ram10[6] , \ram10[5] , \ram10[4] , 
        \ram10[3] , \ram10[2] , \ram10[1] , \ram10[0] , \ram11[7] , \ram11[6] , 
        \ram11[5] , \ram11[4] , \ram11[3] , \ram11[2] , \ram11[1] , \ram11[0] , 
        \ram12[7] , \ram12[6] , \ram12[5] , \ram12[4] , \ram12[3] , \ram12[2] , 
        \ram12[1] , \ram12[0] , \ram13[7] , \ram13[6] , \ram13[5] , \ram13[4] , 
        \ram13[3] , \ram13[2] , \ram13[1] , \ram13[0] , \ram14[7] , \ram14[6] , 
        \ram14[5] , \ram14[4] , \ram14[3] , \ram14[2] , \ram14[1] , \ram14[0] , 
        \ram15[7] , \ram15[6] , \ram15[5] , \ram15[4] , \ram15[3] , \ram15[2] , 
        \ram15[1] , \ram15[0] , N353, N369, N385, N401, N417, N433, N449, N465, 
        N481, N497, N513, N529, N545, N561, N577, N593, n25, n26, n27, n28, 
        n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        n43, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
        n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, 
        n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
        n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
        n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
        n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176;
    tri \_0_ca_[7] , \_0_ca_[6] , \_0_ca_[5] , \_0_ca_[4] , \_0_ca_[3] , 
        \_0_ca_[2] , \_0_ca_[1] , \_0_ca_[0] ;
    tran( \_0_ca_[7] , data[7] );
    tran( \_0_ca_[6] , data[6] );
    tran( \_0_ca_[5] , data[5] );
    tran( \_0_ca_[4] , data[4] );
    tran( \_0_ca_[3] , data[3] );
    tran( \_0_ca_[2] , data[2] );
    tran( \_0_ca_[1] , data[1] );
    tran( \_0_ca_[0] , data[0] );
    inv1a1 U3 ( .A(addr[0]), .Y(n142) );
    ao1d2 U4 ( .A(n126), .B(n125), .C(n147), .Y(n28) );
    ao1d2 U5 ( .A(n128), .B(n127), .C(n151), .Y(n27) );
    ao1d2 U6 ( .A(n130), .B(n129), .C(n149), .Y(n26) );
    ao1d2 U7 ( .A(n132), .B(n131), .C(n153), .Y(n25) );
    ao1d2 U8 ( .A(n118), .B(n117), .C(n147), .Y(n32) );
    ao1d2 U9 ( .A(n120), .B(n119), .C(n151), .Y(n31) );
    ao1d2 U10 ( .A(n122), .B(n121), .C(n149), .Y(n30) );
    ao1d2 U11 ( .A(n124), .B(n123), .C(n153), .Y(n29) );
    ao1d2 U12 ( .A(n110), .B(n109), .C(n147), .Y(n36) );
    ao1d2 U13 ( .A(n112), .B(n111), .C(n151), .Y(n35) );
    ao1d2 U14 ( .A(n114), .B(n113), .C(n149), .Y(n34) );
    ao1d2 U15 ( .A(n116), .B(n115), .C(n153), .Y(n33) );
    ao1d2 U16 ( .A(n102), .B(n101), .C(n147), .Y(n40) );
    ao1d2 U17 ( .A(n104), .B(n103), .C(n151), .Y(n39) );
    ao1d2 U18 ( .A(n106), .B(n105), .C(n149), .Y(n38) );
    ao1d2 U19 ( .A(n108), .B(n107), .C(n153), .Y(n37) );
    ao1d2 U20 ( .A(n94), .B(n93), .C(n147), .Y(n51) );
    ao1d2 U21 ( .A(n96), .B(n95), .C(n151), .Y(n43) );
    ao1d2 U22 ( .A(n98), .B(n97), .C(n149), .Y(n42) );
    ao1d2 U23 ( .A(n100), .B(n99), .C(n153), .Y(n41) );
    ao1d2 U24 ( .A(n86), .B(n85), .C(n147), .Y(n55) );
    ao1d2 U25 ( .A(n88), .B(n87), .C(n151), .Y(n54) );
    ao1d2 U26 ( .A(n90), .B(n89), .C(n149), .Y(n53) );
    ao1d2 U27 ( .A(n92), .B(n91), .C(n153), .Y(n52) );
    ao1d2 U28 ( .A(n78), .B(n77), .C(n147), .Y(n59) );
    ao1d2 U29 ( .A(n80), .B(n79), .C(n151), .Y(n58) );
    ao1d2 U30 ( .A(n82), .B(n81), .C(n149), .Y(n57) );
    ao1d2 U31 ( .A(n84), .B(n83), .C(n153), .Y(n56) );
    ao1d2 U32 ( .A(n70), .B(n69), .C(n147), .Y(n63) );
    clk1b6 U33 ( .A(n65), .Y(n147) );
    ao1d2 U34 ( .A(n72), .B(n71), .C(n151), .Y(n62) );
    clk1b6 U35 ( .A(n66), .Y(n151) );
    ao1d2 U36 ( .A(n74), .B(n73), .C(n149), .Y(n61) );
    clk1b6 U37 ( .A(n67), .Y(n149) );
    ao1d2 U38 ( .A(n76), .B(n75), .C(n153), .Y(n60) );
    clk1b6 U39 ( .A(n68), .Y(n153) );
    or2b2 U40 ( .A(n64), .B(addr[2]), .Y(n68) );
    inv1a1 U41 ( .A(addr[3]), .Y(n64) );
    inv1a3 U42 ( .A(n148), .Y(n169) );
    inv1a3 U43 ( .A(n150), .Y(n164) );
    inv1a3 U44 ( .A(n152), .Y(n159) );
    clk1b15 U45 ( .A(n145), .Y(n157) );
    clk1b15 U46 ( .A(n141), .Y(n154) );
    clk1b15 U47 ( .A(n143), .Y(n155) );
    clk1b15 U48 ( .A(n144), .Y(n156) );
    fdef1a3 \ram11_reg[0]  ( .D(\_0_ca_[0] ), .E(N529), .CLK(clk), .Q(
        \ram11[0] ) );
    fdef1a3 \ram11_reg[1]  ( .D(\_0_ca_[1] ), .E(N529), .CLK(clk), .Q(
        \ram11[1] ) );
    fdef1a3 \ram11_reg[2]  ( .D(\_0_ca_[2] ), .E(N529), .CLK(clk), .Q(
        \ram11[2] ) );
    fdef1a3 \ram11_reg[3]  ( .D(\_0_ca_[3] ), .E(N529), .CLK(clk), .Q(
        \ram11[3] ) );
    fdef1a3 \ram11_reg[4]  ( .D(\_0_ca_[4] ), .E(N529), .CLK(clk), .Q(
        \ram11[4] ) );
    fdef1a3 \ram11_reg[5]  ( .D(\_0_ca_[5] ), .E(N529), .CLK(clk), .Q(
        \ram11[5] ) );
    fdef1a3 \ram11_reg[6]  ( .D(\_0_ca_[6] ), .E(N529), .CLK(clk), .Q(
        \ram11[6] ) );
    fdef1a3 \ram11_reg[7]  ( .D(\_0_ca_[7] ), .E(N529), .CLK(clk), .Q(
        \ram11[7] ) );
    fdef1a3 \ram10_reg[0]  ( .D(\_0_ca_[0] ), .E(N513), .CLK(clk), .Q(
        \ram10[0] ) );
    fdef1a3 \ram10_reg[1]  ( .D(\_0_ca_[1] ), .E(N513), .CLK(clk), .Q(
        \ram10[1] ) );
    fdef1a3 \ram10_reg[2]  ( .D(\_0_ca_[2] ), .E(N513), .CLK(clk), .Q(
        \ram10[2] ) );
    fdef1a3 \ram10_reg[3]  ( .D(\_0_ca_[3] ), .E(N513), .CLK(clk), .Q(
        \ram10[3] ) );
    fdef1a3 \ram10_reg[4]  ( .D(\_0_ca_[4] ), .E(N513), .CLK(clk), .Q(
        \ram10[4] ) );
    fdef1a3 \ram10_reg[5]  ( .D(\_0_ca_[5] ), .E(N513), .CLK(clk), .Q(
        \ram10[5] ) );
    fdef1a3 \ram10_reg[6]  ( .D(\_0_ca_[6] ), .E(N513), .CLK(clk), .Q(
        \ram10[6] ) );
    fdef1a3 \ram10_reg[7]  ( .D(\_0_ca_[7] ), .E(N513), .CLK(clk), .Q(
        \ram10[7] ) );
    fdef1a3 \ram9_reg[0]  ( .D(\_0_ca_[0] ), .E(N497), .CLK(clk), .Q(\ram9[0] 
        ) );
    fdef1a3 \ram9_reg[1]  ( .D(\_0_ca_[1] ), .E(N497), .CLK(clk), .Q(\ram9[1] 
        ) );
    fdef1a3 \ram9_reg[2]  ( .D(\_0_ca_[2] ), .E(N497), .CLK(clk), .Q(\ram9[2] 
        ) );
    fdef1a3 \ram9_reg[3]  ( .D(\_0_ca_[3] ), .E(N497), .CLK(clk), .Q(\ram9[3] 
        ) );
    fdef1a3 \ram9_reg[4]  ( .D(\_0_ca_[4] ), .E(N497), .CLK(clk), .Q(\ram9[4] 
        ) );
    fdef1a3 \ram9_reg[5]  ( .D(\_0_ca_[5] ), .E(N497), .CLK(clk), .Q(\ram9[5] 
        ) );
    fdef1a3 \ram9_reg[6]  ( .D(\_0_ca_[6] ), .E(N497), .CLK(clk), .Q(\ram9[6] 
        ) );
    fdef1a3 \ram9_reg[7]  ( .D(\_0_ca_[7] ), .E(N497), .CLK(clk), .Q(\ram9[7] 
        ) );
    fdef1a3 \ram8_reg[0]  ( .D(\_0_ca_[0] ), .E(N481), .CLK(clk), .Q(\ram8[0] 
        ) );
    fdef1a3 \ram8_reg[1]  ( .D(\_0_ca_[1] ), .E(N481), .CLK(clk), .Q(\ram8[1] 
        ) );
    fdef1a3 \ram8_reg[2]  ( .D(\_0_ca_[2] ), .E(N481), .CLK(clk), .Q(\ram8[2] 
        ) );
    fdef1a3 \ram8_reg[3]  ( .D(\_0_ca_[3] ), .E(N481), .CLK(clk), .Q(\ram8[3] 
        ) );
    fdef1a3 \ram8_reg[4]  ( .D(\_0_ca_[4] ), .E(N481), .CLK(clk), .Q(\ram8[4] 
        ) );
    fdef1a3 \ram8_reg[5]  ( .D(\_0_ca_[5] ), .E(N481), .CLK(clk), .Q(\ram8[5] 
        ) );
    fdef1a3 \ram8_reg[6]  ( .D(\_0_ca_[6] ), .E(N481), .CLK(clk), .Q(\ram8[6] 
        ) );
    fdef1a3 \ram8_reg[7]  ( .D(\_0_ca_[7] ), .E(N481), .CLK(clk), .Q(\ram8[7] 
        ) );
    fdef1a3 \ram7_reg[0]  ( .D(\_0_ca_[0] ), .E(N465), .CLK(clk), .Q(\ram7[0] 
        ) );
    fdef1a3 \ram7_reg[1]  ( .D(\_0_ca_[1] ), .E(N465), .CLK(clk), .Q(\ram7[1] 
        ) );
    fdef1a3 \ram7_reg[2]  ( .D(\_0_ca_[2] ), .E(N465), .CLK(clk), .Q(\ram7[2] 
        ) );
    fdef1a3 \ram7_reg[3]  ( .D(\_0_ca_[3] ), .E(N465), .CLK(clk), .Q(\ram7[3] 
        ) );
    fdef1a3 \ram7_reg[4]  ( .D(\_0_ca_[4] ), .E(N465), .CLK(clk), .Q(\ram7[4] 
        ) );
    fdef1a3 \ram7_reg[5]  ( .D(\_0_ca_[5] ), .E(N465), .CLK(clk), .Q(\ram7[5] 
        ) );
    fdef1a3 \ram7_reg[6]  ( .D(\_0_ca_[6] ), .E(N465), .CLK(clk), .Q(\ram7[6] 
        ) );
    fdef1a3 \ram7_reg[7]  ( .D(\_0_ca_[7] ), .E(N465), .CLK(clk), .Q(\ram7[7] 
        ) );
    fdef1a3 \ram6_reg[0]  ( .D(\_0_ca_[0] ), .E(N449), .CLK(clk), .Q(\ram6[0] 
        ) );
    fdef1a3 \ram6_reg[1]  ( .D(\_0_ca_[1] ), .E(N449), .CLK(clk), .Q(\ram6[1] 
        ) );
    fdef1a3 \ram6_reg[2]  ( .D(\_0_ca_[2] ), .E(N449), .CLK(clk), .Q(\ram6[2] 
        ) );
    fdef1a3 \ram6_reg[3]  ( .D(\_0_ca_[3] ), .E(N449), .CLK(clk), .Q(\ram6[3] 
        ) );
    fdef1a3 \ram6_reg[4]  ( .D(\_0_ca_[4] ), .E(N449), .CLK(clk), .Q(\ram6[4] 
        ) );
    fdef1a3 \ram6_reg[5]  ( .D(\_0_ca_[5] ), .E(N449), .CLK(clk), .Q(\ram6[5] 
        ) );
    fdef1a3 \ram6_reg[6]  ( .D(\_0_ca_[6] ), .E(N449), .CLK(clk), .Q(\ram6[6] 
        ) );
    fdef1a3 \ram6_reg[7]  ( .D(\_0_ca_[7] ), .E(N449), .CLK(clk), .Q(\ram6[7] 
        ) );
    fdef1a3 \ram5_reg[0]  ( .D(\_0_ca_[0] ), .E(N433), .CLK(clk), .Q(\ram5[0] 
        ) );
    fdef1a3 \ram5_reg[1]  ( .D(\_0_ca_[1] ), .E(N433), .CLK(clk), .Q(\ram5[1] 
        ) );
    fdef1a3 \ram5_reg[2]  ( .D(\_0_ca_[2] ), .E(N433), .CLK(clk), .Q(\ram5[2] 
        ) );
    fdef1a3 \ram5_reg[3]  ( .D(\_0_ca_[3] ), .E(N433), .CLK(clk), .Q(\ram5[3] 
        ) );
    fdef1a3 \ram5_reg[4]  ( .D(\_0_ca_[4] ), .E(N433), .CLK(clk), .Q(\ram5[4] 
        ) );
    fdef1a3 \ram5_reg[5]  ( .D(\_0_ca_[5] ), .E(N433), .CLK(clk), .Q(\ram5[5] 
        ) );
    fdef1a3 \ram5_reg[6]  ( .D(\_0_ca_[6] ), .E(N433), .CLK(clk), .Q(\ram5[6] 
        ) );
    fdef1a3 \ram5_reg[7]  ( .D(\_0_ca_[7] ), .E(N433), .CLK(clk), .Q(\ram5[7] 
        ) );
    fdef1a3 \ram4_reg[0]  ( .D(\_0_ca_[0] ), .E(N417), .CLK(clk), .Q(\ram4[0] 
        ) );
    fdef1a3 \ram4_reg[1]  ( .D(\_0_ca_[1] ), .E(N417), .CLK(clk), .Q(\ram4[1] 
        ) );
    fdef1a3 \ram4_reg[2]  ( .D(\_0_ca_[2] ), .E(N417), .CLK(clk), .Q(\ram4[2] 
        ) );
    fdef1a3 \ram4_reg[3]  ( .D(\_0_ca_[3] ), .E(N417), .CLK(clk), .Q(\ram4[3] 
        ) );
    fdef1a3 \ram4_reg[4]  ( .D(\_0_ca_[4] ), .E(N417), .CLK(clk), .Q(\ram4[4] 
        ) );
    fdef1a3 \ram4_reg[5]  ( .D(\_0_ca_[5] ), .E(N417), .CLK(clk), .Q(\ram4[5] 
        ) );
    fdef1a3 \ram4_reg[6]  ( .D(\_0_ca_[6] ), .E(N417), .CLK(clk), .Q(\ram4[6] 
        ) );
    fdef1a3 \ram4_reg[7]  ( .D(\_0_ca_[7] ), .E(N417), .CLK(clk), .Q(\ram4[7] 
        ) );
    fdef1a3 \ram3_reg[0]  ( .D(\_0_ca_[0] ), .E(N401), .CLK(clk), .Q(\ram3[0] 
        ) );
    fdef1a3 \ram3_reg[1]  ( .D(\_0_ca_[1] ), .E(N401), .CLK(clk), .Q(\ram3[1] 
        ) );
    fdef1a3 \ram3_reg[2]  ( .D(\_0_ca_[2] ), .E(N401), .CLK(clk), .Q(\ram3[2] 
        ) );
    fdef1a3 \ram3_reg[3]  ( .D(\_0_ca_[3] ), .E(N401), .CLK(clk), .Q(\ram3[3] 
        ) );
    fdef1a3 \ram3_reg[4]  ( .D(\_0_ca_[4] ), .E(N401), .CLK(clk), .Q(\ram3[4] 
        ) );
    fdef1a3 \ram3_reg[5]  ( .D(\_0_ca_[5] ), .E(N401), .CLK(clk), .Q(\ram3[5] 
        ) );
    fdef1a3 \ram3_reg[6]  ( .D(\_0_ca_[6] ), .E(N401), .CLK(clk), .Q(\ram3[6] 
        ) );
    fdef1a3 \ram3_reg[7]  ( .D(\_0_ca_[7] ), .E(N401), .CLK(clk), .Q(\ram3[7] 
        ) );
    fdef1a3 \ram2_reg[0]  ( .D(\_0_ca_[0] ), .E(N385), .CLK(clk), .Q(\ram2[0] 
        ) );
    fdef1a3 \ram2_reg[1]  ( .D(\_0_ca_[1] ), .E(N385), .CLK(clk), .Q(\ram2[1] 
        ) );
    fdef1a3 \ram2_reg[2]  ( .D(\_0_ca_[2] ), .E(N385), .CLK(clk), .Q(\ram2[2] 
        ) );
    fdef1a3 \ram2_reg[3]  ( .D(\_0_ca_[3] ), .E(N385), .CLK(clk), .Q(\ram2[3] 
        ) );
    fdef1a3 \ram2_reg[4]  ( .D(\_0_ca_[4] ), .E(N385), .CLK(clk), .Q(\ram2[4] 
        ) );
    fdef1a3 \ram2_reg[5]  ( .D(\_0_ca_[5] ), .E(N385), .CLK(clk), .Q(\ram2[5] 
        ) );
    fdef1a3 \ram2_reg[6]  ( .D(\_0_ca_[6] ), .E(N385), .CLK(clk), .Q(\ram2[6] 
        ) );
    fdef1a3 \ram2_reg[7]  ( .D(\_0_ca_[7] ), .E(N385), .CLK(clk), .Q(\ram2[7] 
        ) );
    fdef1a3 \ram1_reg[0]  ( .D(\_0_ca_[0] ), .E(N369), .CLK(clk), .Q(\ram1[0] 
        ) );
    fdef1a3 \ram1_reg[1]  ( .D(\_0_ca_[1] ), .E(N369), .CLK(clk), .Q(\ram1[1] 
        ) );
    fdef1a3 \ram1_reg[2]  ( .D(\_0_ca_[2] ), .E(N369), .CLK(clk), .Q(\ram1[2] 
        ) );
    fdef1a3 \ram1_reg[3]  ( .D(\_0_ca_[3] ), .E(N369), .CLK(clk), .Q(\ram1[3] 
        ) );
    fdef1a3 \ram1_reg[4]  ( .D(\_0_ca_[4] ), .E(N369), .CLK(clk), .Q(\ram1[4] 
        ) );
    fdef1a3 \ram1_reg[5]  ( .D(\_0_ca_[5] ), .E(N369), .CLK(clk), .Q(\ram1[5] 
        ) );
    fdef1a3 \ram1_reg[6]  ( .D(\_0_ca_[6] ), .E(N369), .CLK(clk), .Q(\ram1[6] 
        ) );
    fdef1a3 \ram1_reg[7]  ( .D(\_0_ca_[7] ), .E(N369), .CLK(clk), .Q(\ram1[7] 
        ) );
    fdef1a3 \ram0_reg[0]  ( .D(\_0_ca_[0] ), .E(N353), .CLK(clk), .Q(\ram0[0] 
        ) );
    fdef1a3 \ram0_reg[1]  ( .D(\_0_ca_[1] ), .E(N353), .CLK(clk), .Q(\ram0[1] 
        ) );
    fdef1a3 \ram0_reg[2]  ( .D(\_0_ca_[2] ), .E(N353), .CLK(clk), .Q(\ram0[2] 
        ) );
    fdef1a3 \ram0_reg[3]  ( .D(\_0_ca_[3] ), .E(N353), .CLK(clk), .Q(\ram0[3] 
        ) );
    fdef1a3 \ram0_reg[4]  ( .D(\_0_ca_[4] ), .E(N353), .CLK(clk), .Q(\ram0[4] 
        ) );
    fdef1a3 \ram0_reg[5]  ( .D(\_0_ca_[5] ), .E(N353), .CLK(clk), .Q(\ram0[5] 
        ) );
    fdef1a3 \ram0_reg[6]  ( .D(\_0_ca_[6] ), .E(N353), .CLK(clk), .Q(\ram0[6] 
        ) );
    fdef1a3 \ram0_reg[7]  ( .D(\_0_ca_[7] ), .E(N353), .CLK(clk), .Q(\ram0[7] 
        ) );
    fdef1a3 \ram15_reg[0]  ( .D(\_0_ca_[0] ), .E(N593), .CLK(clk), .Q(
        \ram15[0] ) );
    fdef1a3 \ram15_reg[1]  ( .D(\_0_ca_[1] ), .E(N593), .CLK(clk), .Q(
        \ram15[1] ) );
    fdef1a3 \ram15_reg[2]  ( .D(\_0_ca_[2] ), .E(N593), .CLK(clk), .Q(
        \ram15[2] ) );
    fdef1a3 \ram15_reg[3]  ( .D(\_0_ca_[3] ), .E(N593), .CLK(clk), .Q(
        \ram15[3] ) );
    fdef1a3 \ram15_reg[4]  ( .D(\_0_ca_[4] ), .E(N593), .CLK(clk), .Q(
        \ram15[4] ) );
    fdef1a3 \ram15_reg[5]  ( .D(\_0_ca_[5] ), .E(N593), .CLK(clk), .Q(
        \ram15[5] ) );
    fdef1a3 \ram15_reg[6]  ( .D(\_0_ca_[6] ), .E(N593), .CLK(clk), .Q(
        \ram15[6] ) );
    fdef1a3 \ram15_reg[7]  ( .D(\_0_ca_[7] ), .E(N593), .CLK(clk), .Q(
        \ram15[7] ) );
    fdef1a3 \ram12_reg[0]  ( .D(\_0_ca_[0] ), .E(N545), .CLK(clk), .Q(
        \ram12[0] ) );
    fdef1a3 \ram12_reg[1]  ( .D(\_0_ca_[1] ), .E(N545), .CLK(clk), .Q(
        \ram12[1] ) );
    fdef1a3 \ram12_reg[2]  ( .D(\_0_ca_[2] ), .E(N545), .CLK(clk), .Q(
        \ram12[2] ) );
    fdef1a3 \ram12_reg[3]  ( .D(\_0_ca_[3] ), .E(N545), .CLK(clk), .Q(
        \ram12[3] ) );
    fdef1a3 \ram12_reg[4]  ( .D(\_0_ca_[4] ), .E(N545), .CLK(clk), .Q(
        \ram12[4] ) );
    fdef1a3 \ram12_reg[5]  ( .D(\_0_ca_[5] ), .E(N545), .CLK(clk), .Q(
        \ram12[5] ) );
    fdef1a3 \ram12_reg[6]  ( .D(\_0_ca_[6] ), .E(N545), .CLK(clk), .Q(
        \ram12[6] ) );
    fdef1a3 \ram12_reg[7]  ( .D(\_0_ca_[7] ), .E(N545), .CLK(clk), .Q(
        \ram12[7] ) );
    fdef1a3 \ram13_reg[0]  ( .D(\_0_ca_[0] ), .E(N561), .CLK(clk), .Q(
        \ram13[0] ) );
    fdef1a3 \ram13_reg[1]  ( .D(\_0_ca_[1] ), .E(N561), .CLK(clk), .Q(
        \ram13[1] ) );
    fdef1a3 \ram13_reg[2]  ( .D(\_0_ca_[2] ), .E(N561), .CLK(clk), .Q(
        \ram13[2] ) );
    fdef1a3 \ram13_reg[3]  ( .D(\_0_ca_[3] ), .E(N561), .CLK(clk), .Q(
        \ram13[3] ) );
    fdef1a3 \ram13_reg[4]  ( .D(\_0_ca_[4] ), .E(N561), .CLK(clk), .Q(
        \ram13[4] ) );
    fdef1a3 \ram13_reg[5]  ( .D(\_0_ca_[5] ), .E(N561), .CLK(clk), .Q(
        \ram13[5] ) );
    fdef1a3 \ram13_reg[6]  ( .D(\_0_ca_[6] ), .E(N561), .CLK(clk), .Q(
        \ram13[6] ) );
    fdef1a3 \ram13_reg[7]  ( .D(\_0_ca_[7] ), .E(N561), .CLK(clk), .Q(
        \ram13[7] ) );
    fdef1a3 \ram14_reg[0]  ( .D(\_0_ca_[0] ), .E(N577), .CLK(clk), .Q(
        \ram14[0] ) );
    fdef1a3 \ram14_reg[1]  ( .D(\_0_ca_[1] ), .E(N577), .CLK(clk), .Q(
        \ram14[1] ) );
    fdef1a3 \ram14_reg[2]  ( .D(\_0_ca_[2] ), .E(N577), .CLK(clk), .Q(
        \ram14[2] ) );
    fdef1a3 \ram14_reg[3]  ( .D(\_0_ca_[3] ), .E(N577), .CLK(clk), .Q(
        \ram14[3] ) );
    fdef1a3 \ram14_reg[4]  ( .D(\_0_ca_[4] ), .E(N577), .CLK(clk), .Q(
        \ram14[4] ) );
    fdef1a3 \ram14_reg[5]  ( .D(\_0_ca_[5] ), .E(N577), .CLK(clk), .Q(
        \ram14[5] ) );
    fdef1a3 \ram14_reg[6]  ( .D(\_0_ca_[6] ), .E(N577), .CLK(clk), .Q(
        \ram14[6] ) );
    fdef1a3 \ram14_reg[7]  ( .D(\_0_ca_[7] ), .E(N577), .CLK(clk), .Q(
        \ram14[7] ) );
    tri1a15 \_0_ca__tri[7]  ( .A(n133), .E(oe), .Y(\_0_ca_[7] ) );
    tri1a15 \_0_ca__tri[6]  ( .A(n134), .E(oe), .Y(\_0_ca_[6] ) );
    tri1a15 \_0_ca__tri[5]  ( .A(n135), .E(oe), .Y(\_0_ca_[5] ) );
    tri1a15 \_0_ca__tri[4]  ( .A(n136), .E(oe), .Y(\_0_ca_[4] ) );
    tri1a15 \_0_ca__tri[3]  ( .A(n137), .E(oe), .Y(\_0_ca_[3] ) );
    tri1a15 \_0_ca__tri[2]  ( .A(n138), .E(oe), .Y(\_0_ca_[2] ) );
    tri1a15 \_0_ca__tri[1]  ( .A(n139), .E(oe), .Y(\_0_ca_[1] ) );
    tri1a15 \_0_ca__tri[0]  ( .A(n140), .E(oe), .Y(\_0_ca_[0] ) );
    or4e3 U49 ( .A(n25), .B(n26), .C(n27), .D(n28), .Y(n140) );
    or4e3 U50 ( .A(n29), .B(n30), .C(n31), .D(n32), .Y(n139) );
    or4e3 U51 ( .A(n33), .B(n34), .C(n35), .D(n36), .Y(n138) );
    or4e3 U52 ( .A(n37), .B(n38), .C(n39), .D(n40), .Y(n137) );
    or4e3 U53 ( .A(n41), .B(n42), .C(n43), .D(n51), .Y(n136) );
    or4e3 U54 ( .A(n52), .B(n53), .C(n54), .D(n55), .Y(n135) );
    or4e3 U55 ( .A(n56), .B(n57), .C(n58), .D(n59), .Y(n134) );
    or4e3 U56 ( .A(n60), .B(n61), .C(n62), .D(n63), .Y(n133) );
    or2b2 U57 ( .A(addr[2]), .B(n64), .Y(n65) );
    or2b2 U58 ( .A(addr[2]), .B(addr[3]), .Y(n66) );
    or2b2 U59 ( .A(addr[3]), .B(addr[2]), .Y(n67) );
    oa4f3 U60 ( .A(\ram15[7] ), .B(n157), .C(\ram14[7] ), .D(n156), .Y(n69) );
    oa4f3 U61 ( .A(\ram13[7] ), .B(n155), .C(\ram12[7] ), .D(n154), .Y(n70) );
    oa4f3 U62 ( .A(\ram7[7] ), .B(n157), .C(\ram6[7] ), .D(n156), .Y(n71) );
    oa4f3 U63 ( .A(\ram5[7] ), .B(n155), .C(\ram4[7] ), .D(n154), .Y(n72) );
    oa4f3 U64 ( .A(\ram11[7] ), .B(n157), .C(\ram10[7] ), .D(n156), .Y(n73) );
    oa4f3 U65 ( .A(\ram9[7] ), .B(n155), .C(\ram8[7] ), .D(n154), .Y(n74) );
    oa4f3 U66 ( .A(\ram3[7] ), .B(n157), .C(\ram2[7] ), .D(n156), .Y(n75) );
    oa4f3 U67 ( .A(\ram1[7] ), .B(n155), .C(\ram0[7] ), .D(n154), .Y(n76) );
    oa4f3 U68 ( .A(\ram15[6] ), .B(n157), .C(\ram14[6] ), .D(n156), .Y(n77) );
    oa4f3 U69 ( .A(\ram13[6] ), .B(n155), .C(\ram12[6] ), .D(n154), .Y(n78) );
    oa4f3 U70 ( .A(\ram7[6] ), .B(n157), .C(\ram6[6] ), .D(n156), .Y(n79) );
    oa4f3 U71 ( .A(\ram5[6] ), .B(n155), .C(\ram4[6] ), .D(n154), .Y(n80) );
    oa4f3 U72 ( .A(\ram11[6] ), .B(n157), .C(\ram10[6] ), .D(n156), .Y(n81) );
    oa4f3 U73 ( .A(\ram9[6] ), .B(n155), .C(\ram8[6] ), .D(n154), .Y(n82) );
    oa4f3 U74 ( .A(\ram3[6] ), .B(n157), .C(\ram2[6] ), .D(n156), .Y(n83) );
    oa4f3 U75 ( .A(\ram1[6] ), .B(n155), .C(\ram0[6] ), .D(n154), .Y(n84) );
    oa4f3 U76 ( .A(\ram15[5] ), .B(n157), .C(\ram14[5] ), .D(n156), .Y(n85) );
    oa4f3 U77 ( .A(\ram13[5] ), .B(n155), .C(\ram12[5] ), .D(n154), .Y(n86) );
    oa4f3 U78 ( .A(\ram7[5] ), .B(n157), .C(\ram6[5] ), .D(n156), .Y(n87) );
    oa4f3 U79 ( .A(\ram5[5] ), .B(n155), .C(\ram4[5] ), .D(n154), .Y(n88) );
    oa4f3 U80 ( .A(\ram11[5] ), .B(n157), .C(\ram10[5] ), .D(n156), .Y(n89) );
    oa4f3 U81 ( .A(\ram9[5] ), .B(n155), .C(\ram8[5] ), .D(n154), .Y(n90) );
    oa4f3 U82 ( .A(\ram3[5] ), .B(n157), .C(\ram2[5] ), .D(n156), .Y(n91) );
    oa4f3 U83 ( .A(\ram1[5] ), .B(n155), .C(\ram0[5] ), .D(n154), .Y(n92) );
    oa4f3 U84 ( .A(\ram15[4] ), .B(n157), .C(\ram14[4] ), .D(n156), .Y(n93) );
    oa4f3 U85 ( .A(\ram13[4] ), .B(n155), .C(\ram12[4] ), .D(n154), .Y(n94) );
    oa4f3 U86 ( .A(\ram7[4] ), .B(n157), .C(\ram6[4] ), .D(n156), .Y(n95) );
    oa4f3 U87 ( .A(\ram5[4] ), .B(n155), .C(\ram4[4] ), .D(n154), .Y(n96) );
    oa4f3 U88 ( .A(\ram11[4] ), .B(n157), .C(\ram10[4] ), .D(n156), .Y(n97) );
    oa4f3 U89 ( .A(\ram9[4] ), .B(n155), .C(\ram8[4] ), .D(n154), .Y(n98) );
    oa4f3 U90 ( .A(\ram3[4] ), .B(n157), .C(\ram2[4] ), .D(n156), .Y(n99) );
    oa4f3 U91 ( .A(\ram1[4] ), .B(n155), .C(\ram0[4] ), .D(n154), .Y(n100) );
    oa4f3 U92 ( .A(\ram15[3] ), .B(n157), .C(\ram14[3] ), .D(n156), .Y(n101)
         );
    oa4f3 U93 ( .A(\ram13[3] ), .B(n155), .C(\ram12[3] ), .D(n154), .Y(n102)
         );
    oa4f3 U94 ( .A(\ram7[3] ), .B(n157), .C(\ram6[3] ), .D(n156), .Y(n103) );
    oa4f3 U95 ( .A(\ram5[3] ), .B(n155), .C(\ram4[3] ), .D(n154), .Y(n104) );
    oa4f3 U96 ( .A(\ram11[3] ), .B(n157), .C(\ram10[3] ), .D(n156), .Y(n105)
         );
    oa4f3 U97 ( .A(\ram9[3] ), .B(n155), .C(\ram8[3] ), .D(n154), .Y(n106) );
    oa4f3 U98 ( .A(\ram3[3] ), .B(n157), .C(\ram2[3] ), .D(n156), .Y(n107) );
    oa4f3 U99 ( .A(\ram1[3] ), .B(n155), .C(\ram0[3] ), .D(n154), .Y(n108) );
    oa4f3 U100 ( .A(\ram15[2] ), .B(n157), .C(\ram14[2] ), .D(n156), .Y(n109)
         );
    oa4f3 U101 ( .A(\ram13[2] ), .B(n155), .C(\ram12[2] ), .D(n154), .Y(n110)
         );
    oa4f3 U102 ( .A(\ram7[2] ), .B(n157), .C(\ram6[2] ), .D(n156), .Y(n111) );
    oa4f3 U103 ( .A(\ram5[2] ), .B(n155), .C(\ram4[2] ), .D(n154), .Y(n112) );
    oa4f3 U104 ( .A(\ram11[2] ), .B(n157), .C(\ram10[2] ), .D(n156), .Y(n113)
         );
    oa4f3 U105 ( .A(\ram9[2] ), .B(n155), .C(\ram8[2] ), .D(n154), .Y(n114) );
    oa4f3 U106 ( .A(\ram3[2] ), .B(n157), .C(\ram2[2] ), .D(n156), .Y(n115) );
    oa4f3 U107 ( .A(\ram1[2] ), .B(n155), .C(\ram0[2] ), .D(n154), .Y(n116) );
    oa4f3 U108 ( .A(\ram15[1] ), .B(n157), .C(\ram14[1] ), .D(n156), .Y(n117)
         );
    oa4f3 U109 ( .A(\ram13[1] ), .B(n155), .C(\ram12[1] ), .D(n154), .Y(n118)
         );
    oa4f3 U110 ( .A(\ram7[1] ), .B(n157), .C(\ram6[1] ), .D(n156), .Y(n119) );
    oa4f3 U111 ( .A(\ram5[1] ), .B(n155), .C(\ram4[1] ), .D(n154), .Y(n120) );
    oa4f3 U112 ( .A(\ram11[1] ), .B(n157), .C(\ram10[1] ), .D(n156), .Y(n121)
         );
    oa4f3 U113 ( .A(\ram9[1] ), .B(n155), .C(\ram8[1] ), .D(n154), .Y(n122) );
    oa4f3 U114 ( .A(\ram3[1] ), .B(n157), .C(\ram2[1] ), .D(n156), .Y(n123) );
    oa4f3 U115 ( .A(\ram1[1] ), .B(n155), .C(\ram0[1] ), .D(n154), .Y(n124) );
    oa4f3 U116 ( .A(\ram15[0] ), .B(n157), .C(\ram14[0] ), .D(n156), .Y(n125)
         );
    oa4f3 U117 ( .A(\ram13[0] ), .B(n155), .C(\ram12[0] ), .D(n154), .Y(n126)
         );
    oa4f3 U118 ( .A(\ram7[0] ), .B(n157), .C(\ram6[0] ), .D(n156), .Y(n127) );
    oa4f3 U119 ( .A(\ram5[0] ), .B(n155), .C(\ram4[0] ), .D(n154), .Y(n128) );
    oa4f3 U120 ( .A(\ram11[0] ), .B(n157), .C(\ram10[0] ), .D(n156), .Y(n129)
         );
    oa4f3 U121 ( .A(\ram9[0] ), .B(n155), .C(\ram8[0] ), .D(n154), .Y(n130) );
    oa4f3 U122 ( .A(\ram3[0] ), .B(n157), .C(\ram2[0] ), .D(n156), .Y(n131) );
    oa4f3 U123 ( .A(\ram1[0] ), .B(n155), .C(\ram0[0] ), .D(n154), .Y(n132) );
    or2b2 U124 ( .A(n142), .B(addr[1]), .Y(n141) );
    or2b2 U125 ( .A(addr[0]), .B(addr[1]), .Y(n143) );
    or2b2 U126 ( .A(addr[1]), .B(addr[0]), .Y(n144) );
    or2b2 U127 ( .A(addr[1]), .B(n142), .Y(n145) );
    or2b2 U128 ( .A(n147), .B(wrN), .Y(n146) );
    or2b2 U129 ( .A(n149), .B(wrN), .Y(n148) );
    or2b2 U130 ( .A(n151), .B(wrN), .Y(n150) );
    or2b2 U131 ( .A(n153), .B(wrN), .Y(n152) );
    or2b2 U132 ( .A(n159), .B(n141), .Y(n158) );
    clk1b6 U133 ( .A(n158), .Y(N353) );
    or2b2 U134 ( .A(n159), .B(n143), .Y(n160) );
    clk1b6 U135 ( .A(n160), .Y(N369) );
    or2b2 U136 ( .A(n159), .B(n144), .Y(n161) );
    clk1b6 U137 ( .A(n161), .Y(N385) );
    or2b2 U138 ( .A(n159), .B(n145), .Y(n162) );
    clk1b6 U139 ( .A(n162), .Y(N401) );
    or2b2 U140 ( .A(n164), .B(n141), .Y(n163) );
    clk1b6 U141 ( .A(n163), .Y(N417) );
    or2b2 U142 ( .A(n164), .B(n143), .Y(n165) );
    clk1b6 U143 ( .A(n165), .Y(N433) );
    or2b2 U144 ( .A(n164), .B(n144), .Y(n166) );
    clk1b6 U145 ( .A(n166), .Y(N449) );
    or2b2 U146 ( .A(n164), .B(n145), .Y(n167) );
    clk1b6 U147 ( .A(n167), .Y(N465) );
    or2b2 U148 ( .A(n169), .B(n141), .Y(n168) );
    clk1b6 U149 ( .A(n168), .Y(N481) );
    or2b2 U150 ( .A(n169), .B(n143), .Y(n170) );
    clk1b6 U151 ( .A(n170), .Y(N497) );
    or2b2 U152 ( .A(n169), .B(n144), .Y(n171) );
    clk1b6 U153 ( .A(n171), .Y(N513) );
    or2b2 U154 ( .A(n169), .B(n145), .Y(n172) );
    clk1b6 U155 ( .A(n172), .Y(N529) );
    or2b2 U156 ( .A(n154), .B(n146), .Y(n173) );
    clk1b6 U157 ( .A(n173), .Y(N545) );
    or2b2 U158 ( .A(n155), .B(n146), .Y(n174) );
    clk1b6 U159 ( .A(n174), .Y(N561) );
    or2b2 U160 ( .A(n156), .B(n146), .Y(n175) );
    clk1b6 U161 ( .A(n175), .Y(N577) );
    or2b2 U162 ( .A(n157), .B(n146), .Y(n176) );
    clk1b6 U163 ( .A(n176), .Y(N593) );
endmodule


module fifo_mem_0_DW01_inc_5_1 ( A, SUM );
input  [4:0] A;
output [4:0] SUM;
    wire net4398, net4404, net4407;
    xor2a2 U5 ( .A(net4407), .B(A[4]), .Y(SUM[4]) );
    ha1a2 U6 ( .A(A[3]), .B(net4398), .S(SUM[3]), .CO(net4407) );
    ha1a2 U7 ( .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(net4404) );
    ha1a2 U8 ( .A(A[2]), .B(net4404), .S(SUM[2]), .CO(net4398) );
endmodule


module fifo_mem_0_DW01_inc_5_0 ( A, SUM );
input  [4:0] A;
output [4:0] SUM;
    wire net4379, net4385, net4388;
    xor2a2 U5 ( .A(net4388), .B(A[4]), .Y(SUM[4]) );
    ha1a2 U6 ( .A(A[3]), .B(net4379), .S(SUM[3]), .CO(net4388) );
    ha1a2 U7 ( .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(net4385) );
    ha1a2 U8 ( .A(A[2]), .B(net4385), .S(SUM[2]), .CO(net4379) );
endmodule


module fifo_mem_0_DW01_cmp6_5_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
input  [4:0] A;
input  [4:0] B;
input  TC;
output LT, GT, EQ, LE, GE, NE;
    wire n44, n45, n46, n47, n48, n49, n50;
    or2c1 U10 ( .A(n49), .B(n50), .Y(n45) );
    xor2b2 U11 ( .A(B[4]), .B(A[4]), .Y(n50) );
    or3d1 U12 ( .A(n46), .B(n47), .C(n48), .Y(n44) );
    xor2b2 U13 ( .A(B[1]), .B(A[1]), .Y(n46) );
    xor2b2 U14 ( .A(A[3]), .B(B[3]), .Y(n47) );
    xor2b2 U15 ( .A(B[2]), .B(A[2]), .Y(n48) );
    and2c3 U16 ( .A(n44), .B(n45), .Y(EQ) );
    xor2b2 U17 ( .A(A[0]), .B(B[0]), .Y(n49) );
endmodule


module fifo_mem_0 ( data, clk, rstN, wrN, rdN, empty, full );
inout  [7:0] data;
input  clk, rstN, wrN, rdN;
output empty, full;
    wire \addr[3] , \addr[1] , \addr[0] , \wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] , N10, N20, \rd_cntr[4] , 
        \rd_cntr[3] , \rd_cntr[2] , \rd_cntr[1] , \rd_cntr[0] , N47, N57, 
        \_que_1[2] , N87, N115, N116, N117, N118, N120, N121, N122, N123, n177, 
        n178, n179, n180, n181;
    tri \data[7] , \data[6] , \data[5] , \data[4] , \data[3] , \data[2] , 
        \data[1] , \data[0] ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 ;
    tran( \data[7] , data[7] );
    tran( \data[6] , data[6] );
    tran( \data[5] , data[5] );
    tran( \data[4] , data[4] );
    tran( \data[3] , data[3] );
    tran( \data[2] , data[2] );
    tran( \data[1] , data[1] );
    tran( \data[0] , data[0] );
    ram16X8_0 ram ( .data({\data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .addr({\addr[3] , 
        \_que_1[2] , \addr[1] , \addr[0] }), .oe(wrN), .wrN(wrN), .clk(clk) );
    mx2a3 U4 ( .D0(\wr_cntr[3] ), .D1(\rd_cntr[3] ), .S(wrN), .Y(\addr[3] ) );
    mx2a3 U5 ( .D0(\wr_cntr[2] ), .D1(\rd_cntr[2] ), .S(wrN), .Y(\_que_1[2] )
         );
    mx2d3 U6 ( .D0(N10), .D1(N47), .S(wrN), .Y(\addr[0] ) );
    mx2a3 U7 ( .D0(\wr_cntr[1] ), .D1(\rd_cntr[1] ), .S(wrN), .Y(\addr[1] ) );
    xor2a2 U8 ( .A(\wr_cntr[4] ), .B(\rd_cntr[4] ), .Y(n180) );
    xor2a2 U9 ( .A(N10), .B(wrN), .Y(n178) );
    and2b2 U10 ( .A(n179), .B(N87), .Y(empty) );
    xor2a2 U11 ( .A(\wr_cntr[4] ), .B(\rd_cntr[4] ), .Y(n179) );
    inv1a3 U12 ( .A(wrN), .Y(N20) );
    inv1a3 U13 ( .A(rdN), .Y(N57) );
    inv1a1 U14 ( .A(N87), .Y(n181) );
    inv1a3 U15 ( .A(\rd_cntr[0] ), .Y(N47) );
    fdef2a3 \rd_cntr_reg[1]  ( .D(N115), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[1] ) );
    fdef2a3 \rd_cntr_reg[2]  ( .D(N116), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[2] ) );
    fdef2a3 \rd_cntr_reg[3]  ( .D(N117), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[3] ) );
    fdef2a3 \rd_cntr_reg[4]  ( .D(N118), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[4] ) );
    fdef2a3 \wr_cntr_reg[1]  ( .D(N120), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[1] ) );
    fdef2a3 \wr_cntr_reg[2]  ( .D(N121), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[2] ) );
    fdef2a3 \wr_cntr_reg[3]  ( .D(N122), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[3] ) );
    fdef2a3 \wr_cntr_reg[4]  ( .D(N123), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[4] ) );
    xor2a2 U16 ( .A(N47), .B(rdN), .Y(n177) );
    fdf2a3 \rd_cntr_reg[0]  ( .D(n177), .CLK(clk), .CLR(rstN), .Q(\rd_cntr[0] 
        ) );
    inv1a3 U17 ( .A(\wr_cntr[0] ), .Y(N10) );
    fdf2a3 \wr_cntr_reg[0]  ( .D(n178), .CLK(clk), .CLR(rstN), .Q(\wr_cntr[0] 
        ) );
    fifo_mem_0_DW01_inc_5_1 C99 ( .A({\rd_cntr[4] , \rd_cntr[3] , \rd_cntr[2] , 
        \rd_cntr[1] , \rd_cntr[0] }), .SUM({N118, N117, N116, N115, 
        SYNOPSYS_UNCONNECTED_1}) );
    fifo_mem_0_DW01_inc_5_0 C101 ( .A({\wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] }), .SUM({N123, N122, N121, 
        N120, SYNOPSYS_UNCONNECTED_2}) );
    fifo_mem_0_DW01_cmp6_5_0 r292 ( .A({\wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] }), .B({\rd_cntr[4] , 
        \rd_cntr[3] , \rd_cntr[2] , \rd_cntr[1] , \rd_cntr[0] }), .TC(1'b0), 
        .EQ(N87) );
    and2b2 U18 ( .A(n181), .B(n180), .Y(full) );
endmodule


module ram16X8_1 ( data, addr, oe, wrN, clk );
inout  [7:0] data;
input  [3:0] addr;
input  oe, wrN, clk;
    wire \ram0[7] , \ram0[6] , \ram0[5] , \ram0[4] , \ram0[3] , \ram0[2] , 
        \ram0[1] , \ram0[0] , \ram1[7] , \ram1[6] , \ram1[5] , \ram1[4] , 
        \ram1[3] , \ram1[2] , \ram1[1] , \ram1[0] , \ram2[7] , \ram2[6] , 
        \ram2[5] , \ram2[4] , \ram2[3] , \ram2[2] , \ram2[1] , \ram2[0] , 
        \ram3[7] , \ram3[6] , \ram3[5] , \ram3[4] , \ram3[3] , \ram3[2] , 
        \ram3[1] , \ram3[0] , \ram4[7] , \ram4[6] , \ram4[5] , \ram4[4] , 
        \ram4[3] , \ram4[2] , \ram4[1] , \ram4[0] , \ram5[7] , \ram5[6] , 
        \ram5[5] , \ram5[4] , \ram5[3] , \ram5[2] , \ram5[1] , \ram5[0] , 
        \ram6[7] , \ram6[6] , \ram6[5] , \ram6[4] , \ram6[3] , \ram6[2] , 
        \ram6[1] , \ram6[0] , \ram7[7] , \ram7[6] , \ram7[5] , \ram7[4] , 
        \ram7[3] , \ram7[2] , \ram7[1] , \ram7[0] , \ram8[7] , \ram8[6] , 
        \ram8[5] , \ram8[4] , \ram8[3] , \ram8[2] , \ram8[1] , \ram8[0] , 
        \ram9[7] , \ram9[6] , \ram9[5] , \ram9[4] , \ram9[3] , \ram9[2] , 
        \ram9[1] , \ram9[0] , \ram10[7] , \ram10[6] , \ram10[5] , \ram10[4] , 
        \ram10[3] , \ram10[2] , \ram10[1] , \ram10[0] , \ram11[7] , \ram11[6] , 
        \ram11[5] , \ram11[4] , \ram11[3] , \ram11[2] , \ram11[1] , \ram11[0] , 
        \ram12[7] , \ram12[6] , \ram12[5] , \ram12[4] , \ram12[3] , \ram12[2] , 
        \ram12[1] , \ram12[0] , \ram13[7] , \ram13[6] , \ram13[5] , \ram13[4] , 
        \ram13[3] , \ram13[2] , \ram13[1] , \ram13[0] , \ram14[7] , \ram14[6] , 
        \ram14[5] , \ram14[4] , \ram14[3] , \ram14[2] , \ram14[1] , \ram14[0] , 
        \ram15[7] , \ram15[6] , \ram15[5] , \ram15[4] , \ram15[3] , \ram15[2] , 
        \ram15[1] , \ram15[0] , N353, N369, N385, N401, N417, N433, N449, N465, 
        N481, N497, N513, N529, N545, N561, N577, N593, n190, n191, n192, n193, 
        n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
        n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
        n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334;
    tri \_0_ca_[7] , \_0_ca_[6] , \_0_ca_[5] , \_0_ca_[4] , \_0_ca_[3] , 
        \_0_ca_[2] , \_0_ca_[1] , \_0_ca_[0] ;
    tran( \_0_ca_[7] , data[7] );
    tran( \_0_ca_[6] , data[6] );
    tran( \_0_ca_[5] , data[5] );
    tran( \_0_ca_[4] , data[4] );
    tran( \_0_ca_[3] , data[3] );
    tran( \_0_ca_[2] , data[2] );
    tran( \_0_ca_[1] , data[1] );
    tran( \_0_ca_[0] , data[0] );
    inv1a1 U3 ( .A(addr[0]), .Y(n300) );
    ao1d2 U4 ( .A(n284), .B(n283), .C(n305), .Y(n193) );
    ao1d2 U5 ( .A(n286), .B(n285), .C(n309), .Y(n192) );
    ao1d2 U6 ( .A(n288), .B(n287), .C(n307), .Y(n191) );
    ao1d2 U7 ( .A(n290), .B(n289), .C(n311), .Y(n190) );
    ao1d2 U8 ( .A(n276), .B(n275), .C(n305), .Y(n197) );
    ao1d2 U9 ( .A(n278), .B(n277), .C(n309), .Y(n196) );
    ao1d2 U10 ( .A(n280), .B(n279), .C(n307), .Y(n195) );
    ao1d2 U11 ( .A(n282), .B(n281), .C(n311), .Y(n194) );
    ao1d2 U12 ( .A(n268), .B(n267), .C(n305), .Y(n201) );
    ao1d2 U13 ( .A(n270), .B(n269), .C(n309), .Y(n200) );
    ao1d2 U14 ( .A(n272), .B(n271), .C(n307), .Y(n199) );
    ao1d2 U15 ( .A(n274), .B(n273), .C(n311), .Y(n198) );
    ao1d2 U16 ( .A(n260), .B(n259), .C(n305), .Y(n205) );
    ao1d2 U17 ( .A(n262), .B(n261), .C(n309), .Y(n204) );
    ao1d2 U18 ( .A(n264), .B(n263), .C(n307), .Y(n203) );
    ao1d2 U19 ( .A(n266), .B(n265), .C(n311), .Y(n202) );
    ao1d2 U20 ( .A(n252), .B(n251), .C(n305), .Y(n209) );
    ao1d2 U21 ( .A(n254), .B(n253), .C(n309), .Y(n208) );
    ao1d2 U22 ( .A(n256), .B(n255), .C(n307), .Y(n207) );
    ao1d2 U23 ( .A(n258), .B(n257), .C(n311), .Y(n206) );
    ao1d2 U24 ( .A(n244), .B(n243), .C(n305), .Y(n213) );
    ao1d2 U25 ( .A(n246), .B(n245), .C(n309), .Y(n212) );
    ao1d2 U26 ( .A(n248), .B(n247), .C(n307), .Y(n211) );
    ao1d2 U27 ( .A(n250), .B(n249), .C(n311), .Y(n210) );
    ao1d2 U28 ( .A(n236), .B(n235), .C(n305), .Y(n217) );
    ao1d2 U29 ( .A(n238), .B(n237), .C(n309), .Y(n216) );
    ao1d2 U30 ( .A(n240), .B(n239), .C(n307), .Y(n215) );
    ao1d2 U31 ( .A(n242), .B(n241), .C(n311), .Y(n214) );
    ao1d2 U32 ( .A(n228), .B(n227), .C(n305), .Y(n221) );
    clk1b6 U33 ( .A(n223), .Y(n305) );
    ao1d2 U34 ( .A(n230), .B(n229), .C(n309), .Y(n220) );
    clk1b6 U35 ( .A(n224), .Y(n309) );
    ao1d2 U36 ( .A(n232), .B(n231), .C(n307), .Y(n219) );
    clk1b6 U37 ( .A(n225), .Y(n307) );
    ao1d2 U38 ( .A(n234), .B(n233), .C(n311), .Y(n218) );
    clk1b6 U39 ( .A(n226), .Y(n311) );
    or2b2 U40 ( .A(n222), .B(addr[2]), .Y(n226) );
    inv1a1 U41 ( .A(addr[3]), .Y(n222) );
    inv1a3 U42 ( .A(n306), .Y(n327) );
    inv1a3 U43 ( .A(n308), .Y(n322) );
    inv1a3 U44 ( .A(n310), .Y(n317) );
    clk1b15 U45 ( .A(n303), .Y(n315) );
    clk1b15 U46 ( .A(n299), .Y(n312) );
    clk1b15 U47 ( .A(n301), .Y(n313) );
    clk1b15 U48 ( .A(n302), .Y(n314) );
    fdef1a3 \ram11_reg[0]  ( .D(\_0_ca_[0] ), .E(N529), .CLK(clk), .Q(
        \ram11[0] ) );
    fdef1a3 \ram11_reg[1]  ( .D(\_0_ca_[1] ), .E(N529), .CLK(clk), .Q(
        \ram11[1] ) );
    fdef1a3 \ram11_reg[2]  ( .D(\_0_ca_[2] ), .E(N529), .CLK(clk), .Q(
        \ram11[2] ) );
    fdef1a3 \ram11_reg[3]  ( .D(\_0_ca_[3] ), .E(N529), .CLK(clk), .Q(
        \ram11[3] ) );
    fdef1a3 \ram11_reg[4]  ( .D(\_0_ca_[4] ), .E(N529), .CLK(clk), .Q(
        \ram11[4] ) );
    fdef1a3 \ram11_reg[5]  ( .D(\_0_ca_[5] ), .E(N529), .CLK(clk), .Q(
        \ram11[5] ) );
    fdef1a3 \ram11_reg[6]  ( .D(\_0_ca_[6] ), .E(N529), .CLK(clk), .Q(
        \ram11[6] ) );
    fdef1a3 \ram11_reg[7]  ( .D(\_0_ca_[7] ), .E(N529), .CLK(clk), .Q(
        \ram11[7] ) );
    fdef1a3 \ram10_reg[0]  ( .D(\_0_ca_[0] ), .E(N513), .CLK(clk), .Q(
        \ram10[0] ) );
    fdef1a3 \ram10_reg[1]  ( .D(\_0_ca_[1] ), .E(N513), .CLK(clk), .Q(
        \ram10[1] ) );
    fdef1a3 \ram10_reg[2]  ( .D(\_0_ca_[2] ), .E(N513), .CLK(clk), .Q(
        \ram10[2] ) );
    fdef1a3 \ram10_reg[3]  ( .D(\_0_ca_[3] ), .E(N513), .CLK(clk), .Q(
        \ram10[3] ) );
    fdef1a3 \ram10_reg[4]  ( .D(\_0_ca_[4] ), .E(N513), .CLK(clk), .Q(
        \ram10[4] ) );
    fdef1a3 \ram10_reg[5]  ( .D(\_0_ca_[5] ), .E(N513), .CLK(clk), .Q(
        \ram10[5] ) );
    fdef1a3 \ram10_reg[6]  ( .D(\_0_ca_[6] ), .E(N513), .CLK(clk), .Q(
        \ram10[6] ) );
    fdef1a3 \ram10_reg[7]  ( .D(\_0_ca_[7] ), .E(N513), .CLK(clk), .Q(
        \ram10[7] ) );
    fdef1a3 \ram9_reg[0]  ( .D(\_0_ca_[0] ), .E(N497), .CLK(clk), .Q(\ram9[0] 
        ) );
    fdef1a3 \ram9_reg[1]  ( .D(\_0_ca_[1] ), .E(N497), .CLK(clk), .Q(\ram9[1] 
        ) );
    fdef1a3 \ram9_reg[2]  ( .D(\_0_ca_[2] ), .E(N497), .CLK(clk), .Q(\ram9[2] 
        ) );
    fdef1a3 \ram9_reg[3]  ( .D(\_0_ca_[3] ), .E(N497), .CLK(clk), .Q(\ram9[3] 
        ) );
    fdef1a3 \ram9_reg[4]  ( .D(\_0_ca_[4] ), .E(N497), .CLK(clk), .Q(\ram9[4] 
        ) );
    fdef1a3 \ram9_reg[5]  ( .D(\_0_ca_[5] ), .E(N497), .CLK(clk), .Q(\ram9[5] 
        ) );
    fdef1a3 \ram9_reg[6]  ( .D(\_0_ca_[6] ), .E(N497), .CLK(clk), .Q(\ram9[6] 
        ) );
    fdef1a3 \ram9_reg[7]  ( .D(\_0_ca_[7] ), .E(N497), .CLK(clk), .Q(\ram9[7] 
        ) );
    fdef1a3 \ram8_reg[0]  ( .D(\_0_ca_[0] ), .E(N481), .CLK(clk), .Q(\ram8[0] 
        ) );
    fdef1a3 \ram8_reg[1]  ( .D(\_0_ca_[1] ), .E(N481), .CLK(clk), .Q(\ram8[1] 
        ) );
    fdef1a3 \ram8_reg[2]  ( .D(\_0_ca_[2] ), .E(N481), .CLK(clk), .Q(\ram8[2] 
        ) );
    fdef1a3 \ram8_reg[3]  ( .D(\_0_ca_[3] ), .E(N481), .CLK(clk), .Q(\ram8[3] 
        ) );
    fdef1a3 \ram8_reg[4]  ( .D(\_0_ca_[4] ), .E(N481), .CLK(clk), .Q(\ram8[4] 
        ) );
    fdef1a3 \ram8_reg[5]  ( .D(\_0_ca_[5] ), .E(N481), .CLK(clk), .Q(\ram8[5] 
        ) );
    fdef1a3 \ram8_reg[6]  ( .D(\_0_ca_[6] ), .E(N481), .CLK(clk), .Q(\ram8[6] 
        ) );
    fdef1a3 \ram8_reg[7]  ( .D(\_0_ca_[7] ), .E(N481), .CLK(clk), .Q(\ram8[7] 
        ) );
    fdef1a3 \ram7_reg[0]  ( .D(\_0_ca_[0] ), .E(N465), .CLK(clk), .Q(\ram7[0] 
        ) );
    fdef1a3 \ram7_reg[1]  ( .D(\_0_ca_[1] ), .E(N465), .CLK(clk), .Q(\ram7[1] 
        ) );
    fdef1a3 \ram7_reg[2]  ( .D(\_0_ca_[2] ), .E(N465), .CLK(clk), .Q(\ram7[2] 
        ) );
    fdef1a3 \ram7_reg[3]  ( .D(\_0_ca_[3] ), .E(N465), .CLK(clk), .Q(\ram7[3] 
        ) );
    fdef1a3 \ram7_reg[4]  ( .D(\_0_ca_[4] ), .E(N465), .CLK(clk), .Q(\ram7[4] 
        ) );
    fdef1a3 \ram7_reg[5]  ( .D(\_0_ca_[5] ), .E(N465), .CLK(clk), .Q(\ram7[5] 
        ) );
    fdef1a3 \ram7_reg[6]  ( .D(\_0_ca_[6] ), .E(N465), .CLK(clk), .Q(\ram7[6] 
        ) );
    fdef1a3 \ram7_reg[7]  ( .D(\_0_ca_[7] ), .E(N465), .CLK(clk), .Q(\ram7[7] 
        ) );
    fdef1a3 \ram6_reg[0]  ( .D(\_0_ca_[0] ), .E(N449), .CLK(clk), .Q(\ram6[0] 
        ) );
    fdef1a3 \ram6_reg[1]  ( .D(\_0_ca_[1] ), .E(N449), .CLK(clk), .Q(\ram6[1] 
        ) );
    fdef1a3 \ram6_reg[2]  ( .D(\_0_ca_[2] ), .E(N449), .CLK(clk), .Q(\ram6[2] 
        ) );
    fdef1a3 \ram6_reg[3]  ( .D(\_0_ca_[3] ), .E(N449), .CLK(clk), .Q(\ram6[3] 
        ) );
    fdef1a3 \ram6_reg[4]  ( .D(\_0_ca_[4] ), .E(N449), .CLK(clk), .Q(\ram6[4] 
        ) );
    fdef1a3 \ram6_reg[5]  ( .D(\_0_ca_[5] ), .E(N449), .CLK(clk), .Q(\ram6[5] 
        ) );
    fdef1a3 \ram6_reg[6]  ( .D(\_0_ca_[6] ), .E(N449), .CLK(clk), .Q(\ram6[6] 
        ) );
    fdef1a3 \ram6_reg[7]  ( .D(\_0_ca_[7] ), .E(N449), .CLK(clk), .Q(\ram6[7] 
        ) );
    fdef1a3 \ram5_reg[0]  ( .D(\_0_ca_[0] ), .E(N433), .CLK(clk), .Q(\ram5[0] 
        ) );
    fdef1a3 \ram5_reg[1]  ( .D(\_0_ca_[1] ), .E(N433), .CLK(clk), .Q(\ram5[1] 
        ) );
    fdef1a3 \ram5_reg[2]  ( .D(\_0_ca_[2] ), .E(N433), .CLK(clk), .Q(\ram5[2] 
        ) );
    fdef1a3 \ram5_reg[3]  ( .D(\_0_ca_[3] ), .E(N433), .CLK(clk), .Q(\ram5[3] 
        ) );
    fdef1a3 \ram5_reg[4]  ( .D(\_0_ca_[4] ), .E(N433), .CLK(clk), .Q(\ram5[4] 
        ) );
    fdef1a3 \ram5_reg[5]  ( .D(\_0_ca_[5] ), .E(N433), .CLK(clk), .Q(\ram5[5] 
        ) );
    fdef1a3 \ram5_reg[6]  ( .D(\_0_ca_[6] ), .E(N433), .CLK(clk), .Q(\ram5[6] 
        ) );
    fdef1a3 \ram5_reg[7]  ( .D(\_0_ca_[7] ), .E(N433), .CLK(clk), .Q(\ram5[7] 
        ) );
    fdef1a3 \ram4_reg[0]  ( .D(\_0_ca_[0] ), .E(N417), .CLK(clk), .Q(\ram4[0] 
        ) );
    fdef1a3 \ram4_reg[1]  ( .D(\_0_ca_[1] ), .E(N417), .CLK(clk), .Q(\ram4[1] 
        ) );
    fdef1a3 \ram4_reg[2]  ( .D(\_0_ca_[2] ), .E(N417), .CLK(clk), .Q(\ram4[2] 
        ) );
    fdef1a3 \ram4_reg[3]  ( .D(\_0_ca_[3] ), .E(N417), .CLK(clk), .Q(\ram4[3] 
        ) );
    fdef1a3 \ram4_reg[4]  ( .D(\_0_ca_[4] ), .E(N417), .CLK(clk), .Q(\ram4[4] 
        ) );
    fdef1a3 \ram4_reg[5]  ( .D(\_0_ca_[5] ), .E(N417), .CLK(clk), .Q(\ram4[5] 
        ) );
    fdef1a3 \ram4_reg[6]  ( .D(\_0_ca_[6] ), .E(N417), .CLK(clk), .Q(\ram4[6] 
        ) );
    fdef1a3 \ram4_reg[7]  ( .D(\_0_ca_[7] ), .E(N417), .CLK(clk), .Q(\ram4[7] 
        ) );
    fdef1a3 \ram3_reg[0]  ( .D(\_0_ca_[0] ), .E(N401), .CLK(clk), .Q(\ram3[0] 
        ) );
    fdef1a3 \ram3_reg[1]  ( .D(\_0_ca_[1] ), .E(N401), .CLK(clk), .Q(\ram3[1] 
        ) );
    fdef1a3 \ram3_reg[2]  ( .D(\_0_ca_[2] ), .E(N401), .CLK(clk), .Q(\ram3[2] 
        ) );
    fdef1a3 \ram3_reg[3]  ( .D(\_0_ca_[3] ), .E(N401), .CLK(clk), .Q(\ram3[3] 
        ) );
    fdef1a3 \ram3_reg[4]  ( .D(\_0_ca_[4] ), .E(N401), .CLK(clk), .Q(\ram3[4] 
        ) );
    fdef1a3 \ram3_reg[5]  ( .D(\_0_ca_[5] ), .E(N401), .CLK(clk), .Q(\ram3[5] 
        ) );
    fdef1a3 \ram3_reg[6]  ( .D(\_0_ca_[6] ), .E(N401), .CLK(clk), .Q(\ram3[6] 
        ) );
    fdef1a3 \ram3_reg[7]  ( .D(\_0_ca_[7] ), .E(N401), .CLK(clk), .Q(\ram3[7] 
        ) );
    fdef1a3 \ram2_reg[0]  ( .D(\_0_ca_[0] ), .E(N385), .CLK(clk), .Q(\ram2[0] 
        ) );
    fdef1a3 \ram2_reg[1]  ( .D(\_0_ca_[1] ), .E(N385), .CLK(clk), .Q(\ram2[1] 
        ) );
    fdef1a3 \ram2_reg[2]  ( .D(\_0_ca_[2] ), .E(N385), .CLK(clk), .Q(\ram2[2] 
        ) );
    fdef1a3 \ram2_reg[3]  ( .D(\_0_ca_[3] ), .E(N385), .CLK(clk), .Q(\ram2[3] 
        ) );
    fdef1a3 \ram2_reg[4]  ( .D(\_0_ca_[4] ), .E(N385), .CLK(clk), .Q(\ram2[4] 
        ) );
    fdef1a3 \ram2_reg[5]  ( .D(\_0_ca_[5] ), .E(N385), .CLK(clk), .Q(\ram2[5] 
        ) );
    fdef1a3 \ram2_reg[6]  ( .D(\_0_ca_[6] ), .E(N385), .CLK(clk), .Q(\ram2[6] 
        ) );
    fdef1a3 \ram2_reg[7]  ( .D(\_0_ca_[7] ), .E(N385), .CLK(clk), .Q(\ram2[7] 
        ) );
    fdef1a3 \ram1_reg[0]  ( .D(\_0_ca_[0] ), .E(N369), .CLK(clk), .Q(\ram1[0] 
        ) );
    fdef1a3 \ram1_reg[1]  ( .D(\_0_ca_[1] ), .E(N369), .CLK(clk), .Q(\ram1[1] 
        ) );
    fdef1a3 \ram1_reg[2]  ( .D(\_0_ca_[2] ), .E(N369), .CLK(clk), .Q(\ram1[2] 
        ) );
    fdef1a3 \ram1_reg[3]  ( .D(\_0_ca_[3] ), .E(N369), .CLK(clk), .Q(\ram1[3] 
        ) );
    fdef1a3 \ram1_reg[4]  ( .D(\_0_ca_[4] ), .E(N369), .CLK(clk), .Q(\ram1[4] 
        ) );
    fdef1a3 \ram1_reg[5]  ( .D(\_0_ca_[5] ), .E(N369), .CLK(clk), .Q(\ram1[5] 
        ) );
    fdef1a3 \ram1_reg[6]  ( .D(\_0_ca_[6] ), .E(N369), .CLK(clk), .Q(\ram1[6] 
        ) );
    fdef1a3 \ram1_reg[7]  ( .D(\_0_ca_[7] ), .E(N369), .CLK(clk), .Q(\ram1[7] 
        ) );
    fdef1a3 \ram0_reg[0]  ( .D(\_0_ca_[0] ), .E(N353), .CLK(clk), .Q(\ram0[0] 
        ) );
    fdef1a3 \ram0_reg[1]  ( .D(\_0_ca_[1] ), .E(N353), .CLK(clk), .Q(\ram0[1] 
        ) );
    fdef1a3 \ram0_reg[2]  ( .D(\_0_ca_[2] ), .E(N353), .CLK(clk), .Q(\ram0[2] 
        ) );
    fdef1a3 \ram0_reg[3]  ( .D(\_0_ca_[3] ), .E(N353), .CLK(clk), .Q(\ram0[3] 
        ) );
    fdef1a3 \ram0_reg[4]  ( .D(\_0_ca_[4] ), .E(N353), .CLK(clk), .Q(\ram0[4] 
        ) );
    fdef1a3 \ram0_reg[5]  ( .D(\_0_ca_[5] ), .E(N353), .CLK(clk), .Q(\ram0[5] 
        ) );
    fdef1a3 \ram0_reg[6]  ( .D(\_0_ca_[6] ), .E(N353), .CLK(clk), .Q(\ram0[6] 
        ) );
    fdef1a3 \ram0_reg[7]  ( .D(\_0_ca_[7] ), .E(N353), .CLK(clk), .Q(\ram0[7] 
        ) );
    fdef1a3 \ram15_reg[0]  ( .D(\_0_ca_[0] ), .E(N593), .CLK(clk), .Q(
        \ram15[0] ) );
    fdef1a3 \ram15_reg[1]  ( .D(\_0_ca_[1] ), .E(N593), .CLK(clk), .Q(
        \ram15[1] ) );
    fdef1a3 \ram15_reg[2]  ( .D(\_0_ca_[2] ), .E(N593), .CLK(clk), .Q(
        \ram15[2] ) );
    fdef1a3 \ram15_reg[3]  ( .D(\_0_ca_[3] ), .E(N593), .CLK(clk), .Q(
        \ram15[3] ) );
    fdef1a3 \ram15_reg[4]  ( .D(\_0_ca_[4] ), .E(N593), .CLK(clk), .Q(
        \ram15[4] ) );
    fdef1a3 \ram15_reg[5]  ( .D(\_0_ca_[5] ), .E(N593), .CLK(clk), .Q(
        \ram15[5] ) );
    fdef1a3 \ram15_reg[6]  ( .D(\_0_ca_[6] ), .E(N593), .CLK(clk), .Q(
        \ram15[6] ) );
    fdef1a3 \ram15_reg[7]  ( .D(\_0_ca_[7] ), .E(N593), .CLK(clk), .Q(
        \ram15[7] ) );
    fdef1a3 \ram12_reg[0]  ( .D(\_0_ca_[0] ), .E(N545), .CLK(clk), .Q(
        \ram12[0] ) );
    fdef1a3 \ram12_reg[1]  ( .D(\_0_ca_[1] ), .E(N545), .CLK(clk), .Q(
        \ram12[1] ) );
    fdef1a3 \ram12_reg[2]  ( .D(\_0_ca_[2] ), .E(N545), .CLK(clk), .Q(
        \ram12[2] ) );
    fdef1a3 \ram12_reg[3]  ( .D(\_0_ca_[3] ), .E(N545), .CLK(clk), .Q(
        \ram12[3] ) );
    fdef1a3 \ram12_reg[4]  ( .D(\_0_ca_[4] ), .E(N545), .CLK(clk), .Q(
        \ram12[4] ) );
    fdef1a3 \ram12_reg[5]  ( .D(\_0_ca_[5] ), .E(N545), .CLK(clk), .Q(
        \ram12[5] ) );
    fdef1a3 \ram12_reg[6]  ( .D(\_0_ca_[6] ), .E(N545), .CLK(clk), .Q(
        \ram12[6] ) );
    fdef1a3 \ram12_reg[7]  ( .D(\_0_ca_[7] ), .E(N545), .CLK(clk), .Q(
        \ram12[7] ) );
    fdef1a3 \ram13_reg[0]  ( .D(\_0_ca_[0] ), .E(N561), .CLK(clk), .Q(
        \ram13[0] ) );
    fdef1a3 \ram13_reg[1]  ( .D(\_0_ca_[1] ), .E(N561), .CLK(clk), .Q(
        \ram13[1] ) );
    fdef1a3 \ram13_reg[2]  ( .D(\_0_ca_[2] ), .E(N561), .CLK(clk), .Q(
        \ram13[2] ) );
    fdef1a3 \ram13_reg[3]  ( .D(\_0_ca_[3] ), .E(N561), .CLK(clk), .Q(
        \ram13[3] ) );
    fdef1a3 \ram13_reg[4]  ( .D(\_0_ca_[4] ), .E(N561), .CLK(clk), .Q(
        \ram13[4] ) );
    fdef1a3 \ram13_reg[5]  ( .D(\_0_ca_[5] ), .E(N561), .CLK(clk), .Q(
        \ram13[5] ) );
    fdef1a3 \ram13_reg[6]  ( .D(\_0_ca_[6] ), .E(N561), .CLK(clk), .Q(
        \ram13[6] ) );
    fdef1a3 \ram13_reg[7]  ( .D(\_0_ca_[7] ), .E(N561), .CLK(clk), .Q(
        \ram13[7] ) );
    fdef1a3 \ram14_reg[0]  ( .D(\_0_ca_[0] ), .E(N577), .CLK(clk), .Q(
        \ram14[0] ) );
    fdef1a3 \ram14_reg[1]  ( .D(\_0_ca_[1] ), .E(N577), .CLK(clk), .Q(
        \ram14[1] ) );
    fdef1a3 \ram14_reg[2]  ( .D(\_0_ca_[2] ), .E(N577), .CLK(clk), .Q(
        \ram14[2] ) );
    fdef1a3 \ram14_reg[3]  ( .D(\_0_ca_[3] ), .E(N577), .CLK(clk), .Q(
        \ram14[3] ) );
    fdef1a3 \ram14_reg[4]  ( .D(\_0_ca_[4] ), .E(N577), .CLK(clk), .Q(
        \ram14[4] ) );
    fdef1a3 \ram14_reg[5]  ( .D(\_0_ca_[5] ), .E(N577), .CLK(clk), .Q(
        \ram14[5] ) );
    fdef1a3 \ram14_reg[6]  ( .D(\_0_ca_[6] ), .E(N577), .CLK(clk), .Q(
        \ram14[6] ) );
    fdef1a3 \ram14_reg[7]  ( .D(\_0_ca_[7] ), .E(N577), .CLK(clk), .Q(
        \ram14[7] ) );
    tri1a15 \_0_ca__tri[0]  ( .A(n298), .E(oe), .Y(\_0_ca_[0] ) );
    tri1a15 \_0_ca__tri[1]  ( .A(n297), .E(oe), .Y(\_0_ca_[1] ) );
    tri1a15 \_0_ca__tri[2]  ( .A(n296), .E(oe), .Y(\_0_ca_[2] ) );
    tri1a15 \_0_ca__tri[3]  ( .A(n295), .E(oe), .Y(\_0_ca_[3] ) );
    tri1a15 \_0_ca__tri[4]  ( .A(n294), .E(oe), .Y(\_0_ca_[4] ) );
    tri1a15 \_0_ca__tri[5]  ( .A(n293), .E(oe), .Y(\_0_ca_[5] ) );
    tri1a15 \_0_ca__tri[6]  ( .A(n292), .E(oe), .Y(\_0_ca_[6] ) );
    tri1a15 \_0_ca__tri[7]  ( .A(n291), .E(oe), .Y(\_0_ca_[7] ) );
    or4e3 U49 ( .A(n190), .B(n191), .C(n192), .D(n193), .Y(n298) );
    or4e3 U50 ( .A(n194), .B(n195), .C(n196), .D(n197), .Y(n297) );
    or4e3 U51 ( .A(n198), .B(n199), .C(n200), .D(n201), .Y(n296) );
    or4e3 U52 ( .A(n202), .B(n203), .C(n204), .D(n205), .Y(n295) );
    or4e3 U53 ( .A(n206), .B(n207), .C(n208), .D(n209), .Y(n294) );
    or4e3 U54 ( .A(n210), .B(n211), .C(n212), .D(n213), .Y(n293) );
    or4e3 U55 ( .A(n214), .B(n215), .C(n216), .D(n217), .Y(n292) );
    or4e3 U56 ( .A(n218), .B(n219), .C(n220), .D(n221), .Y(n291) );
    or2b2 U57 ( .A(addr[2]), .B(n222), .Y(n223) );
    or2b2 U58 ( .A(addr[2]), .B(addr[3]), .Y(n224) );
    or2b2 U59 ( .A(addr[3]), .B(addr[2]), .Y(n225) );
    oa4f3 U60 ( .A(\ram15[7] ), .B(n315), .C(\ram14[7] ), .D(n314), .Y(n227)
         );
    oa4f3 U61 ( .A(\ram13[7] ), .B(n313), .C(\ram12[7] ), .D(n312), .Y(n228)
         );
    oa4f3 U62 ( .A(\ram7[7] ), .B(n315), .C(\ram6[7] ), .D(n314), .Y(n229) );
    oa4f3 U63 ( .A(\ram5[7] ), .B(n313), .C(\ram4[7] ), .D(n312), .Y(n230) );
    oa4f3 U64 ( .A(\ram11[7] ), .B(n315), .C(\ram10[7] ), .D(n314), .Y(n231)
         );
    oa4f3 U65 ( .A(\ram9[7] ), .B(n313), .C(\ram8[7] ), .D(n312), .Y(n232) );
    oa4f3 U66 ( .A(\ram3[7] ), .B(n315), .C(\ram2[7] ), .D(n314), .Y(n233) );
    oa4f3 U67 ( .A(\ram1[7] ), .B(n313), .C(\ram0[7] ), .D(n312), .Y(n234) );
    oa4f3 U68 ( .A(\ram15[6] ), .B(n315), .C(\ram14[6] ), .D(n314), .Y(n235)
         );
    oa4f3 U69 ( .A(\ram13[6] ), .B(n313), .C(\ram12[6] ), .D(n312), .Y(n236)
         );
    oa4f3 U70 ( .A(\ram7[6] ), .B(n315), .C(\ram6[6] ), .D(n314), .Y(n237) );
    oa4f3 U71 ( .A(\ram5[6] ), .B(n313), .C(\ram4[6] ), .D(n312), .Y(n238) );
    oa4f3 U72 ( .A(\ram11[6] ), .B(n315), .C(\ram10[6] ), .D(n314), .Y(n239)
         );
    oa4f3 U73 ( .A(\ram9[6] ), .B(n313), .C(\ram8[6] ), .D(n312), .Y(n240) );
    oa4f3 U74 ( .A(\ram3[6] ), .B(n315), .C(\ram2[6] ), .D(n314), .Y(n241) );
    oa4f3 U75 ( .A(\ram1[6] ), .B(n313), .C(\ram0[6] ), .D(n312), .Y(n242) );
    oa4f3 U76 ( .A(\ram15[5] ), .B(n315), .C(\ram14[5] ), .D(n314), .Y(n243)
         );
    oa4f3 U77 ( .A(\ram13[5] ), .B(n313), .C(\ram12[5] ), .D(n312), .Y(n244)
         );
    oa4f3 U78 ( .A(\ram7[5] ), .B(n315), .C(\ram6[5] ), .D(n314), .Y(n245) );
    oa4f3 U79 ( .A(\ram5[5] ), .B(n313), .C(\ram4[5] ), .D(n312), .Y(n246) );
    oa4f3 U80 ( .A(\ram11[5] ), .B(n315), .C(\ram10[5] ), .D(n314), .Y(n247)
         );
    oa4f3 U81 ( .A(\ram9[5] ), .B(n313), .C(\ram8[5] ), .D(n312), .Y(n248) );
    oa4f3 U82 ( .A(\ram3[5] ), .B(n315), .C(\ram2[5] ), .D(n314), .Y(n249) );
    oa4f3 U83 ( .A(\ram1[5] ), .B(n313), .C(\ram0[5] ), .D(n312), .Y(n250) );
    oa4f3 U84 ( .A(\ram15[4] ), .B(n315), .C(\ram14[4] ), .D(n314), .Y(n251)
         );
    oa4f3 U85 ( .A(\ram13[4] ), .B(n313), .C(\ram12[4] ), .D(n312), .Y(n252)
         );
    oa4f3 U86 ( .A(\ram7[4] ), .B(n315), .C(\ram6[4] ), .D(n314), .Y(n253) );
    oa4f3 U87 ( .A(\ram5[4] ), .B(n313), .C(\ram4[4] ), .D(n312), .Y(n254) );
    oa4f3 U88 ( .A(\ram11[4] ), .B(n315), .C(\ram10[4] ), .D(n314), .Y(n255)
         );
    oa4f3 U89 ( .A(\ram9[4] ), .B(n313), .C(\ram8[4] ), .D(n312), .Y(n256) );
    oa4f3 U90 ( .A(\ram3[4] ), .B(n315), .C(\ram2[4] ), .D(n314), .Y(n257) );
    oa4f3 U91 ( .A(\ram1[4] ), .B(n313), .C(\ram0[4] ), .D(n312), .Y(n258) );
    oa4f3 U92 ( .A(\ram15[3] ), .B(n315), .C(\ram14[3] ), .D(n314), .Y(n259)
         );
    oa4f3 U93 ( .A(\ram13[3] ), .B(n313), .C(\ram12[3] ), .D(n312), .Y(n260)
         );
    oa4f3 U94 ( .A(\ram7[3] ), .B(n315), .C(\ram6[3] ), .D(n314), .Y(n261) );
    oa4f3 U95 ( .A(\ram5[3] ), .B(n313), .C(\ram4[3] ), .D(n312), .Y(n262) );
    oa4f3 U96 ( .A(\ram11[3] ), .B(n315), .C(\ram10[3] ), .D(n314), .Y(n263)
         );
    oa4f3 U97 ( .A(\ram9[3] ), .B(n313), .C(\ram8[3] ), .D(n312), .Y(n264) );
    oa4f3 U98 ( .A(\ram3[3] ), .B(n315), .C(\ram2[3] ), .D(n314), .Y(n265) );
    oa4f3 U99 ( .A(\ram1[3] ), .B(n313), .C(\ram0[3] ), .D(n312), .Y(n266) );
    oa4f3 U100 ( .A(\ram15[2] ), .B(n315), .C(\ram14[2] ), .D(n314), .Y(n267)
         );
    oa4f3 U101 ( .A(\ram13[2] ), .B(n313), .C(\ram12[2] ), .D(n312), .Y(n268)
         );
    oa4f3 U102 ( .A(\ram7[2] ), .B(n315), .C(\ram6[2] ), .D(n314), .Y(n269) );
    oa4f3 U103 ( .A(\ram5[2] ), .B(n313), .C(\ram4[2] ), .D(n312), .Y(n270) );
    oa4f3 U104 ( .A(\ram11[2] ), .B(n315), .C(\ram10[2] ), .D(n314), .Y(n271)
         );
    oa4f3 U105 ( .A(\ram9[2] ), .B(n313), .C(\ram8[2] ), .D(n312), .Y(n272) );
    oa4f3 U106 ( .A(\ram3[2] ), .B(n315), .C(\ram2[2] ), .D(n314), .Y(n273) );
    oa4f3 U107 ( .A(\ram1[2] ), .B(n313), .C(\ram0[2] ), .D(n312), .Y(n274) );
    oa4f3 U108 ( .A(\ram15[1] ), .B(n315), .C(\ram14[1] ), .D(n314), .Y(n275)
         );
    oa4f3 U109 ( .A(\ram13[1] ), .B(n313), .C(\ram12[1] ), .D(n312), .Y(n276)
         );
    oa4f3 U110 ( .A(\ram7[1] ), .B(n315), .C(\ram6[1] ), .D(n314), .Y(n277) );
    oa4f3 U111 ( .A(\ram5[1] ), .B(n313), .C(\ram4[1] ), .D(n312), .Y(n278) );
    oa4f3 U112 ( .A(\ram11[1] ), .B(n315), .C(\ram10[1] ), .D(n314), .Y(n279)
         );
    oa4f3 U113 ( .A(\ram9[1] ), .B(n313), .C(\ram8[1] ), .D(n312), .Y(n280) );
    oa4f3 U114 ( .A(\ram3[1] ), .B(n315), .C(\ram2[1] ), .D(n314), .Y(n281) );
    oa4f3 U115 ( .A(\ram1[1] ), .B(n313), .C(\ram0[1] ), .D(n312), .Y(n282) );
    oa4f3 U116 ( .A(\ram15[0] ), .B(n315), .C(\ram14[0] ), .D(n314), .Y(n283)
         );
    oa4f3 U117 ( .A(\ram13[0] ), .B(n313), .C(\ram12[0] ), .D(n312), .Y(n284)
         );
    oa4f3 U118 ( .A(\ram7[0] ), .B(n315), .C(\ram6[0] ), .D(n314), .Y(n285) );
    oa4f3 U119 ( .A(\ram5[0] ), .B(n313), .C(\ram4[0] ), .D(n312), .Y(n286) );
    oa4f3 U120 ( .A(\ram11[0] ), .B(n315), .C(\ram10[0] ), .D(n314), .Y(n287)
         );
    oa4f3 U121 ( .A(\ram9[0] ), .B(n313), .C(\ram8[0] ), .D(n312), .Y(n288) );
    oa4f3 U122 ( .A(\ram3[0] ), .B(n315), .C(\ram2[0] ), .D(n314), .Y(n289) );
    oa4f3 U123 ( .A(\ram1[0] ), .B(n313), .C(\ram0[0] ), .D(n312), .Y(n290) );
    or2b2 U124 ( .A(n300), .B(addr[1]), .Y(n299) );
    or2b2 U125 ( .A(addr[0]), .B(addr[1]), .Y(n301) );
    or2b2 U126 ( .A(addr[1]), .B(addr[0]), .Y(n302) );
    or2b2 U127 ( .A(addr[1]), .B(n300), .Y(n303) );
    or2b2 U128 ( .A(n305), .B(wrN), .Y(n304) );
    or2b2 U129 ( .A(n307), .B(wrN), .Y(n306) );
    or2b2 U130 ( .A(n309), .B(wrN), .Y(n308) );
    or2b2 U131 ( .A(n311), .B(wrN), .Y(n310) );
    or2b2 U132 ( .A(n317), .B(n299), .Y(n316) );
    clk1b6 U133 ( .A(n316), .Y(N353) );
    or2b2 U134 ( .A(n317), .B(n301), .Y(n318) );
    clk1b6 U135 ( .A(n318), .Y(N369) );
    or2b2 U136 ( .A(n317), .B(n302), .Y(n319) );
    clk1b6 U137 ( .A(n319), .Y(N385) );
    or2b2 U138 ( .A(n317), .B(n303), .Y(n320) );
    clk1b6 U139 ( .A(n320), .Y(N401) );
    or2b2 U140 ( .A(n322), .B(n299), .Y(n321) );
    clk1b6 U141 ( .A(n321), .Y(N417) );
    or2b2 U142 ( .A(n322), .B(n301), .Y(n323) );
    clk1b6 U143 ( .A(n323), .Y(N433) );
    or2b2 U144 ( .A(n322), .B(n302), .Y(n324) );
    clk1b6 U145 ( .A(n324), .Y(N449) );
    or2b2 U146 ( .A(n322), .B(n303), .Y(n325) );
    clk1b6 U147 ( .A(n325), .Y(N465) );
    or2b2 U148 ( .A(n327), .B(n299), .Y(n326) );
    clk1b6 U149 ( .A(n326), .Y(N481) );
    or2b2 U150 ( .A(n327), .B(n301), .Y(n328) );
    clk1b6 U151 ( .A(n328), .Y(N497) );
    or2b2 U152 ( .A(n327), .B(n302), .Y(n329) );
    clk1b6 U153 ( .A(n329), .Y(N513) );
    or2b2 U154 ( .A(n327), .B(n303), .Y(n330) );
    clk1b6 U155 ( .A(n330), .Y(N529) );
    or2b2 U156 ( .A(n312), .B(n304), .Y(n331) );
    clk1b6 U157 ( .A(n331), .Y(N545) );
    or2b2 U158 ( .A(n313), .B(n304), .Y(n332) );
    clk1b6 U159 ( .A(n332), .Y(N561) );
    or2b2 U160 ( .A(n314), .B(n304), .Y(n333) );
    clk1b6 U161 ( .A(n333), .Y(N577) );
    or2b2 U162 ( .A(n315), .B(n304), .Y(n334) );
    clk1b6 U163 ( .A(n334), .Y(N593) );
endmodule


module fifo_mem_1_DW01_inc_5_1 ( A, SUM );
input  [4:0] A;
output [4:0] SUM;
    wire \C99/carry[3] , \C99/carry[2] , \C99/carry[4] ;
    xor2a2 U5 ( .A(\C99/carry[4] ), .B(A[4]), .Y(SUM[4]) );
    ha1a2 \C99/U1_1_3  ( .A(A[3]), .B(\C99/carry[3] ), .S(SUM[3]), .CO(
        \C99/carry[4] ) );
    ha1a2 \C99/U1_1_1  ( .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(\C99/carry[2] )
         );
    ha1a2 \C99/U1_1_2  ( .A(A[2]), .B(\C99/carry[2] ), .S(SUM[2]), .CO(
        \C99/carry[3] ) );
endmodule


module fifo_mem_1_DW01_inc_5_0 ( A, SUM );
input  [4:0] A;
output [4:0] SUM;
    wire \C101/carry[3] , \C101/carry[2] , \C101/carry[4] ;
    xor2a2 U5 ( .A(\C101/carry[4] ), .B(A[4]), .Y(SUM[4]) );
    ha1a2 \C101/U1_1_3  ( .A(A[3]), .B(\C101/carry[3] ), .S(SUM[3]), .CO(
        \C101/carry[4] ) );
    ha1a2 \C101/U1_1_1  ( .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(\C101/carry[2] )
         );
    ha1a2 \C101/U1_1_2  ( .A(A[2]), .B(\C101/carry[2] ), .S(SUM[2]), .CO(
        \C101/carry[3] ) );
endmodule


module fifo_mem_1_DW01_cmp6_5_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
input  [4:0] A;
input  [4:0] B;
input  TC;
output LT, GT, EQ, LE, GE, NE;
    wire n183, n184, n185, n186, n187, n188, n189;
    or2c1 U10 ( .A(n188), .B(n189), .Y(n184) );
    xor2b2 U11 ( .A(B[4]), .B(A[4]), .Y(n189) );
    or3d1 U12 ( .A(n185), .B(n186), .C(n187), .Y(n183) );
    xor2b2 U13 ( .A(B[1]), .B(A[1]), .Y(n185) );
    xor2b2 U14 ( .A(A[3]), .B(B[3]), .Y(n186) );
    xor2b2 U15 ( .A(B[2]), .B(A[2]), .Y(n187) );
    and2c3 U16 ( .A(n183), .B(n184), .Y(EQ) );
    xor2b2 U17 ( .A(A[0]), .B(B[0]), .Y(n188) );
endmodule


module fifo_mem_1 ( data, clk, rstN, wrN, rdN, empty, full );
inout  [7:0] data;
input  clk, rstN, wrN, rdN;
output empty, full;
    wire \addr[3] , \addr[1] , \addr[0] , \wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] , N10, N20, \rd_cntr[4] , 
        \rd_cntr[3] , \rd_cntr[2] , \rd_cntr[1] , \rd_cntr[0] , N47, N57, 
        \_que_1[2] , N87, N115, N116, N117, N118, N120, N121, N122, N123, n335, 
        n336, n337, n338, n339;
    tri \data[7] , \data[6] , \data[5] , \data[4] , \data[3] , \data[2] , 
        \data[1] , \data[0] ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 ;
    tran( \data[7] , data[7] );
    tran( \data[6] , data[6] );
    tran( \data[5] , data[5] );
    tran( \data[4] , data[4] );
    tran( \data[3] , data[3] );
    tran( \data[2] , data[2] );
    tran( \data[1] , data[1] );
    tran( \data[0] , data[0] );
    ram16X8_1 ram ( .data({\data[7] , \data[6] , \data[5] , \data[4] , 
        \data[3] , \data[2] , \data[1] , \data[0] }), .addr({\addr[3] , 
        \_que_1[2] , \addr[1] , \addr[0] }), .oe(wrN), .wrN(wrN), .clk(clk) );
    mx2a3 U4 ( .D0(\wr_cntr[3] ), .D1(\rd_cntr[3] ), .S(wrN), .Y(\addr[3] ) );
    mx2a3 U5 ( .D0(\wr_cntr[2] ), .D1(\rd_cntr[2] ), .S(wrN), .Y(\_que_1[2] )
         );
    mx2d3 U6 ( .D0(N10), .D1(N47), .S(wrN), .Y(\addr[0] ) );
    mx2a3 U7 ( .D0(\wr_cntr[1] ), .D1(\rd_cntr[1] ), .S(wrN), .Y(\addr[1] ) );
    xor2a2 U8 ( .A(\wr_cntr[4] ), .B(\rd_cntr[4] ), .Y(n338) );
    xor2a2 U9 ( .A(N10), .B(wrN), .Y(n336) );
    and2b3 U10 ( .A(n337), .B(N87), .Y(empty) );
    xor2a2 U11 ( .A(\wr_cntr[4] ), .B(\rd_cntr[4] ), .Y(n337) );
    inv1a3 U12 ( .A(wrN), .Y(N20) );
    inv1a3 U13 ( .A(rdN), .Y(N57) );
    inv1a1 U14 ( .A(N87), .Y(n339) );
    inv1a3 U15 ( .A(\rd_cntr[0] ), .Y(N47) );
    fdef2a3 \rd_cntr_reg[1]  ( .D(N115), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[1] ) );
    fdef2a3 \rd_cntr_reg[2]  ( .D(N116), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[2] ) );
    fdef2a3 \rd_cntr_reg[3]  ( .D(N117), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[3] ) );
    fdef2a3 \rd_cntr_reg[4]  ( .D(N118), .E(N57), .CLK(clk), .CLR(rstN), .Q(
        \rd_cntr[4] ) );
    fdef2a3 \wr_cntr_reg[1]  ( .D(N120), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[1] ) );
    fdef2a3 \wr_cntr_reg[2]  ( .D(N121), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[2] ) );
    fdef2a3 \wr_cntr_reg[3]  ( .D(N122), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[3] ) );
    fdef2a3 \wr_cntr_reg[4]  ( .D(N123), .E(N20), .CLK(clk), .CLR(rstN), .Q(
        \wr_cntr[4] ) );
    xor2a2 U16 ( .A(N47), .B(rdN), .Y(n335) );
    fdf2a3 \rd_cntr_reg[0]  ( .D(n335), .CLK(clk), .CLR(rstN), .Q(\rd_cntr[0] 
        ) );
    inv1a3 U17 ( .A(\wr_cntr[0] ), .Y(N10) );
    fdf2a3 \wr_cntr_reg[0]  ( .D(n336), .CLK(clk), .CLR(rstN), .Q(\wr_cntr[0] 
        ) );
    fifo_mem_1_DW01_inc_5_1 C99 ( .A({\rd_cntr[4] , \rd_cntr[3] , \rd_cntr[2] , 
        \rd_cntr[1] , \rd_cntr[0] }), .SUM({N118, N117, N116, N115, 
        SYNOPSYS_UNCONNECTED_1}) );
    fifo_mem_1_DW01_inc_5_0 C101 ( .A({\wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] }), .SUM({N123, N122, N121, 
        N120, SYNOPSYS_UNCONNECTED_2}) );
    fifo_mem_1_DW01_cmp6_5_0 r292 ( .A({\wr_cntr[4] , \wr_cntr[3] , 
        \wr_cntr[2] , \wr_cntr[1] , \wr_cntr[0] }), .B({\rd_cntr[4] , 
        \rd_cntr[3] , \rd_cntr[2] , \rd_cntr[1] , \rd_cntr[0] }), .TC(1'b0), 
        .EQ(N87) );
    and2b2 U18 ( .A(n339), .B(n338), .Y(full) );
endmodule


module fifo32X8 ( din, dout, clk, rstN, wrN, rdN, empty, full );
input  [7:0] din;
output [7:0] dout;
input  clk, rstN, wrN, rdN;
output empty, full;
    wire n9, n23, rdN_even, mem_empty_even, mem_full_even, rdN_odd, 
        mem_empty_odd, mem_full_odd, ldN_even, ldN_odd, \din_even[7] , 
        \din_even[6] , \din_even[5] , \din_even[4] , \din_even[3] , 
        \din_even[2] , \din_even[1] , \din_even[0] , N9, \din_odd[7] , 
        \din_odd[6] , \din_odd[5] , \din_odd[4] , \din_odd[3] , \din_odd[2] , 
        \din_odd[1] , \din_odd[0] , N44, \dout_even[7] , \dout_even[6] , 
        \dout_even[5] , \dout_even[4] , \dout_even[3] , \dout_even[2] , 
        \dout_even[1] , \dout_even[0] , N71, \dout_odd[7] , \dout_odd[6] , 
        \dout_odd[5] , \dout_odd[4] , \dout_odd[3] , \dout_odd[2] , 
        \dout_odd[1] , \dout_odd[0] , N98, _if_0, n341, n342;
    tri \data_even[7] , \data_even[6] , \data_even[5] , \data_even[4] , 
        \data_even[3] , \data_even[2] , \data_even[1] , \data_even[0] , 
        \data_odd[7] , \data_odd[6] , \data_odd[5] , \data_odd[4] , 
        \data_odd[3] , \data_odd[2] , \data_odd[1] , \data_odd[0] ;
    fifo_mem_1 mem_even ( .data({\data_even[7] , \data_even[6] , 
        \data_even[5] , \data_even[4] , \data_even[3] , \data_even[2] , 
        \data_even[1] , \data_even[0] }), .clk(clk), .rstN(rstN), .wrN(n9), 
        .rdN(rdN_even), .empty(mem_empty_even), .full(mem_full_even) );
    fifo_mem_0 mem_odd ( .data({\data_odd[7] , \data_odd[6] , \data_odd[5] , 
        \data_odd[4] , \data_odd[3] , \data_odd[2] , \data_odd[1] , 
        \data_odd[0] }), .clk(clk), .rstN(rstN), .wrN(n23), .rdN(rdN_odd), 
        .empty(mem_empty_odd), .full(mem_full_odd) );
    fifo_cntrl cntrl ( .clk(clk), .rstN(rstN), .wrN(wrN), .rdN(rdN), .empty(
        empty), .full(full), .mem_empty_even(mem_empty_even), .mem_empty_odd(
        mem_empty_odd), .mem_full_even(mem_full_even), .mem_full_odd(
        mem_full_odd), .ldN_even(ldN_even), .ldN_odd(ldN_odd), 
        .out_sel_odd_evenN(_if_0), .rdN_even(rdN_even), .wrN_even(n9), 
        .rdN_odd(rdN_odd), .wrN_odd(n23) );
    inv1a9 U3 ( .A(n23), .Y(n342) );
    inv1a9 U4 ( .A(n9), .Y(n341) );
    mx2a1 U5 ( .D0(\dout_even[3] ), .D1(\dout_odd[3] ), .S(_if_0), .Y(dout[3])
         );
    mx2a1 U6 ( .D0(\dout_even[5] ), .D1(\dout_odd[5] ), .S(_if_0), .Y(dout[5])
         );
    fdef1a3 \dout_odd_reg[0]  ( .D(\data_odd[0] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[0] ) );
    fdef1a3 \dout_odd_reg[1]  ( .D(\data_odd[1] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[1] ) );
    fdef1a3 \dout_odd_reg[2]  ( .D(\data_odd[2] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[2] ) );
    fdef1a3 \dout_odd_reg[3]  ( .D(\data_odd[3] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[3] ) );
    fdef1a3 \dout_odd_reg[4]  ( .D(\data_odd[4] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[4] ) );
    fdef1a3 \dout_odd_reg[5]  ( .D(\data_odd[5] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[5] ) );
    fdef1a3 \dout_odd_reg[6]  ( .D(\data_odd[6] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[6] ) );
    fdef1a3 \dout_odd_reg[7]  ( .D(\data_odd[7] ), .E(N98), .CLK(clk), .Q(
        \dout_odd[7] ) );
    fdef1a3 \dout_even_reg[0]  ( .D(\data_even[0] ), .E(N71), .CLK(clk), .Q(
        \dout_even[0] ) );
    fdef1a3 \dout_even_reg[1]  ( .D(\data_even[1] ), .E(N71), .CLK(clk), .Q(
        \dout_even[1] ) );
    fdef1a3 \dout_even_reg[2]  ( .D(\data_even[2] ), .E(N71), .CLK(clk), .Q(
        \dout_even[2] ) );
    fdef1a3 \dout_even_reg[3]  ( .D(\data_even[3] ), .E(N71), .CLK(clk), .Q(
        \dout_even[3] ) );
    fdef1a3 \dout_even_reg[4]  ( .D(\data_even[4] ), .E(N71), .CLK(clk), .Q(
        \dout_even[4] ) );
    fdef1a3 \dout_even_reg[5]  ( .D(\data_even[5] ), .E(N71), .CLK(clk), .Q(
        \dout_even[5] ) );
    fdef1a3 \dout_even_reg[6]  ( .D(\data_even[6] ), .E(N71), .CLK(clk), .Q(
        \dout_even[6] ) );
    fdef1a3 \dout_even_reg[7]  ( .D(\data_even[7] ), .E(N71), .CLK(clk), .Q(
        \dout_even[7] ) );
    fdef1a3 \din_odd_reg[0]  ( .D(din[0]), .E(N44), .CLK(clk), .Q(\din_odd[0] 
        ) );
    fdef1a3 \din_odd_reg[1]  ( .D(din[1]), .E(N44), .CLK(clk), .Q(\din_odd[1] 
        ) );
    fdef1a3 \din_odd_reg[2]  ( .D(din[2]), .E(N44), .CLK(clk), .Q(\din_odd[2] 
        ) );
    fdef1a3 \din_odd_reg[3]  ( .D(din[3]), .E(N44), .CLK(clk), .Q(\din_odd[3] 
        ) );
    fdef1a3 \din_odd_reg[4]  ( .D(din[4]), .E(N44), .CLK(clk), .Q(\din_odd[4] 
        ) );
    fdef1a3 \din_odd_reg[5]  ( .D(din[5]), .E(N44), .CLK(clk), .Q(\din_odd[5] 
        ) );
    fdef1a3 \din_odd_reg[6]  ( .D(din[6]), .E(N44), .CLK(clk), .Q(\din_odd[6] 
        ) );
    fdef1a3 \din_odd_reg[7]  ( .D(din[7]), .E(N44), .CLK(clk), .Q(\din_odd[7] 
        ) );
    fdef1a3 \din_even_reg[0]  ( .D(din[0]), .E(N9), .CLK(clk), .Q(
        \din_even[0] ) );
    fdef1a3 \din_even_reg[1]  ( .D(din[1]), .E(N9), .CLK(clk), .Q(
        \din_even[1] ) );
    fdef1a3 \din_even_reg[2]  ( .D(din[2]), .E(N9), .CLK(clk), .Q(
        \din_even[2] ) );
    fdef1a3 \din_even_reg[3]  ( .D(din[3]), .E(N9), .CLK(clk), .Q(
        \din_even[3] ) );
    fdef1a3 \din_even_reg[4]  ( .D(din[4]), .E(N9), .CLK(clk), .Q(
        \din_even[4] ) );
    fdef1a3 \din_even_reg[5]  ( .D(din[5]), .E(N9), .CLK(clk), .Q(
        \din_even[5] ) );
    fdef1a3 \din_even_reg[6]  ( .D(din[6]), .E(N9), .CLK(clk), .Q(
        \din_even[6] ) );
    fdef1a3 \din_even_reg[7]  ( .D(din[7]), .E(N9), .CLK(clk), .Q(
        \din_even[7] ) );
    mx2a1 U7 ( .D0(\dout_even[6] ), .D1(\dout_odd[6] ), .S(_if_0), .Y(dout[6])
         );
    mx2a1 U8 ( .D0(\dout_even[0] ), .D1(\dout_odd[0] ), .S(_if_0), .Y(dout[0])
         );
    mx2a1 U9 ( .D0(\dout_even[1] ), .D1(\dout_odd[1] ), .S(_if_0), .Y(dout[1])
         );
    mx2a1 U10 ( .D0(\dout_even[7] ), .D1(\dout_odd[7] ), .S(_if_0), .Y(dout[7]
        ) );
    mx2a1 U11 ( .D0(\dout_even[2] ), .D1(\dout_odd[2] ), .S(_if_0), .Y(dout[2]
        ) );
    mx2a1 U12 ( .D0(\dout_even[4] ), .D1(\dout_odd[4] ), .S(_if_0), .Y(dout[4]
        ) );
    tri1a15 \_1_ca__tri[0]  ( .A(\din_even[0] ), .E(n341), .Y(\data_even[0] )
         );
    tri1a15 \_2_ca__tri[7]  ( .A(\din_odd[7] ), .E(n342), .Y(\data_odd[7] ) );
    tri1a15 \_1_ca__tri[1]  ( .A(\din_even[1] ), .E(n341), .Y(\data_even[1] )
         );
    tri1a15 \_2_ca__tri[6]  ( .A(\din_odd[6] ), .E(n342), .Y(\data_odd[6] ) );
    tri1a15 \_1_ca__tri[2]  ( .A(\din_even[2] ), .E(n341), .Y(\data_even[2] )
         );
    tri1a15 \_2_ca__tri[5]  ( .A(\din_odd[5] ), .E(n342), .Y(\data_odd[5] ) );
    tri1a15 \_1_ca__tri[3]  ( .A(\din_even[3] ), .E(n341), .Y(\data_even[3] )
         );
    tri1a15 \_2_ca__tri[4]  ( .A(\din_odd[4] ), .E(n342), .Y(\data_odd[4] ) );
    tri1a15 \_1_ca__tri[4]  ( .A(\din_even[4] ), .E(n341), .Y(\data_even[4] )
         );
    tri1a15 \_2_ca__tri[3]  ( .A(\din_odd[3] ), .E(n342), .Y(\data_odd[3] ) );
    tri1a15 \_1_ca__tri[5]  ( .A(\din_even[5] ), .E(n341), .Y(\data_even[5] )
         );
    tri1a15 \_2_ca__tri[2]  ( .A(\din_odd[2] ), .E(n342), .Y(\data_odd[2] ) );
    tri1a15 \_1_ca__tri[6]  ( .A(\din_even[6] ), .E(n341), .Y(\data_even[6] )
         );
    tri1a15 \_2_ca__tri[1]  ( .A(\din_odd[1] ), .E(n342), .Y(\data_odd[1] ) );
    tri1a15 \_1_ca__tri[7]  ( .A(\din_even[7] ), .E(n341), .Y(\data_even[7] )
         );
    tri1a15 \_2_ca__tri[0]  ( .A(\din_odd[0] ), .E(n342), .Y(\data_odd[0] ) );
    clk1b6 U13 ( .A(ldN_even), .Y(N9) );
    clk1b6 U14 ( .A(ldN_odd), .Y(N44) );
    clk1b6 U15 ( .A(rdN_even), .Y(N71) );
    clk1b6 U16 ( .A(rdN_odd), .Y(N98) );
endmodule

