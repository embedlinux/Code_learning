`timescale 1ns/1ps

module FIFOTop ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, ClkW, Reseter
 );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

initial $sdf_annotate("FIFOTopNetlist.sdf");

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(n85), .WriteReq(n88), .ClkR(ClkR), 
        .ClkW(ClkW), .Reset(n141) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({n187, n186, n185, 
        n184, n183, n182, n181, n180, n179, n178, n177, n176, n175, n174, n173, 
        n172, n171, n170, n169, n168, n167, n166, n165, n164, n163, n162, n161, 
        n160, n159, n158, n157, n156}), .AddrR(SM_ReadAddr), .AddrW(
        SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), .ChipEna(\*Logic1* ), .Read(
        n91), .Write(SM_MemWriteCmd), .Reset(n154) );
  CKBD0 U2 ( .CLK(SM_MemReadCmd), .C(n155) );
  BUFFD0 U3 ( .I(n74), .Z(n158) );
  INVD0 U4 ( .I(n1), .ZN(n2) );
  CKNXD16 U5 ( .I(Din[31]), .ZN(n1) );
  BUFFD0 U6 ( .I(n2), .Z(n3) );
  BUFFD0 U7 ( .I(n3), .Z(n4) );
  BUFFD0 U8 ( .I(n4), .Z(n5) );
  BUFFD0 U9 ( .I(n5), .Z(n6) );
  BUFFD0 U10 ( .I(n6), .Z(n7) );
  BUFFD0 U11 ( .I(n7), .Z(n8) );
  BUFFD0 U12 ( .I(n8), .Z(n9) );
  BUFFD0 U13 ( .I(n9), .Z(n10) );
  BUFFD0 U14 ( .I(n10), .Z(n11) );
  BUFFD0 U15 ( .I(n11), .Z(n12) );
  BUFFD0 U16 ( .I(n12), .Z(n13) );
  BUFFD0 U17 ( .I(n13), .Z(n14) );
  BUFFD0 U18 ( .I(n14), .Z(n15) );
  BUFFD0 U19 ( .I(n15), .Z(n16) );
  BUFFD0 U20 ( .I(n16), .Z(n17) );
  BUFFD0 U21 ( .I(n17), .Z(n18) );
  BUFFD0 U22 ( .I(n18), .Z(n19) );
  BUFFD0 U23 ( .I(n19), .Z(n20) );
  BUFFD0 U24 ( .I(n20), .Z(n21) );
  BUFFD0 U25 ( .I(n21), .Z(n22) );
  BUFFD0 U26 ( .I(n24), .Z(n186) );
  INVD0 U27 ( .I(n23), .ZN(n24) );
  CKNXD16 U28 ( .I(Din[30]), .ZN(n23) );
  BUFFD0 U29 ( .I(n26), .Z(n185) );
  INVD0 U30 ( .I(n25), .ZN(n26) );
  CKNXD16 U31 ( .I(Din[29]), .ZN(n25) );
  INVD0 U32 ( .I(n27), .ZN(n28) );
  CKNXD16 U33 ( .I(Din[28]), .ZN(n27) );
  INVD0 U34 ( .I(n29), .ZN(n30) );
  CKNXD16 U35 ( .I(Din[24]), .ZN(n29) );
  INVD0 U36 ( .I(n31), .ZN(n32) );
  CKNXD16 U37 ( .I(Din[23]), .ZN(n31) );
  BUFFD0 U38 ( .I(n34), .Z(n178) );
  INVD0 U39 ( .I(n33), .ZN(n34) );
  CKNXD16 U40 ( .I(Din[22]), .ZN(n33) );
  BUFFD0 U41 ( .I(n36), .Z(n177) );
  INVD0 U42 ( .I(n35), .ZN(n36) );
  CKNXD16 U43 ( .I(Din[21]), .ZN(n35) );
  INVD0 U44 ( .I(n37), .ZN(n38) );
  CKNXD16 U45 ( .I(Din[20]), .ZN(n37) );
  INVD0 U46 ( .I(n39), .ZN(n40) );
  CKNXD16 U47 ( .I(Din[19]), .ZN(n39) );
  BUFFD0 U48 ( .I(n42), .Z(n174) );
  INVD0 U49 ( .I(n41), .ZN(n42) );
  CKNXD16 U50 ( .I(Din[18]), .ZN(n41) );
  BUFFD0 U51 ( .I(n44), .Z(n173) );
  INVD0 U52 ( .I(n43), .ZN(n44) );
  CKNXD16 U53 ( .I(Din[17]), .ZN(n43) );
  INVD0 U54 ( .I(n45), .ZN(n46) );
  CKNXD16 U55 ( .I(Din[16]), .ZN(n45) );
  BUFFD0 U56 ( .I(n48), .Z(n171) );
  INVD0 U57 ( .I(n47), .ZN(n48) );
  CKNXD16 U58 ( .I(Din[15]), .ZN(n47) );
  BUFFD0 U59 ( .I(n50), .Z(n170) );
  INVD0 U60 ( .I(n49), .ZN(n50) );
  CKNXD16 U61 ( .I(Din[14]), .ZN(n49) );
  INVD0 U62 ( .I(n51), .ZN(n52) );
  CKNXD16 U63 ( .I(Din[13]), .ZN(n51) );
  INVD0 U64 ( .I(n53), .ZN(n54) );
  CKNXD16 U65 ( .I(Din[12]), .ZN(n53) );
  BUFFD0 U66 ( .I(n56), .Z(n167) );
  INVD0 U67 ( .I(n55), .ZN(n56) );
  CKNXD16 U68 ( .I(Din[11]), .ZN(n55) );
  BUFFD0 U69 ( .I(n58), .Z(n166) );
  INVD0 U70 ( .I(n57), .ZN(n58) );
  CKNXD16 U71 ( .I(Din[10]), .ZN(n57) );
  INVD0 U72 ( .I(n59), .ZN(n60) );
  CKNXD16 U73 ( .I(Din[9]), .ZN(n59) );
  BUFFD0 U74 ( .I(n62), .Z(n164) );
  INVD0 U75 ( .I(n61), .ZN(n62) );
  CKNXD16 U76 ( .I(Din[8]), .ZN(n61) );
  BUFFD0 U77 ( .I(n64), .Z(n163) );
  INVD0 U78 ( .I(n63), .ZN(n64) );
  CKNXD16 U79 ( .I(Din[7]), .ZN(n63) );
  INVD0 U80 ( .I(n65), .ZN(n66) );
  CKNXD16 U81 ( .I(Din[6]), .ZN(n65) );
  INVD0 U82 ( .I(n67), .ZN(n68) );
  CKNXD16 U83 ( .I(Din[5]), .ZN(n67) );
  BUFFD0 U84 ( .I(n70), .Z(n160) );
  INVD0 U85 ( .I(n69), .ZN(n70) );
  CKNXD16 U86 ( .I(Din[4]), .ZN(n69) );
  BUFFD0 U87 ( .I(n72), .Z(n159) );
  INVD0 U88 ( .I(n71), .ZN(n72) );
  CKNXD16 U89 ( .I(Din[3]), .ZN(n71) );
  INVD0 U90 ( .I(n73), .ZN(n74) );
  CKNXD16 U91 ( .I(Din[2]), .ZN(n73) );
  BUFFD0 U92 ( .I(n76), .Z(n157) );
  INVD0 U93 ( .I(n75), .ZN(n76) );
  CKNXD16 U94 ( .I(Din[1]), .ZN(n75) );
  INVD0 U95 ( .I(n77), .ZN(n78) );
  CKNXD16 U96 ( .I(Din[0]), .ZN(n77) );
  INVD0 U97 ( .I(n79), .ZN(n80) );
  CKNXD16 U98 ( .I(Din[27]), .ZN(n79) );
  BUFFD0 U99 ( .I(n82), .Z(n181) );
  INVD0 U100 ( .I(n81), .ZN(n82) );
  CKNXD16 U101 ( .I(Din[25]), .ZN(n81) );
  BUFFD0 U102 ( .I(n84), .Z(n182) );
  INVD0 U103 ( .I(n83), .ZN(n84) );
  CKNXD16 U104 ( .I(Din[26]), .ZN(n83) );
  BUFFD0 U105 ( .I(n86), .Z(n85) );
  BUFFD0 U106 ( .I(n87), .Z(n86) );
  BUFFD0 U107 ( .I(n152), .Z(n87) );
  BUFFD0 U108 ( .I(n89), .Z(n88) );
  BUFFD0 U109 ( .I(n90), .Z(n89) );
  BUFFD0 U110 ( .I(n146), .Z(n90) );
  CKNXD0 U111 ( .I(n145), .ZN(n146) );
  BUFFD0 U112 ( .I(n92), .Z(n91) );
  BUFFD0 U113 ( .I(n93), .Z(n92) );
  BUFFD0 U114 ( .I(n94), .Z(n93) );
  BUFFD0 U115 ( .I(n95), .Z(n94) );
  BUFFD0 U116 ( .I(n96), .Z(n95) );
  BUFFD0 U117 ( .I(n97), .Z(n96) );
  BUFFD0 U118 ( .I(n98), .Z(n97) );
  BUFFD0 U119 ( .I(n99), .Z(n98) );
  BUFFD0 U120 ( .I(n100), .Z(n99) );
  BUFFD0 U121 ( .I(n101), .Z(n100) );
  BUFFD0 U122 ( .I(n102), .Z(n101) );
  BUFFD0 U123 ( .I(n103), .Z(n102) );
  BUFFD0 U124 ( .I(n104), .Z(n103) );
  BUFFD0 U125 ( .I(n105), .Z(n104) );
  BUFFD0 U126 ( .I(n106), .Z(n105) );
  BUFFD0 U127 ( .I(n107), .Z(n106) );
  BUFFD0 U128 ( .I(n108), .Z(n107) );
  BUFFD0 U129 ( .I(n109), .Z(n108) );
  BUFFD0 U130 ( .I(n110), .Z(n109) );
  BUFFD0 U131 ( .I(n111), .Z(n110) );
  BUFFD0 U132 ( .I(n112), .Z(n111) );
  BUFFD0 U133 ( .I(n113), .Z(n112) );
  BUFFD0 U134 ( .I(n114), .Z(n113) );
  BUFFD0 U135 ( .I(n115), .Z(n114) );
  BUFFD0 U136 ( .I(n116), .Z(n115) );
  BUFFD0 U137 ( .I(n117), .Z(n116) );
  BUFFD0 U138 ( .I(n118), .Z(n117) );
  BUFFD0 U139 ( .I(n119), .Z(n118) );
  BUFFD0 U140 ( .I(n120), .Z(n119) );
  BUFFD0 U141 ( .I(n121), .Z(n120) );
  BUFFD0 U142 ( .I(n122), .Z(n121) );
  BUFFD0 U143 ( .I(n123), .Z(n122) );
  BUFFD0 U144 ( .I(n124), .Z(n123) );
  BUFFD0 U145 ( .I(n125), .Z(n124) );
  BUFFD0 U146 ( .I(n126), .Z(n125) );
  BUFFD0 U147 ( .I(n127), .Z(n126) );
  BUFFD0 U148 ( .I(n128), .Z(n127) );
  BUFFD0 U149 ( .I(n129), .Z(n128) );
  BUFFD0 U150 ( .I(n130), .Z(n129) );
  BUFFD0 U151 ( .I(n131), .Z(n130) );
  BUFFD0 U152 ( .I(n132), .Z(n131) );
  BUFFD0 U153 ( .I(n133), .Z(n132) );
  BUFFD0 U154 ( .I(n134), .Z(n133) );
  BUFFD0 U155 ( .I(n135), .Z(n134) );
  BUFFD0 U156 ( .I(n136), .Z(n135) );
  BUFFD0 U157 ( .I(n137), .Z(n136) );
  BUFFD0 U158 ( .I(n138), .Z(n137) );
  BUFFD0 U159 ( .I(n139), .Z(n138) );
  BUFFD0 U160 ( .I(n140), .Z(n139) );
  BUFFD0 U161 ( .I(n155), .Z(n140) );
  BUFFD0 U162 ( .I(n142), .Z(n141) );
  BUFFD0 U163 ( .I(n143), .Z(n142) );
  BUFFD0 U164 ( .I(n144), .Z(n143) );
  BUFFD0 U165 ( .I(n147), .Z(n144) );
  CKNXD16 U166 ( .I(WriteIn), .ZN(n145) );
  BUFFD0 U167 ( .I(n148), .Z(n147) );
  BUFFD0 U168 ( .I(n149), .Z(n148) );
  BUFFD0 U169 ( .I(n150), .Z(n149) );
  BUFFD0 U170 ( .I(n153), .Z(n150) );
  INVD0 U171 ( .I(n151), .ZN(n152) );
  CKNXD16 U172 ( .I(ReadIn), .ZN(n151) );
  BUFFD0 U173 ( .I(n154), .Z(n153) );
  BUFFD1 U174 ( .I(Reseter), .Z(n154) );
  BUFFD1 U175 ( .I(n28), .Z(n184) );
  BUFFD1 U176 ( .I(n22), .Z(n187) );
  BUFFD1 U177 ( .I(n78), .Z(n156) );
  BUFFD1 U178 ( .I(n68), .Z(n161) );
  BUFFD1 U179 ( .I(n66), .Z(n162) );
  BUFFD1 U180 ( .I(n60), .Z(n165) );
  BUFFD1 U181 ( .I(n54), .Z(n168) );
  BUFFD1 U182 ( .I(n52), .Z(n169) );
  BUFFD1 U183 ( .I(n46), .Z(n172) );
  BUFFD1 U184 ( .I(n40), .Z(n175) );
  BUFFD1 U185 ( .I(n38), .Z(n176) );
  BUFFD1 U186 ( .I(n32), .Z(n179) );
  BUFFD1 U187 ( .I(n30), .Z(n180) );
  BUFFD1 U188 ( .I(n80), .Z(n183) );
  TIEH U189 ( .Z(\*Logic1* ) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n1777, n1778, n1779, n1780, StateClockRaw, StateClock, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N169, N171, N172, N173, N321, N323, N324,
         N325, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, \add_387/carry[2] ,
         \add_387/carry[3] , \add_387/carry[4] , \add_306/carry[2] ,
         \add_306/carry[3] , \add_306/carry[4] , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n86, n88, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1654, n1656, n1657, n1672, n1674, n1675, n1677, n1679, n1681,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  assign WriteAddr[0] = N321;
  assign WriteAddr[1] = \add_387/carry[2] ;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  FIFOStateM_AWid5_DW01_inc_0 r151 ( .A({WriteAddr[4:2], \add_387/carry[2] , 
        N321}), .SUM({N70, N69, N68, N67, N66}) );
  FIFOStateM_AWid5_DW01_inc_1 r150 ( .A({ReadAddr[4], n981, ReadAddr[2:1], 
        n1023}), .SUM({N47, N46, N45, N44, N43}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n16), .CPN(StateClock), .CDN(n1672), .QN(n89) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n74), .CPN(StateClock), .CDN(n1672), .QN(
        n87) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n153), .CPN(StateClock), .CDN(n1672), .QN(
        n80) );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n210), .CPN(StateClock), .CDN(n106), .QN(n77) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n267), .CPN(StateClock), .CDN(n106), .QN(n75) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n324), .CPN(StateClock), .CDN(n106), .QN(
        n73) );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n381), .CPN(StateClock), .CDN(n1672), .QN(
        n82) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n437), .CPN(StateClock), .CDN(n1672), .QN(
        n81) );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n494), .CPN(StateClock), .CDN(n1672), .QN(
        n79) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n550), .CPN(StateClock), .CDN(n106), .QN(n78) );
  DFNCND1 \NextState_reg[1]  ( .D(n666), .CPN(StateClock), .CDN(n1672), .Q(
        NextState[1]), .QN(n85) );
  DFNCND1 \NextState_reg[2]  ( .D(n714), .CPN(StateClock), .CDN(n1672), .Q(
        NextState[2]), .QN(n84) );
  DFNCND1 \NextState_reg[0]  ( .D(n772), .CPN(StateClock), .CDN(n1672), .Q(
        NextState[0]), .QN(n83) );
  DFNCND1 ReadCmdr_reg ( .D(n832), .CPN(StateClock), .CDN(n1672), .Q(n1779) );
  DFNCND1 WriteCmdr_reg ( .D(n885), .CPN(StateClock), .CDN(n1672), .Q(n1780)
         );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n1672), 
        .Q(CurState[0]) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n106), 
        .Q(CurState[2]) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n1672), 
        .Q(CurState[1]) );
  EDFCNQD1 \ReadAr_reg[3]  ( .D(N51), .E(N52), .CP(StateClock), .CDN(n1672), 
        .Q(n1777) );
  EDFCNQD1 \ReadAr_reg[0]  ( .D(N48), .E(N52), .CP(StateClock), .CDN(n106), 
        .Q(N169) );
  EDFCNQD1 \ReadAr_reg[1]  ( .D(n1024), .E(N52), .CP(StateClock), .CDN(n106), 
        .Q(\add_306/carry[2] ) );
  EDFCND1 \ReadAr_reg[4]  ( .D(n1072), .E(N52), .CP(StateClock), .CDN(n106), 
        .QN(n1683) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n1118), .E(N52), .CP(StateClock), .CDN(n106), 
        .QN(n1679) );
  EDFCND1 \WriteAr_reg[4]  ( .D(n1200), .E(n1515), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[4]), .QN(n1684) );
  EDFCND1 \WriteAr_reg[3]  ( .D(n1262), .E(n1515), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[3]), .QN(n1687) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n1317), .E(n1515), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[2]), .QN(n1686) );
  EDFCND1 \WriteAr_reg[1]  ( .D(n1373), .E(n1515), .CP(StateClock), .CDN(n106), 
        .Q(\add_387/carry[2] ), .QN(n4) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n1423), .E(n1515), .CP(StateClock), .CDN(n106), 
        .Q(N321), .QN(n1706) );
  DFND4 EmptyFIFOr_reg ( .D(n2), .CPN(StateClock), .QN(n6) );
  DFND1 FullFIFOr_reg ( .D(n1594), .CPN(StateClock), .Q(n1778), .QN(n76) );
  BUFFD0 U3 ( .I(n1709), .Z(n1) );
  MUX2ND1 U4 ( .I0(n935), .I1(n1711), .S(n1707), .ZN(n103) );
  BUFFD0 U5 ( .I(n1591), .Z(n1593) );
  BUFFD0 U6 ( .I(n1538), .Z(n2) );
  OAI22D0 U7 ( .A1(n1681), .A2(n1689), .B1(n1711), .B2(n1774), .ZN(N74) );
  AN2D1 U8 ( .A1(n1708), .A2(WriteReq), .Z(n3) );
  INVD1 U9 ( .I(n3), .ZN(n1710) );
  ND2D1 U10 ( .A1(CurState[2]), .A2(CurState[0]), .ZN(n1691) );
  INVD1 U11 ( .I(n1691), .ZN(n1731) );
  OAI21D1 U12 ( .A1(Reset), .A2(n1693), .B(n1657), .ZN(n5) );
  MUX2ND1 U13 ( .I0(n7), .I1(n1674), .S(n1688), .ZN(n107) );
  BUFFD0 U14 ( .I(n8), .Z(n7) );
  BUFFD0 U15 ( .I(n9), .Z(n8) );
  BUFFD0 U16 ( .I(n10), .Z(n9) );
  BUFFD0 U17 ( .I(n11), .Z(n10) );
  BUFFD0 U18 ( .I(n12), .Z(n11) );
  BUFFD0 U19 ( .I(n13), .Z(n12) );
  BUFFD0 U20 ( .I(n14), .Z(n13) );
  BUFFD0 U21 ( .I(n15), .Z(n14) );
  BUFFD0 U22 ( .I(n89), .Z(n15) );
  BUFFD0 U23 ( .I(n17), .Z(n16) );
  BUFFD0 U24 ( .I(n18), .Z(n17) );
  BUFFD0 U25 ( .I(n19), .Z(n18) );
  BUFFD0 U26 ( .I(n20), .Z(n19) );
  BUFFD0 U27 ( .I(n21), .Z(n20) );
  BUFFD0 U28 ( .I(n22), .Z(n21) );
  BUFFD0 U29 ( .I(n23), .Z(n22) );
  BUFFD0 U30 ( .I(n24), .Z(n23) );
  BUFFD0 U31 ( .I(n25), .Z(n24) );
  BUFFD0 U32 ( .I(n26), .Z(n25) );
  BUFFD0 U33 ( .I(n27), .Z(n26) );
  BUFFD0 U34 ( .I(n28), .Z(n27) );
  BUFFD0 U35 ( .I(n29), .Z(n28) );
  BUFFD0 U36 ( .I(n30), .Z(n29) );
  BUFFD0 U37 ( .I(n31), .Z(n30) );
  BUFFD0 U38 ( .I(n32), .Z(n31) );
  BUFFD0 U39 ( .I(n33), .Z(n32) );
  BUFFD0 U40 ( .I(n34), .Z(n33) );
  BUFFD0 U41 ( .I(n35), .Z(n34) );
  BUFFD0 U42 ( .I(n36), .Z(n35) );
  BUFFD0 U43 ( .I(n37), .Z(n36) );
  BUFFD0 U44 ( .I(n38), .Z(n37) );
  BUFFD0 U45 ( .I(n39), .Z(n38) );
  BUFFD0 U46 ( .I(n40), .Z(n39) );
  BUFFD0 U47 ( .I(n41), .Z(n40) );
  BUFFD0 U48 ( .I(n42), .Z(n41) );
  BUFFD0 U49 ( .I(n43), .Z(n42) );
  BUFFD0 U50 ( .I(n44), .Z(n43) );
  BUFFD0 U51 ( .I(n45), .Z(n44) );
  BUFFD0 U52 ( .I(n46), .Z(n45) );
  BUFFD0 U53 ( .I(n47), .Z(n46) );
  BUFFD0 U54 ( .I(n48), .Z(n47) );
  BUFFD0 U55 ( .I(n49), .Z(n48) );
  BUFFD0 U56 ( .I(n50), .Z(n49) );
  BUFFD0 U57 ( .I(n51), .Z(n50) );
  BUFFD0 U58 ( .I(n52), .Z(n51) );
  BUFFD0 U59 ( .I(n53), .Z(n52) );
  BUFFD0 U60 ( .I(n54), .Z(n53) );
  BUFFD0 U61 ( .I(n55), .Z(n54) );
  BUFFD0 U62 ( .I(n56), .Z(n55) );
  BUFFD0 U63 ( .I(n57), .Z(n56) );
  BUFFD0 U64 ( .I(n58), .Z(n57) );
  BUFFD0 U65 ( .I(n59), .Z(n58) );
  BUFFD0 U66 ( .I(n60), .Z(n59) );
  BUFFD0 U67 ( .I(n61), .Z(n60) );
  BUFFD0 U68 ( .I(n62), .Z(n61) );
  BUFFD0 U69 ( .I(n63), .Z(n62) );
  BUFFD0 U70 ( .I(n107), .Z(n63) );
  MUX2ND1 U71 ( .I0(n64), .I1(n1706), .S(n1685), .ZN(n104) );
  BUFFD0 U72 ( .I(n65), .Z(n64) );
  BUFFD0 U73 ( .I(n66), .Z(n65) );
  BUFFD0 U74 ( .I(n67), .Z(n66) );
  BUFFD0 U75 ( .I(n68), .Z(n67) );
  BUFFD0 U76 ( .I(n69), .Z(n68) );
  BUFFD0 U77 ( .I(n70), .Z(n69) );
  BUFFD0 U78 ( .I(n71), .Z(n70) );
  BUFFD0 U79 ( .I(n72), .Z(n71) );
  BUFFD0 U80 ( .I(n87), .Z(n72) );
  BUFFD0 U81 ( .I(n86), .Z(n74) );
  BUFFD0 U82 ( .I(n88), .Z(n86) );
  BUFFD0 U83 ( .I(n108), .Z(n88) );
  BUFFD0 U84 ( .I(n109), .Z(n108) );
  BUFFD0 U85 ( .I(n110), .Z(n109) );
  BUFFD0 U86 ( .I(n111), .Z(n110) );
  BUFFD0 U87 ( .I(n112), .Z(n111) );
  BUFFD0 U88 ( .I(n113), .Z(n112) );
  BUFFD0 U89 ( .I(n114), .Z(n113) );
  BUFFD0 U90 ( .I(n115), .Z(n114) );
  BUFFD0 U91 ( .I(n116), .Z(n115) );
  BUFFD0 U92 ( .I(n117), .Z(n116) );
  BUFFD0 U93 ( .I(n118), .Z(n117) );
  BUFFD0 U94 ( .I(n119), .Z(n118) );
  BUFFD0 U95 ( .I(n120), .Z(n119) );
  BUFFD0 U96 ( .I(n121), .Z(n120) );
  BUFFD0 U97 ( .I(n122), .Z(n121) );
  BUFFD0 U98 ( .I(n123), .Z(n122) );
  BUFFD0 U99 ( .I(n124), .Z(n123) );
  BUFFD0 U100 ( .I(n125), .Z(n124) );
  BUFFD0 U101 ( .I(n126), .Z(n125) );
  BUFFD0 U102 ( .I(n127), .Z(n126) );
  BUFFD0 U103 ( .I(n128), .Z(n127) );
  BUFFD0 U104 ( .I(n129), .Z(n128) );
  BUFFD0 U105 ( .I(n130), .Z(n129) );
  BUFFD0 U106 ( .I(n131), .Z(n130) );
  BUFFD0 U107 ( .I(n132), .Z(n131) );
  BUFFD0 U108 ( .I(n133), .Z(n132) );
  BUFFD0 U109 ( .I(n134), .Z(n133) );
  BUFFD0 U110 ( .I(n135), .Z(n134) );
  BUFFD0 U111 ( .I(n136), .Z(n135) );
  BUFFD0 U112 ( .I(n137), .Z(n136) );
  BUFFD0 U113 ( .I(n138), .Z(n137) );
  BUFFD0 U114 ( .I(n139), .Z(n138) );
  BUFFD0 U115 ( .I(n140), .Z(n139) );
  BUFFD0 U116 ( .I(n141), .Z(n140) );
  BUFFD0 U117 ( .I(n142), .Z(n141) );
  BUFFD0 U118 ( .I(n143), .Z(n142) );
  BUFFD0 U119 ( .I(n144), .Z(n143) );
  BUFFD0 U120 ( .I(n145), .Z(n144) );
  BUFFD0 U121 ( .I(n146), .Z(n145) );
  BUFFD0 U122 ( .I(n147), .Z(n146) );
  BUFFD0 U123 ( .I(n148), .Z(n147) );
  BUFFD0 U124 ( .I(n149), .Z(n148) );
  BUFFD0 U125 ( .I(n150), .Z(n149) );
  BUFFD0 U126 ( .I(n151), .Z(n150) );
  BUFFD0 U127 ( .I(n152), .Z(n151) );
  BUFFD0 U128 ( .I(n104), .Z(n152) );
  BUFFD0 U129 ( .I(n162), .Z(n153) );
  BUFFD0 U130 ( .I(n155), .Z(n154) );
  BUFFD0 U131 ( .I(n156), .Z(n155) );
  BUFFD0 U132 ( .I(n157), .Z(n156) );
  BUFFD0 U133 ( .I(n158), .Z(n157) );
  BUFFD0 U134 ( .I(n159), .Z(n158) );
  BUFFD0 U135 ( .I(n160), .Z(n159) );
  BUFFD0 U136 ( .I(n161), .Z(n160) );
  BUFFD0 U137 ( .I(n80), .Z(n161) );
  BUFFD0 U138 ( .I(n163), .Z(n162) );
  BUFFD0 U139 ( .I(n164), .Z(n163) );
  BUFFD0 U140 ( .I(n165), .Z(n164) );
  BUFFD0 U141 ( .I(n166), .Z(n165) );
  BUFFD0 U142 ( .I(n167), .Z(n166) );
  BUFFD0 U143 ( .I(n168), .Z(n167) );
  BUFFD0 U144 ( .I(n169), .Z(n168) );
  BUFFD0 U145 ( .I(n170), .Z(n169) );
  BUFFD0 U146 ( .I(n171), .Z(n170) );
  BUFFD0 U147 ( .I(n172), .Z(n171) );
  BUFFD0 U148 ( .I(n173), .Z(n172) );
  BUFFD0 U149 ( .I(n174), .Z(n173) );
  BUFFD0 U150 ( .I(n175), .Z(n174) );
  BUFFD0 U151 ( .I(n176), .Z(n175) );
  BUFFD0 U152 ( .I(n177), .Z(n176) );
  BUFFD0 U153 ( .I(n178), .Z(n177) );
  BUFFD0 U154 ( .I(n179), .Z(n178) );
  BUFFD0 U155 ( .I(n180), .Z(n179) );
  BUFFD0 U156 ( .I(n181), .Z(n180) );
  BUFFD0 U157 ( .I(n182), .Z(n181) );
  BUFFD0 U158 ( .I(n183), .Z(n182) );
  BUFFD0 U159 ( .I(n184), .Z(n183) );
  BUFFD0 U160 ( .I(n185), .Z(n184) );
  BUFFD0 U161 ( .I(n186), .Z(n185) );
  BUFFD0 U162 ( .I(n187), .Z(n186) );
  BUFFD0 U163 ( .I(n188), .Z(n187) );
  BUFFD0 U164 ( .I(n189), .Z(n188) );
  BUFFD0 U165 ( .I(n190), .Z(n189) );
  BUFFD0 U166 ( .I(n191), .Z(n190) );
  BUFFD0 U167 ( .I(n192), .Z(n191) );
  BUFFD0 U168 ( .I(n193), .Z(n192) );
  BUFFD0 U169 ( .I(n194), .Z(n193) );
  BUFFD0 U170 ( .I(n195), .Z(n194) );
  BUFFD0 U171 ( .I(n196), .Z(n195) );
  BUFFD0 U172 ( .I(n197), .Z(n196) );
  BUFFD0 U173 ( .I(n198), .Z(n197) );
  BUFFD0 U174 ( .I(n199), .Z(n198) );
  BUFFD0 U175 ( .I(n200), .Z(n199) );
  BUFFD0 U176 ( .I(n201), .Z(n200) );
  BUFFD0 U177 ( .I(n202), .Z(n201) );
  BUFFD0 U178 ( .I(n203), .Z(n202) );
  BUFFD0 U179 ( .I(n204), .Z(n203) );
  BUFFD0 U180 ( .I(n205), .Z(n204) );
  BUFFD0 U181 ( .I(n206), .Z(n205) );
  BUFFD0 U182 ( .I(n207), .Z(n206) );
  BUFFD0 U183 ( .I(n208), .Z(n207) );
  BUFFD0 U184 ( .I(n209), .Z(n208) );
  BUFFD0 U185 ( .I(n97), .Z(n209) );
  BUFFD0 U186 ( .I(n219), .Z(n210) );
  BUFFD0 U187 ( .I(n212), .Z(n211) );
  BUFFD0 U188 ( .I(n213), .Z(n212) );
  BUFFD0 U189 ( .I(n214), .Z(n213) );
  BUFFD0 U190 ( .I(n215), .Z(n214) );
  BUFFD0 U191 ( .I(n216), .Z(n215) );
  BUFFD0 U192 ( .I(n217), .Z(n216) );
  BUFFD0 U193 ( .I(n218), .Z(n217) );
  BUFFD0 U194 ( .I(n77), .Z(n218) );
  BUFFD0 U195 ( .I(n220), .Z(n219) );
  BUFFD0 U196 ( .I(n221), .Z(n220) );
  BUFFD0 U197 ( .I(n222), .Z(n221) );
  BUFFD0 U198 ( .I(n223), .Z(n222) );
  BUFFD0 U199 ( .I(n224), .Z(n223) );
  BUFFD0 U200 ( .I(n225), .Z(n224) );
  BUFFD0 U201 ( .I(n226), .Z(n225) );
  BUFFD0 U202 ( .I(n227), .Z(n226) );
  BUFFD0 U203 ( .I(n228), .Z(n227) );
  BUFFD0 U204 ( .I(n229), .Z(n228) );
  BUFFD0 U205 ( .I(n230), .Z(n229) );
  BUFFD0 U206 ( .I(n231), .Z(n230) );
  BUFFD0 U207 ( .I(n232), .Z(n231) );
  BUFFD0 U208 ( .I(n233), .Z(n232) );
  BUFFD0 U209 ( .I(n234), .Z(n233) );
  BUFFD0 U210 ( .I(n235), .Z(n234) );
  BUFFD0 U211 ( .I(n236), .Z(n235) );
  BUFFD0 U212 ( .I(n237), .Z(n236) );
  BUFFD0 U213 ( .I(n238), .Z(n237) );
  BUFFD0 U214 ( .I(n239), .Z(n238) );
  BUFFD0 U215 ( .I(n240), .Z(n239) );
  BUFFD0 U216 ( .I(n241), .Z(n240) );
  BUFFD0 U217 ( .I(n242), .Z(n241) );
  BUFFD0 U218 ( .I(n243), .Z(n242) );
  BUFFD0 U219 ( .I(n244), .Z(n243) );
  BUFFD0 U220 ( .I(n245), .Z(n244) );
  BUFFD0 U221 ( .I(n246), .Z(n245) );
  BUFFD0 U222 ( .I(n247), .Z(n246) );
  BUFFD0 U223 ( .I(n248), .Z(n247) );
  BUFFD0 U224 ( .I(n249), .Z(n248) );
  BUFFD0 U225 ( .I(n250), .Z(n249) );
  BUFFD0 U226 ( .I(n251), .Z(n250) );
  BUFFD0 U227 ( .I(n252), .Z(n251) );
  BUFFD0 U228 ( .I(n253), .Z(n252) );
  BUFFD0 U229 ( .I(n254), .Z(n253) );
  BUFFD0 U230 ( .I(n255), .Z(n254) );
  BUFFD0 U231 ( .I(n256), .Z(n255) );
  BUFFD0 U232 ( .I(n257), .Z(n256) );
  BUFFD0 U233 ( .I(n258), .Z(n257) );
  BUFFD0 U234 ( .I(n259), .Z(n258) );
  BUFFD0 U235 ( .I(n260), .Z(n259) );
  BUFFD0 U236 ( .I(n261), .Z(n260) );
  BUFFD0 U237 ( .I(n262), .Z(n261) );
  BUFFD0 U238 ( .I(n263), .Z(n262) );
  BUFFD0 U239 ( .I(n264), .Z(n263) );
  BUFFD0 U240 ( .I(n265), .Z(n264) );
  BUFFD0 U241 ( .I(n266), .Z(n265) );
  BUFFD0 U242 ( .I(n94), .Z(n266) );
  BUFFD0 U243 ( .I(n276), .Z(n267) );
  BUFFD0 U244 ( .I(n269), .Z(n268) );
  BUFFD0 U245 ( .I(n270), .Z(n269) );
  BUFFD0 U246 ( .I(n271), .Z(n270) );
  BUFFD0 U247 ( .I(n272), .Z(n271) );
  BUFFD0 U248 ( .I(n273), .Z(n272) );
  BUFFD0 U249 ( .I(n274), .Z(n273) );
  BUFFD0 U250 ( .I(n275), .Z(n274) );
  BUFFD0 U251 ( .I(n75), .Z(n275) );
  BUFFD0 U252 ( .I(n277), .Z(n276) );
  BUFFD0 U253 ( .I(n278), .Z(n277) );
  BUFFD0 U254 ( .I(n279), .Z(n278) );
  BUFFD0 U255 ( .I(n280), .Z(n279) );
  BUFFD0 U256 ( .I(n281), .Z(n280) );
  BUFFD0 U257 ( .I(n282), .Z(n281) );
  BUFFD0 U258 ( .I(n283), .Z(n282) );
  BUFFD0 U259 ( .I(n284), .Z(n283) );
  BUFFD0 U260 ( .I(n285), .Z(n284) );
  BUFFD0 U261 ( .I(n286), .Z(n285) );
  BUFFD0 U262 ( .I(n287), .Z(n286) );
  BUFFD0 U263 ( .I(n288), .Z(n287) );
  BUFFD0 U264 ( .I(n289), .Z(n288) );
  BUFFD0 U265 ( .I(n290), .Z(n289) );
  BUFFD0 U266 ( .I(n291), .Z(n290) );
  BUFFD0 U267 ( .I(n292), .Z(n291) );
  BUFFD0 U268 ( .I(n293), .Z(n292) );
  BUFFD0 U269 ( .I(n294), .Z(n293) );
  BUFFD0 U270 ( .I(n295), .Z(n294) );
  BUFFD0 U271 ( .I(n296), .Z(n295) );
  BUFFD0 U272 ( .I(n297), .Z(n296) );
  BUFFD0 U273 ( .I(n298), .Z(n297) );
  BUFFD0 U274 ( .I(n299), .Z(n298) );
  BUFFD0 U275 ( .I(n300), .Z(n299) );
  BUFFD0 U276 ( .I(n301), .Z(n300) );
  BUFFD0 U277 ( .I(n302), .Z(n301) );
  BUFFD0 U278 ( .I(n303), .Z(n302) );
  BUFFD0 U279 ( .I(n304), .Z(n303) );
  BUFFD0 U280 ( .I(n305), .Z(n304) );
  BUFFD0 U281 ( .I(n306), .Z(n305) );
  BUFFD0 U282 ( .I(n307), .Z(n306) );
  BUFFD0 U283 ( .I(n308), .Z(n307) );
  BUFFD0 U284 ( .I(n309), .Z(n308) );
  BUFFD0 U285 ( .I(n310), .Z(n309) );
  BUFFD0 U286 ( .I(n311), .Z(n310) );
  BUFFD0 U287 ( .I(n312), .Z(n311) );
  BUFFD0 U288 ( .I(n313), .Z(n312) );
  BUFFD0 U289 ( .I(n314), .Z(n313) );
  BUFFD0 U290 ( .I(n315), .Z(n314) );
  BUFFD0 U291 ( .I(n316), .Z(n315) );
  BUFFD0 U292 ( .I(n317), .Z(n316) );
  BUFFD0 U293 ( .I(n318), .Z(n317) );
  BUFFD0 U294 ( .I(n319), .Z(n318) );
  BUFFD0 U295 ( .I(n320), .Z(n319) );
  BUFFD0 U296 ( .I(n321), .Z(n320) );
  BUFFD0 U297 ( .I(n322), .Z(n321) );
  BUFFD0 U298 ( .I(n323), .Z(n322) );
  BUFFD0 U299 ( .I(n92), .Z(n323) );
  BUFFD0 U300 ( .I(n333), .Z(n324) );
  BUFFD0 U301 ( .I(n326), .Z(n325) );
  BUFFD0 U302 ( .I(n327), .Z(n326) );
  BUFFD0 U303 ( .I(n328), .Z(n327) );
  BUFFD0 U304 ( .I(n329), .Z(n328) );
  BUFFD0 U305 ( .I(n330), .Z(n329) );
  BUFFD0 U306 ( .I(n331), .Z(n330) );
  BUFFD0 U307 ( .I(n332), .Z(n331) );
  BUFFD0 U308 ( .I(n73), .Z(n332) );
  BUFFD0 U309 ( .I(n334), .Z(n333) );
  BUFFD0 U310 ( .I(n335), .Z(n334) );
  BUFFD0 U311 ( .I(n336), .Z(n335) );
  BUFFD0 U312 ( .I(n337), .Z(n336) );
  BUFFD0 U313 ( .I(n338), .Z(n337) );
  BUFFD0 U314 ( .I(n339), .Z(n338) );
  BUFFD0 U315 ( .I(n340), .Z(n339) );
  BUFFD0 U316 ( .I(n341), .Z(n340) );
  BUFFD0 U317 ( .I(n342), .Z(n341) );
  BUFFD0 U318 ( .I(n343), .Z(n342) );
  BUFFD0 U319 ( .I(n344), .Z(n343) );
  BUFFD0 U320 ( .I(n345), .Z(n344) );
  BUFFD0 U321 ( .I(n346), .Z(n345) );
  BUFFD0 U322 ( .I(n347), .Z(n346) );
  BUFFD0 U323 ( .I(n348), .Z(n347) );
  BUFFD0 U324 ( .I(n349), .Z(n348) );
  BUFFD0 U325 ( .I(n350), .Z(n349) );
  BUFFD0 U326 ( .I(n351), .Z(n350) );
  BUFFD0 U327 ( .I(n352), .Z(n351) );
  BUFFD0 U328 ( .I(n353), .Z(n352) );
  BUFFD0 U329 ( .I(n354), .Z(n353) );
  BUFFD0 U330 ( .I(n355), .Z(n354) );
  BUFFD0 U331 ( .I(n356), .Z(n355) );
  BUFFD0 U332 ( .I(n357), .Z(n356) );
  BUFFD0 U333 ( .I(n358), .Z(n357) );
  BUFFD0 U334 ( .I(n359), .Z(n358) );
  BUFFD0 U335 ( .I(n360), .Z(n359) );
  BUFFD0 U336 ( .I(n361), .Z(n360) );
  BUFFD0 U337 ( .I(n362), .Z(n361) );
  BUFFD0 U338 ( .I(n363), .Z(n362) );
  BUFFD0 U339 ( .I(n364), .Z(n363) );
  BUFFD0 U340 ( .I(n365), .Z(n364) );
  BUFFD0 U341 ( .I(n366), .Z(n365) );
  BUFFD0 U342 ( .I(n367), .Z(n366) );
  BUFFD0 U343 ( .I(n368), .Z(n367) );
  BUFFD0 U344 ( .I(n369), .Z(n368) );
  BUFFD0 U345 ( .I(n370), .Z(n369) );
  BUFFD0 U346 ( .I(n371), .Z(n370) );
  BUFFD0 U347 ( .I(n372), .Z(n371) );
  BUFFD0 U348 ( .I(n373), .Z(n372) );
  BUFFD0 U349 ( .I(n374), .Z(n373) );
  BUFFD0 U350 ( .I(n375), .Z(n374) );
  BUFFD0 U351 ( .I(n376), .Z(n375) );
  BUFFD0 U352 ( .I(n377), .Z(n376) );
  BUFFD0 U353 ( .I(n378), .Z(n377) );
  BUFFD0 U354 ( .I(n379), .Z(n378) );
  BUFFD0 U355 ( .I(n380), .Z(n379) );
  BUFFD0 U356 ( .I(n90), .Z(n380) );
  BUFFD0 U357 ( .I(n389), .Z(n381) );
  BUFFD0 U358 ( .I(n383), .Z(n382) );
  BUFFD0 U359 ( .I(n384), .Z(n383) );
  BUFFD0 U360 ( .I(n385), .Z(n384) );
  BUFFD0 U361 ( .I(n386), .Z(n385) );
  BUFFD0 U362 ( .I(n387), .Z(n386) );
  BUFFD0 U363 ( .I(n388), .Z(n387) );
  BUFFD0 U364 ( .I(n884), .Z(n388) );
  BUFFD0 U365 ( .I(n390), .Z(n389) );
  BUFFD0 U366 ( .I(n391), .Z(n390) );
  BUFFD0 U367 ( .I(n392), .Z(n391) );
  BUFFD0 U368 ( .I(n393), .Z(n392) );
  BUFFD0 U369 ( .I(n394), .Z(n393) );
  BUFFD0 U370 ( .I(n395), .Z(n394) );
  BUFFD0 U371 ( .I(n396), .Z(n395) );
  BUFFD0 U372 ( .I(n397), .Z(n396) );
  BUFFD0 U373 ( .I(n398), .Z(n397) );
  BUFFD0 U374 ( .I(n399), .Z(n398) );
  BUFFD0 U375 ( .I(n400), .Z(n399) );
  BUFFD0 U376 ( .I(n401), .Z(n400) );
  BUFFD0 U377 ( .I(n402), .Z(n401) );
  BUFFD0 U378 ( .I(n403), .Z(n402) );
  BUFFD0 U379 ( .I(n404), .Z(n403) );
  BUFFD0 U380 ( .I(n405), .Z(n404) );
  BUFFD0 U381 ( .I(n406), .Z(n405) );
  BUFFD0 U382 ( .I(n407), .Z(n406) );
  BUFFD0 U383 ( .I(n408), .Z(n407) );
  BUFFD0 U384 ( .I(n409), .Z(n408) );
  BUFFD0 U385 ( .I(n410), .Z(n409) );
  BUFFD0 U386 ( .I(n411), .Z(n410) );
  BUFFD0 U387 ( .I(n412), .Z(n411) );
  BUFFD0 U388 ( .I(n413), .Z(n412) );
  BUFFD0 U389 ( .I(n414), .Z(n413) );
  BUFFD0 U390 ( .I(n415), .Z(n414) );
  BUFFD0 U391 ( .I(n416), .Z(n415) );
  BUFFD0 U392 ( .I(n417), .Z(n416) );
  BUFFD0 U393 ( .I(n418), .Z(n417) );
  BUFFD0 U394 ( .I(n419), .Z(n418) );
  BUFFD0 U395 ( .I(n420), .Z(n419) );
  BUFFD0 U396 ( .I(n421), .Z(n420) );
  BUFFD0 U397 ( .I(n422), .Z(n421) );
  BUFFD0 U398 ( .I(n423), .Z(n422) );
  BUFFD0 U399 ( .I(n424), .Z(n423) );
  BUFFD0 U400 ( .I(n425), .Z(n424) );
  BUFFD0 U401 ( .I(n426), .Z(n425) );
  BUFFD0 U402 ( .I(n427), .Z(n426) );
  BUFFD0 U403 ( .I(n428), .Z(n427) );
  BUFFD0 U404 ( .I(n429), .Z(n428) );
  BUFFD0 U405 ( .I(n430), .Z(n429) );
  BUFFD0 U406 ( .I(n431), .Z(n430) );
  BUFFD0 U407 ( .I(n432), .Z(n431) );
  BUFFD0 U408 ( .I(n433), .Z(n432) );
  BUFFD0 U409 ( .I(n434), .Z(n433) );
  BUFFD0 U410 ( .I(n435), .Z(n434) );
  BUFFD0 U411 ( .I(n436), .Z(n435) );
  BUFFD0 U412 ( .I(n99), .Z(n436) );
  BUFFD0 U413 ( .I(n446), .Z(n437) );
  BUFFD0 U414 ( .I(n439), .Z(n438) );
  BUFFD0 U415 ( .I(n440), .Z(n439) );
  BUFFD0 U416 ( .I(n441), .Z(n440) );
  BUFFD0 U417 ( .I(n442), .Z(n441) );
  BUFFD0 U418 ( .I(n443), .Z(n442) );
  BUFFD0 U419 ( .I(n444), .Z(n443) );
  BUFFD0 U420 ( .I(n445), .Z(n444) );
  BUFFD0 U421 ( .I(n81), .Z(n445) );
  BUFFD0 U422 ( .I(n447), .Z(n446) );
  BUFFD0 U423 ( .I(n448), .Z(n447) );
  BUFFD0 U424 ( .I(n449), .Z(n448) );
  BUFFD0 U425 ( .I(n450), .Z(n449) );
  BUFFD0 U426 ( .I(n451), .Z(n450) );
  BUFFD0 U427 ( .I(n452), .Z(n451) );
  BUFFD0 U428 ( .I(n453), .Z(n452) );
  BUFFD0 U429 ( .I(n454), .Z(n453) );
  BUFFD0 U430 ( .I(n455), .Z(n454) );
  BUFFD0 U431 ( .I(n456), .Z(n455) );
  BUFFD0 U432 ( .I(n457), .Z(n456) );
  BUFFD0 U433 ( .I(n458), .Z(n457) );
  BUFFD0 U434 ( .I(n459), .Z(n458) );
  BUFFD0 U435 ( .I(n460), .Z(n459) );
  BUFFD0 U436 ( .I(n461), .Z(n460) );
  BUFFD0 U437 ( .I(n462), .Z(n461) );
  BUFFD0 U438 ( .I(n463), .Z(n462) );
  BUFFD0 U439 ( .I(n464), .Z(n463) );
  BUFFD0 U440 ( .I(n465), .Z(n464) );
  BUFFD0 U441 ( .I(n466), .Z(n465) );
  BUFFD0 U442 ( .I(n467), .Z(n466) );
  BUFFD0 U443 ( .I(n468), .Z(n467) );
  BUFFD0 U444 ( .I(n469), .Z(n468) );
  BUFFD0 U445 ( .I(n470), .Z(n469) );
  BUFFD0 U446 ( .I(n471), .Z(n470) );
  BUFFD0 U447 ( .I(n472), .Z(n471) );
  BUFFD0 U448 ( .I(n473), .Z(n472) );
  BUFFD0 U449 ( .I(n474), .Z(n473) );
  BUFFD0 U450 ( .I(n475), .Z(n474) );
  BUFFD0 U451 ( .I(n476), .Z(n475) );
  BUFFD0 U452 ( .I(n477), .Z(n476) );
  BUFFD0 U453 ( .I(n478), .Z(n477) );
  BUFFD0 U454 ( .I(n479), .Z(n478) );
  BUFFD0 U455 ( .I(n480), .Z(n479) );
  BUFFD0 U456 ( .I(n481), .Z(n480) );
  BUFFD0 U457 ( .I(n482), .Z(n481) );
  BUFFD0 U458 ( .I(n483), .Z(n482) );
  BUFFD0 U459 ( .I(n484), .Z(n483) );
  BUFFD0 U460 ( .I(n485), .Z(n484) );
  BUFFD0 U461 ( .I(n486), .Z(n485) );
  BUFFD0 U462 ( .I(n487), .Z(n486) );
  BUFFD0 U463 ( .I(n488), .Z(n487) );
  BUFFD0 U464 ( .I(n489), .Z(n488) );
  BUFFD0 U465 ( .I(n490), .Z(n489) );
  BUFFD0 U466 ( .I(n491), .Z(n490) );
  BUFFD0 U467 ( .I(n492), .Z(n491) );
  BUFFD0 U468 ( .I(n493), .Z(n492) );
  BUFFD0 U469 ( .I(n98), .Z(n493) );
  BUFFD0 U470 ( .I(n502), .Z(n494) );
  BUFFD0 U471 ( .I(n496), .Z(n495) );
  BUFFD0 U472 ( .I(n497), .Z(n496) );
  BUFFD0 U473 ( .I(n498), .Z(n497) );
  BUFFD0 U474 ( .I(n499), .Z(n498) );
  BUFFD0 U475 ( .I(n500), .Z(n499) );
  BUFFD0 U476 ( .I(n501), .Z(n500) );
  BUFFD0 U477 ( .I(n831), .Z(n501) );
  BUFFD0 U478 ( .I(n503), .Z(n502) );
  BUFFD0 U479 ( .I(n504), .Z(n503) );
  BUFFD0 U480 ( .I(n505), .Z(n504) );
  BUFFD0 U481 ( .I(n506), .Z(n505) );
  BUFFD0 U482 ( .I(n507), .Z(n506) );
  BUFFD0 U483 ( .I(n508), .Z(n507) );
  BUFFD0 U484 ( .I(n509), .Z(n508) );
  BUFFD0 U485 ( .I(n510), .Z(n509) );
  BUFFD0 U486 ( .I(n511), .Z(n510) );
  BUFFD0 U487 ( .I(n512), .Z(n511) );
  BUFFD0 U488 ( .I(n513), .Z(n512) );
  BUFFD0 U489 ( .I(n514), .Z(n513) );
  BUFFD0 U490 ( .I(n515), .Z(n514) );
  BUFFD0 U491 ( .I(n516), .Z(n515) );
  BUFFD0 U492 ( .I(n517), .Z(n516) );
  BUFFD0 U493 ( .I(n518), .Z(n517) );
  BUFFD0 U494 ( .I(n519), .Z(n518) );
  BUFFD0 U495 ( .I(n520), .Z(n519) );
  BUFFD0 U496 ( .I(n521), .Z(n520) );
  BUFFD0 U497 ( .I(n522), .Z(n521) );
  BUFFD0 U498 ( .I(n523), .Z(n522) );
  BUFFD0 U499 ( .I(n524), .Z(n523) );
  BUFFD0 U500 ( .I(n525), .Z(n524) );
  BUFFD0 U501 ( .I(n526), .Z(n525) );
  BUFFD0 U502 ( .I(n527), .Z(n526) );
  BUFFD0 U503 ( .I(n528), .Z(n527) );
  BUFFD0 U504 ( .I(n529), .Z(n528) );
  BUFFD0 U505 ( .I(n530), .Z(n529) );
  BUFFD0 U506 ( .I(n531), .Z(n530) );
  BUFFD0 U507 ( .I(n532), .Z(n531) );
  BUFFD0 U508 ( .I(n533), .Z(n532) );
  BUFFD0 U509 ( .I(n534), .Z(n533) );
  BUFFD0 U510 ( .I(n535), .Z(n534) );
  BUFFD0 U511 ( .I(n536), .Z(n535) );
  BUFFD0 U512 ( .I(n537), .Z(n536) );
  BUFFD0 U513 ( .I(n538), .Z(n537) );
  BUFFD0 U514 ( .I(n539), .Z(n538) );
  BUFFD0 U515 ( .I(n540), .Z(n539) );
  BUFFD0 U516 ( .I(n541), .Z(n540) );
  BUFFD0 U517 ( .I(n542), .Z(n541) );
  BUFFD0 U518 ( .I(n543), .Z(n542) );
  BUFFD0 U519 ( .I(n544), .Z(n543) );
  BUFFD0 U520 ( .I(n545), .Z(n544) );
  BUFFD0 U521 ( .I(n546), .Z(n545) );
  BUFFD0 U522 ( .I(n547), .Z(n546) );
  BUFFD0 U523 ( .I(n548), .Z(n547) );
  BUFFD0 U524 ( .I(n549), .Z(n548) );
  BUFFD0 U525 ( .I(n96), .Z(n549) );
  BUFFD0 U526 ( .I(n558), .Z(n550) );
  BUFFD0 U527 ( .I(n552), .Z(n551) );
  BUFFD0 U528 ( .I(n553), .Z(n552) );
  BUFFD0 U529 ( .I(n554), .Z(n553) );
  BUFFD0 U530 ( .I(n555), .Z(n554) );
  BUFFD0 U531 ( .I(n556), .Z(n555) );
  BUFFD0 U532 ( .I(n557), .Z(n556) );
  BUFFD0 U533 ( .I(n830), .Z(n557) );
  BUFFD0 U534 ( .I(n559), .Z(n558) );
  BUFFD0 U535 ( .I(n560), .Z(n559) );
  BUFFD0 U536 ( .I(n561), .Z(n560) );
  BUFFD0 U537 ( .I(n562), .Z(n561) );
  BUFFD0 U538 ( .I(n563), .Z(n562) );
  BUFFD0 U539 ( .I(n564), .Z(n563) );
  BUFFD0 U540 ( .I(n565), .Z(n564) );
  BUFFD0 U541 ( .I(n566), .Z(n565) );
  BUFFD0 U542 ( .I(n567), .Z(n566) );
  BUFFD0 U543 ( .I(n568), .Z(n567) );
  BUFFD0 U544 ( .I(n569), .Z(n568) );
  BUFFD0 U545 ( .I(n570), .Z(n569) );
  BUFFD0 U546 ( .I(n571), .Z(n570) );
  BUFFD0 U547 ( .I(n572), .Z(n571) );
  BUFFD0 U548 ( .I(n573), .Z(n572) );
  BUFFD0 U549 ( .I(n574), .Z(n573) );
  BUFFD0 U550 ( .I(n575), .Z(n574) );
  BUFFD0 U551 ( .I(n576), .Z(n575) );
  BUFFD0 U552 ( .I(n577), .Z(n576) );
  BUFFD0 U553 ( .I(n578), .Z(n577) );
  BUFFD0 U554 ( .I(n579), .Z(n578) );
  BUFFD0 U555 ( .I(n580), .Z(n579) );
  BUFFD0 U556 ( .I(n581), .Z(n580) );
  BUFFD0 U557 ( .I(n582), .Z(n581) );
  BUFFD0 U558 ( .I(n583), .Z(n582) );
  BUFFD0 U559 ( .I(n584), .Z(n583) );
  BUFFD0 U560 ( .I(n585), .Z(n584) );
  BUFFD0 U561 ( .I(n586), .Z(n585) );
  BUFFD0 U562 ( .I(n587), .Z(n586) );
  BUFFD0 U563 ( .I(n588), .Z(n587) );
  BUFFD0 U564 ( .I(n589), .Z(n588) );
  BUFFD0 U565 ( .I(n590), .Z(n589) );
  BUFFD0 U566 ( .I(n591), .Z(n590) );
  BUFFD0 U567 ( .I(n592), .Z(n591) );
  BUFFD0 U568 ( .I(n593), .Z(n592) );
  BUFFD0 U569 ( .I(n594), .Z(n593) );
  BUFFD0 U570 ( .I(n595), .Z(n594) );
  BUFFD0 U571 ( .I(n596), .Z(n595) );
  BUFFD0 U572 ( .I(n597), .Z(n596) );
  BUFFD0 U573 ( .I(n598), .Z(n597) );
  BUFFD0 U574 ( .I(n599), .Z(n598) );
  BUFFD0 U575 ( .I(n600), .Z(n599) );
  BUFFD0 U576 ( .I(n601), .Z(n600) );
  BUFFD0 U577 ( .I(n602), .Z(n601) );
  BUFFD0 U578 ( .I(n603), .Z(n602) );
  BUFFD0 U579 ( .I(n604), .Z(n603) );
  BUFFD0 U580 ( .I(n605), .Z(n604) );
  BUFFD0 U581 ( .I(n95), .Z(n605) );
  BUFFD0 U582 ( .I(n934), .Z(n606) );
  BUFFD0 U583 ( .I(n606), .Z(n607) );
  BUFFD0 U584 ( .I(n607), .Z(n608) );
  BUFFD0 U585 ( .I(n608), .Z(n609) );
  BUFFD0 U586 ( .I(n609), .Z(n610) );
  BUFFD0 U587 ( .I(n610), .Z(n611) );
  BUFFD0 U588 ( .I(n611), .Z(n612) );
  BUFFD0 U589 ( .I(n612), .Z(n613) );
  BUFFD0 U590 ( .I(n613), .Z(n614) );
  BUFFD0 U591 ( .I(n614), .Z(n615) );
  BUFFD0 U592 ( .I(n615), .Z(n616) );
  BUFFD0 U593 ( .I(n616), .Z(n617) );
  BUFFD0 U594 ( .I(n617), .Z(n618) );
  BUFFD0 U595 ( .I(n618), .Z(n619) );
  BUFFD0 U596 ( .I(n619), .Z(n620) );
  BUFFD0 U597 ( .I(n620), .Z(n621) );
  BUFFD0 U598 ( .I(n621), .Z(n622) );
  BUFFD0 U599 ( .I(n622), .Z(n623) );
  BUFFD0 U600 ( .I(n623), .Z(n624) );
  BUFFD0 U601 ( .I(n624), .Z(n625) );
  BUFFD0 U602 ( .I(n625), .Z(n626) );
  BUFFD0 U603 ( .I(n626), .Z(n627) );
  BUFFD0 U604 ( .I(n627), .Z(n628) );
  BUFFD0 U605 ( .I(n628), .Z(n629) );
  BUFFD0 U606 ( .I(n629), .Z(n630) );
  BUFFD0 U607 ( .I(n630), .Z(n631) );
  BUFFD0 U608 ( .I(n631), .Z(n632) );
  BUFFD0 U609 ( .I(n632), .Z(n633) );
  BUFFD0 U610 ( .I(n633), .Z(n634) );
  BUFFD0 U611 ( .I(n634), .Z(n635) );
  BUFFD0 U612 ( .I(n635), .Z(n636) );
  BUFFD0 U613 ( .I(n636), .Z(n637) );
  BUFFD0 U614 ( .I(n637), .Z(n638) );
  BUFFD0 U615 ( .I(n638), .Z(n639) );
  BUFFD0 U616 ( .I(n639), .Z(n640) );
  BUFFD0 U617 ( .I(n640), .Z(n641) );
  BUFFD0 U618 ( .I(n641), .Z(n642) );
  BUFFD0 U619 ( .I(n642), .Z(n643) );
  BUFFD0 U620 ( .I(n643), .Z(n644) );
  BUFFD0 U621 ( .I(n644), .Z(n645) );
  BUFFD0 U622 ( .I(n645), .Z(n646) );
  BUFFD0 U623 ( .I(n646), .Z(n647) );
  BUFFD0 U624 ( .I(n1780), .Z(n648) );
  BUFFD0 U625 ( .I(n647), .Z(n649) );
  BUFFD0 U626 ( .I(n649), .Z(n650) );
  BUFFD0 U627 ( .I(n650), .Z(n651) );
  BUFFD0 U628 ( .I(n651), .Z(n652) );
  BUFFD0 U629 ( .I(n652), .Z(n653) );
  BUFFD0 U630 ( .I(n648), .Z(n654) );
  BUFFD0 U631 ( .I(n654), .Z(n655) );
  CKBD0 U632 ( .CLK(n653), .C(WriteCmd) );
  MUX2ND1 U633 ( .I0(n1719), .I1(n657), .S(n1720), .ZN(n102) );
  BUFFD0 U634 ( .I(n658), .Z(n657) );
  BUFFD0 U635 ( .I(n659), .Z(n658) );
  BUFFD0 U636 ( .I(n660), .Z(n659) );
  BUFFD0 U637 ( .I(n661), .Z(n660) );
  BUFFD0 U638 ( .I(n662), .Z(n661) );
  BUFFD0 U639 ( .I(n663), .Z(n662) );
  BUFFD0 U640 ( .I(n664), .Z(n663) );
  BUFFD0 U641 ( .I(n665), .Z(n664) );
  BUFFD0 U642 ( .I(n85), .Z(n665) );
  BUFFD0 U643 ( .I(n667), .Z(n666) );
  BUFFD0 U644 ( .I(n668), .Z(n667) );
  BUFFD0 U645 ( .I(n669), .Z(n668) );
  BUFFD0 U646 ( .I(n670), .Z(n669) );
  BUFFD0 U647 ( .I(n671), .Z(n670) );
  BUFFD0 U648 ( .I(n672), .Z(n671) );
  BUFFD0 U649 ( .I(n673), .Z(n672) );
  BUFFD0 U650 ( .I(n674), .Z(n673) );
  BUFFD0 U651 ( .I(n675), .Z(n674) );
  BUFFD0 U652 ( .I(n676), .Z(n675) );
  BUFFD0 U653 ( .I(n677), .Z(n676) );
  BUFFD0 U654 ( .I(n678), .Z(n677) );
  BUFFD0 U655 ( .I(n679), .Z(n678) );
  BUFFD0 U656 ( .I(n680), .Z(n679) );
  BUFFD0 U657 ( .I(n681), .Z(n680) );
  BUFFD0 U658 ( .I(n682), .Z(n681) );
  BUFFD0 U659 ( .I(n683), .Z(n682) );
  BUFFD0 U660 ( .I(n684), .Z(n683) );
  BUFFD0 U661 ( .I(n685), .Z(n684) );
  BUFFD0 U662 ( .I(n686), .Z(n685) );
  BUFFD0 U663 ( .I(n687), .Z(n686) );
  BUFFD0 U664 ( .I(n688), .Z(n687) );
  BUFFD0 U665 ( .I(n689), .Z(n688) );
  BUFFD0 U666 ( .I(n690), .Z(n689) );
  BUFFD0 U667 ( .I(n691), .Z(n690) );
  BUFFD0 U668 ( .I(n692), .Z(n691) );
  BUFFD0 U669 ( .I(n693), .Z(n692) );
  BUFFD0 U670 ( .I(n694), .Z(n693) );
  BUFFD0 U671 ( .I(n695), .Z(n694) );
  BUFFD0 U672 ( .I(n696), .Z(n695) );
  BUFFD0 U673 ( .I(n697), .Z(n696) );
  BUFFD0 U674 ( .I(n698), .Z(n697) );
  BUFFD0 U675 ( .I(n699), .Z(n698) );
  BUFFD0 U676 ( .I(n700), .Z(n699) );
  BUFFD0 U677 ( .I(n701), .Z(n700) );
  BUFFD0 U678 ( .I(n702), .Z(n701) );
  BUFFD0 U679 ( .I(n703), .Z(n702) );
  BUFFD0 U680 ( .I(n704), .Z(n703) );
  BUFFD0 U681 ( .I(n705), .Z(n704) );
  BUFFD0 U682 ( .I(n706), .Z(n705) );
  BUFFD0 U683 ( .I(n707), .Z(n706) );
  BUFFD0 U684 ( .I(n708), .Z(n707) );
  BUFFD0 U685 ( .I(n709), .Z(n708) );
  BUFFD0 U686 ( .I(n710), .Z(n709) );
  BUFFD0 U687 ( .I(n711), .Z(n710) );
  BUFFD0 U688 ( .I(n712), .Z(n711) );
  BUFFD0 U689 ( .I(n713), .Z(n712) );
  BUFFD0 U690 ( .I(n102), .Z(n713) );
  BUFFD0 U691 ( .I(n724), .Z(n714) );
  BUFFD0 U692 ( .I(n716), .Z(n715) );
  BUFFD0 U693 ( .I(n717), .Z(n716) );
  BUFFD0 U694 ( .I(n718), .Z(n717) );
  BUFFD0 U695 ( .I(n719), .Z(n718) );
  BUFFD0 U696 ( .I(n720), .Z(n719) );
  BUFFD0 U697 ( .I(n721), .Z(n720) );
  BUFFD0 U698 ( .I(n722), .Z(n721) );
  BUFFD0 U699 ( .I(n723), .Z(n722) );
  BUFFD0 U700 ( .I(n84), .Z(n723) );
  BUFFD0 U701 ( .I(n725), .Z(n724) );
  BUFFD0 U702 ( .I(n726), .Z(n725) );
  BUFFD0 U703 ( .I(n727), .Z(n726) );
  BUFFD0 U704 ( .I(n728), .Z(n727) );
  BUFFD0 U705 ( .I(n729), .Z(n728) );
  BUFFD0 U706 ( .I(n730), .Z(n729) );
  BUFFD0 U707 ( .I(n731), .Z(n730) );
  BUFFD0 U708 ( .I(n732), .Z(n731) );
  BUFFD0 U709 ( .I(n733), .Z(n732) );
  BUFFD0 U710 ( .I(n734), .Z(n733) );
  BUFFD0 U711 ( .I(n735), .Z(n734) );
  BUFFD0 U712 ( .I(n736), .Z(n735) );
  BUFFD0 U713 ( .I(n737), .Z(n736) );
  BUFFD0 U714 ( .I(n738), .Z(n737) );
  BUFFD0 U715 ( .I(n739), .Z(n738) );
  BUFFD0 U716 ( .I(n740), .Z(n739) );
  BUFFD0 U717 ( .I(n741), .Z(n740) );
  BUFFD0 U718 ( .I(n742), .Z(n741) );
  BUFFD0 U719 ( .I(n743), .Z(n742) );
  BUFFD0 U720 ( .I(n744), .Z(n743) );
  BUFFD0 U721 ( .I(n745), .Z(n744) );
  BUFFD0 U722 ( .I(n746), .Z(n745) );
  BUFFD0 U723 ( .I(n747), .Z(n746) );
  BUFFD0 U724 ( .I(n748), .Z(n747) );
  BUFFD0 U725 ( .I(n749), .Z(n748) );
  BUFFD0 U726 ( .I(n750), .Z(n749) );
  BUFFD0 U727 ( .I(n751), .Z(n750) );
  BUFFD0 U728 ( .I(n752), .Z(n751) );
  BUFFD0 U729 ( .I(n753), .Z(n752) );
  BUFFD0 U730 ( .I(n754), .Z(n753) );
  BUFFD0 U731 ( .I(n755), .Z(n754) );
  BUFFD0 U732 ( .I(n756), .Z(n755) );
  BUFFD0 U733 ( .I(n757), .Z(n756) );
  BUFFD0 U734 ( .I(n758), .Z(n757) );
  BUFFD0 U735 ( .I(n759), .Z(n758) );
  BUFFD0 U736 ( .I(n760), .Z(n759) );
  BUFFD0 U737 ( .I(n761), .Z(n760) );
  BUFFD0 U738 ( .I(n762), .Z(n761) );
  BUFFD0 U739 ( .I(n763), .Z(n762) );
  BUFFD0 U740 ( .I(n764), .Z(n763) );
  BUFFD0 U741 ( .I(n765), .Z(n764) );
  BUFFD0 U742 ( .I(n766), .Z(n765) );
  BUFFD0 U743 ( .I(n767), .Z(n766) );
  BUFFD0 U744 ( .I(n768), .Z(n767) );
  BUFFD0 U745 ( .I(n769), .Z(n768) );
  BUFFD0 U746 ( .I(n770), .Z(n769) );
  BUFFD0 U747 ( .I(n771), .Z(n770) );
  BUFFD0 U748 ( .I(n101), .Z(n771) );
  BUFFD0 U749 ( .I(n782), .Z(n772) );
  BUFFD0 U750 ( .I(n774), .Z(n773) );
  BUFFD0 U751 ( .I(n775), .Z(n774) );
  BUFFD0 U752 ( .I(n776), .Z(n775) );
  BUFFD0 U753 ( .I(n777), .Z(n776) );
  BUFFD0 U754 ( .I(n778), .Z(n777) );
  BUFFD0 U755 ( .I(n779), .Z(n778) );
  BUFFD0 U756 ( .I(n780), .Z(n779) );
  BUFFD0 U757 ( .I(n781), .Z(n780) );
  BUFFD0 U758 ( .I(n83), .Z(n781) );
  BUFFD0 U759 ( .I(n783), .Z(n782) );
  BUFFD0 U760 ( .I(n784), .Z(n783) );
  BUFFD0 U761 ( .I(n785), .Z(n784) );
  BUFFD0 U762 ( .I(n786), .Z(n785) );
  BUFFD0 U763 ( .I(n787), .Z(n786) );
  BUFFD0 U764 ( .I(n788), .Z(n787) );
  BUFFD0 U765 ( .I(n789), .Z(n788) );
  BUFFD0 U766 ( .I(n790), .Z(n789) );
  BUFFD0 U767 ( .I(n791), .Z(n790) );
  BUFFD0 U768 ( .I(n792), .Z(n791) );
  BUFFD0 U769 ( .I(n793), .Z(n792) );
  BUFFD0 U770 ( .I(n794), .Z(n793) );
  BUFFD0 U771 ( .I(n795), .Z(n794) );
  BUFFD0 U772 ( .I(n796), .Z(n795) );
  BUFFD0 U773 ( .I(n797), .Z(n796) );
  BUFFD0 U774 ( .I(n798), .Z(n797) );
  BUFFD0 U775 ( .I(n799), .Z(n798) );
  BUFFD0 U776 ( .I(n800), .Z(n799) );
  BUFFD0 U777 ( .I(n801), .Z(n800) );
  BUFFD0 U778 ( .I(n802), .Z(n801) );
  BUFFD0 U779 ( .I(n803), .Z(n802) );
  BUFFD0 U780 ( .I(n804), .Z(n803) );
  BUFFD0 U781 ( .I(n805), .Z(n804) );
  BUFFD0 U782 ( .I(n806), .Z(n805) );
  BUFFD0 U783 ( .I(n807), .Z(n806) );
  BUFFD0 U784 ( .I(n808), .Z(n807) );
  BUFFD0 U785 ( .I(n809), .Z(n808) );
  BUFFD0 U786 ( .I(n810), .Z(n809) );
  BUFFD0 U787 ( .I(n811), .Z(n810) );
  BUFFD0 U788 ( .I(n812), .Z(n811) );
  BUFFD0 U789 ( .I(n813), .Z(n812) );
  BUFFD0 U790 ( .I(n814), .Z(n813) );
  BUFFD0 U791 ( .I(n815), .Z(n814) );
  BUFFD0 U792 ( .I(n816), .Z(n815) );
  BUFFD0 U793 ( .I(n817), .Z(n816) );
  BUFFD0 U794 ( .I(n818), .Z(n817) );
  BUFFD0 U795 ( .I(n819), .Z(n818) );
  BUFFD0 U796 ( .I(n820), .Z(n819) );
  BUFFD0 U797 ( .I(n821), .Z(n820) );
  BUFFD0 U798 ( .I(n822), .Z(n821) );
  BUFFD0 U799 ( .I(n823), .Z(n822) );
  BUFFD0 U800 ( .I(n824), .Z(n823) );
  BUFFD0 U801 ( .I(n825), .Z(n824) );
  BUFFD0 U802 ( .I(n826), .Z(n825) );
  BUFFD0 U803 ( .I(n827), .Z(n826) );
  BUFFD0 U804 ( .I(n828), .Z(n827) );
  BUFFD0 U805 ( .I(n829), .Z(n828) );
  BUFFD0 U806 ( .I(n100), .Z(n829) );
  BUFFD0 U807 ( .I(n78), .Z(n830) );
  BUFFD0 U808 ( .I(n79), .Z(n831) );
  BUFFD0 U809 ( .I(n833), .Z(n832) );
  BUFFD0 U810 ( .I(n834), .Z(n833) );
  BUFFD0 U811 ( .I(n835), .Z(n834) );
  BUFFD0 U812 ( .I(n836), .Z(n835) );
  BUFFD0 U813 ( .I(n837), .Z(n836) );
  BUFFD0 U814 ( .I(n838), .Z(n837) );
  BUFFD0 U815 ( .I(n839), .Z(n838) );
  BUFFD0 U816 ( .I(n840), .Z(n839) );
  BUFFD0 U817 ( .I(n841), .Z(n840) );
  BUFFD0 U818 ( .I(n842), .Z(n841) );
  BUFFD0 U819 ( .I(n843), .Z(n842) );
  BUFFD0 U820 ( .I(n844), .Z(n843) );
  BUFFD0 U821 ( .I(n845), .Z(n844) );
  BUFFD0 U822 ( .I(n846), .Z(n845) );
  BUFFD0 U823 ( .I(n847), .Z(n846) );
  BUFFD0 U824 ( .I(n848), .Z(n847) );
  BUFFD0 U825 ( .I(n849), .Z(n848) );
  BUFFD0 U826 ( .I(n850), .Z(n849) );
  BUFFD0 U827 ( .I(n851), .Z(n850) );
  BUFFD0 U828 ( .I(n852), .Z(n851) );
  BUFFD0 U829 ( .I(n853), .Z(n852) );
  BUFFD0 U830 ( .I(n854), .Z(n853) );
  BUFFD0 U831 ( .I(n855), .Z(n854) );
  BUFFD0 U832 ( .I(n856), .Z(n855) );
  BUFFD0 U833 ( .I(n857), .Z(n856) );
  BUFFD0 U834 ( .I(n858), .Z(n857) );
  BUFFD0 U835 ( .I(n859), .Z(n858) );
  BUFFD0 U836 ( .I(n860), .Z(n859) );
  BUFFD0 U837 ( .I(n861), .Z(n860) );
  BUFFD0 U838 ( .I(n862), .Z(n861) );
  BUFFD0 U839 ( .I(n863), .Z(n862) );
  BUFFD0 U840 ( .I(n864), .Z(n863) );
  BUFFD0 U841 ( .I(n865), .Z(n864) );
  BUFFD0 U842 ( .I(n866), .Z(n865) );
  BUFFD0 U843 ( .I(n867), .Z(n866) );
  BUFFD0 U844 ( .I(n868), .Z(n867) );
  BUFFD0 U845 ( .I(n869), .Z(n868) );
  BUFFD0 U846 ( .I(n870), .Z(n869) );
  BUFFD0 U847 ( .I(n871), .Z(n870) );
  BUFFD0 U848 ( .I(n872), .Z(n871) );
  BUFFD0 U849 ( .I(n873), .Z(n872) );
  BUFFD0 U850 ( .I(n874), .Z(n873) );
  BUFFD0 U851 ( .I(n875), .Z(n874) );
  BUFFD0 U852 ( .I(n876), .Z(n875) );
  BUFFD0 U853 ( .I(n877), .Z(n876) );
  BUFFD0 U854 ( .I(n878), .Z(n877) );
  BUFFD0 U855 ( .I(n879), .Z(n878) );
  BUFFD0 U856 ( .I(n880), .Z(n879) );
  BUFFD0 U857 ( .I(n881), .Z(n880) );
  BUFFD0 U858 ( .I(n882), .Z(n881) );
  BUFFD0 U859 ( .I(n883), .Z(n882) );
  BUFFD0 U860 ( .I(n105), .Z(n883) );
  ND2D8 U861 ( .A1(n1695), .A2(ReadReq), .ZN(n1696) );
  BUFFD0 U862 ( .I(n82), .Z(n884) );
  BUFFD0 U863 ( .I(n886), .Z(n885) );
  BUFFD0 U864 ( .I(n887), .Z(n886) );
  BUFFD0 U865 ( .I(n888), .Z(n887) );
  BUFFD0 U866 ( .I(n889), .Z(n888) );
  BUFFD0 U867 ( .I(n890), .Z(n889) );
  BUFFD0 U868 ( .I(n891), .Z(n890) );
  BUFFD0 U869 ( .I(n892), .Z(n891) );
  BUFFD0 U870 ( .I(n893), .Z(n892) );
  BUFFD0 U871 ( .I(n894), .Z(n893) );
  BUFFD0 U872 ( .I(n895), .Z(n894) );
  BUFFD0 U873 ( .I(n896), .Z(n895) );
  BUFFD0 U874 ( .I(n897), .Z(n896) );
  BUFFD0 U875 ( .I(n898), .Z(n897) );
  BUFFD0 U876 ( .I(n899), .Z(n898) );
  BUFFD0 U877 ( .I(n900), .Z(n899) );
  BUFFD0 U878 ( .I(n901), .Z(n900) );
  BUFFD0 U879 ( .I(n902), .Z(n901) );
  BUFFD0 U880 ( .I(n903), .Z(n902) );
  BUFFD0 U881 ( .I(n904), .Z(n903) );
  BUFFD0 U882 ( .I(n905), .Z(n904) );
  BUFFD0 U883 ( .I(n906), .Z(n905) );
  BUFFD0 U884 ( .I(n907), .Z(n906) );
  BUFFD0 U885 ( .I(n908), .Z(n907) );
  BUFFD0 U886 ( .I(n909), .Z(n908) );
  BUFFD0 U887 ( .I(n910), .Z(n909) );
  BUFFD0 U888 ( .I(n911), .Z(n910) );
  BUFFD0 U889 ( .I(n912), .Z(n911) );
  BUFFD0 U890 ( .I(n913), .Z(n912) );
  BUFFD0 U891 ( .I(n914), .Z(n913) );
  BUFFD0 U892 ( .I(n915), .Z(n914) );
  BUFFD0 U893 ( .I(n916), .Z(n915) );
  BUFFD0 U894 ( .I(n917), .Z(n916) );
  BUFFD0 U895 ( .I(n918), .Z(n917) );
  BUFFD0 U896 ( .I(n919), .Z(n918) );
  BUFFD0 U897 ( .I(n920), .Z(n919) );
  BUFFD0 U898 ( .I(n921), .Z(n920) );
  BUFFD0 U899 ( .I(n922), .Z(n921) );
  BUFFD0 U900 ( .I(n923), .Z(n922) );
  BUFFD0 U901 ( .I(n924), .Z(n923) );
  BUFFD0 U902 ( .I(n925), .Z(n924) );
  BUFFD0 U903 ( .I(n926), .Z(n925) );
  BUFFD0 U904 ( .I(n927), .Z(n926) );
  BUFFD0 U905 ( .I(n928), .Z(n927) );
  BUFFD0 U906 ( .I(n929), .Z(n928) );
  BUFFD0 U907 ( .I(n930), .Z(n929) );
  BUFFD0 U908 ( .I(n931), .Z(n930) );
  BUFFD0 U909 ( .I(n932), .Z(n931) );
  BUFFD0 U910 ( .I(n936), .Z(n932) );
  BUFFD0 U911 ( .I(n1710), .Z(n933) );
  CKBXD0 U912 ( .I(n655), .Z(n934) );
  CKBD0 U913 ( .CLK(n933), .C(n935) );
  BUFFD0 U914 ( .I(n103), .Z(n936) );
  BUFFD0 U915 ( .I(n938), .Z(n937) );
  BUFFD0 U916 ( .I(n939), .Z(n938) );
  BUFFD0 U917 ( .I(n940), .Z(n939) );
  BUFFD0 U918 ( .I(n941), .Z(n940) );
  BUFFD0 U919 ( .I(n942), .Z(n941) );
  BUFFD0 U920 ( .I(n943), .Z(n942) );
  BUFFD0 U921 ( .I(n944), .Z(n943) );
  BUFFD0 U922 ( .I(n945), .Z(n944) );
  BUFFD0 U923 ( .I(n946), .Z(n945) );
  BUFFD0 U924 ( .I(n947), .Z(n946) );
  BUFFD0 U925 ( .I(n948), .Z(n947) );
  BUFFD0 U926 ( .I(n949), .Z(n948) );
  BUFFD0 U927 ( .I(n950), .Z(n949) );
  BUFFD0 U928 ( .I(n951), .Z(n950) );
  BUFFD0 U929 ( .I(n952), .Z(n951) );
  BUFFD0 U930 ( .I(n953), .Z(n952) );
  BUFFD0 U931 ( .I(n954), .Z(n953) );
  BUFFD0 U932 ( .I(n955), .Z(n954) );
  BUFFD0 U933 ( .I(n956), .Z(n955) );
  BUFFD0 U934 ( .I(n957), .Z(n956) );
  BUFFD0 U935 ( .I(n958), .Z(n957) );
  BUFFD0 U936 ( .I(n959), .Z(n958) );
  BUFFD0 U937 ( .I(n960), .Z(n959) );
  BUFFD0 U938 ( .I(n961), .Z(n960) );
  BUFFD0 U939 ( .I(n962), .Z(n961) );
  BUFFD0 U940 ( .I(n963), .Z(n962) );
  BUFFD0 U941 ( .I(n964), .Z(n963) );
  BUFFD0 U942 ( .I(n965), .Z(n964) );
  BUFFD0 U943 ( .I(n966), .Z(n965) );
  BUFFD0 U944 ( .I(n967), .Z(n966) );
  BUFFD0 U945 ( .I(n968), .Z(n967) );
  BUFFD0 U946 ( .I(n969), .Z(n968) );
  BUFFD0 U947 ( .I(n970), .Z(n969) );
  BUFFD0 U948 ( .I(n971), .Z(n970) );
  BUFFD0 U949 ( .I(n972), .Z(n971) );
  BUFFD0 U950 ( .I(n973), .Z(n972) );
  BUFFD0 U951 ( .I(n974), .Z(n973) );
  BUFFD0 U952 ( .I(n975), .Z(n974) );
  BUFFD0 U953 ( .I(n976), .Z(n975) );
  BUFFD0 U954 ( .I(n977), .Z(n976) );
  BUFFD0 U955 ( .I(n978), .Z(n977) );
  BUFFD0 U956 ( .I(n979), .Z(n978) );
  BUFFD0 U957 ( .I(n980), .Z(n979) );
  BUFFD0 U958 ( .I(n1767), .Z(n980) );
  BUFFD0 U959 ( .I(ReadAddr[3]), .Z(n981) );
  CKBD0 U960 ( .CLK(N169), .C(n1018) );
  BUFFD0 U961 ( .I(ReadAddr[0]), .Z(n982) );
  BUFFD0 U962 ( .I(n982), .Z(n983) );
  BUFFD0 U963 ( .I(n983), .Z(n984) );
  BUFFD0 U964 ( .I(n984), .Z(n985) );
  BUFFD0 U965 ( .I(n985), .Z(n986) );
  BUFFD0 U966 ( .I(n986), .Z(n987) );
  BUFFD0 U967 ( .I(n987), .Z(n988) );
  BUFFD0 U968 ( .I(n988), .Z(n989) );
  BUFFD0 U969 ( .I(n989), .Z(n990) );
  BUFFD0 U970 ( .I(n990), .Z(n991) );
  BUFFD0 U971 ( .I(n991), .Z(n992) );
  BUFFD0 U972 ( .I(n992), .Z(n993) );
  BUFFD0 U973 ( .I(n993), .Z(n994) );
  BUFFD0 U974 ( .I(n994), .Z(n995) );
  BUFFD0 U975 ( .I(n995), .Z(n996) );
  BUFFD0 U976 ( .I(n996), .Z(n997) );
  BUFFD0 U977 ( .I(n997), .Z(n998) );
  BUFFD0 U978 ( .I(n998), .Z(n999) );
  BUFFD0 U979 ( .I(n999), .Z(n1000) );
  BUFFD0 U980 ( .I(n1000), .Z(n1001) );
  BUFFD0 U981 ( .I(n1001), .Z(n1002) );
  BUFFD0 U982 ( .I(n1002), .Z(n1003) );
  BUFFD0 U983 ( .I(n1003), .Z(n1004) );
  BUFFD0 U984 ( .I(n1004), .Z(n1005) );
  BUFFD0 U985 ( .I(n1005), .Z(n1006) );
  BUFFD0 U986 ( .I(n1006), .Z(n1007) );
  BUFFD0 U987 ( .I(n1007), .Z(n1008) );
  BUFFD0 U988 ( .I(n1008), .Z(n1009) );
  BUFFD0 U989 ( .I(n1009), .Z(n1010) );
  BUFFD0 U990 ( .I(n1010), .Z(n1011) );
  BUFFD0 U991 ( .I(n1011), .Z(n1012) );
  BUFFD0 U992 ( .I(n1012), .Z(n1013) );
  BUFFD0 U993 ( .I(n1013), .Z(n1014) );
  BUFFD0 U994 ( .I(n1014), .Z(n1015) );
  BUFFD0 U995 ( .I(n1015), .Z(n1016) );
  BUFFD0 U996 ( .I(n1016), .Z(n1017) );
  BUFFD0 U997 ( .I(n1017), .Z(n1019) );
  BUFFD0 U998 ( .I(n1019), .Z(n1020) );
  BUFFD0 U999 ( .I(n1020), .Z(n1021) );
  BUFFD0 U1000 ( .I(n1021), .Z(n1022) );
  BUFFD0 U1001 ( .I(n1022), .Z(n1023) );
  BUFFD0 U1002 ( .I(N49), .Z(n1024) );
  BUFFD0 U1003 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1004 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1005 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1006 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1007 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1008 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1009 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1010 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1011 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1012 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1013 ( .I(n1036), .Z(n1035) );
  BUFFD0 U1014 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1015 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1016 ( .I(n1039), .Z(n1038) );
  BUFFD0 U1017 ( .I(n1040), .Z(n1039) );
  BUFFD0 U1018 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1019 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1020 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1021 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1022 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1023 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1024 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1025 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1026 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1027 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1028 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1029 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1030 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1031 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1032 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1033 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1034 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1035 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1036 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1037 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1038 ( .I(n1061), .Z(n1060) );
  BUFFD0 U1039 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1040 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1041 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1042 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1043 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1044 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1045 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1046 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1047 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1048 ( .I(n1766), .Z(n1070) );
  BUFFD0 U1049 ( .I(n1779), .Z(ReadCmd) );
  INR2XD4 U1050 ( .A1(N47), .B1(n1697), .ZN(N53) );
  BUFFD0 U1051 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1052 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1053 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1054 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1055 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1056 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1057 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1058 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1059 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1060 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1061 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1062 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1063 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1064 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1065 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1066 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1067 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1068 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1069 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1070 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1071 ( .I(n1093), .Z(n1092) );
  BUFFD0 U1072 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1073 ( .I(n1095), .Z(n1094) );
  BUFFD0 U1074 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1075 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1076 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1077 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1078 ( .I(n1100), .Z(n1099) );
  BUFFD0 U1079 ( .I(n1101), .Z(n1100) );
  BUFFD0 U1080 ( .I(n1102), .Z(n1101) );
  BUFFD0 U1081 ( .I(n1103), .Z(n1102) );
  BUFFD0 U1082 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1083 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1084 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1085 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1086 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1087 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1088 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1089 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1090 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1091 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1092 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1093 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1094 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1095 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1096 ( .I(N53), .Z(n1117) );
  BUFFD0 U1097 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1098 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1099 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1100 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1101 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1102 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1103 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1104 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1105 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1106 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1107 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1108 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1109 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1110 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1111 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1112 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1113 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1114 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1115 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1116 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1117 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1118 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1119 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1120 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1121 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1122 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1123 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1124 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1125 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1126 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1127 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1128 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1129 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1130 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1131 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1132 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1133 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1134 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1135 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1136 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1137 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1138 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1139 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1140 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1141 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1142 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1143 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1144 ( .I(N50), .Z(n1165) );
  BUFFD0 U1145 ( .I(n1517), .Z(n1166) );
  BUFFD0 U1146 ( .I(n1692), .Z(n1167) );
  BUFFD0 U1147 ( .I(n1167), .Z(n1168) );
  BUFFD0 U1148 ( .I(n1168), .Z(n1169) );
  BUFFD0 U1149 ( .I(n1169), .Z(n1170) );
  BUFFD0 U1150 ( .I(n1170), .Z(n1171) );
  BUFFD0 U1151 ( .I(n1171), .Z(n1172) );
  BUFFD0 U1152 ( .I(n1172), .Z(n1173) );
  BUFFD0 U1153 ( .I(n1173), .Z(n1174) );
  BUFFD0 U1154 ( .I(n1174), .Z(n1175) );
  BUFFD0 U1155 ( .I(n1175), .Z(n1176) );
  BUFFD0 U1156 ( .I(n1176), .Z(n1177) );
  BUFFD0 U1157 ( .I(n1177), .Z(n1178) );
  BUFFD0 U1158 ( .I(n1178), .Z(n1179) );
  BUFFD0 U1159 ( .I(n1179), .Z(n1180) );
  BUFFD0 U1160 ( .I(n1180), .Z(n1181) );
  BUFFD0 U1161 ( .I(n1181), .Z(n1182) );
  BUFFD0 U1162 ( .I(n1182), .Z(n1183) );
  BUFFD0 U1163 ( .I(n1183), .Z(n1184) );
  BUFFD0 U1164 ( .I(n1184), .Z(n1185) );
  BUFFD0 U1165 ( .I(n1185), .Z(n1186) );
  BUFFD0 U1166 ( .I(n1186), .Z(n1187) );
  BUFFD0 U1167 ( .I(n1187), .Z(n1188) );
  BUFFD0 U1168 ( .I(n1188), .Z(n1189) );
  BUFFD0 U1169 ( .I(n1189), .Z(n1190) );
  BUFFD0 U1170 ( .I(n1190), .Z(n1191) );
  BUFFD0 U1171 ( .I(n1191), .Z(n1192) );
  BUFFD0 U1172 ( .I(n1192), .Z(n1193) );
  BUFFD0 U1173 ( .I(n1193), .Z(n1194) );
  BUFFD0 U1174 ( .I(n1194), .Z(n1195) );
  BUFFD0 U1175 ( .I(n1195), .Z(n1196) );
  BUFFD0 U1176 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1177 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1178 ( .I(n1693), .Z(n1199) );
  BUFFD0 U1179 ( .I(n1206), .Z(n1200) );
  BUFFD0 U1180 ( .I(N75), .Z(n1201) );
  BUFFD0 U1181 ( .I(n1201), .Z(n1202) );
  BUFFD0 U1182 ( .I(n1202), .Z(n1203) );
  BUFFD0 U1183 ( .I(n1203), .Z(n1204) );
  BUFFD0 U1184 ( .I(n1204), .Z(n1205) );
  BUFFD0 U1185 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1186 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1187 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1188 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1189 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1190 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1191 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1192 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1193 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1194 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1195 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1196 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1197 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1198 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1199 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1200 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1201 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1202 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1203 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1204 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1205 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1206 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1207 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1208 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1209 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1210 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1211 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1212 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1213 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1214 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1215 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1216 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1217 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1218 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1219 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1220 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1221 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1222 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1223 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1224 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1225 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1226 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1227 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1228 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1229 ( .I(n1251), .Z(n1250) );
  BUFFD0 U1230 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1231 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1232 ( .I(n1205), .Z(n1253) );
  BUFFD0 U1233 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1234 ( .I(n1683), .Z(n1255) );
  BUFFD0 U1235 ( .I(N74), .Z(n1256) );
  BUFFD0 U1236 ( .I(n1256), .Z(n1257) );
  BUFFD0 U1237 ( .I(n1257), .Z(n1258) );
  BUFFD0 U1238 ( .I(n1258), .Z(n1259) );
  BUFFD0 U1239 ( .I(n1259), .Z(n1260) );
  BUFFD0 U1240 ( .I(n1260), .Z(n1261) );
  BUFFD0 U1241 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1242 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1243 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1244 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1245 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1246 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1247 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1248 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1249 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1250 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1251 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1252 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1253 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1254 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1255 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1256 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1257 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1258 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1259 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1260 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1261 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1262 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1263 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1264 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1265 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1266 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1267 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1268 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1269 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1270 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1271 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1272 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1273 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1274 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1275 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1276 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1277 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1278 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1279 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1280 ( .I(n1302), .Z(n1301) );
  BUFFD0 U1281 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1282 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1283 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1284 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1285 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1286 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1287 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1288 ( .I(n1261), .Z(n1309) );
  BUFFD0 U1289 ( .I(n1777), .Z(n1310) );
  BUFFD0 U1290 ( .I(n1310), .Z(n1311) );
  INVD0 U1291 ( .I(n1311), .ZN(n1681) );
  INVD0 U1292 ( .I(N68), .ZN(n1748) );
  BUFFD0 U1293 ( .I(N73), .Z(n1312) );
  BUFFD0 U1294 ( .I(n1312), .Z(n1313) );
  BUFFD0 U1295 ( .I(n1313), .Z(n1314) );
  BUFFD0 U1296 ( .I(n1314), .Z(n1315) );
  BUFFD0 U1297 ( .I(n1315), .Z(n1316) );
  BUFFD0 U1298 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1299 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1300 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1301 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1302 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1303 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1304 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1305 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1306 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1307 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1308 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1309 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1310 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1311 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1312 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1313 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1314 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1315 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1316 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1317 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1318 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1319 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1320 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1321 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1322 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1323 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1324 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1325 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1326 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1327 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1328 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1329 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1330 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1331 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1332 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1333 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1334 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1335 ( .I(n1355), .Z(n1354) );
  BUFFD0 U1336 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1337 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1338 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1339 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1340 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1341 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1342 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1343 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1344 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1345 ( .I(n1316), .Z(n1364) );
  BUFFD0 U1346 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1347 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1348 ( .I(n1679), .Z(n1367) );
  INVD4 U1349 ( .I(N67), .ZN(n1775) );
  BUFFD0 U1350 ( .I(N72), .Z(n1368) );
  BUFFD0 U1351 ( .I(n1368), .Z(n1369) );
  BUFFD0 U1352 ( .I(n1369), .Z(n1370) );
  BUFFD0 U1353 ( .I(n1370), .Z(n1371) );
  BUFFD0 U1354 ( .I(n1371), .Z(n1372) );
  BUFFD0 U1355 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1356 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1357 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1358 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1359 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1360 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1361 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1362 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1363 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1364 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1365 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1366 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1367 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1368 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1369 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1370 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1371 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1372 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1373 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1374 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1375 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1376 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1377 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1378 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1379 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1380 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1381 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1382 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1383 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1384 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1385 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1386 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1387 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1388 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1389 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1390 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1391 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1392 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1393 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1394 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1395 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1396 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1397 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1398 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1399 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1400 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1401 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1402 ( .I(n1372), .Z(n1420) );
  BUFFD0 U1403 ( .I(\add_306/carry[2] ), .Z(n1421) );
  BUFFD0 U1404 ( .I(n1421), .Z(n1422) );
  INVD0 U1405 ( .I(n1422), .ZN(n1677) );
  BUFFD0 U1406 ( .I(n1427), .Z(n1423) );
  BUFFD0 U1407 ( .I(N71), .Z(n1424) );
  BUFFD0 U1408 ( .I(n1424), .Z(n1425) );
  BUFFD0 U1409 ( .I(n1425), .Z(n1426) );
  BUFFD0 U1410 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1411 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1412 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1413 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1414 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1415 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1416 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1417 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1418 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1419 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1420 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1421 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1422 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1423 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1424 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1425 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1426 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1427 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1428 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1429 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1430 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1431 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1432 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1433 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1434 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1435 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1436 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1437 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1438 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1439 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1440 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1441 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1442 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1443 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1444 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1445 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1446 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1447 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1448 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1449 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1450 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1451 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1452 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1453 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1454 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1455 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1456 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1457 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1458 ( .I(n1426), .Z(n1475) );
  BUFFD0 U1459 ( .I(n1018), .Z(n1476) );
  BUFFD0 U1460 ( .I(n1476), .Z(n1477) );
  BUFFD0 U1461 ( .I(n1477), .Z(n1478) );
  INVD0 U1462 ( .I(n1478), .ZN(n1674) );
  BUFFD0 U1463 ( .I(N76), .Z(n1479) );
  BUFFD0 U1464 ( .I(n1479), .Z(n1480) );
  BUFFD0 U1465 ( .I(n1480), .Z(n1481) );
  BUFFD0 U1466 ( .I(n1481), .Z(n1482) );
  BUFFD0 U1467 ( .I(n1482), .Z(n1483) );
  BUFFD0 U1468 ( .I(n1483), .Z(n1484) );
  BUFFD0 U1469 ( .I(n1484), .Z(n1485) );
  BUFFD0 U1470 ( .I(n1485), .Z(n1486) );
  BUFFD0 U1471 ( .I(n1486), .Z(n1487) );
  BUFFD0 U1472 ( .I(n1487), .Z(n1488) );
  BUFFD0 U1473 ( .I(n1488), .Z(n1489) );
  BUFFD0 U1474 ( .I(n1489), .Z(n1490) );
  BUFFD0 U1475 ( .I(n1490), .Z(n1491) );
  BUFFD0 U1476 ( .I(n1491), .Z(n1492) );
  BUFFD0 U1477 ( .I(n1492), .Z(n1493) );
  BUFFD0 U1478 ( .I(n1493), .Z(n1494) );
  BUFFD0 U1479 ( .I(n1494), .Z(n1495) );
  BUFFD0 U1480 ( .I(n1495), .Z(n1496) );
  BUFFD0 U1481 ( .I(n1496), .Z(n1497) );
  BUFFD0 U1482 ( .I(n1497), .Z(n1498) );
  BUFFD0 U1483 ( .I(n1498), .Z(n1499) );
  BUFFD0 U1484 ( .I(n1499), .Z(n1500) );
  BUFFD0 U1485 ( .I(n1500), .Z(n1501) );
  BUFFD0 U1486 ( .I(n1501), .Z(n1502) );
  BUFFD0 U1487 ( .I(n1502), .Z(n1503) );
  BUFFD0 U1488 ( .I(n1503), .Z(n1504) );
  BUFFD0 U1489 ( .I(n1504), .Z(n1505) );
  BUFFD0 U1490 ( .I(n1505), .Z(n1506) );
  BUFFD0 U1491 ( .I(n1506), .Z(n1507) );
  BUFFD0 U1492 ( .I(n1507), .Z(n1508) );
  BUFFD0 U1493 ( .I(n1508), .Z(n1509) );
  BUFFD0 U1494 ( .I(n1509), .Z(n1510) );
  BUFFD0 U1495 ( .I(n1510), .Z(n1511) );
  BUFFD0 U1496 ( .I(n1511), .Z(n1512) );
  BUFFD0 U1497 ( .I(n1512), .Z(n1513) );
  BUFFD0 U1498 ( .I(n1513), .Z(n1514) );
  CKBD0 U1499 ( .CLK(n1514), .C(n1515) );
  ND3D8 U1500 ( .A1(n1689), .A2(n1517), .A3(n1711), .ZN(N76) );
  BUFFD0 U1501 ( .I(n1518), .Z(n1516) );
  BUFFD0 U1502 ( .I(n1519), .Z(n1517) );
  BUFFD0 U1503 ( .I(n1520), .Z(n1518) );
  BUFFD0 U1504 ( .I(n1521), .Z(n1519) );
  BUFFD0 U1505 ( .I(n1522), .Z(n1520) );
  BUFFD0 U1506 ( .I(n1523), .Z(n1521) );
  BUFFD0 U1507 ( .I(n1524), .Z(n1522) );
  BUFFD0 U1508 ( .I(n1529), .Z(n1523) );
  BUFFD0 U1509 ( .I(n1527), .Z(n1524) );
  CKNXD16 U1510 ( .I(n1525), .ZN(n1526) );
  INVD0 U1511 ( .I(n1731), .ZN(n1525) );
  BUFFD0 U1512 ( .I(n1530), .Z(n1527) );
  BUFFD0 U1513 ( .I(n1526), .Z(n1528) );
  BUFFD0 U1514 ( .I(n1531), .Z(n1529) );
  BUFFD0 U1515 ( .I(n1532), .Z(n1530) );
  BUFFD0 U1516 ( .I(n1533), .Z(n1531) );
  BUFFD0 U1517 ( .I(n1534), .Z(n1532) );
  BUFFD0 U1518 ( .I(n1535), .Z(n1533) );
  BUFFD0 U1519 ( .I(n1536), .Z(n1534) );
  BUFFD0 U1520 ( .I(n1537), .Z(n1535) );
  BUFFD0 U1521 ( .I(CurState[1]), .Z(n1536) );
  BUFFD0 U1522 ( .I(n1196), .Z(n1537) );
  CKND2D0 U1523 ( .A1(n1516), .A2(n1528), .ZN(n1689) );
  BUFFD0 U1524 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1525 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1526 ( .I(n1543), .Z(n1540) );
  BUFFD0 U1527 ( .I(n91), .Z(n1541) );
  BUFFD0 U1528 ( .I(n1541), .Z(n1542) );
  BUFFD0 U1529 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1530 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1531 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1532 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1533 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1534 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1535 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1536 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1537 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1538 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1539 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1540 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1541 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1542 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1543 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1544 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1545 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1546 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1547 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1548 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1549 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1550 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1551 ( .I(n1566), .Z(n1565) );
  BUFFD0 U1552 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1553 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1554 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1555 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1556 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1557 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1558 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1559 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1560 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1561 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1562 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1563 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1564 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1565 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1566 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1567 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1568 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1569 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1570 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1571 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1572 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1573 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1574 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1575 ( .I(n1592), .Z(n1589) );
  BUFFD0 U1576 ( .I(n1542), .Z(n1590) );
  BUFFD0 U1577 ( .I(n1590), .Z(n1591) );
  CKBD0 U1578 ( .CLK(n1593), .C(n1592) );
  OAI31D4 U1579 ( .A1(n1692), .A2(WriteReq), .A3(Reset), .B(n5), .ZN(n91) );
  BUFFD0 U1580 ( .I(n1599), .Z(n1594) );
  OAI32XD4 U1581 ( .A1(n1689), .A2(Reset), .A3(ReadReq), .B1(n76), .B2(n1690), 
        .ZN(n93) );
  BUFFD0 U1582 ( .I(n93), .Z(n1595) );
  BUFFD0 U1583 ( .I(n1595), .Z(n1596) );
  BUFFD0 U1584 ( .I(n1596), .Z(n1597) );
  BUFFD0 U1585 ( .I(n1597), .Z(n1598) );
  BUFFD0 U1586 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1587 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1588 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1589 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1590 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1591 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1592 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1593 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1594 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1595 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1596 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1597 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1598 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1599 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1600 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1601 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1602 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1603 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1604 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1605 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1606 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1607 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1608 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1609 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1610 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1611 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1612 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1613 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1614 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1615 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1616 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1617 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1618 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1619 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1620 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1621 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1622 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1623 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1624 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1625 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1626 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1627 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1628 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1629 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1630 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1631 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1632 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1633 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1634 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1635 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1636 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1637 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1638 ( .I(n1598), .Z(n1651) );
  CKBXD0 U1639 ( .I(n6), .Z(n1652) );
  CKNXD16 U1640 ( .I(n1652), .ZN(EmptyFIFO) );
  CKBD0 U1641 ( .CLK(n1656), .C(n1654) );
  CKNXD16 U1642 ( .I(n1654), .ZN(FullFIFO) );
  CKND0 U1643 ( .CLK(n1778), .CN(n1656) );
  CKNXD4 U1644 ( .I(n6), .ZN(n1657) );
  INVD1 U1645 ( .I(N43), .ZN(n1675) );
  INVD1 U1646 ( .I(Reset), .ZN(n1672) );
  INVD1 U1647 ( .I(n1674), .ZN(ReadAddr[0]) );
  INVD1 U1648 ( .I(n1677), .ZN(ReadAddr[1]) );
  INVD1 U1649 ( .I(n1681), .ZN(ReadAddr[3]) );
  INVD1 U1650 ( .I(n1365), .ZN(ReadAddr[2]) );
  INVD1 U1651 ( .I(n1254), .ZN(ReadAddr[4]) );
  CKXOR2D0 U1652 ( .A1(ReadAddr[4]), .A2(\add_306/carry[4] ), .Z(N173) );
  AN2D0 U1653 ( .A1(ReadAddr[3]), .A2(\add_306/carry[3] ), .Z(
        \add_306/carry[4] ) );
  CKXOR2D0 U1654 ( .A1(\add_306/carry[3] ), .A2(ReadAddr[3]), .Z(N172) );
  AN2D0 U1655 ( .A1(ReadAddr[2]), .A2(ReadAddr[1]), .Z(\add_306/carry[3] ) );
  CKXOR2D0 U1656 ( .A1(ReadAddr[1]), .A2(ReadAddr[2]), .Z(N171) );
  CKXOR2D0 U1657 ( .A1(WriteAddr[4]), .A2(\add_387/carry[4] ), .Z(N325) );
  AN2D0 U1658 ( .A1(WriteAddr[3]), .A2(\add_387/carry[3] ), .Z(
        \add_387/carry[4] ) );
  CKXOR2D0 U1659 ( .A1(\add_387/carry[3] ), .A2(WriteAddr[3]), .Z(N324) );
  AN2D0 U1660 ( .A1(WriteAddr[2]), .A2(\add_387/carry[2] ), .Z(
        \add_387/carry[3] ) );
  CKXOR2D0 U1661 ( .A1(\add_387/carry[2] ), .A2(WriteAddr[2]), .Z(N323) );
  MUX2ND0 U1662 ( .I0(n382), .I1(n1684), .S(n1685), .ZN(n99) );
  MUX2ND0 U1663 ( .I0(n438), .I1(n1686), .S(n1685), .ZN(n98) );
  MUX2ND0 U1664 ( .I0(n154), .I1(n1687), .S(n1685), .ZN(n97) );
  MUX2ND0 U1665 ( .I0(n495), .I1(n1683), .S(n1688), .ZN(n96) );
  MUX2ND0 U1666 ( .I0(n551), .I1(n1679), .S(n1688), .ZN(n95) );
  MUX2ND0 U1667 ( .I0(n211), .I1(n1681), .S(n1688), .ZN(n94) );
  AOI21D0 U1668 ( .A1(n1691), .A2(n1692), .B(Reset), .ZN(n1690) );
  MUX2ND0 U1669 ( .I0(n268), .I1(n1677), .S(n1688), .ZN(n92) );
  MUX2ND0 U1670 ( .I0(n325), .I1(n4), .S(n1685), .ZN(n90) );
  INR3D0 U1671 ( .A1(ReadReq), .B1(n1694), .B2(n1695), .ZN(n1688) );
  CKND0 U1672 ( .CLK(Reset), .CN(n106) );
  MUX2ND0 U1673 ( .I0(n1696), .I1(n1697), .S(n1694), .ZN(n105) );
  NR2D0 U1674 ( .A1(n1698), .A2(n1699), .ZN(n1694) );
  AN3D0 U1675 ( .A1(n1700), .A2(n1701), .A3(n1702), .Z(n1695) );
  NR3D0 U1676 ( .A1(n1703), .A2(n1704), .A3(n1705), .ZN(n1702) );
  CKXOR2D0 U1677 ( .A1(n1681), .A2(n211), .Z(n1705) );
  CKXOR2D0 U1678 ( .A1(n1677), .A2(n268), .Z(n1704) );
  CKXOR2D0 U1679 ( .A1(n1674), .A2(n89), .Z(n1703) );
  CKXOR2D0 U1680 ( .A1(n551), .A2(ReadAddr[2]), .Z(n1701) );
  CKXOR2D0 U1681 ( .A1(n495), .A2(ReadAddr[4]), .Z(n1700) );
  NR3D0 U1682 ( .A1(n1707), .A2(n1708), .A3(n1), .ZN(n1685) );
  NR2D0 U1683 ( .A1(n1698), .A2(n1712), .ZN(n1707) );
  AN3D0 U1684 ( .A1(n1713), .A2(n1714), .A3(n1715), .Z(n1708) );
  NR3D0 U1685 ( .A1(n1716), .A2(n1717), .A3(n1718), .ZN(n1715) );
  CKXOR2D0 U1686 ( .A1(n1687), .A2(n154), .Z(n1718) );
  CKXOR2D0 U1687 ( .A1(n4), .A2(n325), .Z(n1717) );
  CKXOR2D0 U1688 ( .A1(n1706), .A2(n87), .Z(n1716) );
  CKXOR2D0 U1689 ( .A1(n438), .A2(WriteAddr[2]), .Z(n1714) );
  CKXOR2D0 U1690 ( .A1(n382), .A2(WriteAddr[4]), .Z(n1713) );
  NR2D0 U1691 ( .A1(n1712), .A2(n1721), .ZN(n1719) );
  MUX2ND0 U1692 ( .I0(n1722), .I1(n1723), .S(CurState[1]), .ZN(n1721) );
  OAI21D0 U1693 ( .A1(n1724), .A2(n1725), .B(n1726), .ZN(n1723) );
  AOI31D0 U1694 ( .A1(n1727), .A2(n1728), .A3(n1729), .B(CurState[2]), .ZN(
        n1726) );
  OAI21D0 U1695 ( .A1(n1729), .A2(n1730), .B(n1731), .ZN(n1722) );
  CKND0 U1696 ( .CLK(n1732), .CN(n1730) );
  AN3D0 U1697 ( .A1(n1733), .A2(n1734), .A3(n1735), .Z(n1729) );
  NR3D0 U1698 ( .A1(n1736), .A2(n1737), .A3(n1738), .ZN(n1735) );
  CKXOR2D0 U1699 ( .A1(WriteAddr[3]), .A2(ReadAddr[3]), .Z(n1738) );
  CKXOR2D0 U1700 ( .A1(\add_387/carry[2] ), .A2(ReadAddr[1]), .Z(n1737) );
  CKXOR2D0 U1701 ( .A1(N321), .A2(ReadAddr[0]), .Z(n1736) );
  CKXOR2D0 U1702 ( .A1(ReadAddr[2]), .A2(n1686), .Z(n1734) );
  CKXOR2D0 U1703 ( .A1(ReadAddr[4]), .A2(n1684), .Z(n1733) );
  MUX2ND0 U1704 ( .I0(n1739), .I1(n715), .S(n1720), .ZN(n101) );
  AOI211D0 U1705 ( .A1(n1731), .A2(n1732), .B(n1699), .C(n1740), .ZN(n1739) );
  NR3D0 U1706 ( .A1(n1725), .A2(n1741), .A3(n1724), .ZN(n1740) );
  ND3D0 U1707 ( .A1(n1742), .A2(n1743), .A3(n1744), .ZN(n1725) );
  NR3D0 U1708 ( .A1(n1745), .A2(n1746), .A3(n1747), .ZN(n1744) );
  CKXOR2D0 U1709 ( .A1(ReadAddr[3]), .A2(N69), .Z(n1747) );
  CKXOR2D0 U1710 ( .A1(ReadAddr[1]), .A2(N67), .Z(n1746) );
  CKXOR2D0 U1711 ( .A1(ReadAddr[0]), .A2(N66), .Z(n1745) );
  CKXOR2D0 U1712 ( .A1(ReadAddr[2]), .A2(n1748), .Z(n1743) );
  CKXOR2D0 U1713 ( .A1(ReadAddr[4]), .A2(n1749), .Z(n1742) );
  CKND0 U1714 ( .CLK(n1689), .CN(n1699) );
  ND3D0 U1715 ( .A1(n1750), .A2(n1751), .A3(n1752), .ZN(n1732) );
  NR3D0 U1716 ( .A1(n1753), .A2(n1754), .A3(n1755), .ZN(n1752) );
  CKXOR2D0 U1717 ( .A1(ReadAddr[3]), .A2(N324), .Z(n1755) );
  CKXOR2D0 U1718 ( .A1(ReadAddr[1]), .A2(n4), .Z(n1754) );
  CKXOR2D0 U1719 ( .A1(ReadAddr[0]), .A2(N321), .Z(n1753) );
  CKXOR2D0 U1720 ( .A1(N323), .A2(n1679), .Z(n1751) );
  CKXOR2D0 U1721 ( .A1(N325), .A2(n1683), .Z(n1750) );
  MUX2ND0 U1722 ( .I0(n1756), .I1(n773), .S(n1720), .ZN(n100) );
  OA211D0 U1723 ( .A1(n1), .A2(n1692), .B(n1757), .C(n1758), .Z(n1720) );
  AOI21D0 U1724 ( .A1(CurState[0]), .A2(n1741), .B(n1698), .ZN(n1758) );
  MUX2ND0 U1725 ( .I0(CurState[2]), .I1(n1691), .S(n1741), .ZN(n1698) );
  CKND0 U1726 ( .CLK(CurState[1]), .CN(n1741) );
  OAI21D0 U1727 ( .A1(ReadReq), .A2(n1728), .B(CurState[2]), .ZN(n1757) );
  CKND0 U1728 ( .CLK(WriteReq), .CN(n1709) );
  AOI21D0 U1729 ( .A1(CurState[1]), .A2(n1759), .B(n1731), .ZN(n1756) );
  OAI21D0 U1730 ( .A1(n1693), .A2(n1727), .B(n1724), .ZN(n1759) );
  OAI31D0 U1731 ( .A1(n1760), .A2(n1761), .A3(n1762), .B(CurState[0]), .ZN(
        n1724) );
  CKXOR2D0 U1732 ( .A1(WriteAddr[4]), .A2(N47), .Z(n1762) );
  CKXOR2D0 U1733 ( .A1(WriteAddr[2]), .A2(N45), .Z(n1761) );
  ND3D0 U1734 ( .A1(n1763), .A2(n1764), .A3(n1765), .ZN(n1760) );
  CKXOR2D0 U1735 ( .A1(N321), .A2(n1675), .Z(n1765) );
  CKXOR2D0 U1736 ( .A1(\add_387/carry[2] ), .A2(n1766), .Z(n1764) );
  CKXOR2D0 U1737 ( .A1(WriteAddr[3]), .A2(n1767), .Z(n1763) );
  ND3D0 U1738 ( .A1(n1768), .A2(n1769), .A3(n1770), .ZN(n1727) );
  NR3D0 U1739 ( .A1(n1771), .A2(n1772), .A3(n1773), .ZN(n1770) );
  CKXOR2D0 U1740 ( .A1(WriteAddr[3]), .A2(N172), .Z(n1773) );
  CKXOR2D0 U1741 ( .A1(\add_387/carry[2] ), .A2(n1677), .Z(n1772) );
  CKXOR2D0 U1742 ( .A1(N321), .A2(ReadAddr[0]), .Z(n1771) );
  CKXOR2D0 U1743 ( .A1(N171), .A2(n1686), .Z(n1769) );
  CKXOR2D0 U1744 ( .A1(N173), .A2(n1684), .Z(n1768) );
  CKND2D0 U1745 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  OAI22D0 U1746 ( .A1(n1254), .A2(n1689), .B1(n1711), .B2(n1749), .ZN(N75) );
  CKND0 U1747 ( .CLK(N70), .CN(n1749) );
  CKND0 U1748 ( .CLK(N69), .CN(n1774) );
  OAI22D0 U1749 ( .A1(n1365), .A2(n1689), .B1(n1711), .B2(n1748), .ZN(N73) );
  OAI22D0 U1750 ( .A1(n1677), .A2(n1689), .B1(n1711), .B2(n1775), .ZN(N72) );
  OAI22D0 U1751 ( .A1(n1674), .A2(n1689), .B1(n1711), .B2(n1776), .ZN(N71) );
  CKND0 U1752 ( .CLK(N66), .CN(n1776) );
  CKND2D0 U1753 ( .A1(n934), .A2(n1689), .ZN(n1711) );
  CKND2D0 U1754 ( .A1(n1166), .A2(n1697), .ZN(N52) );
  NR2D0 U1755 ( .A1(n1697), .A2(n937), .ZN(N51) );
  CKND0 U1756 ( .CLK(N46), .CN(n1767) );
  INR2D0 U1757 ( .A1(N45), .B1(n1697), .ZN(N50) );
  NR2D0 U1758 ( .A1(n1697), .A2(n1025), .ZN(N49) );
  CKND0 U1759 ( .CLK(N44), .CN(n1766) );
  NR2D0 U1760 ( .A1(n1697), .A2(n1675), .ZN(N48) );
  CKND2D0 U1761 ( .A1(ReadCmd), .A2(n1166), .ZN(n1697) );
  CKND0 U1762 ( .CLK(n1712), .CN(n1692) );
  NR2D0 U1763 ( .A1(n1197), .A2(n1516), .ZN(n1712) );
  IND2D0 U1764 ( .A1(CurState[2]), .B1(n1728), .ZN(n1693) );
  CKND0 U1765 ( .CLK(CurState[0]), .CN(n1728) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, ClockR, ClockW, Dreadyr, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N85, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n107,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  XNR4D1 U18 ( .A1(n4706), .A2(n4704), .A3(n4711), .A4(n4708), .ZN(n84) );
  XOR4D1 U19 ( .A1(n4716), .A2(n4714), .A3(n4721), .A4(n4718), .Z(n83) );
  XOR4D1 U20 ( .A1(n4696), .A2(n4694), .A3(n4701), .A4(n4698), .Z(n80) );
  XOR4D1 U21 ( .A1(n4678), .A2(n4676), .A3(n4683), .A4(n4680), .Z(n77) );
  XNR4D1 U22 ( .A1(n4660), .A2(n4658), .A3(n4665), .A4(n4662), .ZN(n74) );
  XOR4D1 U27 ( .A1(n90), .A2(n3172), .A3(n91), .A4(n3798), .Z(n89) );
  XNR4D1 U28 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n91) );
  XNR4D1 U33 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n97) );
  XOR4D1 U34 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n96) );
  XNR4D1 U35 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .ZN(n93) );
  XNR4D1 U36 ( .A1(n3800), .A2(n3821), .A3(n3819), .A4(n3801), .ZN(n87) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(N85), .E(n4523), .CP(n4596), .CDN(n4476), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(n10), .E(n4523), .CP(n4596), .CDN(n4475), 
        .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(n45), .E(n4522), .CP(n4596), .CDN(n4475), 
        .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(n139), .E(n4523), .CP(n4596), .CDN(n4475), .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(n191), .E(n4522), .CP(n4596), .CDN(n4475), .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(n1565), .E(n4523), .CP(n4597), .CDN(
        n4475), .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(n1671), .E(n4522), .CP(n4597), .CDN(
        n4475), .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(n1619), .E(n4523), .CP(n4597), .CDN(
        n4475), .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(n245), .E(n4522), .CP(n4597), .CDN(n4475), .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(n299), .E(n4523), .CP(n4597), .CDN(n4475), .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n353), .E(n4522), .CP(n4597), .CDN(n4475), .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(n405), .E(n4522), .CP(n4597), .CDN(n4475), .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(n457), .E(n4522), .CP(n4597), .CDN(n4474), .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(n1), .E(n4522), .CP(n4597), .CDN(n4474), 
        .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(n4689), .E(n4522), .CP(n4597), .CDN(
        n4474), .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(n4686), .E(n4522), .CP(n4598), .CDN(
        n4474), .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(n669), .E(n4522), .CP(n4598), .CDN(n4474), .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n723), .E(n4522), .CP(n4598), .CDN(n4474), .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n775), .E(n4522), .CP(n4598), .CDN(n4474), .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(n827), .E(n4522), .CP(n4598), .CDN(n4474), .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n2), .E(n4522), .CP(n4598), .CDN(n4474), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(n4671), .E(n4522), .CP(n4598), .CDN(
        n4474), .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(n4668), .E(n4523), .CP(n4598), .CDN(
        n4474), .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n1039), .E(n4523), .CP(n4598), .CDN(n4473), .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(n1093), .E(n4523), .CP(n4598), .CDN(n4473), .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n1145), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n1197), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n3), .E(n4523), .CP(n4599), .CDN(n4473), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n4653), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(n4650), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n1428), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(n4645), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n1532), .E(n4523), .CP(n4599), .CDN(n4473), .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(n4576), .E(n4527), .CP(n4603), .CDN(
        n4470), .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(n10), .E(n4527), .CP(n4603), .CDN(n4469), 
        .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(n45), .E(n4526), .CP(n4603), .CDN(n4469), 
        .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(n139), .E(n4527), .CP(n4603), .CDN(n4469), .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(n191), .E(n4526), .CP(n4603), .CDN(n4469), .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(n1565), .E(n4527), .CP(n4603), .CDN(
        n4469), .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(n1671), .E(n4526), .CP(n4603), .CDN(
        n4469), .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(n1619), .E(n4527), .CP(n4603), .CDN(
        n4469), .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(n245), .E(n4526), .CP(n4603), .CDN(n4469), .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(n299), .E(n4527), .CP(n4604), .CDN(n4469), .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n353), .E(n4526), .CP(n4604), .CDN(n4469), .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(n405), .E(n4526), .CP(n4604), .CDN(n4469), .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(n457), .E(n4526), .CP(n4604), .CDN(n4468), .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(n5), .E(n4526), .CP(n4604), .CDN(n4468), 
        .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(n4689), .E(n4526), .CP(n4604), .CDN(
        n4468), .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(n4686), .E(n4526), .CP(n4604), .CDN(
        n4468), .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(n669), .E(n4526), .CP(n4604), .CDN(n4468), .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n723), .E(n4526), .CP(n4604), .CDN(n4468), .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n775), .E(n4526), .CP(n4604), .CDN(n4468), .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(n827), .E(n4526), .CP(n4605), .CDN(n4468), .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n6), .E(n4526), .CP(n4605), .CDN(n4468), 
        .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(n4671), .E(n4526), .CP(n4605), .CDN(
        n4468), .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(n4668), .E(n4527), .CP(n4605), .CDN(
        n4468), .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n1039), .E(n4527), .CP(n4605), .CDN(n4467), .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(n1093), .E(n4527), .CP(n4605), .CDN(n4467), .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n1145), .E(n4527), .CP(n4605), .CDN(n4467), .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n1197), .E(n4527), .CP(n4605), .CDN(n4467), .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n7), .E(n4527), .CP(n4605), .CDN(n4467), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n4653), .E(n4527), .CP(n4605), .CDN(n4467), .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(n4650), .E(n4527), .CP(n4606), .CDN(n4467), .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n1428), .E(n4527), .CP(n4606), .CDN(n4467), .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(n4645), .E(n4527), .CP(n4606), .CDN(n4467), .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n1532), .E(n4527), .CP(n4606), .CDN(n4467), .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(n4576), .E(n4515), .CP(n4583), .CDN(
        n4488), .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(n10), .E(n4515), .CP(n4583), .CDN(n4487), 
        .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(n45), .E(n4514), .CP(n4583), .CDN(n4487), 
        .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(n139), .E(n4515), .CP(n4583), .CDN(n4487), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(n191), .E(n4514), .CP(n4583), .CDN(n4487), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(n1565), .E(n4515), .CP(n4583), .CDN(
        n4487), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(n245), .E(n4514), .CP(n4584), .CDN(n4487), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(n299), .E(n4515), .CP(n4584), .CDN(n4487), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(n353), .E(n4514), .CP(n4584), .CDN(n4487), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(n405), .E(n4514), .CP(n4584), .CDN(n4487), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(n457), .E(n4514), .CP(n4584), .CDN(n4486), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(n5), .E(n4514), .CP(n4584), .CDN(n4486), 
        .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(n4689), .E(n4514), .CP(n4584), .CDN(
        n4486), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(n4686), .E(n4514), .CP(n4584), .CDN(
        n4486), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(n669), .E(n4514), .CP(n4584), .CDN(n4486), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(n723), .E(n4514), .CP(n4585), .CDN(n4486), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(n775), .E(n4514), .CP(n4585), .CDN(n4486), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(n827), .E(n4514), .CP(n4585), .CDN(n4486), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(n6), .E(n4514), .CP(n4585), .CDN(n4486), 
        .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(n4671), .E(n4514), .CP(n4585), .CDN(
        n4486), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(n4668), .E(n4515), .CP(n4585), .CDN(
        n4486), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(n1039), .E(n4515), .CP(n4585), .CDN(n4485), .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(n1093), .E(n4515), .CP(n4585), .CDN(n4485), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(n1145), .E(n4515), .CP(n4585), .CDN(n4485), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(n1197), .E(n4515), .CP(n4585), .CDN(n4485), .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(n7), .E(n4515), .CP(n4586), .CDN(n4485), 
        .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(n4653), .E(n4515), .CP(n4586), .CDN(n4485), .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(n4650), .E(n4515), .CP(n4586), .CDN(n4485), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(n1428), .E(n4515), .CP(n4586), .CDN(n4485), .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(n4645), .E(n4515), .CP(n4586), .CDN(n4485), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(n1532), .E(n4515), .CP(n4586), .CDN(n4485), .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n4576), .E(n4517), .CP(n4586), .CDN(
        n4485), .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(n10), .E(n4517), .CP(n4586), .CDN(n4484), 
        .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(n45), .E(n4516), .CP(n4586), .CDN(n4484), 
        .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(n139), .E(n4517), .CP(n4586), .CDN(n4484), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(n191), .E(n4516), .CP(n4587), .CDN(n4484), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(n1565), .E(n4517), .CP(n4587), .CDN(
        n4484), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(n245), .E(n4516), .CP(n4587), .CDN(n4484), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(n299), .E(n4517), .CP(n4587), .CDN(n4484), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(n353), .E(n4516), .CP(n4587), .CDN(n4484), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(n405), .E(n4516), .CP(n4587), .CDN(n4484), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(n457), .E(n4516), .CP(n4587), .CDN(n4483), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(n5), .E(n4516), .CP(n4587), .CDN(n4483), 
        .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(n4689), .E(n4516), .CP(n4588), .CDN(
        n4483), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(n4686), .E(n4516), .CP(n4588), .CDN(
        n4483), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(n669), .E(n4516), .CP(n4588), .CDN(n4483), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(n723), .E(n4516), .CP(n4588), .CDN(n4483), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(n775), .E(n4516), .CP(n4588), .CDN(n4483), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(n827), .E(n4516), .CP(n4588), .CDN(n4483), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(n6), .E(n4516), .CP(n4588), .CDN(n4483), 
        .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(n4671), .E(n4516), .CP(n4588), .CDN(
        n4483), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(n4668), .E(n4517), .CP(n4588), .CDN(
        n4483), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(n1039), .E(n4517), .CP(n4588), .CDN(n4482), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(n1093), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(n1145), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(n1197), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(n7), .E(n4517), .CP(n4589), .CDN(n4482), 
        .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(n4653), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(n4650), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(n1428), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(n4645), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(n1532), .E(n4517), .CP(n4589), .CDN(n4482), .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(n4576), .E(n4519), .CP(n4589), .CDN(
        n4482), .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(n10), .E(n4519), .CP(n4590), .CDN(n4481), 
        .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(n45), .E(n4518), .CP(n4590), .CDN(n4481), 
        .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(n139), .E(n4519), .CP(n4590), .CDN(n4481), .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(n191), .E(n4518), .CP(n4590), .CDN(n4481), .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(n245), .E(n4519), .CP(n4590), .CDN(n4481), .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(n299), .E(n4518), .CP(n4590), .CDN(n4481), .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n353), .E(n4519), .CP(n4590), .CDN(n4481), .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(n405), .E(n4518), .CP(n4591), .CDN(n4481), .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(n457), .E(n4518), .CP(n4591), .CDN(n4480), .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(n5), .E(n4518), .CP(n4591), .CDN(n4480), 
        .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(n4689), .E(n4518), .CP(n4591), .CDN(
        n4480), .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(n4686), .E(n4518), .CP(n4591), .CDN(
        n4480), .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(n669), .E(n4518), .CP(n4591), .CDN(n4480), .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(n723), .E(n4518), .CP(n4591), .CDN(n4480), .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(n775), .E(n4518), .CP(n4591), .CDN(n4480), .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(n827), .E(n4518), .CP(n4591), .CDN(n4480), .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n6), .E(n4518), .CP(n4591), .CDN(n4480), 
        .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(n4671), .E(n4518), .CP(n4592), .CDN(
        n4480), .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(n4668), .E(n4519), .CP(n4592), .CDN(
        n4480), .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n1039), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(n1093), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(n1145), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n1197), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n7), .E(n4519), .CP(n4592), .CDN(n4479), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n4653), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(n4650), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n1428), .E(n4519), .CP(n4592), .CDN(n4479), .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(n4645), .E(n4519), .CP(n4593), .CDN(n4479), .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n1532), .E(n4519), .CP(n4593), .CDN(n4479), .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n4576), .E(n4521), .CP(n4593), .CDN(
        n4479), .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(n10), .E(n4521), .CP(n4593), .CDN(n4478), 
        .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(n46), .E(n4520), .CP(n4593), .CDN(n4478), 
        .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(n140), .E(n4521), .CP(n4593), .CDN(n4478), .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(n191), .E(n4520), .CP(n4593), .CDN(n4478), .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(n1565), .E(n4521), .CP(n4593), .CDN(
        n4478), .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(n1672), .E(n4520), .CP(n4593), .CDN(
        n4478), .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(n1620), .E(n4521), .CP(n4593), .CDN(
        n4478), .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(n245), .E(n4520), .CP(n4594), .CDN(n4478), .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(n299), .E(n4521), .CP(n4594), .CDN(n4478), .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n354), .E(n4520), .CP(n4594), .CDN(n4478), .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(n406), .E(n4520), .CP(n4594), .CDN(n4478), .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(n457), .E(n4520), .CP(n4594), .CDN(n4477), .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(n5), .E(n4520), .CP(n4594), .CDN(n4477), 
        .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(n4689), .E(n4520), .CP(n4594), .CDN(
        n4477), .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(n4686), .E(n4520), .CP(n4594), .CDN(
        n4477), .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(n669), .E(n4520), .CP(n4594), .CDN(n4477), .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n724), .E(n4520), .CP(n4594), .CDN(n4477), .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n776), .E(n4520), .CP(n4595), .CDN(n4477), .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(n827), .E(n4520), .CP(n4595), .CDN(n4477), .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n6), .E(n4520), .CP(n4595), .CDN(n4477), 
        .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(n4671), .E(n4520), .CP(n4595), .CDN(
        n4477), .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(n4668), .E(n4521), .CP(n4595), .CDN(
        n4477), .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n1039), .E(n4521), .CP(n4595), .CDN(n4476), .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(n1094), .E(n4521), .CP(n4595), .CDN(n4476), .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n1146), .E(n4521), .CP(n4595), .CDN(n4476), .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n1197), .E(n4521), .CP(n4595), .CDN(n4476), .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n7), .E(n4521), .CP(n4595), .CDN(n4476), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n4653), .E(n4521), .CP(n4596), .CDN(n4476), .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(n4650), .E(n4521), .CP(n4596), .CDN(n4476), .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n1428), .E(n4521), .CP(n4596), .CDN(n4476), .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(n4645), .E(n4521), .CP(n4596), .CDN(n4476), .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n1532), .E(n4521), .CP(n4596), .CDN(n4476), .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n4576), .E(n4525), .CP(n4599), .CDN(
        n4473), .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(n10), .E(n4525), .CP(n4599), .CDN(n4472), 
        .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(n45), .E(n4524), .CP(n4600), .CDN(n4472), 
        .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(n139), .E(n4525), .CP(n4600), .CDN(n4472), .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(n191), .E(n4524), .CP(n4600), .CDN(n4472), .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(n1565), .E(n4525), .CP(n4600), .CDN(
        n4472), .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(n1671), .E(n4524), .CP(n4600), .CDN(
        n4472), .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(n1619), .E(n4525), .CP(n4600), .CDN(
        n4472), .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(n245), .E(n4524), .CP(n4600), .CDN(n4472), .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(n299), .E(n4525), .CP(n4600), .CDN(n4472), .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n353), .E(n4524), .CP(n4600), .CDN(n4472), .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(n405), .E(n4524), .CP(n4600), .CDN(n4472), .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(n457), .E(n4524), .CP(n4601), .CDN(n4471), .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(n1), .E(n4524), .CP(n4601), .CDN(n4471), 
        .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(n4689), .E(n4524), .CP(n4601), .CDN(
        n4471), .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(n4686), .E(n4524), .CP(n4601), .CDN(
        n4471), .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(n669), .E(n4524), .CP(n4601), .CDN(n4471), .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(n723), .E(n4524), .CP(n4601), .CDN(n4471), .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(n775), .E(n4524), .CP(n4601), .CDN(n4471), .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(n827), .E(n4524), .CP(n4601), .CDN(n4471), .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n2), .E(n4524), .CP(n4601), .CDN(n4471), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(n4671), .E(n4524), .CP(n4601), .CDN(
        n4471), .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(n4668), .E(n4525), .CP(n4602), .CDN(
        n4471), .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n1039), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(n1093), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(n1145), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n1197), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n3), .E(n4525), .CP(n4602), .CDN(n4470), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n4653), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(n4650), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n1428), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(n4645), .E(n4525), .CP(n4602), .CDN(n4470), .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n1532), .E(n4525), .CP(n4603), .CDN(n4470), .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(n4576), .E(n4531), .CP(n4609), .CDN(
        n4464), .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n4720), .E(n4531), .CP(n4609), .CDN(
        n4463), .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n46), .E(n4530), .CP(n4609), .CDN(n4463), 
        .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(n140), .E(n4531), .CP(n4628), .CDN(n4463), .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(n4713), .E(n4530), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(n4710), .E(n4531), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n1672), .E(n4530), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(n1620), .E(n4531), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(n4703), .E(n4530), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(n4700), .E(n4531), .CP(n4579), .CDN(
        n4463), .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(n354), .E(n4530), .CP(n4579), .CDN(n4463), .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(n406), .E(n4530), .CP(n4579), .CDN(n4463), .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(n4693), .E(n4530), .CP(n4627), .CDN(
        n4462), .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(n5), .E(n4530), .CP(n4626), .CDN(n4462), 
        .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(n4689), .E(n4530), .CP(n4579), .CDN(
        n4462), .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n4686), .E(n4530), .CP(n4623), .CDN(
        n4462), .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(n4682), .E(n4530), .CP(n4622), .CDN(
        n4462), .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(n724), .E(n4530), .CP(n4579), .CDN(n4462), .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(n776), .E(n4530), .CP(n4623), .CDN(n4462), .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n4675), .E(n4530), .CP(n4622), .CDN(
        n4462), .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(n6), .E(n4530), .CP(n4627), .CDN(n4462), 
        .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(n4671), .E(n4530), .CP(n4626), .CDN(
        n4462), .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(n4668), .E(n4531), .CP(n4625), .CDN(
        n4462), .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(n4664), .E(n4531), .CP(n4624), .CDN(n4461), .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(n1094), .E(n4531), .CP(n4624), .CDN(n4461), .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(n1146), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n4657), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n7), .E(n4531), .CP(ClockW), .CDN(n4461), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(n4653), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(n4650), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(n1428), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(n4645), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n1532), .E(n4531), .CP(ClockW), .CDN(
        n4461), .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(N85), .E(n4533), .CP(n4610), .CDN(n4461), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n4720), .E(n4533), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n46), .E(n4532), .CP(n4610), .CDN(n4460), 
        .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n140), .E(n4533), .CP(n4610), .CDN(n4460), .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n4713), .E(n4532), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(n4710), .E(n4533), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n1672), .E(n4532), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n1620), .E(n4533), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n4703), .E(n4532), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(n4700), .E(n4533), .CP(n4610), .CDN(
        n4460), .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n354), .E(n4532), .CP(n4611), .CDN(n4460), .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n406), .E(n4532), .CP(n4611), .CDN(n4460), .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n4693), .E(n4532), .CP(n4611), .CDN(
        n4459), .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n1), .E(n4532), .CP(n4611), .CDN(n4459), 
        .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(n4689), .E(n4532), .CP(n4611), .CDN(
        n4459), .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n4686), .E(n4532), .CP(n4611), .CDN(
        n4459), .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n4682), .E(n4532), .CP(n4611), .CDN(
        n4459), .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n724), .E(n4532), .CP(n4611), .CDN(n4459), .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n776), .E(n4532), .CP(n4611), .CDN(n4459), .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n4675), .E(n4532), .CP(n4611), .CDN(
        n4459), .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n2), .E(n4532), .CP(n4621), .CDN(n4459), 
        .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n4671), .E(n4532), .CP(n4620), .CDN(
        n4459), .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n4668), .E(n4533), .CP(n4619), .CDN(
        n4459), .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n4664), .E(n4533), .CP(n4629), .CDN(n4458), .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n1094), .E(n4533), .CP(n4627), .CDN(n4458), .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n1146), .E(n4533), .CP(n4626), .CDN(n4458), .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n4657), .E(n4533), .CP(n4625), .CDN(n4458), .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n3), .E(n4533), .CP(n4578), .CDN(n4458), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n4653), .E(n4533), .CP(n4628), .CDN(n4458), .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(n4650), .E(n4533), .CP(n4623), .CDN(n4458), .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n8), .E(n4533), .CP(n4631), .CDN(n4458), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n4645), .E(n4533), .CP(n4618), .CDN(n4458), .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n9), .E(n4533), .CP(n4631), .CDN(n4458), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(N85), .E(n4539), .CP(n4632), .CDN(n4452), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(n4720), .E(n4539), .CP(n4627), .CDN(
        n4451), .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(n46), .E(n4538), .CP(n4626), .CDN(n4451), 
        .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(n140), .E(n4539), .CP(n4615), .CDN(n4451), .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(n4713), .E(n4538), .CP(n4621), .CDN(
        n4451), .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(n4710), .E(n4539), .CP(n4620), .CDN(
        n4451), .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(n1672), .E(n4538), .CP(n4619), .CDN(
        n4451), .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(n1620), .E(n4539), .CP(n4625), .CDN(
        n4451), .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(n4703), .E(n4538), .CP(n4626), .CDN(
        n4451), .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(n4700), .E(n4539), .CP(ClockW), .CDN(
        n4451), .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n354), .E(n4538), .CP(n4629), .CDN(n4451), .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(n406), .E(n4538), .CP(n4623), .CDN(n4451), .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(n4693), .E(n4538), .CP(n4630), .CDN(
        n4450), .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(n1), .E(n4538), .CP(n4632), .CDN(n4450), 
        .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(n4689), .E(n4538), .CP(n4629), .CDN(
        n4450), .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(n4686), .E(n4538), .CP(n4625), .CDN(
        n4450), .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(n4682), .E(n4538), .CP(n4626), .CDN(
        n4450), .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(n724), .E(n4538), .CP(n4622), .CDN(n4450), .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(n776), .E(n4538), .CP(n4617), .CDN(n4450), .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n4675), .E(n4538), .CP(n4630), .CDN(
        n4450), .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n2), .E(n4538), .CP(n4613), .CDN(n4450), 
        .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(n4671), .E(n4538), .CP(n4632), .CDN(
        n4450), .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(n4668), .E(n4539), .CP(n4579), .CDN(
        n4450), .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n4664), .E(n4539), .CP(n4621), .CDN(n4449), .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(n1094), .E(n4539), .CP(n4620), .CDN(n4449), .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(n1146), .E(n4539), .CP(n4619), .CDN(n4449), .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n4657), .E(n4539), .CP(n4627), .CDN(n4449), .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n3), .E(n4539), .CP(n4626), .CDN(n4449), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n4653), .E(n4539), .CP(n4625), .CDN(n4449), .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(n4650), .E(n4539), .CP(n4578), .CDN(n4449), .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n1428), .E(n4539), .CP(n4621), .CDN(n4449), .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(n4645), .E(n4539), .CP(n4614), .CDN(n4449), .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n1532), .E(n4539), .CP(n4613), .CDN(n4449), .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n4576), .E(n4541), .CP(n4629), .CDN(
        n4449), .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n4720), .E(n4541), .CP(n4627), .CDN(
        n4448), .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n46), .E(n4540), .CP(n4627), .CDN(n4448), 
        .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(n140), .E(n4541), .CP(n4621), .CDN(n4448), .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(n4713), .E(n4540), .CP(n4628), .CDN(
        n4448), .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n4710), .E(n4541), .CP(n4620), .CDN(
        n4448), .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n1672), .E(n4540), .CP(n4578), .CDN(
        n4448), .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(n1620), .E(n4541), .CP(n4619), .CDN(
        n4448), .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(n4703), .E(n4540), .CP(n4622), .CDN(
        n4448), .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n4700), .E(n4541), .CP(n4623), .CDN(
        n4448), .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n354), .E(n4540), .CP(n4615), .CDN(n4448), .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(n406), .E(n4540), .CP(n4617), .CDN(n4448), .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(n4693), .E(n4540), .CP(n4616), .CDN(
        n4447), .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(n1), .E(n4540), .CP(n4621), .CDN(n4447), 
        .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n4689), .E(n4540), .CP(n4620), .CDN(
        n4447), .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n4686), .E(n4540), .CP(n4624), .CDN(
        n4447), .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(n4682), .E(n4540), .CP(n4596), .CDN(
        n4447), .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(n724), .E(n4540), .CP(n4597), .CDN(n4447), .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(n776), .E(n4540), .CP(n4601), .CDN(n4447), .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n4675), .E(n4540), .CP(n4615), .CDN(
        n4447), .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n2), .E(n4540), .CP(n4614), .CDN(n4447), 
        .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(n4671), .E(n4540), .CP(n4613), .CDN(
        n4447), .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(n4668), .E(n4541), .CP(n4632), .CDN(
        n4447), .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n4664), .E(n4541), .CP(n4626), .CDN(n4444), .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(n1094), .E(n4541), .CP(n4627), .CDN(n4446), .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(n1146), .E(n4541), .CP(n4622), .CDN(n4437), .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n4657), .E(n4541), .CP(n4624), .CDN(n4402), .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n3), .E(n4541), .CP(n4623), .CDN(n4446), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n4653), .E(n4541), .CP(n4615), .CDN(n4444), .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n4650), .E(n4541), .CP(n4618), .CDN(n4401), .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n1428), .E(n4541), .CP(n4599), .CDN(n4446), .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(n4645), .E(n4541), .CP(n4599), .CDN(n4478), .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n1532), .E(n4541), .CP(n4599), .CDN(n4400), .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n4576), .E(n4547), .CP(n4630), .CDN(
        n4443), .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n4720), .E(n4547), .CP(n4603), .CDN(
        n4475), .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n46), .E(n4546), .CP(n4616), .CDN(n4464), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n140), .E(n4547), .CP(n4616), .CDN(n4458), .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n4713), .E(n4546), .CP(n4616), .CDN(
        n4457), .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n4710), .E(n4547), .CP(n4616), .CDN(
        n4456), .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n1672), .E(n4546), .CP(n4616), .CDN(
        n4455), .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n1620), .E(n4547), .CP(n4616), .CDN(
        n4466), .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n4703), .E(n4546), .CP(n4616), .CDN(
        n4463), .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n4700), .E(n4547), .CP(n4602), .CDN(
        n4443), .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n354), .E(n4546), .CP(n4602), .CDN(n4465), .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n406), .E(n4546), .CP(n4602), .CDN(n4444), .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n4693), .E(n4546), .CP(n4584), .CDN(
        n4442), .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n1), .E(n4546), .CP(n4586), .CDN(n4442), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n4689), .E(n4546), .CP(n4587), .CDN(
        n4442), .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n4686), .E(n4546), .CP(n4588), .CDN(
        n4442), .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n4682), .E(n4546), .CP(n4589), .CDN(
        n4442), .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n724), .E(n4546), .CP(n4590), .CDN(n4442), .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n776), .E(n4546), .CP(n4591), .CDN(n4442), .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n4675), .E(n4546), .CP(n4606), .CDN(
        n4442), .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n2), .E(n4546), .CP(n4607), .CDN(n4442), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n4671), .E(n4546), .CP(n4608), .CDN(
        n4442), .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n4668), .E(n4547), .CP(n4609), .CDN(
        n4442), .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n4664), .E(n4547), .CP(n4623), .CDN(n4441), .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n1094), .E(n4547), .CP(n4579), .CDN(n4441), .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n1146), .E(n4547), .CP(n4624), .CDN(n4441), .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n4657), .E(n4547), .CP(n4610), .CDN(n4441), .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n3), .E(n4547), .CP(n4613), .CDN(n4441), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n4653), .E(n4547), .CP(n4625), .CDN(n4441), .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n4650), .E(n4547), .CP(n4613), .CDN(n4441), .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n1428), .E(n4547), .CP(n4623), .CDN(n4441), .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n4645), .E(n4547), .CP(n4619), .CDN(n4441), .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n1532), .E(n4547), .CP(n4617), .CDN(n4441), .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n4576), .E(n4549), .CP(n4627), .CDN(
        n4441), .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n4720), .E(n4549), .CP(n4626), .CDN(
        n4440), .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n46), .E(n4548), .CP(n4623), .CDN(n4440), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n140), .E(n4549), .CP(n4625), .CDN(n4440), .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n4713), .E(n4548), .CP(n4624), .CDN(
        n4440), .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n4710), .E(n4549), .CP(n4622), .CDN(
        n4440), .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n1672), .E(n4548), .CP(n4628), .CDN(
        n4440), .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n1620), .E(n4549), .CP(n4617), .CDN(
        n4440), .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n4703), .E(n4548), .CP(n4622), .CDN(
        n4440), .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n4700), .E(n4549), .CP(n4614), .CDN(
        n4440), .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n354), .E(n4548), .CP(n4621), .CDN(n4440), .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n406), .E(n4548), .CP(n4620), .CDN(n4440), .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n4693), .E(n4548), .CP(n4610), .CDN(
        n4439), .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n1), .E(n4548), .CP(n4624), .CDN(n4439), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n4689), .E(n4548), .CP(n4613), .CDN(
        n4439), .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n4686), .E(n4548), .CP(n4623), .CDN(
        n4439), .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n4682), .E(n4548), .CP(n4630), .CDN(
        n4439), .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n724), .E(n4548), .CP(n4605), .CDN(n4439), .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n776), .E(n4548), .CP(n4615), .CDN(n4439), .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n4675), .E(n4548), .CP(n4615), .CDN(
        n4439), .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n2), .E(n4548), .CP(n4615), .CDN(n4439), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n4671), .E(n4548), .CP(n4627), .CDN(
        n4439), .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n4668), .E(n4549), .CP(n4622), .CDN(
        n4439), .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n4664), .E(n4549), .CP(n4608), .CDN(n4475), .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n1094), .E(n4549), .CP(n4609), .CDN(n4475), .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n1146), .E(n4549), .CP(n4613), .CDN(n4477), .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n4657), .E(n4549), .CP(n4594), .CDN(n4478), .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n3), .E(n4549), .CP(n4580), .CDN(n4476), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n4653), .E(n4549), .CP(n4581), .CDN(n4475), .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n4650), .E(n4549), .CP(n4582), .CDN(n4477), .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n8), .E(n4549), .CP(n4583), .CDN(n4478), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n4645), .E(n4549), .CP(n4584), .CDN(n4476), .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n1532), .E(n4549), .CP(n4585), .CDN(n4444), .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(n4576), .E(n4555), .CP(n4593), .CDN(
        n4433), .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n10), .E(n4555), .CP(n4592), .CDN(n4432), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n46), .E(n4554), .CP(n4591), .CDN(n4432), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n140), .E(n4555), .CP(n4590), .CDN(n4432), .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n191), .E(n4554), .CP(n4589), .CDN(n4432), .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n1565), .E(n4555), .CP(n4588), .CDN(
        n4432), .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n1672), .E(n4554), .CP(n4587), .CDN(
        n4432), .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n1620), .E(n4555), .CP(n4608), .CDN(
        n4432), .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n245), .E(n4554), .CP(n4607), .CDN(n4432), .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n299), .E(n4555), .CP(n4604), .CDN(n4432), .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n354), .E(n4554), .CP(n4625), .CDN(n4432), .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n406), .E(n4554), .CP(n4600), .CDN(n4432), .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n457), .E(n4554), .CP(n4601), .CDN(n4431), .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n1), .E(n4554), .CP(n4622), .CDN(n4431), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n4688), .E(n4554), .CP(n4603), .CDN(
        n4431), .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n4685), .E(n4554), .CP(ClockW), .CDN(
        n4431), .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n669), .E(n4554), .CP(n4610), .CDN(n4431), .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n724), .E(n4554), .CP(n4605), .CDN(n4431), .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n776), .E(n4554), .CP(n4591), .CDN(n4431), .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n827), .E(n4554), .CP(n4625), .CDN(n4431), .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n2), .E(n4554), .CP(n4616), .CDN(n4431), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n4670), .E(n4554), .CP(n4595), .CDN(
        n4431), .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n4667), .E(n4555), .CP(n4607), .CDN(
        n4431), .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n1039), .E(n4555), .CP(n4578), .CDN(n4430), .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n1094), .E(n4555), .CP(n4632), .CDN(n4430), .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n1146), .E(n4555), .CP(n4615), .CDN(n4430), .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n1197), .E(n4555), .CP(n4593), .CDN(n4430), .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n3), .E(n4555), .CP(n4610), .CDN(n4430), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n4652), .E(n4555), .CP(n4597), .CDN(n4430), .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n4649), .E(n4555), .CP(n4609), .CDN(n4430), .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n1428), .E(n4555), .CP(n4604), .CDN(n4430), .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n4644), .E(n4555), .CP(n4607), .CDN(n4430), .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n1532), .E(n4555), .CP(n4606), .CDN(n4430), .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n4576), .E(n4557), .CP(n4608), .CDN(n4430), .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n4720), .E(n4557), .CP(n4609), .CDN(n4429), .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n46), .E(n4556), .CP(n4628), .CDN(n4429), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n140), .E(n4557), .CP(n4623), .CDN(n4429), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n4713), .E(n4556), .CP(n4594), .CDN(n4429), .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n4710), .E(n4557), .CP(n4594), .CDN(n4429), .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n1672), .E(n4556), .CP(n4613), .CDN(n4429), .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n1620), .E(n4557), .CP(n4593), .CDN(n4429), .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n4703), .E(n4556), .CP(n4582), .CDN(n4429), .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n4700), .E(n4557), .CP(n4581), .CDN(n4429), .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n354), .E(n4556), .CP(n4595), .CDN(n4429), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n406), .E(n4556), .CP(n4631), .CDN(n4429), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n4693), .E(n4556), .CP(n4581), .CDN(n4428), .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n5), .E(n4556), .CP(n4602), .CDN(n4428), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n4688), .E(n4556), .CP(n4588), .CDN(n4428), .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n4685), .E(n4556), .CP(n4625), .CDN(n4428), .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n4682), .E(n4556), .CP(n4580), .CDN(n4428), .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n724), .E(n4556), .CP(n4581), .CDN(n4428), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n776), .E(n4556), .CP(n4582), .CDN(n4428), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n4675), .E(n4556), .CP(n4583), .CDN(n4428), .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n6), .E(n4556), .CP(n4584), .CDN(n4428), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n4670), .E(n4556), .CP(n4585), .CDN(n4428), .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n4667), .E(n4557), .CP(n4586), .CDN(n4428), .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n4664), .E(n4557), .CP(n4587), .CDN(n4427), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n1094), .E(n4557), .CP(n4599), .CDN(n4427), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n1146), .E(n4557), .CP(n4589), .CDN(n4427), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n4657), .E(n4557), .CP(n4590), .CDN(n4427), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n7), .E(n4557), .CP(n4592), .CDN(n4427), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n4652), .E(n4557), .CP(n4593), .CDN(n4427), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n4649), .E(n4557), .CP(n4594), .CDN(n4427), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n8), .E(n4557), .CP(n4595), .CDN(n4427), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n4644), .E(n4557), .CP(n4596), .CDN(n4427), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n9), .E(n4557), .CP(n4597), .CDN(n4427), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n4576), .E(n4563), .CP(n4617), .CDN(n4421), .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n10), .E(n4563), .CP(ClockW), .CDN(n4420), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n46), .E(n4562), .CP(n4610), .CDN(n4420), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n140), .E(n4563), .CP(n4611), .CDN(n4420), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n191), .E(n4562), .CP(n4615), .CDN(n4420), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n1565), .E(n4563), .CP(n4580), .CDN(n4420), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n1672), .E(n4562), .CP(n4617), .CDN(n4420), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n1620), .E(n4563), .CP(n4622), .CDN(n4420), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n245), .E(n4562), .CP(n4616), .CDN(n4420), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n299), .E(n4563), .CP(n4594), .CDN(n4420), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n354), .E(n4562), .CP(n4620), .CDN(n4420), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n406), .E(n4562), .CP(n4614), .CDN(n4420), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n457), .E(n4562), .CP(n4614), .CDN(n4419), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n5), .E(n4562), .CP(n4619), .CDN(n4419), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n4688), .E(n4562), .CP(n4592), .CDN(n4419), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n4685), .E(n4562), .CP(n4606), .CDN(n4419), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n669), .E(n4562), .CP(n4597), .CDN(n4419), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n724), .E(n4562), .CP(n4598), .CDN(n4419), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n776), .E(n4562), .CP(n4599), .CDN(n4419), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n827), .E(n4562), .CP(n4600), .CDN(n4419), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n6), .E(n4562), .CP(n4601), .CDN(n4419), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n4670), .E(n4562), .CP(n4602), .CDN(n4419), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n4667), .E(n4563), .CP(n4603), .CDN(n4419), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n1039), .E(n4563), .CP(n4604), .CDN(n4418), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n1094), .E(n4563), .CP(n4605), .CDN(n4418), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n1146), .E(n4563), .CP(n4629), .CDN(n4418), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n1197), .E(n4563), .CP(n4607), .CDN(n4418), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n7), .E(n4563), .CP(n4608), .CDN(n4418), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n4652), .E(n4563), .CP(n4609), .CDN(n4418), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n4649), .E(n4563), .CP(n4628), .CDN(n4418), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n8), .E(n4563), .CP(n4579), .CDN(n4418), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n4644), .E(n4563), .CP(ClockW), .CDN(n4418), .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n9), .E(n4563), .CP(n4610), .CDN(n4418), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N85), .E(n4565), .CP(n4611), .CDN(n4418), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n4720), .E(n4565), .CP(n4628), .CDN(n4417), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n45), .E(n4564), .CP(n4621), .CDN(n4417), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n139), .E(n4565), .CP(n4616), .CDN(n4417), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n4713), .E(n4564), .CP(n4612), .CDN(n4417), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n4710), .E(n4565), .CP(n4615), .CDN(n4417), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n1671), .E(n4564), .CP(n4596), .CDN(n4417), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n1619), .E(n4565), .CP(n4613), .CDN(n4417), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n4703), .E(n4564), .CP(n4613), .CDN(n4417), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n4700), .E(n4565), .CP(n4628), .CDN(n4417), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n353), .E(n4564), .CP(n4616), .CDN(n4417), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n405), .E(n4564), .CP(n4593), .CDN(n4417), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n4693), .E(n4564), .CP(n4580), .CDN(n4416), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n5), .E(n4564), .CP(n4630), .CDN(n4416), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n4688), .E(n4564), .CP(n4630), .CDN(n4416), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n4685), .E(n4564), .CP(n4628), .CDN(n4416), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n4682), .E(n4564), .CP(n4591), .CDN(n4416), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n723), .E(n4564), .CP(n4622), .CDN(n4416), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n775), .E(n4564), .CP(n4595), .CDN(n4416), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n4675), .E(n4564), .CP(n4614), .CDN(n4416), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n6), .E(n4564), .CP(n4592), .CDN(n4416), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n4670), .E(n4564), .CP(n4581), .CDN(n4416), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n4667), .E(n4565), .CP(n4625), .CDN(n4416), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n4664), .E(n4565), .CP(n4583), .CDN(n4415), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n1093), .E(n4565), .CP(n4615), .CDN(n4415), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n1145), .E(n4565), .CP(n4625), .CDN(n4415), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n4657), .E(n4565), .CP(n4625), .CDN(n4415), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n7), .E(n4565), .CP(n4614), .CDN(n4415), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n4652), .E(n4565), .CP(n4623), .CDN(n4415), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n4649), .E(n4565), .CP(n4626), .CDN(n4415), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n8), .E(n4565), .CP(n4619), .CDN(n4415), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n4644), .E(n4565), .CP(n4624), .CDN(n4415), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n9), .E(n4565), .CP(n4580), .CDN(n4415), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N85), .E(n4571), .CP(n4596), .CDN(n4409), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n4720), .E(n4571), .CP(n4587), .CDN(n4408), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n45), .E(n4570), .CP(n4588), .CDN(n4408), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n139), .E(n4571), .CP(n4614), .CDN(n4408), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n4713), .E(n4570), .CP(n4623), .CDN(n4408), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n4710), .E(n4571), .CP(ClockW), .CDN(
        n4408), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n1671), .E(n4570), .CP(n4610), .CDN(n4408), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n1619), .E(n4571), .CP(n4611), .CDN(n4408), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n4703), .E(n4570), .CP(n4578), .CDN(n4408), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n4700), .E(n4571), .CP(n4625), .CDN(n4408), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n353), .E(n4570), .CP(n4624), .CDN(n4408), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n405), .E(n4570), .CP(n4622), .CDN(n4408), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n4693), .E(n4570), .CP(n4629), .CDN(n4407), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n5), .E(n4570), .CP(n4592), .CDN(n4407), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n4688), .E(n4570), .CP(n4588), .CDN(n4407), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n4685), .E(n4570), .CP(n4628), .CDN(n4407), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n4682), .E(n4570), .CP(n4630), .CDN(n4407), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n723), .E(n4570), .CP(n4630), .CDN(n4407), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n775), .E(n4570), .CP(n4578), .CDN(n4407), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n4675), .E(n4570), .CP(n4617), .CDN(n4407), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n6), .E(n4570), .CP(n4621), .CDN(n4407), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n4670), .E(n4570), .CP(n4612), .CDN(n4407), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n4667), .E(n4571), .CP(n4578), .CDN(n4407), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n4664), .E(n4571), .CP(n4626), .CDN(n4406), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n1093), .E(n4571), .CP(n4588), .CDN(n4406), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n1145), .E(n4571), .CP(n4586), .CDN(n4406), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n4657), .E(n4571), .CP(n4587), .CDN(n4406), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n7), .E(n4571), .CP(n4620), .CDN(n4406), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n4652), .E(n4571), .CP(n4583), .CDN(n4406), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n4649), .E(n4571), .CP(n4589), .CDN(n4406), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n8), .E(n4571), .CP(n4599), .CDN(n4406), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n4644), .E(n4571), .CP(n4608), .CDN(n4406), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n9), .E(n4571), .CP(n4587), .CDN(n4406), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(n4576), .E(n4572), .CP(n4609), .CDN(n4406), .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n4720), .E(n4572), .CP(n4600), .CDN(n4405), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n45), .E(n4573), .CP(n4592), .CDN(n4405), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n139), .E(n4572), .CP(n4619), .CDN(n4405), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n4713), .E(n4573), .CP(n4580), .CDN(n4405), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n4710), .E(n4572), .CP(n4581), .CDN(n4405), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n1671), .E(n4573), .CP(n4582), .CDN(n4405), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n1619), .E(n4572), .CP(n4583), .CDN(n4405), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n4703), .E(n4573), .CP(n4584), .CDN(n4405), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n4700), .E(n4572), .CP(n4585), .CDN(n4405), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n353), .E(n4573), .CP(n4598), .CDN(n4405), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n405), .E(n4572), .CP(n4597), .CDN(n4405), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n4693), .E(n4572), .CP(n4596), .CDN(n4404), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n5), .E(n4572), .CP(n4595), .CDN(n4404), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n4688), .E(n4572), .CP(n4594), .CDN(n4404), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n4685), .E(n4572), .CP(n4593), .CDN(n4404), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n4682), .E(n4572), .CP(n4592), .CDN(n4404), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n723), .E(n4572), .CP(n4591), .CDN(n4404), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n775), .E(n4572), .CP(n4590), .CDN(n4404), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n4675), .E(n4572), .CP(n4589), .CDN(n4404), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n6), .E(n4572), .CP(n4607), .CDN(n4404), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n4670), .E(n4572), .CP(n4606), .CDN(n4404), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n4667), .E(n4573), .CP(n4605), .CDN(n4404), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n4664), .E(n4573), .CP(n4604), .CDN(n4403), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n1093), .E(n4573), .CP(n4603), .CDN(n4403), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n1145), .E(n4573), .CP(n4602), .CDN(n4403), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n4657), .E(n4573), .CP(n4601), .CDN(n4403), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n7), .E(n4573), .CP(n4586), .CDN(n4403), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n4652), .E(n4573), .CP(n4630), .CDN(n4403), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n4649), .E(n4573), .CP(n4584), .CDN(n4403), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n8), .E(n4573), .CP(n4630), .CDN(n4403), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n4644), .E(n4573), .CP(n4591), .CDN(n4403), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n9), .E(n4573), .CP(n4628), .CDN(n4403), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n4576), .E(n4529), .CP(n4606), .CDN(
        n4467), .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(n10), .E(n4529), .CP(n4606), .CDN(n4466), 
        .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(n45), .E(n4528), .CP(n4606), .CDN(n4466), 
        .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(n139), .E(n4529), .CP(n4606), .CDN(n4466), .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(n191), .E(n4528), .CP(n4606), .CDN(n4466), .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(n1565), .E(n4529), .CP(n4606), .CDN(
        n4466), .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(n1671), .E(n4528), .CP(n4607), .CDN(
        n4466), .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(n1619), .E(n4529), .CP(n4607), .CDN(
        n4466), .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(n245), .E(n4528), .CP(n4607), .CDN(n4466), .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(n299), .E(n4529), .CP(n4607), .CDN(n4466), .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n353), .E(n4528), .CP(n4607), .CDN(n4466), .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(n405), .E(n4528), .CP(n4607), .CDN(n4466), .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(n457), .E(n4528), .CP(n4607), .CDN(n4465), .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(n5), .E(n4528), .CP(n4607), .CDN(n4465), 
        .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(n4689), .E(n4528), .CP(n4607), .CDN(
        n4465), .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(n4686), .E(n4528), .CP(n4607), .CDN(
        n4465), .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(n669), .E(n4528), .CP(n4608), .CDN(n4465), .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(n723), .E(n4528), .CP(n4608), .CDN(n4465), .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(n775), .E(n4528), .CP(n4608), .CDN(n4465), .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n827), .E(n4528), .CP(n4608), .CDN(n4465), .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n6), .E(n4528), .CP(n4608), .CDN(n4465), 
        .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(n4671), .E(n4528), .CP(n4608), .CDN(
        n4465), .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(n4668), .E(n4529), .CP(n4608), .CDN(
        n4465), .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n1039), .E(n4529), .CP(n4608), .CDN(n4464), .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(n1093), .E(n4529), .CP(n4608), .CDN(n4464), .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(n1145), .E(n4529), .CP(n4608), .CDN(n4464), .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n1197), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n7), .E(n4529), .CP(n4609), .CDN(n4464), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n4653), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(n4650), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n1428), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(n4645), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n1532), .E(n4529), .CP(n4609), .CDN(n4464), .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(N85), .E(n4535), .CP(n4618), .CDN(n4458), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(n4720), .E(n4535), .CP(n4618), .CDN(
        n4457), .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(n45), .E(n4534), .CP(n4618), .CDN(n4457), 
        .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(n139), .E(n4535), .CP(n4618), .CDN(n4457), .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(n4713), .E(n4534), .CP(n4618), .CDN(
        n4457), .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(n4710), .E(n4535), .CP(n4618), .CDN(
        n4457), .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(n1671), .E(n4534), .CP(n4618), .CDN(
        n4457), .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(n1619), .E(n4535), .CP(n4613), .CDN(
        n4457), .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(n4703), .E(n4534), .CP(n4629), .CDN(
        n4457), .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(n4700), .E(n4535), .CP(n4611), .CDN(
        n4457), .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n353), .E(n4534), .CP(n4623), .CDN(n4457), .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(n405), .E(n4534), .CP(n4627), .CDN(n4457), .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(n4693), .E(n4534), .CP(n4626), .CDN(
        n4456), .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(n1), .E(n4534), .CP(n4625), .CDN(n4456), 
        .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(n4689), .E(n4534), .CP(n4578), .CDN(
        n4456), .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(n4686), .E(n4534), .CP(n4621), .CDN(
        n4456), .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(n4682), .E(n4534), .CP(n4620), .CDN(
        n4456), .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(n723), .E(n4534), .CP(n4631), .CDN(n4456), .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(n775), .E(n4534), .CP(n4617), .CDN(n4456), .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(n4675), .E(n4534), .CP(n4579), .CDN(
        n4456), .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n2), .E(n4534), .CP(n4615), .CDN(n4456), 
        .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(n4671), .E(n4534), .CP(n4614), .CDN(
        n4456), .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(n4668), .E(n4535), .CP(n4613), .CDN(
        n4456), .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n4664), .E(n4535), .CP(n4632), .CDN(n4455), .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(n1093), .E(n4535), .CP(n4622), .CDN(n4455), .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(n1145), .E(n4535), .CP(n4621), .CDN(n4455), .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n4657), .E(n4535), .CP(n4620), .CDN(n4455), .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n3), .E(n4535), .CP(n4631), .CDN(n4455), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n4653), .E(n4535), .CP(n4631), .CDN(n4455), .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(n4650), .E(n4535), .CP(n4631), .CDN(n4455), .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n8), .E(n4535), .CP(n4631), .CDN(n4455), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(n4645), .E(n4535), .CP(n4631), .CDN(n4455), .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n1532), .E(n4535), .CP(n4631), .CDN(n4455), .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(N85), .E(n4537), .CP(n4631), .CDN(n4455), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(n4720), .E(n4537), .CP(n4631), .CDN(
        n4454), .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(n45), .E(n4536), .CP(n4631), .CDN(n4454), 
        .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(n139), .E(n4537), .CP(n4631), .CDN(n4454), .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(n4713), .E(n4536), .CP(n4627), .CDN(
        n4454), .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(n4710), .E(n4537), .CP(n4623), .CDN(
        n4454), .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(n1671), .E(n4536), .CP(n4632), .CDN(
        n4454), .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(n1619), .E(n4537), .CP(n4629), .CDN(
        n4454), .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(n4703), .E(n4536), .CP(n4630), .CDN(
        n4454), .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(n4700), .E(n4537), .CP(n4628), .CDN(
        n4454), .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n353), .E(n4536), .CP(n4620), .CDN(n4454), .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(n405), .E(n4536), .CP(n4629), .CDN(n4454), .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(n4693), .E(n4536), .CP(n4631), .CDN(
        n4453), .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(n1), .E(n4536), .CP(n4619), .CDN(n4453), 
        .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(n4689), .E(n4536), .CP(n4619), .CDN(
        n4453), .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(n4686), .E(n4536), .CP(n4626), .CDN(
        n4453), .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(n4682), .E(n4536), .CP(n4629), .CDN(
        n4453), .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(n723), .E(n4536), .CP(n4624), .CDN(n4453), .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(n775), .E(n4536), .CP(n4632), .CDN(n4453), .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(n4675), .E(n4536), .CP(n4579), .CDN(
        n4453), .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n2), .E(n4536), .CP(n4622), .CDN(n4453), 
        .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(n4671), .E(n4536), .CP(n4612), .CDN(
        n4453), .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(n4668), .E(n4537), .CP(n4613), .CDN(
        n4453), .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n4664), .E(n4537), .CP(n4630), .CDN(n4452), .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(n1093), .E(n4537), .CP(n4629), .CDN(n4452), .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(n1145), .E(n4537), .CP(n4618), .CDN(n4452), .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n4657), .E(n4537), .CP(n4619), .CDN(n4452), .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n3), .E(n4537), .CP(n4620), .CDN(n4452), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n4653), .E(n4537), .CP(n4621), .CDN(n4452), .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(n4650), .E(n4537), .CP(n4627), .CDN(n4452), .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n1428), .E(n4537), .CP(n4598), .CDN(n4452), .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(n4645), .E(n4537), .CP(n4618), .CDN(n4452), .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n9), .E(n4537), .CP(n4618), .CDN(n4452), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(N85), .E(n4543), .CP(n4599), .CDN(n4446), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(n4720), .E(n4543), .CP(n4599), .CDN(
        n4400), .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(n45), .E(n4542), .CP(n4600), .CDN(n4401), 
        .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(n139), .E(n4543), .CP(n4613), .CDN(n4403), .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(n4713), .E(n4542), .CP(n4630), .CDN(
        n4402), .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(n4710), .E(n4543), .CP(n4617), .CDN(
        n4477), .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(n1671), .E(n4542), .CP(n4621), .CDN(
        n4400), .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(n1619), .E(n4543), .CP(n4612), .CDN(
        n4475), .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(n4703), .E(n4542), .CP(n4578), .CDN(
        n4476), .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(n4700), .E(n4543), .CP(n4629), .CDN(
        n4478), .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n353), .E(n4542), .CP(n4628), .CDN(n4402), .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(n405), .E(n4542), .CP(n4627), .CDN(n4403), .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(n4693), .E(n4542), .CP(n4626), .CDN(
        n4477), .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(n1), .E(n4542), .CP(n4616), .CDN(n4476), 
        .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(n4689), .E(n4542), .CP(n4632), .CDN(
        n4453), .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(n4686), .E(n4542), .CP(n4617), .CDN(
        n4452), .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(n4682), .E(n4542), .CP(n4605), .CDN(
        n4451), .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(n723), .E(n4542), .CP(n4605), .CDN(n4489), .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(n775), .E(n4542), .CP(n4605), .CDN(n4488), .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(n4675), .E(n4542), .CP(n4632), .CDN(
        n4436), .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n2), .E(n4542), .CP(n4615), .CDN(n4454), 
        .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(n4671), .E(n4542), .CP(n4614), .CDN(
        n4437), .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(n4668), .E(n4543), .CP(n4621), .CDN(
        n4444), .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n4664), .E(n4543), .CP(n4620), .CDN(n4446), .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(n1093), .E(n4543), .CP(n4628), .CDN(n4446), .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(n1145), .E(n4543), .CP(n4579), .CDN(n4446), .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n4657), .E(n4543), .CP(n4615), .CDN(n4446), .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n3), .E(n4543), .CP(n4614), .CDN(n4446), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n4653), .E(n4543), .CP(n4613), .CDN(n4446), .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(n4650), .E(n4543), .CP(n4627), .CDN(n4446), .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n8), .E(n4543), .CP(n4632), .CDN(n4446), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(n4645), .E(n4543), .CP(n4611), .CDN(n4446), .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n9), .E(n4543), .CP(n4628), .CDN(n4446), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N85), .E(n4545), .CP(n4600), .CDN(n4446), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n4720), .E(n4545), .CP(n4601), .CDN(
        n4445), .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n45), .E(n4544), .CP(n4578), .CDN(n4445), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n139), .E(n4545), .CP(n4619), .CDN(n4445), .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n4713), .E(n4544), .CP(n4626), .CDN(
        n4445), .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n4710), .E(n4545), .CP(n4620), .CDN(
        n4445), .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n1671), .E(n4544), .CP(n4621), .CDN(
        n4445), .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n1619), .E(n4545), .CP(n4628), .CDN(
        n4445), .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n4703), .E(n4544), .CP(n4629), .CDN(
        n4445), .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n4700), .E(n4545), .CP(n4578), .CDN(
        n4445), .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n353), .E(n4544), .CP(n4578), .CDN(n4445), .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n405), .E(n4544), .CP(n4615), .CDN(n4445), .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n4693), .E(n4544), .CP(n4598), .CDN(
        n4444), .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n1), .E(n4544), .CP(n4632), .CDN(n4444), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n4689), .E(n4544), .CP(n4620), .CDN(
        n4444), .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n4686), .E(n4544), .CP(n4621), .CDN(
        n4444), .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n4682), .E(n4544), .CP(n4619), .CDN(
        n4444), .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n723), .E(n4544), .CP(n4630), .CDN(n4444), .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n775), .E(n4544), .CP(n4615), .CDN(n4444), .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n4675), .E(n4544), .CP(n4617), .CDN(
        n4444), .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n2), .E(n4544), .CP(n4624), .CDN(n4444), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n4671), .E(n4544), .CP(n4632), .CDN(
        n4444), .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n4668), .E(n4545), .CP(n4612), .CDN(
        n4444), .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n4664), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n1093), .E(n4545), .CP(n4617), .CDN(n4443), .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n1145), .E(n4545), .CP(n4615), .CDN(n4443), .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n4657), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n3), .E(n4545), .CP(n4612), .CDN(n4443), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n4653), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n4650), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n1428), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n4645), .E(n4545), .CP(n4612), .CDN(n4443), .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n1532), .E(n4545), .CP(n4616), .CDN(n4443), .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N85), .E(n4551), .CP(n4586), .CDN(n4437), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n4720), .E(n4551), .CP(n4587), .CDN(
        n4438), .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n46), .E(n4550), .CP(n4588), .CDN(n4438), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n140), .E(n4551), .CP(n4582), .CDN(n4438), .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n4713), .E(n4550), .CP(n4595), .CDN(
        n4438), .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n4710), .E(n4551), .CP(n4596), .CDN(
        n4438), .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n1672), .E(n4550), .CP(n4597), .CDN(
        n4438), .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n1620), .E(n4551), .CP(n4600), .CDN(
        n4438), .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n4703), .E(n4550), .CP(n4601), .CDN(
        n4438), .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n4700), .E(n4551), .CP(n4603), .CDN(
        n4438), .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n354), .E(n4550), .CP(n4624), .CDN(n4438), .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n406), .E(n4550), .CP(n4611), .CDN(n4438), .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n4693), .E(n4550), .CP(n4631), .CDN(
        n4437), .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n1), .E(n4550), .CP(n4603), .CDN(n4437), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n4688), .E(n4550), .CP(n4583), .CDN(
        n4437), .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n4685), .E(n4550), .CP(n4584), .CDN(
        n4437), .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n4682), .E(n4550), .CP(n4585), .CDN(
        n4437), .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n724), .E(n4550), .CP(n4586), .CDN(n4437), .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n776), .E(n4550), .CP(n4587), .CDN(n4437), .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n4675), .E(n4550), .CP(n4588), .CDN(
        n4437), .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n2), .E(n4550), .CP(n4589), .CDN(n4437), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n4670), .E(n4550), .CP(n4590), .CDN(
        n4437), .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n4667), .E(n4551), .CP(n4591), .CDN(
        n4437), .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n4664), .E(n4551), .CP(n4580), .CDN(n4436), .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n1094), .E(n4551), .CP(n4579), .CDN(n4436), .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n1146), .E(n4551), .CP(n4622), .CDN(n4436), .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n4657), .E(n4551), .CP(n4624), .CDN(n4436), .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n3), .E(n4551), .CP(n4610), .CDN(n4436), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n4652), .E(n4551), .CP(n4606), .CDN(n4436), .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n4649), .E(n4551), .CP(n4607), .CDN(n4436), .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n8), .E(n4551), .CP(n4608), .CDN(n4436), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n4644), .E(n4551), .CP(n4609), .CDN(n4436), .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n9), .E(n4551), .CP(n4604), .CDN(n4436), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N85), .E(n4553), .CP(n4594), .CDN(n4436), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n4720), .E(n4553), .CP(n4582), .CDN(
        n4435), .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n46), .E(n4552), .CP(n4583), .CDN(n4435), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n140), .E(n4553), .CP(n4585), .CDN(n4435), .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n4713), .E(n4552), .CP(n4584), .CDN(
        n4435), .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n4710), .E(n4553), .CP(n4587), .CDN(
        n4435), .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n1672), .E(n4552), .CP(n4586), .CDN(
        n4435), .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n1620), .E(n4553), .CP(n4588), .CDN(
        n4435), .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n4703), .E(n4552), .CP(n4589), .CDN(
        n4435), .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n4700), .E(n4553), .CP(n4590), .CDN(
        n4435), .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n354), .E(n4552), .CP(n4585), .CDN(n4435), .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n406), .E(n4552), .CP(n4603), .CDN(n4435), .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n4693), .E(n4552), .CP(n4611), .CDN(
        n4434), .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n1), .E(n4552), .CP(n4629), .CDN(n4434), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n4688), .E(n4552), .CP(n4597), .CDN(
        n4434), .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n4685), .E(n4552), .CP(n4596), .CDN(
        n4434), .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n4682), .E(n4552), .CP(n4600), .CDN(
        n4434), .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n724), .E(n4552), .CP(n4601), .CDN(n4434), .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n776), .E(n4552), .CP(n4619), .CDN(n4434), .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n4675), .E(n4552), .CP(n4617), .CDN(
        n4434), .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n2), .E(n4552), .CP(n4582), .CDN(n4434), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n4670), .E(n4552), .CP(n4596), .CDN(
        n4434), .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n4667), .E(n4553), .CP(n4595), .CDN(
        n4434), .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n4664), .E(n4553), .CP(n4627), .CDN(n4433), .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n1094), .E(n4553), .CP(n4578), .CDN(n4433), .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n1146), .E(n4553), .CP(n4626), .CDN(n4433), .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n4657), .E(n4553), .CP(n4615), .CDN(n4433), .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n3), .E(n4553), .CP(ClockW), .CDN(n4433), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n4652), .E(n4553), .CP(n4624), .CDN(n4433), .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n4649), .E(n4553), .CP(n4612), .CDN(n4433), .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n1428), .E(n4553), .CP(n4586), .CDN(n4433), .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n4644), .E(n4553), .CP(n4585), .CDN(n4433), .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n1532), .E(n4553), .CP(n4584), .CDN(n4433), .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N85), .E(n4559), .CP(n4598), .CDN(n4427), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n4720), .E(n4559), .CP(n4609), .CDN(n4426), .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n46), .E(n4558), .CP(n4600), .CDN(n4426), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n140), .E(n4559), .CP(n4601), .CDN(n4426), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n4713), .E(n4558), .CP(n4602), .CDN(n4426), .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n4710), .E(n4559), .CP(n4603), .CDN(n4426), .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n1672), .E(n4558), .CP(n4604), .CDN(n4426), .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n1620), .E(n4559), .CP(n4605), .CDN(n4426), .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n4703), .E(n4558), .CP(n4606), .CDN(n4426), .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n4700), .E(n4559), .CP(n4607), .CDN(n4426), .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n354), .E(n4558), .CP(n4608), .CDN(n4426), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n406), .E(n4558), .CP(n4614), .CDN(n4426), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n4693), .E(n4558), .CP(n4619), .CDN(n4425), .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n5), .E(n4558), .CP(n4624), .CDN(n4425), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n4688), .E(n4558), .CP(n4578), .CDN(n4425), .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n4685), .E(n4558), .CP(n4621), .CDN(n4425), .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n4682), .E(n4558), .CP(n4623), .CDN(n4425), .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n724), .E(n4558), .CP(n4626), .CDN(n4425), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n776), .E(n4558), .CP(ClockW), .CDN(n4425), .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n4675), .E(n4558), .CP(n4610), .CDN(n4425), .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n6), .E(n4558), .CP(n4611), .CDN(n4425), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n4670), .E(n4558), .CP(n4623), .CDN(n4425), .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n4667), .E(n4559), .CP(n4591), .CDN(n4425), .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n4664), .E(n4559), .CP(n4598), .CDN(n4424), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n1094), .E(n4559), .CP(n4620), .CDN(n4424), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n1146), .E(n4559), .CP(n4616), .CDN(n4424), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n4657), .E(n4559), .CP(n4617), .CDN(n4424), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n7), .E(n4559), .CP(n4632), .CDN(n4424), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n4652), .E(n4559), .CP(n4630), .CDN(n4424), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n4649), .E(n4559), .CP(n4619), .CDN(n4424), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n8), .E(n4559), .CP(n4632), .CDN(n4424), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n4644), .E(n4559), .CP(n4590), .CDN(n4424), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n9), .E(n4559), .CP(n4581), .CDN(n4424), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N85), .E(n4561), .CP(n4582), .CDN(n4424), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n4720), .E(n4561), .CP(n4583), .CDN(n4423), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n46), .E(n4560), .CP(n4584), .CDN(n4423), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n140), .E(n4561), .CP(n4585), .CDN(n4423), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n4713), .E(n4560), .CP(n4586), .CDN(n4423), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n4710), .E(n4561), .CP(n4587), .CDN(n4423), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n1672), .E(n4560), .CP(n4588), .CDN(n4423), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n1620), .E(n4561), .CP(n4589), .CDN(n4423), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n4703), .E(n4560), .CP(n4601), .CDN(n4423), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n4700), .E(n4561), .CP(n4592), .CDN(n4423), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n354), .E(n4560), .CP(n4593), .CDN(n4423), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n406), .E(n4560), .CP(n4594), .CDN(n4423), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n4693), .E(n4560), .CP(n4595), .CDN(n4422), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n5), .E(n4560), .CP(n4596), .CDN(n4422), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n4688), .E(n4560), .CP(n4597), .CDN(n4422), .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n4685), .E(n4560), .CP(n4598), .CDN(n4422), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n4682), .E(n4560), .CP(n4599), .CDN(n4422), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n724), .E(n4560), .CP(n4600), .CDN(n4422), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n776), .E(n4560), .CP(n4627), .CDN(n4422), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n4675), .E(n4560), .CP(n4602), .CDN(n4422), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n6), .E(n4560), .CP(n4603), .CDN(n4422), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n4670), .E(n4560), .CP(n4604), .CDN(n4422), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n4667), .E(n4561), .CP(n4605), .CDN(n4422), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n4664), .E(n4561), .CP(n4606), .CDN(n4421), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n1094), .E(n4561), .CP(n4607), .CDN(n4421), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n1146), .E(n4561), .CP(n4608), .CDN(n4421), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n4657), .E(n4561), .CP(n4609), .CDN(n4421), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n7), .E(n4561), .CP(n4579), .CDN(n4421), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n4652), .E(n4561), .CP(n4578), .CDN(n4421), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n4649), .E(n4561), .CP(n4620), .CDN(n4421), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n8), .E(n4561), .CP(n4616), .CDN(n4421), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n4644), .E(n4561), .CP(n4617), .CDN(n4421), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n9), .E(n4561), .CP(n4597), .CDN(n4421), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N85), .E(n4567), .CP(n4618), .CDN(n4415), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n4720), .E(n4567), .CP(n4618), .CDN(n4414), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n46), .E(n4566), .CP(n4629), .CDN(n4414), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n140), .E(n4567), .CP(n4598), .CDN(n4414), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n4713), .E(n4566), .CP(n4618), .CDN(n4414), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n4710), .E(n4567), .CP(n4626), .CDN(n4414), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n1672), .E(n4566), .CP(n4578), .CDN(n4414), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n1620), .E(n4567), .CP(n4578), .CDN(n4414), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n4703), .E(n4566), .CP(n4618), .CDN(n4414), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n4700), .E(n4567), .CP(n4598), .CDN(n4414), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n354), .E(n4566), .CP(n4589), .CDN(n4414), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n406), .E(n4566), .CP(n4590), .CDN(n4414), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n4693), .E(n4566), .CP(n4591), .CDN(n4413), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n5), .E(n4566), .CP(n4592), .CDN(n4413), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n4688), .E(n4566), .CP(n4593), .CDN(n4413), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n4685), .E(n4566), .CP(n4594), .CDN(n4413), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n4682), .E(n4566), .CP(n4595), .CDN(n4413), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n724), .E(n4566), .CP(n4596), .CDN(n4413), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n776), .E(n4566), .CP(n4597), .CDN(n4413), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n4675), .E(n4566), .CP(n4608), .CDN(n4413), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n6), .E(n4566), .CP(n4599), .CDN(n4413), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n4670), .E(n4566), .CP(n4600), .CDN(n4413), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n4667), .E(n4567), .CP(n4601), .CDN(n4413), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n4664), .E(n4567), .CP(n4602), .CDN(n4412), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n1094), .E(n4567), .CP(n4603), .CDN(n4412), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n1146), .E(n4567), .CP(n4604), .CDN(n4412), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n4657), .E(n4567), .CP(n4605), .CDN(n4412), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n7), .E(n4567), .CP(n4606), .CDN(n4412), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n4652), .E(n4567), .CP(n4607), .CDN(n4412), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n4649), .E(n4567), .CP(n4629), .CDN(n4412), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n8), .E(n4567), .CP(n4609), .CDN(n4412), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n4644), .E(n4567), .CP(n4625), .CDN(n4412), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n9), .E(n4567), .CP(n4622), .CDN(n4412), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N85), .E(n4569), .CP(ClockW), .CDN(n4412), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n10), .E(n4569), .CP(n4610), .CDN(n4411), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n46), .E(n4568), .CP(n4611), .CDN(n4411), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n140), .E(n4569), .CP(n4613), .CDN(n4411), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n191), .E(n4568), .CP(n4616), .CDN(n4411), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n1565), .E(n4569), .CP(n4578), .CDN(n4411), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n1672), .E(n4568), .CP(n4602), .CDN(n4411), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n1620), .E(n4569), .CP(ClockW), .CDN(
        n4411), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n245), .E(n4568), .CP(n4617), .CDN(n4411), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n299), .E(n4569), .CP(n4590), .CDN(n4411), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n354), .E(n4568), .CP(n4617), .CDN(n4411), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n406), .E(n4568), .CP(n4593), .CDN(n4411), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n457), .E(n4568), .CP(n4612), .CDN(n4410), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n5), .E(n4568), .CP(n4604), .CDN(n4410), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n4688), .E(n4568), .CP(n4580), .CDN(n4410), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n4685), .E(n4568), .CP(n4625), .CDN(n4410), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n669), .E(n4568), .CP(n4586), .CDN(n4410), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n724), .E(n4568), .CP(n4613), .CDN(n4410), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n776), .E(n4568), .CP(n4606), .CDN(n4410), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n827), .E(n4568), .CP(n4606), .CDN(n4410), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n6), .E(n4568), .CP(n4580), .CDN(n4410), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n4670), .E(n4568), .CP(n4581), .CDN(n4410), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n4667), .E(n4569), .CP(n4582), .CDN(n4410), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n1039), .E(n4569), .CP(n4583), .CDN(n4409), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n1094), .E(n4569), .CP(n4584), .CDN(n4409), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n1146), .E(n4569), .CP(n4585), .CDN(n4409), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n1197), .E(n4569), .CP(n4589), .CDN(n4409), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n7), .E(n4569), .CP(n4591), .CDN(n4409), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n4652), .E(n4569), .CP(n4590), .CDN(n4409), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n4649), .E(n4569), .CP(n4593), .CDN(n4409), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n8), .E(n4569), .CP(n4592), .CDN(n4409), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n4644), .E(n4569), .CP(n4594), .CDN(n4409), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n9), .E(n4569), .CP(n4595), .CDN(n4409), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(n4576), .E(n4574), .CP(n4630), .CDN(n4403), .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n4720), .E(n4574), .CP(n4583), .CDN(n4402), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n46), .E(n4574), .CP(n4611), .CDN(n4402), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n140), .E(n4574), .CP(n4581), .CDN(n4402), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n4713), .E(n4575), .CP(n4618), .CDN(n4402), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n4710), .E(n4574), .CP(n4623), .CDN(n4402), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n1672), .E(n4575), .CP(n4624), .CDN(n4402), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n1620), .E(n4574), .CP(n4585), .CDN(n4402), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n4703), .E(n4575), .CP(n4619), .CDN(n4402), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n4700), .E(n4574), .CP(n4631), .CDN(n4402), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n354), .E(n4575), .CP(n4598), .CDN(n4402), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n406), .E(n4574), .CP(n4625), .CDN(n4402), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n4693), .E(n4574), .CP(n4612), .CDN(n4401), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n5), .E(n4574), .CP(n4621), .CDN(n4401), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n4688), .E(n4574), .CP(n4580), .CDN(n4401), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n4685), .E(n4574), .CP(n4581), .CDN(n4401), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n4682), .E(n4574), .CP(n4582), .CDN(n4401), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n724), .E(n4574), .CP(n4613), .CDN(n4401), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n776), .E(n4574), .CP(n4620), .CDN(n4401), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n4675), .E(n4574), .CP(n4630), .CDN(n4401), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n6), .E(n4574), .CP(n4612), .CDN(n4401), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n4670), .E(n4574), .CP(n4616), .CDN(n4401), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n4667), .E(n4575), .CP(n4604), .CDN(n4401), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n4664), .E(n4575), .CP(n4612), .CDN(n4400), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n1094), .E(n4575), .CP(n4628), .CDN(n4400), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n1146), .E(n4575), .CP(n4617), .CDN(n4400), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n4657), .E(n4575), .CP(n4622), .CDN(n4400), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n7), .E(n4575), .CP(n4622), .CDN(n4400), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n4652), .E(n4575), .CP(n4619), .CDN(n4400), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n4649), .E(n4575), .CP(n4632), .CDN(n4400), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n8), .E(n4575), .CP(n4618), .CDN(n4400), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n4644), .E(n4575), .CP(n4612), .CDN(n4400), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n9), .E(n4575), .CP(n4627), .CDN(n4400), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(N85), .E(n4513), .CP(n4580), .CDN(n4490), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(n10), .E(n4512), .CP(n4580), .CDN(n4446), 
        .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(n45), .E(n4513), .CP(n4580), .CDN(n4403), 
        .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(n139), .E(n4512), .CP(n4580), .CDN(n4446), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(n191), .E(n4513), .CP(n4580), .CDN(n4477), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(n1565), .E(n4512), .CP(n4580), .CDN(
        n4446), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(n1619), .E(n4513), .CP(n4580), .CDN(
        n4478), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(n245), .E(n4512), .CP(n4580), .CDN(n4446), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(n299), .E(n4513), .CP(n4580), .CDN(n4476), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(n353), .E(n4512), .CP(n4581), .CDN(n4446), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(n405), .E(n4512), .CP(n4581), .CDN(n4475), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(n457), .E(n4512), .CP(n4581), .CDN(n4489), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(n1), .E(n4512), .CP(n4581), .CDN(n4489), 
        .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(n4688), .E(n4512), .CP(n4581), .CDN(
        n4489), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(n4685), .E(n4512), .CP(n4581), .CDN(
        n4489), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(n669), .E(n4512), .CP(n4581), .CDN(n4489), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(n723), .E(n4512), .CP(n4581), .CDN(n4489), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(n775), .E(n4512), .CP(n4581), .CDN(n4489), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(n827), .E(n4512), .CP(n4581), .CDN(n4489), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(n2), .E(n4512), .CP(n4582), .CDN(n4489), 
        .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(n4670), .E(n4512), .CP(n4582), .CDN(
        n4489), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(n4667), .E(n4513), .CP(n4582), .CDN(
        n4489), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(n1039), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(n1093), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(n1145), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(n1197), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(n3), .E(n4513), .CP(n4582), .CDN(n4488), 
        .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(n4652), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(n4649), .E(n4513), .CP(n4582), .CDN(n4488), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(n1428), .E(n4513), .CP(n4583), .CDN(n4488), .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(n4644), .E(n4513), .CP(n4583), .CDN(n4488), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(n1532), .E(n4513), .CP(n4583), .CDN(n4488), .Q(\Storage[31][0] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(n1671), .E(n4515), .CP(n4583), .CDN(
        n4487), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(n1619), .E(n4514), .CP(n4584), .CDN(
        n4487), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(n1671), .E(n4517), .CP(n4587), .CDN(
        n4484), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(n1619), .E(n4516), .CP(n4587), .CDN(
        n4484), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(n1565), .E(n4518), .CP(n4590), .CDN(
        n4481), .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(n1671), .E(n4519), .CP(n4590), .CDN(
        n4481), .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(n1619), .E(n4518), .CP(n4590), .CDN(
        n4481), .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(n1671), .E(n4512), .CP(n4580), .CDN(
        n4437), .Q(\Storage[31][26] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(n1723), .E(n4637), .CP(n4633), .CDN(n4478), 
        .Q(DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(n1789), .E(n4637), .CP(ClockR), .CDN(n4454), 
        .Q(DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(n1855), .E(n4637), .CP(ClockR), .CDN(n4494), 
        .Q(DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(n1921), .E(n4637), .CP(ClockR), .CDN(n4452), 
        .Q(DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(n1987), .E(n4637), .CP(ClockR), .CDN(n4453), 
        .Q(DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(n2053), .E(n4637), .CP(ClockR), .CDN(n4451), 
        .Q(DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(n2119), .E(n4637), .CP(n4633), .CDN(n4436), 
        .Q(DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(n2185), .E(n4637), .CP(ClockR), .CDN(n4488), 
        .Q(DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(n2251), .E(n4637), .CP(ClockR), .CDN(n4489), 
        .Q(DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(n2317), .E(n4637), .CP(n4633), .CDN(n4488), 
        .Q(DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(n2383), .E(n4637), .CP(n4633), .CDN(n4401), 
        .Q(DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(n2449), .E(n4638), .CP(ClockR), .CDN(n4437), 
        .Q(DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(n2515), .E(n4638), .CP(n4633), .CDN(n4444), 
        .Q(DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(n2581), .E(n4638), .CP(ClockR), .CDN(n4437), 
        .Q(DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(n2647), .E(n4638), .CP(n4633), .CDN(n4489), 
        .Q(DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(n2713), .E(n4638), .CP(ClockR), .CDN(n4488), 
        .Q(DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(n2779), .E(n4638), .CP(n4633), .CDN(n4436), 
        .Q(DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(n2845), .E(n4638), .CP(ClockR), .CDN(n4451), 
        .Q(DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(n2911), .E(n4638), .CP(n4633), .CDN(n4453), 
        .Q(DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(n2977), .E(n4638), .CP(ClockR), .CDN(n4454), 
        .Q(DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(n3043), .E(n4638), .CP(n4633), .CDN(n4452), 
        .Q(DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(n3109), .E(n4638), .CP(n4633), .CDN(n4476), 
        .Q(DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(n3174), .E(n4639), .CP(n4633), .CDN(n4477), 
        .Q(DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(n3236), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(n3301), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(n3360), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(n3423), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(n3486), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(n3550), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(n3614), .E(n4639), .CP(n4633), .CDN(n4490), 
        .Q(DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(n3677), .E(n4639), .CP(ClockR), .CDN(n4490), 
        .Q(DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(n3735), .E(n4639), .CP(ClockR), .CDN(n4490), 
        .Q(DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(n3802), .E(n4639), .CP(ClockR), .CDN(n4490), .Q(
        ParityErr) );
  BUFTD16 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  BUFTD16 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD16 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD16 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD16 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD16 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD16 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD16 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD16 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD16 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD16 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD16 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD16 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD16 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD16 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD16 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD16 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD16 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD16 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD16 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD16 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD16 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD16 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD16 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD16 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD16 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD16 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD16 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD16 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD16 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD16 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD16 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  EDFCNQD1 Dreadyr_reg ( .D(n3889), .E(n3887), .CP(ClockR), .CDN(n108), .Q(
        Dreadyr) );
  TIEH U3 ( .Z(n3889) );
  XOR3D0 U4 ( .A1(n3799), .A2(n3864), .A3(n86), .Z(N83) );
  CKBD0 U5 ( .CLK(n1409), .C(n4) );
  INVD0 U6 ( .I(n4), .ZN(n4647) );
  CKBD0 U7 ( .CLK(n1514), .C(n1513) );
  CKBD0 U8 ( .CLK(n4642), .C(n9) );
  INVD0 U9 ( .I(n1513), .ZN(n4642) );
  CKBXD0 U10 ( .I(n1460), .Z(n1459) );
  CKNXD0 U11 ( .I(n1459), .ZN(n4645) );
  CKBXD0 U12 ( .I(n1356), .Z(n1355) );
  CKNXD0 U13 ( .I(n1355), .ZN(n4650) );
  CKBXD0 U14 ( .I(n1302), .Z(n1301) );
  CKNXD0 U15 ( .I(n1301), .ZN(n4653) );
  CKBXD0 U16 ( .I(n986), .Z(n985) );
  CKNXD0 U17 ( .I(n985), .ZN(n4668) );
  CKBXD0 U23 ( .I(n932), .Z(n931) );
  CKNXD0 U24 ( .I(n931), .ZN(n4671) );
  CKBXD0 U25 ( .I(n616), .Z(n615) );
  CKNXD0 U26 ( .I(n615), .ZN(n4686) );
  CKBXD0 U29 ( .I(n562), .Z(n561) );
  CKNXD0 U30 ( .I(n561), .ZN(n4689) );
  BUFFD0 U31 ( .I(n5), .Z(n1) );
  BUFFD0 U32 ( .I(n6), .Z(n2) );
  BUFFD0 U37 ( .I(n7), .Z(n3) );
  XOR3D0 U38 ( .A1(n4647), .A2(n4644), .A3(n73), .Z(N85) );
  BUFFD0 U39 ( .I(n4691), .Z(n5) );
  BUFFD0 U40 ( .I(n4673), .Z(n6) );
  BUFFD0 U41 ( .I(n4655), .Z(n7) );
  BUFFD0 U42 ( .I(n4647), .Z(n8) );
  BUFFD0 U43 ( .I(n4721), .Z(n10) );
  BUFFD0 U44 ( .I(n12), .Z(n11) );
  BUFFD0 U45 ( .I(n13), .Z(n12) );
  BUFFD0 U46 ( .I(n14), .Z(n13) );
  BUFFD0 U47 ( .I(n15), .Z(n14) );
  BUFFD0 U48 ( .I(n16), .Z(n15) );
  BUFFD0 U49 ( .I(n17), .Z(n16) );
  BUFFD0 U50 ( .I(n18), .Z(n17) );
  BUFFD0 U51 ( .I(n19), .Z(n18) );
  BUFFD0 U52 ( .I(n20), .Z(n19) );
  BUFFD0 U53 ( .I(n21), .Z(n20) );
  BUFFD0 U54 ( .I(n22), .Z(n21) );
  BUFFD0 U55 ( .I(n23), .Z(n22) );
  BUFFD0 U56 ( .I(n24), .Z(n23) );
  BUFFD0 U57 ( .I(n25), .Z(n24) );
  BUFFD0 U58 ( .I(n26), .Z(n25) );
  BUFFD0 U59 ( .I(n27), .Z(n26) );
  BUFFD0 U60 ( .I(n28), .Z(n27) );
  BUFFD0 U61 ( .I(n29), .Z(n28) );
  BUFFD0 U62 ( .I(n30), .Z(n29) );
  BUFFD0 U63 ( .I(n31), .Z(n30) );
  BUFFD0 U64 ( .I(n32), .Z(n31) );
  BUFFD0 U65 ( .I(n33), .Z(n32) );
  BUFFD0 U66 ( .I(n34), .Z(n33) );
  BUFFD0 U67 ( .I(n35), .Z(n34) );
  BUFFD0 U68 ( .I(n36), .Z(n35) );
  BUFFD0 U69 ( .I(n37), .Z(n36) );
  BUFFD0 U70 ( .I(n38), .Z(n37) );
  BUFFD0 U71 ( .I(n39), .Z(n38) );
  BUFFD0 U72 ( .I(n40), .Z(n39) );
  BUFFD0 U73 ( .I(n41), .Z(n40) );
  BUFFD0 U74 ( .I(n42), .Z(n41) );
  BUFFD0 U75 ( .I(n43), .Z(n42) );
  BUFFD0 U76 ( .I(n44), .Z(n43) );
  BUFFD0 U77 ( .I(n4722), .Z(n44) );
  BUFFD0 U78 ( .I(n46), .Z(n45) );
  BUFFD0 U79 ( .I(n4718), .Z(n46) );
  BUFFD0 U80 ( .I(n48), .Z(n47) );
  BUFFD0 U81 ( .I(n49), .Z(n48) );
  BUFFD0 U82 ( .I(n50), .Z(n49) );
  BUFFD0 U83 ( .I(n51), .Z(n50) );
  BUFFD0 U84 ( .I(n52), .Z(n51) );
  BUFFD0 U85 ( .I(n53), .Z(n52) );
  BUFFD0 U86 ( .I(n54), .Z(n53) );
  BUFFD0 U87 ( .I(n55), .Z(n54) );
  BUFFD0 U88 ( .I(n56), .Z(n55) );
  BUFFD0 U89 ( .I(n57), .Z(n56) );
  BUFFD0 U90 ( .I(n58), .Z(n57) );
  BUFFD0 U91 ( .I(n59), .Z(n58) );
  BUFFD0 U92 ( .I(n60), .Z(n59) );
  BUFFD0 U93 ( .I(n61), .Z(n60) );
  BUFFD0 U94 ( .I(n62), .Z(n61) );
  BUFFD0 U95 ( .I(n63), .Z(n62) );
  BUFFD0 U96 ( .I(n64), .Z(n63) );
  BUFFD0 U97 ( .I(n65), .Z(n64) );
  BUFFD0 U98 ( .I(n107), .Z(n65) );
  BUFFD0 U99 ( .I(n109), .Z(n107) );
  BUFFD0 U100 ( .I(n110), .Z(n109) );
  BUFFD0 U101 ( .I(n111), .Z(n110) );
  BUFFD0 U102 ( .I(n112), .Z(n111) );
  BUFFD0 U103 ( .I(n113), .Z(n112) );
  BUFFD0 U104 ( .I(n114), .Z(n113) );
  BUFFD0 U105 ( .I(n115), .Z(n114) );
  BUFFD0 U106 ( .I(n116), .Z(n115) );
  BUFFD0 U107 ( .I(n117), .Z(n116) );
  BUFFD0 U108 ( .I(n118), .Z(n117) );
  BUFFD0 U109 ( .I(n119), .Z(n118) );
  BUFFD0 U110 ( .I(n120), .Z(n119) );
  BUFFD0 U111 ( .I(n121), .Z(n120) );
  BUFFD0 U112 ( .I(n122), .Z(n121) );
  BUFFD0 U113 ( .I(n123), .Z(n122) );
  BUFFD0 U114 ( .I(n124), .Z(n123) );
  BUFFD0 U115 ( .I(n125), .Z(n124) );
  BUFFD0 U116 ( .I(n126), .Z(n125) );
  BUFFD0 U117 ( .I(n127), .Z(n126) );
  BUFFD0 U118 ( .I(n128), .Z(n127) );
  BUFFD0 U119 ( .I(n129), .Z(n128) );
  BUFFD0 U120 ( .I(n130), .Z(n129) );
  BUFFD0 U121 ( .I(n131), .Z(n130) );
  BUFFD0 U122 ( .I(n132), .Z(n131) );
  BUFFD0 U123 ( .I(n133), .Z(n132) );
  BUFFD0 U124 ( .I(n134), .Z(n133) );
  BUFFD0 U125 ( .I(n135), .Z(n134) );
  BUFFD0 U126 ( .I(n136), .Z(n135) );
  BUFFD0 U127 ( .I(n137), .Z(n136) );
  BUFFD0 U128 ( .I(n138), .Z(n137) );
  BUFFD0 U129 ( .I(n4719), .Z(n138) );
  BUFFD0 U130 ( .I(n140), .Z(n139) );
  BUFFD0 U131 ( .I(n4716), .Z(n140) );
  BUFFD0 U132 ( .I(n142), .Z(n141) );
  BUFFD0 U133 ( .I(n143), .Z(n142) );
  BUFFD0 U134 ( .I(n144), .Z(n143) );
  BUFFD0 U135 ( .I(n145), .Z(n144) );
  BUFFD0 U136 ( .I(n146), .Z(n145) );
  BUFFD0 U137 ( .I(n147), .Z(n146) );
  BUFFD0 U138 ( .I(n148), .Z(n147) );
  BUFFD0 U139 ( .I(n149), .Z(n148) );
  BUFFD0 U140 ( .I(n150), .Z(n149) );
  BUFFD0 U141 ( .I(n151), .Z(n150) );
  BUFFD0 U142 ( .I(n152), .Z(n151) );
  BUFFD0 U143 ( .I(n153), .Z(n152) );
  BUFFD0 U144 ( .I(n154), .Z(n153) );
  BUFFD0 U145 ( .I(n155), .Z(n154) );
  BUFFD0 U146 ( .I(n156), .Z(n155) );
  BUFFD0 U147 ( .I(n157), .Z(n156) );
  BUFFD0 U148 ( .I(n158), .Z(n157) );
  BUFFD0 U149 ( .I(n159), .Z(n158) );
  BUFFD0 U150 ( .I(n160), .Z(n159) );
  BUFFD0 U151 ( .I(n161), .Z(n160) );
  BUFFD0 U152 ( .I(n162), .Z(n161) );
  BUFFD0 U153 ( .I(n163), .Z(n162) );
  BUFFD0 U154 ( .I(n164), .Z(n163) );
  BUFFD0 U155 ( .I(n165), .Z(n164) );
  BUFFD0 U156 ( .I(n166), .Z(n165) );
  BUFFD0 U157 ( .I(n167), .Z(n166) );
  BUFFD0 U158 ( .I(n168), .Z(n167) );
  BUFFD0 U159 ( .I(n169), .Z(n168) );
  BUFFD0 U160 ( .I(n170), .Z(n169) );
  BUFFD0 U161 ( .I(n171), .Z(n170) );
  BUFFD0 U162 ( .I(n172), .Z(n171) );
  BUFFD0 U163 ( .I(n173), .Z(n172) );
  BUFFD0 U164 ( .I(n174), .Z(n173) );
  BUFFD0 U165 ( .I(n175), .Z(n174) );
  BUFFD0 U166 ( .I(n176), .Z(n175) );
  BUFFD0 U167 ( .I(n177), .Z(n176) );
  BUFFD0 U168 ( .I(n178), .Z(n177) );
  BUFFD0 U169 ( .I(n179), .Z(n178) );
  BUFFD0 U170 ( .I(n180), .Z(n179) );
  BUFFD0 U171 ( .I(n181), .Z(n180) );
  BUFFD0 U172 ( .I(n182), .Z(n181) );
  BUFFD0 U173 ( .I(n183), .Z(n182) );
  BUFFD0 U174 ( .I(n184), .Z(n183) );
  BUFFD0 U175 ( .I(n185), .Z(n184) );
  BUFFD0 U176 ( .I(n186), .Z(n185) );
  BUFFD0 U177 ( .I(n187), .Z(n186) );
  BUFFD0 U178 ( .I(n188), .Z(n187) );
  BUFFD0 U179 ( .I(n189), .Z(n188) );
  BUFFD0 U180 ( .I(n190), .Z(n189) );
  BUFFD0 U181 ( .I(n4717), .Z(n190) );
  BUFFD0 U182 ( .I(n4714), .Z(n191) );
  BUFFD0 U183 ( .I(n193), .Z(n192) );
  BUFFD0 U184 ( .I(n194), .Z(n193) );
  BUFFD0 U185 ( .I(n195), .Z(n194) );
  BUFFD0 U186 ( .I(n196), .Z(n195) );
  BUFFD0 U187 ( .I(n197), .Z(n196) );
  BUFFD0 U188 ( .I(n198), .Z(n197) );
  BUFFD0 U189 ( .I(n199), .Z(n198) );
  BUFFD0 U190 ( .I(n200), .Z(n199) );
  BUFFD0 U191 ( .I(n201), .Z(n200) );
  BUFFD0 U192 ( .I(n202), .Z(n201) );
  BUFFD0 U193 ( .I(n203), .Z(n202) );
  BUFFD0 U194 ( .I(n204), .Z(n203) );
  BUFFD0 U195 ( .I(n205), .Z(n204) );
  BUFFD0 U196 ( .I(n206), .Z(n205) );
  BUFFD0 U197 ( .I(n207), .Z(n206) );
  BUFFD0 U198 ( .I(n208), .Z(n207) );
  BUFFD0 U199 ( .I(n209), .Z(n208) );
  BUFFD0 U200 ( .I(n210), .Z(n209) );
  BUFFD0 U201 ( .I(n211), .Z(n210) );
  BUFFD0 U202 ( .I(n212), .Z(n211) );
  BUFFD0 U203 ( .I(n213), .Z(n212) );
  BUFFD0 U204 ( .I(n214), .Z(n213) );
  BUFFD0 U205 ( .I(n215), .Z(n214) );
  BUFFD0 U206 ( .I(n216), .Z(n215) );
  BUFFD0 U207 ( .I(n217), .Z(n216) );
  BUFFD0 U208 ( .I(n218), .Z(n217) );
  BUFFD0 U209 ( .I(n219), .Z(n218) );
  BUFFD0 U210 ( .I(n220), .Z(n219) );
  BUFFD0 U211 ( .I(n221), .Z(n220) );
  BUFFD0 U212 ( .I(n222), .Z(n221) );
  BUFFD0 U213 ( .I(n223), .Z(n222) );
  BUFFD0 U214 ( .I(n224), .Z(n223) );
  BUFFD0 U215 ( .I(n225), .Z(n224) );
  BUFFD0 U216 ( .I(n226), .Z(n225) );
  BUFFD0 U217 ( .I(n227), .Z(n226) );
  BUFFD0 U218 ( .I(n228), .Z(n227) );
  BUFFD0 U219 ( .I(n229), .Z(n228) );
  BUFFD0 U220 ( .I(n230), .Z(n229) );
  BUFFD0 U221 ( .I(n231), .Z(n230) );
  BUFFD0 U222 ( .I(n232), .Z(n231) );
  BUFFD0 U223 ( .I(n233), .Z(n232) );
  BUFFD0 U224 ( .I(n234), .Z(n233) );
  BUFFD0 U225 ( .I(n235), .Z(n234) );
  BUFFD0 U226 ( .I(n236), .Z(n235) );
  BUFFD0 U227 ( .I(n237), .Z(n236) );
  BUFFD0 U228 ( .I(n238), .Z(n237) );
  BUFFD0 U229 ( .I(n239), .Z(n238) );
  BUFFD0 U230 ( .I(n240), .Z(n239) );
  BUFFD0 U231 ( .I(n241), .Z(n240) );
  BUFFD0 U232 ( .I(n242), .Z(n241) );
  BUFFD0 U233 ( .I(n243), .Z(n242) );
  BUFFD0 U234 ( .I(n244), .Z(n243) );
  BUFFD0 U235 ( .I(n4715), .Z(n244) );
  BUFFD0 U236 ( .I(n4704), .Z(n245) );
  BUFFD0 U237 ( .I(n247), .Z(n246) );
  BUFFD0 U238 ( .I(n248), .Z(n247) );
  BUFFD0 U239 ( .I(n249), .Z(n248) );
  BUFFD0 U240 ( .I(n250), .Z(n249) );
  BUFFD0 U241 ( .I(n251), .Z(n250) );
  BUFFD0 U242 ( .I(n252), .Z(n251) );
  BUFFD0 U243 ( .I(n253), .Z(n252) );
  BUFFD0 U244 ( .I(n254), .Z(n253) );
  BUFFD0 U245 ( .I(n255), .Z(n254) );
  BUFFD0 U246 ( .I(n256), .Z(n255) );
  BUFFD0 U247 ( .I(n257), .Z(n256) );
  BUFFD0 U248 ( .I(n258), .Z(n257) );
  BUFFD0 U249 ( .I(n259), .Z(n258) );
  BUFFD0 U250 ( .I(n260), .Z(n259) );
  BUFFD0 U251 ( .I(n261), .Z(n260) );
  BUFFD0 U252 ( .I(n262), .Z(n261) );
  BUFFD0 U253 ( .I(n263), .Z(n262) );
  BUFFD0 U254 ( .I(n264), .Z(n263) );
  BUFFD0 U255 ( .I(n265), .Z(n264) );
  BUFFD0 U256 ( .I(n266), .Z(n265) );
  BUFFD0 U257 ( .I(n267), .Z(n266) );
  BUFFD0 U258 ( .I(n268), .Z(n267) );
  BUFFD0 U259 ( .I(n269), .Z(n268) );
  BUFFD0 U260 ( .I(n270), .Z(n269) );
  BUFFD0 U261 ( .I(n271), .Z(n270) );
  BUFFD0 U262 ( .I(n272), .Z(n271) );
  BUFFD0 U263 ( .I(n273), .Z(n272) );
  BUFFD0 U264 ( .I(n274), .Z(n273) );
  BUFFD0 U265 ( .I(n275), .Z(n274) );
  BUFFD0 U266 ( .I(n276), .Z(n275) );
  BUFFD0 U267 ( .I(n277), .Z(n276) );
  BUFFD0 U268 ( .I(n278), .Z(n277) );
  BUFFD0 U269 ( .I(n279), .Z(n278) );
  BUFFD0 U270 ( .I(n280), .Z(n279) );
  BUFFD0 U271 ( .I(n281), .Z(n280) );
  BUFFD0 U272 ( .I(n282), .Z(n281) );
  BUFFD0 U273 ( .I(n283), .Z(n282) );
  BUFFD0 U274 ( .I(n284), .Z(n283) );
  BUFFD0 U275 ( .I(n285), .Z(n284) );
  BUFFD0 U276 ( .I(n286), .Z(n285) );
  BUFFD0 U277 ( .I(n287), .Z(n286) );
  BUFFD0 U278 ( .I(n288), .Z(n287) );
  BUFFD0 U279 ( .I(n289), .Z(n288) );
  BUFFD0 U280 ( .I(n290), .Z(n289) );
  BUFFD0 U281 ( .I(n291), .Z(n290) );
  BUFFD0 U282 ( .I(n292), .Z(n291) );
  BUFFD0 U283 ( .I(n293), .Z(n292) );
  BUFFD0 U284 ( .I(n294), .Z(n293) );
  BUFFD0 U285 ( .I(n295), .Z(n294) );
  BUFFD0 U286 ( .I(n296), .Z(n295) );
  BUFFD0 U287 ( .I(n297), .Z(n296) );
  BUFFD0 U288 ( .I(n298), .Z(n297) );
  BUFFD0 U289 ( .I(n4705), .Z(n298) );
  BUFFD0 U290 ( .I(n4701), .Z(n299) );
  BUFFD0 U291 ( .I(n301), .Z(n300) );
  BUFFD0 U292 ( .I(n302), .Z(n301) );
  BUFFD0 U293 ( .I(n303), .Z(n302) );
  BUFFD0 U294 ( .I(n304), .Z(n303) );
  BUFFD0 U295 ( .I(n305), .Z(n304) );
  BUFFD0 U296 ( .I(n306), .Z(n305) );
  BUFFD0 U297 ( .I(n307), .Z(n306) );
  BUFFD0 U298 ( .I(n308), .Z(n307) );
  BUFFD0 U299 ( .I(n309), .Z(n308) );
  BUFFD0 U300 ( .I(n310), .Z(n309) );
  BUFFD0 U301 ( .I(n311), .Z(n310) );
  BUFFD0 U302 ( .I(n312), .Z(n311) );
  BUFFD0 U303 ( .I(n313), .Z(n312) );
  BUFFD0 U304 ( .I(n314), .Z(n313) );
  BUFFD0 U305 ( .I(n315), .Z(n314) );
  BUFFD0 U306 ( .I(n316), .Z(n315) );
  BUFFD0 U307 ( .I(n317), .Z(n316) );
  BUFFD0 U308 ( .I(n318), .Z(n317) );
  BUFFD0 U309 ( .I(n319), .Z(n318) );
  BUFFD0 U310 ( .I(n320), .Z(n319) );
  BUFFD0 U311 ( .I(n321), .Z(n320) );
  BUFFD0 U312 ( .I(n322), .Z(n321) );
  BUFFD0 U313 ( .I(n323), .Z(n322) );
  BUFFD0 U314 ( .I(n324), .Z(n323) );
  BUFFD0 U315 ( .I(n325), .Z(n324) );
  BUFFD0 U316 ( .I(n326), .Z(n325) );
  BUFFD0 U317 ( .I(n327), .Z(n326) );
  BUFFD0 U318 ( .I(n328), .Z(n327) );
  BUFFD0 U319 ( .I(n329), .Z(n328) );
  BUFFD0 U320 ( .I(n330), .Z(n329) );
  BUFFD0 U321 ( .I(n331), .Z(n330) );
  BUFFD0 U322 ( .I(n332), .Z(n331) );
  BUFFD0 U323 ( .I(n333), .Z(n332) );
  BUFFD0 U324 ( .I(n334), .Z(n333) );
  BUFFD0 U325 ( .I(n335), .Z(n334) );
  BUFFD0 U326 ( .I(n336), .Z(n335) );
  BUFFD0 U327 ( .I(n337), .Z(n336) );
  BUFFD0 U328 ( .I(n338), .Z(n337) );
  BUFFD0 U329 ( .I(n339), .Z(n338) );
  BUFFD0 U330 ( .I(n340), .Z(n339) );
  BUFFD0 U331 ( .I(n341), .Z(n340) );
  BUFFD0 U332 ( .I(n342), .Z(n341) );
  BUFFD0 U333 ( .I(n343), .Z(n342) );
  BUFFD0 U334 ( .I(n344), .Z(n343) );
  BUFFD0 U335 ( .I(n345), .Z(n344) );
  BUFFD0 U336 ( .I(n346), .Z(n345) );
  BUFFD0 U337 ( .I(n347), .Z(n346) );
  BUFFD0 U338 ( .I(n348), .Z(n347) );
  BUFFD0 U339 ( .I(n349), .Z(n348) );
  BUFFD0 U340 ( .I(n350), .Z(n349) );
  BUFFD0 U341 ( .I(n351), .Z(n350) );
  BUFFD0 U342 ( .I(n352), .Z(n351) );
  BUFFD0 U343 ( .I(n4702), .Z(n352) );
  BUFFD0 U344 ( .I(n354), .Z(n353) );
  BUFFD0 U345 ( .I(n4698), .Z(n354) );
  BUFFD0 U346 ( .I(n356), .Z(n355) );
  BUFFD0 U347 ( .I(n357), .Z(n356) );
  BUFFD0 U348 ( .I(n358), .Z(n357) );
  BUFFD0 U349 ( .I(n359), .Z(n358) );
  BUFFD0 U350 ( .I(n360), .Z(n359) );
  BUFFD0 U351 ( .I(n361), .Z(n360) );
  BUFFD0 U352 ( .I(n362), .Z(n361) );
  BUFFD0 U353 ( .I(n363), .Z(n362) );
  BUFFD0 U354 ( .I(n364), .Z(n363) );
  BUFFD0 U355 ( .I(n365), .Z(n364) );
  BUFFD0 U356 ( .I(n366), .Z(n365) );
  BUFFD0 U357 ( .I(n367), .Z(n366) );
  BUFFD0 U358 ( .I(n368), .Z(n367) );
  BUFFD0 U359 ( .I(n369), .Z(n368) );
  BUFFD0 U360 ( .I(n370), .Z(n369) );
  BUFFD0 U361 ( .I(n371), .Z(n370) );
  BUFFD0 U362 ( .I(n372), .Z(n371) );
  BUFFD0 U363 ( .I(n373), .Z(n372) );
  BUFFD0 U364 ( .I(n374), .Z(n373) );
  BUFFD0 U365 ( .I(n375), .Z(n374) );
  BUFFD0 U366 ( .I(n376), .Z(n375) );
  BUFFD0 U367 ( .I(n377), .Z(n376) );
  BUFFD0 U368 ( .I(n378), .Z(n377) );
  BUFFD0 U369 ( .I(n379), .Z(n378) );
  BUFFD0 U370 ( .I(n380), .Z(n379) );
  BUFFD0 U371 ( .I(n381), .Z(n380) );
  BUFFD0 U372 ( .I(n382), .Z(n381) );
  BUFFD0 U373 ( .I(n383), .Z(n382) );
  BUFFD0 U374 ( .I(n384), .Z(n383) );
  BUFFD0 U375 ( .I(n385), .Z(n384) );
  BUFFD0 U376 ( .I(n386), .Z(n385) );
  BUFFD0 U377 ( .I(n387), .Z(n386) );
  BUFFD0 U378 ( .I(n388), .Z(n387) );
  BUFFD0 U379 ( .I(n389), .Z(n388) );
  BUFFD0 U380 ( .I(n390), .Z(n389) );
  BUFFD0 U381 ( .I(n391), .Z(n390) );
  BUFFD0 U382 ( .I(n392), .Z(n391) );
  BUFFD0 U383 ( .I(n393), .Z(n392) );
  BUFFD0 U384 ( .I(n394), .Z(n393) );
  BUFFD0 U385 ( .I(n395), .Z(n394) );
  BUFFD0 U386 ( .I(n396), .Z(n395) );
  BUFFD0 U387 ( .I(n397), .Z(n396) );
  BUFFD0 U388 ( .I(n398), .Z(n397) );
  BUFFD0 U389 ( .I(n399), .Z(n398) );
  BUFFD0 U390 ( .I(n400), .Z(n399) );
  BUFFD0 U391 ( .I(n401), .Z(n400) );
  BUFFD0 U392 ( .I(n402), .Z(n401) );
  BUFFD0 U393 ( .I(n403), .Z(n402) );
  BUFFD0 U394 ( .I(n404), .Z(n403) );
  BUFFD0 U395 ( .I(n4699), .Z(n404) );
  BUFFD0 U396 ( .I(n406), .Z(n405) );
  BUFFD0 U397 ( .I(n4696), .Z(n406) );
  BUFFD0 U398 ( .I(n408), .Z(n407) );
  BUFFD0 U399 ( .I(n409), .Z(n408) );
  BUFFD0 U400 ( .I(n410), .Z(n409) );
  BUFFD0 U401 ( .I(n411), .Z(n410) );
  BUFFD0 U402 ( .I(n412), .Z(n411) );
  BUFFD0 U403 ( .I(n413), .Z(n412) );
  BUFFD0 U404 ( .I(n414), .Z(n413) );
  BUFFD0 U405 ( .I(n415), .Z(n414) );
  BUFFD0 U406 ( .I(n416), .Z(n415) );
  BUFFD0 U407 ( .I(n417), .Z(n416) );
  BUFFD0 U408 ( .I(n418), .Z(n417) );
  BUFFD0 U409 ( .I(n419), .Z(n418) );
  BUFFD0 U410 ( .I(n420), .Z(n419) );
  BUFFD0 U411 ( .I(n421), .Z(n420) );
  BUFFD0 U412 ( .I(n422), .Z(n421) );
  BUFFD0 U413 ( .I(n423), .Z(n422) );
  BUFFD0 U414 ( .I(n424), .Z(n423) );
  BUFFD0 U415 ( .I(n425), .Z(n424) );
  BUFFD0 U416 ( .I(n426), .Z(n425) );
  BUFFD0 U417 ( .I(n427), .Z(n426) );
  BUFFD0 U418 ( .I(n428), .Z(n427) );
  BUFFD0 U419 ( .I(n429), .Z(n428) );
  BUFFD0 U420 ( .I(n430), .Z(n429) );
  BUFFD0 U421 ( .I(n431), .Z(n430) );
  BUFFD0 U422 ( .I(n432), .Z(n431) );
  BUFFD0 U423 ( .I(n433), .Z(n432) );
  BUFFD0 U424 ( .I(n434), .Z(n433) );
  BUFFD0 U425 ( .I(n435), .Z(n434) );
  BUFFD0 U426 ( .I(n436), .Z(n435) );
  BUFFD0 U427 ( .I(n437), .Z(n436) );
  BUFFD0 U428 ( .I(n438), .Z(n437) );
  BUFFD0 U429 ( .I(n439), .Z(n438) );
  BUFFD0 U430 ( .I(n440), .Z(n439) );
  BUFFD0 U431 ( .I(n441), .Z(n440) );
  BUFFD0 U432 ( .I(n442), .Z(n441) );
  BUFFD0 U433 ( .I(n443), .Z(n442) );
  BUFFD0 U434 ( .I(n444), .Z(n443) );
  BUFFD0 U435 ( .I(n445), .Z(n444) );
  BUFFD0 U436 ( .I(n446), .Z(n445) );
  BUFFD0 U437 ( .I(n447), .Z(n446) );
  BUFFD0 U438 ( .I(n448), .Z(n447) );
  BUFFD0 U439 ( .I(n449), .Z(n448) );
  BUFFD0 U440 ( .I(n450), .Z(n449) );
  BUFFD0 U441 ( .I(n451), .Z(n450) );
  BUFFD0 U442 ( .I(n452), .Z(n451) );
  BUFFD0 U443 ( .I(n453), .Z(n452) );
  BUFFD0 U444 ( .I(n454), .Z(n453) );
  BUFFD0 U445 ( .I(n455), .Z(n454) );
  BUFFD0 U446 ( .I(n456), .Z(n455) );
  BUFFD0 U447 ( .I(n4697), .Z(n456) );
  BUFFD0 U448 ( .I(n4694), .Z(n457) );
  BUFFD0 U449 ( .I(n459), .Z(n458) );
  BUFFD0 U450 ( .I(n460), .Z(n459) );
  BUFFD0 U451 ( .I(n461), .Z(n460) );
  BUFFD0 U452 ( .I(n462), .Z(n461) );
  BUFFD0 U453 ( .I(n463), .Z(n462) );
  BUFFD0 U454 ( .I(n464), .Z(n463) );
  BUFFD0 U455 ( .I(n465), .Z(n464) );
  BUFFD0 U456 ( .I(n466), .Z(n465) );
  BUFFD0 U457 ( .I(n467), .Z(n466) );
  BUFFD0 U458 ( .I(n468), .Z(n467) );
  BUFFD0 U459 ( .I(n469), .Z(n468) );
  BUFFD0 U460 ( .I(n470), .Z(n469) );
  BUFFD0 U461 ( .I(n471), .Z(n470) );
  BUFFD0 U462 ( .I(n472), .Z(n471) );
  BUFFD0 U463 ( .I(n473), .Z(n472) );
  BUFFD0 U464 ( .I(n474), .Z(n473) );
  BUFFD0 U465 ( .I(n475), .Z(n474) );
  BUFFD0 U466 ( .I(n476), .Z(n475) );
  BUFFD0 U467 ( .I(n477), .Z(n476) );
  BUFFD0 U468 ( .I(n478), .Z(n477) );
  BUFFD0 U469 ( .I(n479), .Z(n478) );
  BUFFD0 U470 ( .I(n480), .Z(n479) );
  BUFFD0 U471 ( .I(n481), .Z(n480) );
  BUFFD0 U472 ( .I(n482), .Z(n481) );
  BUFFD0 U473 ( .I(n483), .Z(n482) );
  BUFFD0 U474 ( .I(n484), .Z(n483) );
  BUFFD0 U475 ( .I(n485), .Z(n484) );
  BUFFD0 U476 ( .I(n486), .Z(n485) );
  BUFFD0 U477 ( .I(n487), .Z(n486) );
  BUFFD0 U478 ( .I(n488), .Z(n487) );
  BUFFD0 U479 ( .I(n489), .Z(n488) );
  BUFFD0 U480 ( .I(n490), .Z(n489) );
  BUFFD0 U481 ( .I(n491), .Z(n490) );
  BUFFD0 U482 ( .I(n492), .Z(n491) );
  BUFFD0 U483 ( .I(n493), .Z(n492) );
  BUFFD0 U484 ( .I(n494), .Z(n493) );
  BUFFD0 U485 ( .I(n495), .Z(n494) );
  BUFFD0 U486 ( .I(n496), .Z(n495) );
  BUFFD0 U487 ( .I(n497), .Z(n496) );
  BUFFD0 U488 ( .I(n498), .Z(n497) );
  BUFFD0 U489 ( .I(n499), .Z(n498) );
  BUFFD0 U490 ( .I(n500), .Z(n499) );
  BUFFD0 U491 ( .I(n501), .Z(n500) );
  BUFFD0 U492 ( .I(n502), .Z(n501) );
  BUFFD0 U493 ( .I(n503), .Z(n502) );
  BUFFD0 U494 ( .I(n504), .Z(n503) );
  BUFFD0 U495 ( .I(n505), .Z(n504) );
  BUFFD0 U496 ( .I(n506), .Z(n505) );
  BUFFD0 U497 ( .I(n507), .Z(n506) );
  BUFFD0 U498 ( .I(n508), .Z(n507) );
  BUFFD0 U499 ( .I(n509), .Z(n508) );
  BUFFD0 U500 ( .I(n510), .Z(n509) );
  BUFFD0 U501 ( .I(n4695), .Z(n510) );
  BUFFD0 U502 ( .I(n512), .Z(n511) );
  BUFFD0 U503 ( .I(n513), .Z(n512) );
  BUFFD0 U504 ( .I(n514), .Z(n513) );
  BUFFD0 U505 ( .I(n515), .Z(n514) );
  BUFFD0 U506 ( .I(n516), .Z(n515) );
  BUFFD0 U507 ( .I(n517), .Z(n516) );
  BUFFD0 U508 ( .I(n518), .Z(n517) );
  BUFFD0 U509 ( .I(n519), .Z(n518) );
  BUFFD0 U510 ( .I(n520), .Z(n519) );
  BUFFD0 U511 ( .I(n521), .Z(n520) );
  BUFFD0 U512 ( .I(n522), .Z(n521) );
  BUFFD0 U513 ( .I(n523), .Z(n522) );
  BUFFD0 U514 ( .I(n524), .Z(n523) );
  BUFFD0 U515 ( .I(n525), .Z(n524) );
  BUFFD0 U516 ( .I(n526), .Z(n525) );
  BUFFD0 U517 ( .I(n527), .Z(n526) );
  BUFFD0 U518 ( .I(n528), .Z(n527) );
  BUFFD0 U519 ( .I(n529), .Z(n528) );
  BUFFD0 U520 ( .I(n530), .Z(n529) );
  BUFFD0 U521 ( .I(n531), .Z(n530) );
  BUFFD0 U522 ( .I(n532), .Z(n531) );
  BUFFD0 U523 ( .I(n533), .Z(n532) );
  BUFFD0 U524 ( .I(n534), .Z(n533) );
  BUFFD0 U525 ( .I(n535), .Z(n534) );
  BUFFD0 U526 ( .I(n536), .Z(n535) );
  BUFFD0 U527 ( .I(n537), .Z(n536) );
  BUFFD0 U528 ( .I(n538), .Z(n537) );
  BUFFD0 U529 ( .I(n539), .Z(n538) );
  BUFFD0 U530 ( .I(n540), .Z(n539) );
  BUFFD0 U531 ( .I(n541), .Z(n540) );
  BUFFD0 U532 ( .I(n542), .Z(n541) );
  BUFFD0 U533 ( .I(n543), .Z(n542) );
  BUFFD0 U534 ( .I(n544), .Z(n543) );
  BUFFD0 U535 ( .I(n545), .Z(n544) );
  BUFFD0 U536 ( .I(n546), .Z(n545) );
  BUFFD0 U537 ( .I(n547), .Z(n546) );
  BUFFD0 U538 ( .I(n548), .Z(n547) );
  BUFFD0 U539 ( .I(n549), .Z(n548) );
  BUFFD0 U540 ( .I(n550), .Z(n549) );
  BUFFD0 U541 ( .I(n551), .Z(n550) );
  BUFFD0 U542 ( .I(n552), .Z(n551) );
  BUFFD0 U543 ( .I(n553), .Z(n552) );
  BUFFD0 U544 ( .I(n554), .Z(n553) );
  BUFFD0 U545 ( .I(n555), .Z(n554) );
  BUFFD0 U546 ( .I(n556), .Z(n555) );
  BUFFD0 U547 ( .I(n557), .Z(n556) );
  BUFFD0 U548 ( .I(n558), .Z(n557) );
  BUFFD0 U549 ( .I(n559), .Z(n558) );
  BUFFD0 U550 ( .I(n560), .Z(n559) );
  BUFFD0 U551 ( .I(n4692), .Z(n560) );
  BUFFD0 U552 ( .I(n563), .Z(n562) );
  BUFFD0 U553 ( .I(n564), .Z(n563) );
  BUFFD0 U554 ( .I(n565), .Z(n564) );
  BUFFD0 U555 ( .I(n566), .Z(n565) );
  BUFFD0 U556 ( .I(n567), .Z(n566) );
  BUFFD0 U557 ( .I(n568), .Z(n567) );
  BUFFD0 U558 ( .I(n569), .Z(n568) );
  BUFFD0 U559 ( .I(n570), .Z(n569) );
  BUFFD0 U560 ( .I(n571), .Z(n570) );
  BUFFD0 U561 ( .I(n572), .Z(n571) );
  BUFFD0 U562 ( .I(n573), .Z(n572) );
  BUFFD0 U563 ( .I(n574), .Z(n573) );
  BUFFD0 U564 ( .I(n575), .Z(n574) );
  BUFFD0 U565 ( .I(n576), .Z(n575) );
  BUFFD0 U566 ( .I(n577), .Z(n576) );
  BUFFD0 U567 ( .I(n578), .Z(n577) );
  BUFFD0 U568 ( .I(n579), .Z(n578) );
  BUFFD0 U569 ( .I(n580), .Z(n579) );
  BUFFD0 U570 ( .I(n581), .Z(n580) );
  BUFFD0 U571 ( .I(n582), .Z(n581) );
  BUFFD0 U572 ( .I(n583), .Z(n582) );
  BUFFD0 U573 ( .I(n584), .Z(n583) );
  BUFFD0 U574 ( .I(n585), .Z(n584) );
  BUFFD0 U575 ( .I(n586), .Z(n585) );
  BUFFD0 U576 ( .I(n587), .Z(n586) );
  BUFFD0 U577 ( .I(n588), .Z(n587) );
  BUFFD0 U578 ( .I(n589), .Z(n588) );
  BUFFD0 U579 ( .I(n590), .Z(n589) );
  BUFFD0 U580 ( .I(n591), .Z(n590) );
  BUFFD0 U581 ( .I(n592), .Z(n591) );
  BUFFD0 U582 ( .I(n593), .Z(n592) );
  BUFFD0 U583 ( .I(n594), .Z(n593) );
  BUFFD0 U584 ( .I(n595), .Z(n594) );
  BUFFD0 U585 ( .I(n596), .Z(n595) );
  BUFFD0 U586 ( .I(n597), .Z(n596) );
  BUFFD0 U587 ( .I(n598), .Z(n597) );
  BUFFD0 U588 ( .I(n599), .Z(n598) );
  BUFFD0 U589 ( .I(n600), .Z(n599) );
  BUFFD0 U590 ( .I(n601), .Z(n600) );
  BUFFD0 U591 ( .I(n602), .Z(n601) );
  BUFFD0 U592 ( .I(n603), .Z(n602) );
  BUFFD0 U593 ( .I(n604), .Z(n603) );
  BUFFD0 U594 ( .I(n605), .Z(n604) );
  BUFFD0 U595 ( .I(n606), .Z(n605) );
  BUFFD0 U596 ( .I(n607), .Z(n606) );
  BUFFD0 U597 ( .I(n608), .Z(n607) );
  BUFFD0 U598 ( .I(n609), .Z(n608) );
  BUFFD0 U599 ( .I(n610), .Z(n609) );
  BUFFD0 U600 ( .I(n611), .Z(n610) );
  BUFFD0 U601 ( .I(n612), .Z(n611) );
  BUFFD0 U602 ( .I(n613), .Z(n612) );
  BUFFD0 U603 ( .I(n614), .Z(n613) );
  BUFFD0 U604 ( .I(n4690), .Z(n614) );
  BUFFD0 U605 ( .I(n617), .Z(n616) );
  BUFFD0 U606 ( .I(n618), .Z(n617) );
  BUFFD0 U607 ( .I(n619), .Z(n618) );
  BUFFD0 U608 ( .I(n620), .Z(n619) );
  BUFFD0 U609 ( .I(n621), .Z(n620) );
  BUFFD0 U610 ( .I(n622), .Z(n621) );
  BUFFD0 U611 ( .I(n623), .Z(n622) );
  BUFFD0 U612 ( .I(n624), .Z(n623) );
  BUFFD0 U613 ( .I(n625), .Z(n624) );
  BUFFD0 U614 ( .I(n626), .Z(n625) );
  BUFFD0 U615 ( .I(n627), .Z(n626) );
  BUFFD0 U616 ( .I(n628), .Z(n627) );
  BUFFD0 U617 ( .I(n629), .Z(n628) );
  BUFFD0 U618 ( .I(n630), .Z(n629) );
  BUFFD0 U619 ( .I(n631), .Z(n630) );
  BUFFD0 U620 ( .I(n632), .Z(n631) );
  BUFFD0 U621 ( .I(n633), .Z(n632) );
  BUFFD0 U622 ( .I(n634), .Z(n633) );
  BUFFD0 U623 ( .I(n635), .Z(n634) );
  BUFFD0 U624 ( .I(n636), .Z(n635) );
  BUFFD0 U625 ( .I(n637), .Z(n636) );
  BUFFD0 U626 ( .I(n638), .Z(n637) );
  BUFFD0 U627 ( .I(n639), .Z(n638) );
  BUFFD0 U628 ( .I(n640), .Z(n639) );
  BUFFD0 U629 ( .I(n641), .Z(n640) );
  BUFFD0 U630 ( .I(n642), .Z(n641) );
  BUFFD0 U631 ( .I(n643), .Z(n642) );
  BUFFD0 U632 ( .I(n644), .Z(n643) );
  BUFFD0 U633 ( .I(n645), .Z(n644) );
  BUFFD0 U634 ( .I(n646), .Z(n645) );
  BUFFD0 U635 ( .I(n647), .Z(n646) );
  BUFFD0 U636 ( .I(n648), .Z(n647) );
  BUFFD0 U637 ( .I(n649), .Z(n648) );
  BUFFD0 U638 ( .I(n650), .Z(n649) );
  BUFFD0 U639 ( .I(n651), .Z(n650) );
  BUFFD0 U640 ( .I(n652), .Z(n651) );
  BUFFD0 U641 ( .I(n653), .Z(n652) );
  BUFFD0 U642 ( .I(n654), .Z(n653) );
  BUFFD0 U643 ( .I(n655), .Z(n654) );
  BUFFD0 U644 ( .I(n656), .Z(n655) );
  BUFFD0 U645 ( .I(n657), .Z(n656) );
  BUFFD0 U646 ( .I(n658), .Z(n657) );
  BUFFD0 U647 ( .I(n659), .Z(n658) );
  BUFFD0 U648 ( .I(n660), .Z(n659) );
  BUFFD0 U649 ( .I(n661), .Z(n660) );
  BUFFD0 U650 ( .I(n662), .Z(n661) );
  BUFFD0 U651 ( .I(n663), .Z(n662) );
  BUFFD0 U652 ( .I(n664), .Z(n663) );
  BUFFD0 U653 ( .I(n665), .Z(n664) );
  BUFFD0 U654 ( .I(n666), .Z(n665) );
  BUFFD0 U655 ( .I(n667), .Z(n666) );
  BUFFD0 U656 ( .I(n668), .Z(n667) );
  BUFFD0 U657 ( .I(n4687), .Z(n668) );
  BUFFD0 U658 ( .I(n4683), .Z(n669) );
  BUFFD0 U659 ( .I(n671), .Z(n670) );
  BUFFD0 U660 ( .I(n672), .Z(n671) );
  BUFFD0 U661 ( .I(n673), .Z(n672) );
  BUFFD0 U662 ( .I(n674), .Z(n673) );
  BUFFD0 U663 ( .I(n675), .Z(n674) );
  BUFFD0 U664 ( .I(n676), .Z(n675) );
  BUFFD0 U665 ( .I(n677), .Z(n676) );
  BUFFD0 U666 ( .I(n678), .Z(n677) );
  BUFFD0 U667 ( .I(n679), .Z(n678) );
  BUFFD0 U668 ( .I(n680), .Z(n679) );
  BUFFD0 U669 ( .I(n681), .Z(n680) );
  BUFFD0 U670 ( .I(n682), .Z(n681) );
  BUFFD0 U671 ( .I(n683), .Z(n682) );
  BUFFD0 U672 ( .I(n684), .Z(n683) );
  BUFFD0 U673 ( .I(n685), .Z(n684) );
  BUFFD0 U674 ( .I(n686), .Z(n685) );
  BUFFD0 U675 ( .I(n687), .Z(n686) );
  BUFFD0 U676 ( .I(n688), .Z(n687) );
  BUFFD0 U677 ( .I(n689), .Z(n688) );
  BUFFD0 U678 ( .I(n690), .Z(n689) );
  BUFFD0 U679 ( .I(n691), .Z(n690) );
  BUFFD0 U680 ( .I(n692), .Z(n691) );
  BUFFD0 U681 ( .I(n693), .Z(n692) );
  BUFFD0 U682 ( .I(n694), .Z(n693) );
  BUFFD0 U683 ( .I(n695), .Z(n694) );
  BUFFD0 U684 ( .I(n696), .Z(n695) );
  BUFFD0 U685 ( .I(n697), .Z(n696) );
  BUFFD0 U686 ( .I(n698), .Z(n697) );
  BUFFD0 U687 ( .I(n699), .Z(n698) );
  BUFFD0 U688 ( .I(n700), .Z(n699) );
  BUFFD0 U689 ( .I(n701), .Z(n700) );
  BUFFD0 U690 ( .I(n702), .Z(n701) );
  BUFFD0 U691 ( .I(n703), .Z(n702) );
  BUFFD0 U692 ( .I(n704), .Z(n703) );
  BUFFD0 U693 ( .I(n705), .Z(n704) );
  BUFFD0 U694 ( .I(n706), .Z(n705) );
  BUFFD0 U695 ( .I(n707), .Z(n706) );
  BUFFD0 U696 ( .I(n708), .Z(n707) );
  BUFFD0 U697 ( .I(n709), .Z(n708) );
  BUFFD0 U698 ( .I(n710), .Z(n709) );
  BUFFD0 U699 ( .I(n711), .Z(n710) );
  BUFFD0 U700 ( .I(n712), .Z(n711) );
  BUFFD0 U701 ( .I(n713), .Z(n712) );
  BUFFD0 U702 ( .I(n714), .Z(n713) );
  BUFFD0 U703 ( .I(n715), .Z(n714) );
  BUFFD0 U704 ( .I(n716), .Z(n715) );
  BUFFD0 U705 ( .I(n717), .Z(n716) );
  BUFFD0 U706 ( .I(n718), .Z(n717) );
  BUFFD0 U707 ( .I(n719), .Z(n718) );
  BUFFD0 U708 ( .I(n720), .Z(n719) );
  BUFFD0 U709 ( .I(n721), .Z(n720) );
  BUFFD0 U710 ( .I(n722), .Z(n721) );
  BUFFD0 U711 ( .I(n4684), .Z(n722) );
  BUFFD0 U712 ( .I(n724), .Z(n723) );
  BUFFD0 U713 ( .I(n4680), .Z(n724) );
  BUFFD0 U714 ( .I(n726), .Z(n725) );
  BUFFD0 U715 ( .I(n727), .Z(n726) );
  BUFFD0 U716 ( .I(n728), .Z(n727) );
  BUFFD0 U717 ( .I(n729), .Z(n728) );
  BUFFD0 U718 ( .I(n730), .Z(n729) );
  BUFFD0 U719 ( .I(n731), .Z(n730) );
  BUFFD0 U720 ( .I(n732), .Z(n731) );
  BUFFD0 U721 ( .I(n733), .Z(n732) );
  BUFFD0 U722 ( .I(n734), .Z(n733) );
  BUFFD0 U723 ( .I(n735), .Z(n734) );
  BUFFD0 U724 ( .I(n736), .Z(n735) );
  BUFFD0 U725 ( .I(n737), .Z(n736) );
  BUFFD0 U726 ( .I(n738), .Z(n737) );
  BUFFD0 U727 ( .I(n739), .Z(n738) );
  BUFFD0 U728 ( .I(n740), .Z(n739) );
  BUFFD0 U729 ( .I(n741), .Z(n740) );
  BUFFD0 U730 ( .I(n742), .Z(n741) );
  BUFFD0 U731 ( .I(n743), .Z(n742) );
  BUFFD0 U732 ( .I(n744), .Z(n743) );
  BUFFD0 U733 ( .I(n745), .Z(n744) );
  BUFFD0 U734 ( .I(n746), .Z(n745) );
  BUFFD0 U735 ( .I(n747), .Z(n746) );
  BUFFD0 U736 ( .I(n748), .Z(n747) );
  BUFFD0 U737 ( .I(n749), .Z(n748) );
  BUFFD0 U738 ( .I(n750), .Z(n749) );
  BUFFD0 U739 ( .I(n751), .Z(n750) );
  BUFFD0 U740 ( .I(n752), .Z(n751) );
  BUFFD0 U741 ( .I(n753), .Z(n752) );
  BUFFD0 U742 ( .I(n754), .Z(n753) );
  BUFFD0 U743 ( .I(n755), .Z(n754) );
  BUFFD0 U744 ( .I(n756), .Z(n755) );
  BUFFD0 U745 ( .I(n757), .Z(n756) );
  BUFFD0 U746 ( .I(n758), .Z(n757) );
  BUFFD0 U747 ( .I(n759), .Z(n758) );
  BUFFD0 U748 ( .I(n760), .Z(n759) );
  BUFFD0 U749 ( .I(n761), .Z(n760) );
  BUFFD0 U750 ( .I(n762), .Z(n761) );
  BUFFD0 U751 ( .I(n763), .Z(n762) );
  BUFFD0 U752 ( .I(n764), .Z(n763) );
  BUFFD0 U753 ( .I(n765), .Z(n764) );
  BUFFD0 U754 ( .I(n766), .Z(n765) );
  BUFFD0 U755 ( .I(n767), .Z(n766) );
  BUFFD0 U756 ( .I(n768), .Z(n767) );
  BUFFD0 U757 ( .I(n769), .Z(n768) );
  BUFFD0 U758 ( .I(n770), .Z(n769) );
  BUFFD0 U759 ( .I(n771), .Z(n770) );
  BUFFD0 U760 ( .I(n772), .Z(n771) );
  BUFFD0 U761 ( .I(n773), .Z(n772) );
  BUFFD0 U762 ( .I(n774), .Z(n773) );
  BUFFD0 U763 ( .I(n4681), .Z(n774) );
  BUFFD0 U764 ( .I(n776), .Z(n775) );
  BUFFD0 U765 ( .I(n4678), .Z(n776) );
  BUFFD0 U766 ( .I(n778), .Z(n777) );
  BUFFD0 U767 ( .I(n779), .Z(n778) );
  BUFFD0 U768 ( .I(n780), .Z(n779) );
  BUFFD0 U769 ( .I(n781), .Z(n780) );
  BUFFD0 U770 ( .I(n782), .Z(n781) );
  BUFFD0 U771 ( .I(n783), .Z(n782) );
  BUFFD0 U772 ( .I(n784), .Z(n783) );
  BUFFD0 U773 ( .I(n785), .Z(n784) );
  BUFFD0 U774 ( .I(n786), .Z(n785) );
  BUFFD0 U775 ( .I(n787), .Z(n786) );
  BUFFD0 U776 ( .I(n788), .Z(n787) );
  BUFFD0 U777 ( .I(n789), .Z(n788) );
  BUFFD0 U778 ( .I(n790), .Z(n789) );
  BUFFD0 U779 ( .I(n791), .Z(n790) );
  BUFFD0 U780 ( .I(n792), .Z(n791) );
  BUFFD0 U781 ( .I(n793), .Z(n792) );
  BUFFD0 U782 ( .I(n794), .Z(n793) );
  BUFFD0 U783 ( .I(n795), .Z(n794) );
  BUFFD0 U784 ( .I(n796), .Z(n795) );
  BUFFD0 U785 ( .I(n797), .Z(n796) );
  BUFFD0 U786 ( .I(n798), .Z(n797) );
  BUFFD0 U787 ( .I(n799), .Z(n798) );
  BUFFD0 U788 ( .I(n800), .Z(n799) );
  BUFFD0 U789 ( .I(n801), .Z(n800) );
  BUFFD0 U790 ( .I(n802), .Z(n801) );
  BUFFD0 U791 ( .I(n803), .Z(n802) );
  BUFFD0 U792 ( .I(n804), .Z(n803) );
  BUFFD0 U793 ( .I(n805), .Z(n804) );
  BUFFD0 U794 ( .I(n806), .Z(n805) );
  BUFFD0 U795 ( .I(n807), .Z(n806) );
  BUFFD0 U796 ( .I(n808), .Z(n807) );
  BUFFD0 U797 ( .I(n809), .Z(n808) );
  BUFFD0 U798 ( .I(n810), .Z(n809) );
  BUFFD0 U799 ( .I(n811), .Z(n810) );
  BUFFD0 U800 ( .I(n812), .Z(n811) );
  BUFFD0 U801 ( .I(n813), .Z(n812) );
  BUFFD0 U802 ( .I(n814), .Z(n813) );
  BUFFD0 U803 ( .I(n815), .Z(n814) );
  BUFFD0 U804 ( .I(n816), .Z(n815) );
  BUFFD0 U805 ( .I(n817), .Z(n816) );
  BUFFD0 U806 ( .I(n818), .Z(n817) );
  BUFFD0 U807 ( .I(n819), .Z(n818) );
  BUFFD0 U808 ( .I(n820), .Z(n819) );
  BUFFD0 U809 ( .I(n821), .Z(n820) );
  BUFFD0 U810 ( .I(n822), .Z(n821) );
  BUFFD0 U811 ( .I(n823), .Z(n822) );
  BUFFD0 U812 ( .I(n824), .Z(n823) );
  BUFFD0 U813 ( .I(n825), .Z(n824) );
  BUFFD0 U814 ( .I(n826), .Z(n825) );
  BUFFD0 U815 ( .I(n4679), .Z(n826) );
  BUFFD0 U816 ( .I(n4676), .Z(n827) );
  BUFFD0 U817 ( .I(n829), .Z(n828) );
  BUFFD0 U818 ( .I(n830), .Z(n829) );
  BUFFD0 U819 ( .I(n831), .Z(n830) );
  BUFFD0 U820 ( .I(n832), .Z(n831) );
  BUFFD0 U821 ( .I(n833), .Z(n832) );
  BUFFD0 U822 ( .I(n834), .Z(n833) );
  BUFFD0 U823 ( .I(n835), .Z(n834) );
  BUFFD0 U824 ( .I(n836), .Z(n835) );
  BUFFD0 U825 ( .I(n837), .Z(n836) );
  BUFFD0 U826 ( .I(n838), .Z(n837) );
  BUFFD0 U827 ( .I(n839), .Z(n838) );
  BUFFD0 U828 ( .I(n840), .Z(n839) );
  BUFFD0 U829 ( .I(n841), .Z(n840) );
  BUFFD0 U830 ( .I(n842), .Z(n841) );
  BUFFD0 U831 ( .I(n843), .Z(n842) );
  BUFFD0 U832 ( .I(n844), .Z(n843) );
  BUFFD0 U833 ( .I(n845), .Z(n844) );
  BUFFD0 U834 ( .I(n846), .Z(n845) );
  BUFFD0 U835 ( .I(n847), .Z(n846) );
  BUFFD0 U836 ( .I(n848), .Z(n847) );
  BUFFD0 U837 ( .I(n849), .Z(n848) );
  BUFFD0 U838 ( .I(n850), .Z(n849) );
  BUFFD0 U839 ( .I(n851), .Z(n850) );
  BUFFD0 U840 ( .I(n852), .Z(n851) );
  BUFFD0 U841 ( .I(n853), .Z(n852) );
  BUFFD0 U842 ( .I(n854), .Z(n853) );
  BUFFD0 U843 ( .I(n855), .Z(n854) );
  BUFFD0 U844 ( .I(n856), .Z(n855) );
  BUFFD0 U845 ( .I(n857), .Z(n856) );
  BUFFD0 U846 ( .I(n858), .Z(n857) );
  BUFFD0 U847 ( .I(n859), .Z(n858) );
  BUFFD0 U848 ( .I(n860), .Z(n859) );
  BUFFD0 U849 ( .I(n861), .Z(n860) );
  BUFFD0 U850 ( .I(n862), .Z(n861) );
  BUFFD0 U851 ( .I(n863), .Z(n862) );
  BUFFD0 U852 ( .I(n864), .Z(n863) );
  BUFFD0 U853 ( .I(n865), .Z(n864) );
  BUFFD0 U854 ( .I(n866), .Z(n865) );
  BUFFD0 U855 ( .I(n867), .Z(n866) );
  BUFFD0 U856 ( .I(n868), .Z(n867) );
  BUFFD0 U857 ( .I(n869), .Z(n868) );
  BUFFD0 U858 ( .I(n870), .Z(n869) );
  BUFFD0 U859 ( .I(n871), .Z(n870) );
  BUFFD0 U860 ( .I(n872), .Z(n871) );
  BUFFD0 U861 ( .I(n873), .Z(n872) );
  BUFFD0 U862 ( .I(n874), .Z(n873) );
  BUFFD0 U863 ( .I(n875), .Z(n874) );
  BUFFD0 U864 ( .I(n876), .Z(n875) );
  BUFFD0 U865 ( .I(n877), .Z(n876) );
  BUFFD0 U866 ( .I(n878), .Z(n877) );
  BUFFD0 U867 ( .I(n879), .Z(n878) );
  BUFFD0 U868 ( .I(n880), .Z(n879) );
  BUFFD0 U869 ( .I(n4677), .Z(n880) );
  BUFFD0 U870 ( .I(n882), .Z(n881) );
  BUFFD0 U871 ( .I(n883), .Z(n882) );
  BUFFD0 U872 ( .I(n884), .Z(n883) );
  BUFFD0 U873 ( .I(n885), .Z(n884) );
  BUFFD0 U874 ( .I(n886), .Z(n885) );
  BUFFD0 U875 ( .I(n887), .Z(n886) );
  BUFFD0 U876 ( .I(n888), .Z(n887) );
  BUFFD0 U877 ( .I(n889), .Z(n888) );
  BUFFD0 U878 ( .I(n890), .Z(n889) );
  BUFFD0 U879 ( .I(n891), .Z(n890) );
  BUFFD0 U880 ( .I(n892), .Z(n891) );
  BUFFD0 U881 ( .I(n893), .Z(n892) );
  BUFFD0 U882 ( .I(n894), .Z(n893) );
  BUFFD0 U883 ( .I(n895), .Z(n894) );
  BUFFD0 U884 ( .I(n896), .Z(n895) );
  BUFFD0 U885 ( .I(n897), .Z(n896) );
  BUFFD0 U886 ( .I(n898), .Z(n897) );
  BUFFD0 U887 ( .I(n899), .Z(n898) );
  BUFFD0 U888 ( .I(n900), .Z(n899) );
  BUFFD0 U889 ( .I(n901), .Z(n900) );
  BUFFD0 U890 ( .I(n902), .Z(n901) );
  BUFFD0 U891 ( .I(n903), .Z(n902) );
  BUFFD0 U892 ( .I(n904), .Z(n903) );
  BUFFD0 U893 ( .I(n905), .Z(n904) );
  BUFFD0 U894 ( .I(n906), .Z(n905) );
  BUFFD0 U895 ( .I(n907), .Z(n906) );
  BUFFD0 U896 ( .I(n908), .Z(n907) );
  BUFFD0 U897 ( .I(n909), .Z(n908) );
  BUFFD0 U898 ( .I(n910), .Z(n909) );
  BUFFD0 U899 ( .I(n911), .Z(n910) );
  BUFFD0 U900 ( .I(n912), .Z(n911) );
  BUFFD0 U901 ( .I(n913), .Z(n912) );
  BUFFD0 U902 ( .I(n914), .Z(n913) );
  BUFFD0 U903 ( .I(n915), .Z(n914) );
  BUFFD0 U904 ( .I(n916), .Z(n915) );
  BUFFD0 U905 ( .I(n917), .Z(n916) );
  BUFFD0 U906 ( .I(n918), .Z(n917) );
  BUFFD0 U907 ( .I(n919), .Z(n918) );
  BUFFD0 U908 ( .I(n920), .Z(n919) );
  BUFFD0 U909 ( .I(n921), .Z(n920) );
  BUFFD0 U910 ( .I(n922), .Z(n921) );
  BUFFD0 U911 ( .I(n923), .Z(n922) );
  BUFFD0 U912 ( .I(n924), .Z(n923) );
  BUFFD0 U913 ( .I(n925), .Z(n924) );
  BUFFD0 U914 ( .I(n926), .Z(n925) );
  BUFFD0 U915 ( .I(n927), .Z(n926) );
  BUFFD0 U916 ( .I(n928), .Z(n927) );
  BUFFD0 U917 ( .I(n929), .Z(n928) );
  BUFFD0 U918 ( .I(n930), .Z(n929) );
  BUFFD0 U919 ( .I(n4674), .Z(n930) );
  BUFFD0 U920 ( .I(n933), .Z(n932) );
  BUFFD0 U921 ( .I(n934), .Z(n933) );
  BUFFD0 U922 ( .I(n935), .Z(n934) );
  BUFFD0 U923 ( .I(n936), .Z(n935) );
  BUFFD0 U924 ( .I(n937), .Z(n936) );
  BUFFD0 U925 ( .I(n938), .Z(n937) );
  BUFFD0 U926 ( .I(n939), .Z(n938) );
  BUFFD0 U927 ( .I(n940), .Z(n939) );
  BUFFD0 U928 ( .I(n941), .Z(n940) );
  BUFFD0 U929 ( .I(n942), .Z(n941) );
  BUFFD0 U930 ( .I(n943), .Z(n942) );
  BUFFD0 U931 ( .I(n944), .Z(n943) );
  BUFFD0 U932 ( .I(n945), .Z(n944) );
  BUFFD0 U933 ( .I(n946), .Z(n945) );
  BUFFD0 U934 ( .I(n947), .Z(n946) );
  BUFFD0 U935 ( .I(n948), .Z(n947) );
  BUFFD0 U936 ( .I(n949), .Z(n948) );
  BUFFD0 U937 ( .I(n950), .Z(n949) );
  BUFFD0 U938 ( .I(n951), .Z(n950) );
  BUFFD0 U939 ( .I(n952), .Z(n951) );
  BUFFD0 U940 ( .I(n953), .Z(n952) );
  BUFFD0 U941 ( .I(n954), .Z(n953) );
  BUFFD0 U942 ( .I(n955), .Z(n954) );
  BUFFD0 U943 ( .I(n956), .Z(n955) );
  BUFFD0 U944 ( .I(n957), .Z(n956) );
  BUFFD0 U945 ( .I(n958), .Z(n957) );
  BUFFD0 U946 ( .I(n959), .Z(n958) );
  BUFFD0 U947 ( .I(n960), .Z(n959) );
  BUFFD0 U948 ( .I(n961), .Z(n960) );
  BUFFD0 U949 ( .I(n962), .Z(n961) );
  BUFFD0 U950 ( .I(n963), .Z(n962) );
  BUFFD0 U951 ( .I(n964), .Z(n963) );
  BUFFD0 U952 ( .I(n965), .Z(n964) );
  BUFFD0 U953 ( .I(n966), .Z(n965) );
  BUFFD0 U954 ( .I(n967), .Z(n966) );
  BUFFD0 U955 ( .I(n968), .Z(n967) );
  BUFFD0 U956 ( .I(n969), .Z(n968) );
  BUFFD0 U957 ( .I(n970), .Z(n969) );
  BUFFD0 U958 ( .I(n971), .Z(n970) );
  BUFFD0 U959 ( .I(n972), .Z(n971) );
  BUFFD0 U960 ( .I(n973), .Z(n972) );
  BUFFD0 U961 ( .I(n974), .Z(n973) );
  BUFFD0 U962 ( .I(n975), .Z(n974) );
  BUFFD0 U963 ( .I(n976), .Z(n975) );
  BUFFD0 U964 ( .I(n977), .Z(n976) );
  BUFFD0 U965 ( .I(n978), .Z(n977) );
  BUFFD0 U966 ( .I(n979), .Z(n978) );
  BUFFD0 U967 ( .I(n980), .Z(n979) );
  BUFFD0 U968 ( .I(n981), .Z(n980) );
  BUFFD0 U969 ( .I(n982), .Z(n981) );
  BUFFD0 U970 ( .I(n983), .Z(n982) );
  BUFFD0 U971 ( .I(n984), .Z(n983) );
  BUFFD0 U972 ( .I(n4672), .Z(n984) );
  BUFFD0 U973 ( .I(n987), .Z(n986) );
  BUFFD0 U974 ( .I(n988), .Z(n987) );
  BUFFD0 U975 ( .I(n989), .Z(n988) );
  BUFFD0 U976 ( .I(n990), .Z(n989) );
  BUFFD0 U977 ( .I(n991), .Z(n990) );
  BUFFD0 U978 ( .I(n992), .Z(n991) );
  BUFFD0 U979 ( .I(n993), .Z(n992) );
  BUFFD0 U980 ( .I(n994), .Z(n993) );
  BUFFD0 U981 ( .I(n995), .Z(n994) );
  BUFFD0 U982 ( .I(n996), .Z(n995) );
  BUFFD0 U983 ( .I(n997), .Z(n996) );
  BUFFD0 U984 ( .I(n998), .Z(n997) );
  BUFFD0 U985 ( .I(n999), .Z(n998) );
  BUFFD0 U986 ( .I(n1000), .Z(n999) );
  BUFFD0 U987 ( .I(n1001), .Z(n1000) );
  BUFFD0 U988 ( .I(n1002), .Z(n1001) );
  BUFFD0 U989 ( .I(n1003), .Z(n1002) );
  BUFFD0 U990 ( .I(n1004), .Z(n1003) );
  BUFFD0 U991 ( .I(n1005), .Z(n1004) );
  BUFFD0 U992 ( .I(n1006), .Z(n1005) );
  BUFFD0 U993 ( .I(n1007), .Z(n1006) );
  BUFFD0 U994 ( .I(n1008), .Z(n1007) );
  BUFFD0 U995 ( .I(n1009), .Z(n1008) );
  BUFFD0 U996 ( .I(n1010), .Z(n1009) );
  BUFFD0 U997 ( .I(n1011), .Z(n1010) );
  BUFFD0 U998 ( .I(n1012), .Z(n1011) );
  BUFFD0 U999 ( .I(n1013), .Z(n1012) );
  BUFFD0 U1000 ( .I(n1014), .Z(n1013) );
  BUFFD0 U1001 ( .I(n1015), .Z(n1014) );
  BUFFD0 U1002 ( .I(n1016), .Z(n1015) );
  BUFFD0 U1003 ( .I(n1017), .Z(n1016) );
  BUFFD0 U1004 ( .I(n1018), .Z(n1017) );
  BUFFD0 U1005 ( .I(n1019), .Z(n1018) );
  BUFFD0 U1006 ( .I(n1020), .Z(n1019) );
  BUFFD0 U1007 ( .I(n1021), .Z(n1020) );
  BUFFD0 U1008 ( .I(n1022), .Z(n1021) );
  BUFFD0 U1009 ( .I(n1023), .Z(n1022) );
  BUFFD0 U1010 ( .I(n1024), .Z(n1023) );
  BUFFD0 U1011 ( .I(n1025), .Z(n1024) );
  BUFFD0 U1012 ( .I(n1026), .Z(n1025) );
  BUFFD0 U1013 ( .I(n1027), .Z(n1026) );
  BUFFD0 U1014 ( .I(n1028), .Z(n1027) );
  BUFFD0 U1015 ( .I(n1029), .Z(n1028) );
  BUFFD0 U1016 ( .I(n1030), .Z(n1029) );
  BUFFD0 U1017 ( .I(n1031), .Z(n1030) );
  BUFFD0 U1018 ( .I(n1032), .Z(n1031) );
  BUFFD0 U1019 ( .I(n1033), .Z(n1032) );
  BUFFD0 U1020 ( .I(n1034), .Z(n1033) );
  BUFFD0 U1021 ( .I(n1035), .Z(n1034) );
  BUFFD0 U1022 ( .I(n1036), .Z(n1035) );
  BUFFD0 U1023 ( .I(n1037), .Z(n1036) );
  BUFFD0 U1024 ( .I(n1038), .Z(n1037) );
  BUFFD0 U1025 ( .I(n4669), .Z(n1038) );
  BUFFD0 U1026 ( .I(n4665), .Z(n1039) );
  BUFFD0 U1027 ( .I(n1041), .Z(n1040) );
  BUFFD0 U1028 ( .I(n1042), .Z(n1041) );
  BUFFD0 U1029 ( .I(n1043), .Z(n1042) );
  BUFFD0 U1030 ( .I(n1044), .Z(n1043) );
  BUFFD0 U1031 ( .I(n1045), .Z(n1044) );
  BUFFD0 U1032 ( .I(n1046), .Z(n1045) );
  BUFFD0 U1033 ( .I(n1047), .Z(n1046) );
  BUFFD0 U1034 ( .I(n1048), .Z(n1047) );
  BUFFD0 U1035 ( .I(n1049), .Z(n1048) );
  BUFFD0 U1036 ( .I(n1050), .Z(n1049) );
  BUFFD0 U1037 ( .I(n1051), .Z(n1050) );
  BUFFD0 U1038 ( .I(n1052), .Z(n1051) );
  BUFFD0 U1039 ( .I(n1053), .Z(n1052) );
  BUFFD0 U1040 ( .I(n1054), .Z(n1053) );
  BUFFD0 U1041 ( .I(n1055), .Z(n1054) );
  BUFFD0 U1042 ( .I(n1056), .Z(n1055) );
  BUFFD0 U1043 ( .I(n1057), .Z(n1056) );
  BUFFD0 U1044 ( .I(n1058), .Z(n1057) );
  BUFFD0 U1045 ( .I(n1059), .Z(n1058) );
  BUFFD0 U1046 ( .I(n1060), .Z(n1059) );
  BUFFD0 U1047 ( .I(n1061), .Z(n1060) );
  BUFFD0 U1048 ( .I(n1062), .Z(n1061) );
  BUFFD0 U1049 ( .I(n1063), .Z(n1062) );
  BUFFD0 U1050 ( .I(n1064), .Z(n1063) );
  BUFFD0 U1051 ( .I(n1065), .Z(n1064) );
  BUFFD0 U1052 ( .I(n1066), .Z(n1065) );
  BUFFD0 U1053 ( .I(n1067), .Z(n1066) );
  BUFFD0 U1054 ( .I(n1068), .Z(n1067) );
  BUFFD0 U1055 ( .I(n1069), .Z(n1068) );
  BUFFD0 U1056 ( .I(n1070), .Z(n1069) );
  BUFFD0 U1057 ( .I(n1071), .Z(n1070) );
  BUFFD0 U1058 ( .I(n1072), .Z(n1071) );
  BUFFD0 U1059 ( .I(n1073), .Z(n1072) );
  BUFFD0 U1060 ( .I(n1074), .Z(n1073) );
  BUFFD0 U1061 ( .I(n1075), .Z(n1074) );
  BUFFD0 U1062 ( .I(n1076), .Z(n1075) );
  BUFFD0 U1063 ( .I(n1077), .Z(n1076) );
  BUFFD0 U1064 ( .I(n1078), .Z(n1077) );
  BUFFD0 U1065 ( .I(n1079), .Z(n1078) );
  BUFFD0 U1066 ( .I(n1080), .Z(n1079) );
  BUFFD0 U1067 ( .I(n1081), .Z(n1080) );
  BUFFD0 U1068 ( .I(n1082), .Z(n1081) );
  BUFFD0 U1069 ( .I(n1083), .Z(n1082) );
  BUFFD0 U1070 ( .I(n1084), .Z(n1083) );
  BUFFD0 U1071 ( .I(n1085), .Z(n1084) );
  BUFFD0 U1072 ( .I(n1086), .Z(n1085) );
  BUFFD0 U1073 ( .I(n1087), .Z(n1086) );
  BUFFD0 U1074 ( .I(n1088), .Z(n1087) );
  BUFFD0 U1075 ( .I(n1089), .Z(n1088) );
  BUFFD0 U1076 ( .I(n1090), .Z(n1089) );
  BUFFD0 U1077 ( .I(n1091), .Z(n1090) );
  BUFFD0 U1078 ( .I(n1092), .Z(n1091) );
  BUFFD0 U1079 ( .I(n4666), .Z(n1092) );
  BUFFD0 U1080 ( .I(n1094), .Z(n1093) );
  BUFFD0 U1081 ( .I(n4662), .Z(n1094) );
  BUFFD0 U1082 ( .I(n1096), .Z(n1095) );
  BUFFD0 U1083 ( .I(n1097), .Z(n1096) );
  BUFFD0 U1084 ( .I(n1098), .Z(n1097) );
  BUFFD0 U1085 ( .I(n1099), .Z(n1098) );
  BUFFD0 U1086 ( .I(n1100), .Z(n1099) );
  BUFFD0 U1087 ( .I(n1101), .Z(n1100) );
  BUFFD0 U1088 ( .I(n1102), .Z(n1101) );
  BUFFD0 U1089 ( .I(n1103), .Z(n1102) );
  BUFFD0 U1090 ( .I(n1104), .Z(n1103) );
  BUFFD0 U1091 ( .I(n1105), .Z(n1104) );
  BUFFD0 U1092 ( .I(n1106), .Z(n1105) );
  BUFFD0 U1093 ( .I(n1107), .Z(n1106) );
  BUFFD0 U1094 ( .I(n1108), .Z(n1107) );
  BUFFD0 U1095 ( .I(n1109), .Z(n1108) );
  BUFFD0 U1096 ( .I(n1110), .Z(n1109) );
  BUFFD0 U1097 ( .I(n1111), .Z(n1110) );
  BUFFD0 U1098 ( .I(n1112), .Z(n1111) );
  BUFFD0 U1099 ( .I(n1113), .Z(n1112) );
  BUFFD0 U1100 ( .I(n1114), .Z(n1113) );
  BUFFD0 U1101 ( .I(n1115), .Z(n1114) );
  BUFFD0 U1102 ( .I(n1116), .Z(n1115) );
  BUFFD0 U1103 ( .I(n1117), .Z(n1116) );
  BUFFD0 U1104 ( .I(n1118), .Z(n1117) );
  BUFFD0 U1105 ( .I(n1119), .Z(n1118) );
  BUFFD0 U1106 ( .I(n1120), .Z(n1119) );
  BUFFD0 U1107 ( .I(n1121), .Z(n1120) );
  BUFFD0 U1108 ( .I(n1122), .Z(n1121) );
  BUFFD0 U1109 ( .I(n1123), .Z(n1122) );
  BUFFD0 U1110 ( .I(n1124), .Z(n1123) );
  BUFFD0 U1111 ( .I(n1125), .Z(n1124) );
  BUFFD0 U1112 ( .I(n1126), .Z(n1125) );
  BUFFD0 U1113 ( .I(n1127), .Z(n1126) );
  BUFFD0 U1114 ( .I(n1128), .Z(n1127) );
  BUFFD0 U1115 ( .I(n1129), .Z(n1128) );
  BUFFD0 U1116 ( .I(n1130), .Z(n1129) );
  BUFFD0 U1117 ( .I(n1131), .Z(n1130) );
  BUFFD0 U1118 ( .I(n1132), .Z(n1131) );
  BUFFD0 U1119 ( .I(n1133), .Z(n1132) );
  BUFFD0 U1120 ( .I(n1134), .Z(n1133) );
  BUFFD0 U1121 ( .I(n1135), .Z(n1134) );
  BUFFD0 U1122 ( .I(n1136), .Z(n1135) );
  BUFFD0 U1123 ( .I(n1137), .Z(n1136) );
  BUFFD0 U1124 ( .I(n1138), .Z(n1137) );
  BUFFD0 U1125 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1126 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1127 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1128 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1129 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1130 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1131 ( .I(n4663), .Z(n1144) );
  BUFFD0 U1132 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1133 ( .I(n4660), .Z(n1146) );
  BUFFD0 U1134 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1135 ( .I(n1149), .Z(n1148) );
  BUFFD0 U1136 ( .I(n1150), .Z(n1149) );
  BUFFD0 U1137 ( .I(n1151), .Z(n1150) );
  BUFFD0 U1138 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1139 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1140 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1141 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1142 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1143 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1144 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1145 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1146 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1147 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1148 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1149 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1150 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1151 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1152 ( .I(n1166), .Z(n1165) );
  BUFFD0 U1153 ( .I(n1167), .Z(n1166) );
  BUFFD0 U1154 ( .I(n1168), .Z(n1167) );
  BUFFD0 U1155 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1156 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1157 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1158 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1159 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1160 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1161 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1162 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1163 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1164 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1165 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1166 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1167 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1168 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1169 ( .I(n1183), .Z(n1182) );
  BUFFD0 U1170 ( .I(n1184), .Z(n1183) );
  BUFFD0 U1171 ( .I(n1185), .Z(n1184) );
  BUFFD0 U1172 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1173 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1174 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1175 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1176 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1177 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1178 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1179 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1180 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1181 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1182 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1183 ( .I(n4661), .Z(n1196) );
  BUFFD0 U1184 ( .I(n4658), .Z(n1197) );
  BUFFD0 U1185 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1186 ( .I(n1200), .Z(n1199) );
  BUFFD0 U1187 ( .I(n1201), .Z(n1200) );
  BUFFD0 U1188 ( .I(n1202), .Z(n1201) );
  BUFFD0 U1189 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1190 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1191 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1192 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1193 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1194 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1195 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1196 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1197 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1198 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1199 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1200 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1201 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1202 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1203 ( .I(n1217), .Z(n1216) );
  BUFFD0 U1204 ( .I(n1218), .Z(n1217) );
  BUFFD0 U1205 ( .I(n1219), .Z(n1218) );
  BUFFD0 U1206 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1207 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1208 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1209 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1210 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1211 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1212 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1213 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1214 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1215 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1216 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1217 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1218 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1219 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1220 ( .I(n1234), .Z(n1233) );
  BUFFD0 U1221 ( .I(n1235), .Z(n1234) );
  BUFFD0 U1222 ( .I(n1236), .Z(n1235) );
  BUFFD0 U1223 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1224 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1225 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1226 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1227 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1228 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1229 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1230 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1231 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1232 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1233 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1234 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1235 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1236 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1237 ( .I(n4659), .Z(n1250) );
  BUFFD0 U1238 ( .I(n1252), .Z(n1251) );
  BUFFD0 U1239 ( .I(n1253), .Z(n1252) );
  BUFFD0 U1240 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1241 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1242 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1243 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1244 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1245 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1246 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1247 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1248 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1249 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1250 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1251 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1252 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1253 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1254 ( .I(n1268), .Z(n1267) );
  BUFFD0 U1255 ( .I(n1269), .Z(n1268) );
  BUFFD0 U1256 ( .I(n1270), .Z(n1269) );
  BUFFD0 U1257 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1258 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1259 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1260 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1261 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1262 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1263 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1264 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1265 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1266 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1267 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1268 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1269 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1270 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1271 ( .I(n1285), .Z(n1284) );
  BUFFD0 U1272 ( .I(n1286), .Z(n1285) );
  BUFFD0 U1273 ( .I(n1287), .Z(n1286) );
  BUFFD0 U1274 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1275 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1276 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1277 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1278 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1279 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1280 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1281 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1282 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1283 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1284 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1285 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1286 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1287 ( .I(n4656), .Z(n1300) );
  BUFFD0 U1288 ( .I(n1303), .Z(n1302) );
  BUFFD0 U1289 ( .I(n1304), .Z(n1303) );
  BUFFD0 U1290 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1291 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1292 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1293 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1294 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1295 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1296 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1297 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1298 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1299 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1300 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1301 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1302 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1303 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1304 ( .I(n1319), .Z(n1318) );
  BUFFD0 U1305 ( .I(n1320), .Z(n1319) );
  BUFFD0 U1306 ( .I(n1321), .Z(n1320) );
  BUFFD0 U1307 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1308 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1309 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1310 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1311 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1312 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1313 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1314 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1315 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1316 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1317 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1318 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1319 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1320 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1321 ( .I(n1336), .Z(n1335) );
  BUFFD0 U1322 ( .I(n1337), .Z(n1336) );
  BUFFD0 U1323 ( .I(n1338), .Z(n1337) );
  BUFFD0 U1324 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1325 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1326 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1327 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1328 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1329 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1330 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1331 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1332 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1333 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1334 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1335 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1336 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1337 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1338 ( .I(n1353), .Z(n1352) );
  BUFFD0 U1339 ( .I(n1354), .Z(n1353) );
  BUFFD0 U1340 ( .I(n4654), .Z(n1354) );
  BUFFD0 U1341 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1342 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1343 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1344 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1345 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1346 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1347 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1348 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1349 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1350 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1351 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1352 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1353 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1354 ( .I(n1370), .Z(n1369) );
  BUFFD0 U1355 ( .I(n1371), .Z(n1370) );
  BUFFD0 U1356 ( .I(n1372), .Z(n1371) );
  BUFFD0 U1357 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1358 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1359 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1360 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1361 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1362 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1363 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1364 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1365 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1366 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1367 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1368 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1369 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1370 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1371 ( .I(n1387), .Z(n1386) );
  BUFFD0 U1372 ( .I(n1388), .Z(n1387) );
  BUFFD0 U1373 ( .I(n1389), .Z(n1388) );
  BUFFD0 U1374 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1375 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1376 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1377 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1378 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1379 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1380 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1381 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1382 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1383 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1384 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1385 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1386 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1387 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1388 ( .I(n1404), .Z(n1403) );
  BUFFD0 U1389 ( .I(n1405), .Z(n1404) );
  BUFFD0 U1390 ( .I(n1406), .Z(n1405) );
  BUFFD0 U1391 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1392 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1393 ( .I(n4651), .Z(n1408) );
  BUFFD0 U1394 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1395 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1396 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1397 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1398 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1399 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1400 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1401 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1402 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1403 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1404 ( .I(n1420), .Z(n1419) );
  BUFFD0 U1405 ( .I(n1421), .Z(n1420) );
  BUFFD0 U1406 ( .I(n1422), .Z(n1421) );
  BUFFD0 U1407 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1408 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1409 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1410 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1411 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1412 ( .I(n1429), .Z(n1427) );
  BUFFD0 U1413 ( .I(n4647), .Z(n1428) );
  BUFFD0 U1414 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1415 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1416 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1417 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1418 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1419 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1420 ( .I(n1436), .Z(n1435) );
  BUFFD0 U1421 ( .I(n1437), .Z(n1436) );
  BUFFD0 U1422 ( .I(n1438), .Z(n1437) );
  BUFFD0 U1423 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1424 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1425 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1426 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1427 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1428 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1429 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1430 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1431 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1432 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1433 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1434 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1435 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1436 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1437 ( .I(n1453), .Z(n1452) );
  BUFFD0 U1438 ( .I(n1454), .Z(n1453) );
  BUFFD0 U1439 ( .I(n1455), .Z(n1454) );
  BUFFD0 U1440 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1441 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1442 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1443 ( .I(n4648), .Z(n1458) );
  BUFFD0 U1444 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1445 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1446 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1447 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1448 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1449 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1450 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1451 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1452 ( .I(n1469), .Z(n1468) );
  BUFFD0 U1453 ( .I(n1470), .Z(n1469) );
  BUFFD0 U1454 ( .I(n1471), .Z(n1470) );
  BUFFD0 U1455 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1456 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1457 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1458 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1459 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1460 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1461 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1462 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1463 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1464 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1465 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1466 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1467 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1468 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1469 ( .I(n1486), .Z(n1485) );
  BUFFD0 U1470 ( .I(n1487), .Z(n1486) );
  BUFFD0 U1471 ( .I(n1488), .Z(n1487) );
  BUFFD0 U1472 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1473 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1474 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1475 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1476 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1477 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1478 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1479 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1480 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1481 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1482 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1483 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1484 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1485 ( .I(n1502), .Z(n1501) );
  BUFFD0 U1486 ( .I(n1503), .Z(n1502) );
  BUFFD0 U1487 ( .I(n1504), .Z(n1503) );
  BUFFD0 U1488 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1489 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1490 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1491 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1492 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1493 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1494 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1495 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1496 ( .I(n4646), .Z(n1512) );
  BUFFD0 U1497 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1498 ( .I(n1516), .Z(n1515) );
  BUFFD0 U1499 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1500 ( .I(n1518), .Z(n1517) );
  BUFFD0 U1501 ( .I(n1519), .Z(n1518) );
  BUFFD0 U1502 ( .I(n1520), .Z(n1519) );
  BUFFD0 U1503 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1504 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1505 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1506 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1507 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1508 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1509 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1510 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1511 ( .I(n1529), .Z(n1528) );
  BUFFD0 U1512 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1513 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1514 ( .I(n1533), .Z(n1531) );
  BUFFD0 U1515 ( .I(n4642), .Z(n1532) );
  BUFFD0 U1516 ( .I(n1534), .Z(n1533) );
  BUFFD0 U1517 ( .I(n1535), .Z(n1534) );
  BUFFD0 U1518 ( .I(n1536), .Z(n1535) );
  BUFFD0 U1519 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1520 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1521 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1522 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1523 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1524 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1525 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1526 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1527 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1528 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1529 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1530 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1531 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1532 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1533 ( .I(n1551), .Z(n1550) );
  BUFFD0 U1534 ( .I(n1552), .Z(n1551) );
  BUFFD0 U1535 ( .I(n1553), .Z(n1552) );
  BUFFD0 U1536 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1537 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1538 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1539 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1540 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1541 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1542 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1543 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1544 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1545 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1546 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1547 ( .I(n4643), .Z(n1564) );
  BUFFD0 U1548 ( .I(n4711), .Z(n1565) );
  BUFFD0 U1549 ( .I(n1567), .Z(n1566) );
  BUFFD0 U1550 ( .I(n1568), .Z(n1567) );
  BUFFD0 U1551 ( .I(n1569), .Z(n1568) );
  BUFFD0 U1552 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1553 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1554 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1555 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1556 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1557 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1558 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1559 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1560 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1561 ( .I(n1579), .Z(n1578) );
  BUFFD0 U1562 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1563 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1564 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1565 ( .I(n1583), .Z(n1582) );
  BUFFD0 U1566 ( .I(n1584), .Z(n1583) );
  BUFFD0 U1567 ( .I(n1585), .Z(n1584) );
  BUFFD0 U1568 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1569 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1570 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1571 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1572 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1573 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1574 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1575 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1576 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1577 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1578 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1579 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1580 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1581 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1582 ( .I(n1600), .Z(n1599) );
  BUFFD0 U1583 ( .I(n1601), .Z(n1600) );
  BUFFD0 U1584 ( .I(n1602), .Z(n1601) );
  BUFFD0 U1585 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1586 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1587 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1588 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1589 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1590 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1591 ( .I(n1609), .Z(n1608) );
  BUFFD0 U1592 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1593 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1594 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1595 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1596 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1597 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1598 ( .I(n1616), .Z(n1615) );
  BUFFD0 U1599 ( .I(n1617), .Z(n1616) );
  BUFFD0 U1600 ( .I(n1618), .Z(n1617) );
  BUFFD0 U1601 ( .I(n4712), .Z(n1618) );
  BUFFD0 U1602 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1603 ( .I(n4706), .Z(n1620) );
  BUFFD0 U1604 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1605 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1606 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1607 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1608 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1609 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1610 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1611 ( .I(n1629), .Z(n1628) );
  BUFFD0 U1612 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1613 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1614 ( .I(n1632), .Z(n1631) );
  BUFFD0 U1615 ( .I(n1633), .Z(n1632) );
  BUFFD0 U1616 ( .I(n1634), .Z(n1633) );
  BUFFD0 U1617 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1618 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1619 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1620 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1621 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1622 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1623 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1624 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1625 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1626 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1627 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1628 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1629 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1630 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1631 ( .I(n1649), .Z(n1648) );
  BUFFD0 U1632 ( .I(n1650), .Z(n1649) );
  BUFFD0 U1633 ( .I(n1651), .Z(n1650) );
  BUFFD0 U1634 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1635 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1636 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1637 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1638 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1639 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1640 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1641 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1642 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1643 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1644 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1645 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1646 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1647 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1648 ( .I(n1666), .Z(n1665) );
  BUFFD0 U1649 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1650 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1651 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1652 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1653 ( .I(n4707), .Z(n1670) );
  BUFFD0 U1654 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1655 ( .I(n4708), .Z(n1672) );
  BUFFD0 U1656 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1657 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1658 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1659 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1660 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1661 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1662 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1663 ( .I(n1681), .Z(n1680) );
  BUFFD0 U1664 ( .I(n1682), .Z(n1681) );
  BUFFD0 U1665 ( .I(n1683), .Z(n1682) );
  BUFFD0 U1666 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1667 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1668 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1669 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1670 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1671 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1672 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1673 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1674 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1675 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1676 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1677 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1678 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1679 ( .I(n1697), .Z(n1696) );
  BUFFD0 U1680 ( .I(n1698), .Z(n1697) );
  BUFFD0 U1681 ( .I(n1699), .Z(n1698) );
  BUFFD0 U1682 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1683 ( .I(n1701), .Z(n1700) );
  BUFFD0 U1684 ( .I(n1702), .Z(n1701) );
  BUFFD0 U1685 ( .I(n1703), .Z(n1702) );
  BUFFD0 U1686 ( .I(n1704), .Z(n1703) );
  BUFFD0 U1687 ( .I(n1705), .Z(n1704) );
  BUFFD0 U1688 ( .I(n1706), .Z(n1705) );
  BUFFD0 U1689 ( .I(n1707), .Z(n1706) );
  BUFFD0 U1690 ( .I(n1708), .Z(n1707) );
  BUFFD0 U1691 ( .I(n1709), .Z(n1708) );
  BUFFD0 U1692 ( .I(n1710), .Z(n1709) );
  BUFFD0 U1693 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1694 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1695 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1696 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1697 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1698 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1699 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1700 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1701 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1702 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1703 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1704 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1705 ( .I(n4709), .Z(n1722) );
  BUFFD0 U1706 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1707 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1708 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1709 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1710 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1711 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1712 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1713 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1714 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1715 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1716 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1717 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1718 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1719 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1720 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1721 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1722 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1723 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1724 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1725 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1726 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1727 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1728 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1729 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1730 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1731 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1732 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1733 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1734 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1735 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1736 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1737 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1738 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1739 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1740 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1741 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1742 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1743 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1744 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1745 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1746 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1747 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1748 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1749 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1750 ( .I(n1768), .Z(n1767) );
  BUFFD0 U1751 ( .I(n1769), .Z(n1768) );
  BUFFD0 U1752 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1753 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1754 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1755 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1756 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1757 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1758 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1759 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1760 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1761 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1762 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1763 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1764 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1765 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1766 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1767 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1768 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1769 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1770 ( .I(N51), .Z(n1787) );
  BUFFD0 U1771 ( .I(n4337), .Z(n1788) );
  BUFFD0 U1772 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1773 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1774 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1775 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1776 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1777 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1778 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1779 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1780 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1781 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1782 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1783 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1784 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1785 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1786 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1787 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1788 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1789 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1790 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1791 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1792 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1793 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1794 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1795 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1796 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1797 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1798 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1799 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1800 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1801 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1802 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1803 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1804 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1805 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1806 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1807 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1808 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1809 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1810 ( .I(n1828), .Z(n1827) );
  BUFFD0 U1811 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1812 ( .I(n1830), .Z(n1829) );
  BUFFD0 U1813 ( .I(n1831), .Z(n1830) );
  BUFFD0 U1814 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1815 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1816 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1817 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1818 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1819 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1820 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1821 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1822 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1823 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1824 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1825 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1826 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1827 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1828 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1829 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1830 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1831 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1832 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1833 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1834 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1835 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1836 ( .I(N52), .Z(n1853) );
  BUFFD0 U1837 ( .I(n4324), .Z(n1854) );
  BUFFD0 U1838 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1839 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1840 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1841 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1842 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1843 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1844 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1845 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1846 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1847 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1848 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1849 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1850 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1851 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1852 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1853 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1854 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1855 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1856 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1857 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1858 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1859 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1860 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1861 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1862 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1863 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1864 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1865 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1866 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1867 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1868 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1869 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1870 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1871 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1872 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1873 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1874 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1875 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1876 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1877 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1878 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1879 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1880 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1881 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1882 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1883 ( .I(n1901), .Z(n1900) );
  BUFFD0 U1884 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1885 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1886 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1887 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1888 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1889 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1890 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1891 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1892 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1893 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1894 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1895 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1896 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1897 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1898 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1899 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1900 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1901 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1902 ( .I(N53), .Z(n1919) );
  BUFFD0 U1903 ( .I(n4311), .Z(n1920) );
  BUFFD0 U1904 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1905 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1906 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1907 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1908 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1909 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1910 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1911 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1912 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1913 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1914 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1915 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1916 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1917 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1918 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1919 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1920 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1921 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1922 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1923 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1924 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1925 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1926 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1927 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1928 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1929 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1930 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1931 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1932 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1933 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1934 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1935 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1936 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1937 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1938 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1939 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1940 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1941 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1942 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1943 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1944 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1945 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1946 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1947 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1948 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1949 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1950 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1951 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1952 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1953 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1954 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1955 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1956 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1957 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1958 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1959 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1960 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1961 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1962 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1963 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1964 ( .I(n1982), .Z(n1981) );
  BUFFD0 U1965 ( .I(n1983), .Z(n1982) );
  BUFFD0 U1966 ( .I(n1984), .Z(n1983) );
  BUFFD0 U1967 ( .I(n1985), .Z(n1984) );
  BUFFD0 U1968 ( .I(N54), .Z(n1985) );
  BUFFD0 U1969 ( .I(n4298), .Z(n1986) );
  BUFFD0 U1970 ( .I(n1988), .Z(n1987) );
  BUFFD0 U1971 ( .I(n1989), .Z(n1988) );
  BUFFD0 U1972 ( .I(n1990), .Z(n1989) );
  BUFFD0 U1973 ( .I(n1991), .Z(n1990) );
  BUFFD0 U1974 ( .I(n1992), .Z(n1991) );
  BUFFD0 U1975 ( .I(n1993), .Z(n1992) );
  BUFFD0 U1976 ( .I(n1994), .Z(n1993) );
  BUFFD0 U1977 ( .I(n1995), .Z(n1994) );
  BUFFD0 U1978 ( .I(n1996), .Z(n1995) );
  BUFFD0 U1979 ( .I(n1997), .Z(n1996) );
  BUFFD0 U1980 ( .I(n1998), .Z(n1997) );
  BUFFD0 U1981 ( .I(n1999), .Z(n1998) );
  BUFFD0 U1982 ( .I(n2000), .Z(n1999) );
  BUFFD0 U1983 ( .I(n2001), .Z(n2000) );
  BUFFD0 U1984 ( .I(n2002), .Z(n2001) );
  BUFFD0 U1985 ( .I(n2003), .Z(n2002) );
  BUFFD0 U1986 ( .I(n2004), .Z(n2003) );
  BUFFD0 U1987 ( .I(n2005), .Z(n2004) );
  BUFFD0 U1988 ( .I(n2006), .Z(n2005) );
  BUFFD0 U1989 ( .I(n2007), .Z(n2006) );
  BUFFD0 U1990 ( .I(n2008), .Z(n2007) );
  BUFFD0 U1991 ( .I(n2009), .Z(n2008) );
  BUFFD0 U1992 ( .I(n2010), .Z(n2009) );
  BUFFD0 U1993 ( .I(n2011), .Z(n2010) );
  BUFFD0 U1994 ( .I(n2012), .Z(n2011) );
  BUFFD0 U1995 ( .I(n2013), .Z(n2012) );
  BUFFD0 U1996 ( .I(n2014), .Z(n2013) );
  BUFFD0 U1997 ( .I(n2015), .Z(n2014) );
  BUFFD0 U1998 ( .I(n2016), .Z(n2015) );
  BUFFD0 U1999 ( .I(n2017), .Z(n2016) );
  BUFFD0 U2000 ( .I(n2018), .Z(n2017) );
  BUFFD0 U2001 ( .I(n2019), .Z(n2018) );
  BUFFD0 U2002 ( .I(n2020), .Z(n2019) );
  BUFFD0 U2003 ( .I(n2021), .Z(n2020) );
  BUFFD0 U2004 ( .I(n2022), .Z(n2021) );
  BUFFD0 U2005 ( .I(n2023), .Z(n2022) );
  BUFFD0 U2006 ( .I(n2024), .Z(n2023) );
  BUFFD0 U2007 ( .I(n2025), .Z(n2024) );
  BUFFD0 U2008 ( .I(n2026), .Z(n2025) );
  BUFFD0 U2009 ( .I(n2027), .Z(n2026) );
  BUFFD0 U2010 ( .I(n2028), .Z(n2027) );
  BUFFD0 U2011 ( .I(n2029), .Z(n2028) );
  BUFFD0 U2012 ( .I(n2030), .Z(n2029) );
  BUFFD0 U2013 ( .I(n2031), .Z(n2030) );
  BUFFD0 U2014 ( .I(n2032), .Z(n2031) );
  BUFFD0 U2015 ( .I(n2033), .Z(n2032) );
  BUFFD0 U2016 ( .I(n2034), .Z(n2033) );
  BUFFD0 U2017 ( .I(n2035), .Z(n2034) );
  BUFFD0 U2018 ( .I(n2036), .Z(n2035) );
  BUFFD0 U2019 ( .I(n2037), .Z(n2036) );
  BUFFD0 U2020 ( .I(n2038), .Z(n2037) );
  BUFFD0 U2021 ( .I(n2039), .Z(n2038) );
  BUFFD0 U2022 ( .I(n2040), .Z(n2039) );
  BUFFD0 U2023 ( .I(n2041), .Z(n2040) );
  BUFFD0 U2024 ( .I(n2042), .Z(n2041) );
  BUFFD0 U2025 ( .I(n2043), .Z(n2042) );
  BUFFD0 U2026 ( .I(n2044), .Z(n2043) );
  BUFFD0 U2027 ( .I(n2045), .Z(n2044) );
  BUFFD0 U2028 ( .I(n2046), .Z(n2045) );
  BUFFD0 U2029 ( .I(n2047), .Z(n2046) );
  BUFFD0 U2030 ( .I(n2048), .Z(n2047) );
  BUFFD0 U2031 ( .I(n2049), .Z(n2048) );
  BUFFD0 U2032 ( .I(n2050), .Z(n2049) );
  BUFFD0 U2033 ( .I(n2051), .Z(n2050) );
  BUFFD0 U2034 ( .I(N55), .Z(n2051) );
  BUFFD0 U2035 ( .I(n4285), .Z(n2052) );
  BUFFD0 U2036 ( .I(n2054), .Z(n2053) );
  BUFFD0 U2037 ( .I(n2055), .Z(n2054) );
  BUFFD0 U2038 ( .I(n2056), .Z(n2055) );
  BUFFD0 U2039 ( .I(n2057), .Z(n2056) );
  BUFFD0 U2040 ( .I(n2058), .Z(n2057) );
  BUFFD0 U2041 ( .I(n2059), .Z(n2058) );
  BUFFD0 U2042 ( .I(n2060), .Z(n2059) );
  BUFFD0 U2043 ( .I(n2061), .Z(n2060) );
  BUFFD0 U2044 ( .I(n2062), .Z(n2061) );
  BUFFD0 U2045 ( .I(n2063), .Z(n2062) );
  BUFFD0 U2046 ( .I(n2064), .Z(n2063) );
  BUFFD0 U2047 ( .I(n2065), .Z(n2064) );
  BUFFD0 U2048 ( .I(n2066), .Z(n2065) );
  BUFFD0 U2049 ( .I(n2067), .Z(n2066) );
  BUFFD0 U2050 ( .I(n2068), .Z(n2067) );
  BUFFD0 U2051 ( .I(n2069), .Z(n2068) );
  BUFFD0 U2052 ( .I(n2070), .Z(n2069) );
  BUFFD0 U2053 ( .I(n2071), .Z(n2070) );
  BUFFD0 U2054 ( .I(n2072), .Z(n2071) );
  BUFFD0 U2055 ( .I(n2073), .Z(n2072) );
  BUFFD0 U2056 ( .I(n2074), .Z(n2073) );
  BUFFD0 U2057 ( .I(n2075), .Z(n2074) );
  BUFFD0 U2058 ( .I(n2076), .Z(n2075) );
  BUFFD0 U2059 ( .I(n2077), .Z(n2076) );
  BUFFD0 U2060 ( .I(n2078), .Z(n2077) );
  BUFFD0 U2061 ( .I(n2079), .Z(n2078) );
  BUFFD0 U2062 ( .I(n2080), .Z(n2079) );
  BUFFD0 U2063 ( .I(n2081), .Z(n2080) );
  BUFFD0 U2064 ( .I(n2082), .Z(n2081) );
  BUFFD0 U2065 ( .I(n2083), .Z(n2082) );
  BUFFD0 U2066 ( .I(n2084), .Z(n2083) );
  BUFFD0 U2067 ( .I(n2085), .Z(n2084) );
  BUFFD0 U2068 ( .I(n2086), .Z(n2085) );
  BUFFD0 U2069 ( .I(n2087), .Z(n2086) );
  BUFFD0 U2070 ( .I(n2088), .Z(n2087) );
  BUFFD0 U2071 ( .I(n2089), .Z(n2088) );
  BUFFD0 U2072 ( .I(n2090), .Z(n2089) );
  BUFFD0 U2073 ( .I(n2091), .Z(n2090) );
  BUFFD0 U2074 ( .I(n2092), .Z(n2091) );
  BUFFD0 U2075 ( .I(n2093), .Z(n2092) );
  BUFFD0 U2076 ( .I(n2094), .Z(n2093) );
  BUFFD0 U2077 ( .I(n2095), .Z(n2094) );
  BUFFD0 U2078 ( .I(n2096), .Z(n2095) );
  BUFFD0 U2079 ( .I(n2097), .Z(n2096) );
  BUFFD0 U2080 ( .I(n2098), .Z(n2097) );
  BUFFD0 U2081 ( .I(n2099), .Z(n2098) );
  BUFFD0 U2082 ( .I(n2100), .Z(n2099) );
  BUFFD0 U2083 ( .I(n2101), .Z(n2100) );
  BUFFD0 U2084 ( .I(n2102), .Z(n2101) );
  BUFFD0 U2085 ( .I(n2103), .Z(n2102) );
  BUFFD0 U2086 ( .I(n2104), .Z(n2103) );
  BUFFD0 U2087 ( .I(n2105), .Z(n2104) );
  BUFFD0 U2088 ( .I(n2106), .Z(n2105) );
  BUFFD0 U2089 ( .I(n2107), .Z(n2106) );
  BUFFD0 U2090 ( .I(n2108), .Z(n2107) );
  BUFFD0 U2091 ( .I(n2109), .Z(n2108) );
  BUFFD0 U2092 ( .I(n2110), .Z(n2109) );
  BUFFD0 U2093 ( .I(n2111), .Z(n2110) );
  BUFFD0 U2094 ( .I(n2112), .Z(n2111) );
  BUFFD0 U2095 ( .I(n2113), .Z(n2112) );
  BUFFD0 U2096 ( .I(n2114), .Z(n2113) );
  BUFFD0 U2097 ( .I(n2115), .Z(n2114) );
  BUFFD0 U2098 ( .I(n2116), .Z(n2115) );
  BUFFD0 U2099 ( .I(n2117), .Z(n2116) );
  BUFFD0 U2100 ( .I(N56), .Z(n2117) );
  BUFFD0 U2101 ( .I(n4272), .Z(n2118) );
  BUFFD0 U2102 ( .I(n2120), .Z(n2119) );
  BUFFD0 U2103 ( .I(n2121), .Z(n2120) );
  BUFFD0 U2104 ( .I(n2122), .Z(n2121) );
  BUFFD0 U2105 ( .I(n2123), .Z(n2122) );
  BUFFD0 U2106 ( .I(n2124), .Z(n2123) );
  BUFFD0 U2107 ( .I(n2125), .Z(n2124) );
  BUFFD0 U2108 ( .I(n2126), .Z(n2125) );
  BUFFD0 U2109 ( .I(n2127), .Z(n2126) );
  BUFFD0 U2110 ( .I(n2128), .Z(n2127) );
  BUFFD0 U2111 ( .I(n2129), .Z(n2128) );
  BUFFD0 U2112 ( .I(n2130), .Z(n2129) );
  BUFFD0 U2113 ( .I(n2131), .Z(n2130) );
  BUFFD0 U2114 ( .I(n2132), .Z(n2131) );
  BUFFD0 U2115 ( .I(n2133), .Z(n2132) );
  BUFFD0 U2116 ( .I(n2134), .Z(n2133) );
  BUFFD0 U2117 ( .I(n2135), .Z(n2134) );
  BUFFD0 U2118 ( .I(n2136), .Z(n2135) );
  BUFFD0 U2119 ( .I(n2137), .Z(n2136) );
  BUFFD0 U2120 ( .I(n2138), .Z(n2137) );
  BUFFD0 U2121 ( .I(n2139), .Z(n2138) );
  BUFFD0 U2122 ( .I(n2140), .Z(n2139) );
  BUFFD0 U2123 ( .I(n2141), .Z(n2140) );
  BUFFD0 U2124 ( .I(n2142), .Z(n2141) );
  BUFFD0 U2125 ( .I(n2143), .Z(n2142) );
  BUFFD0 U2126 ( .I(n2144), .Z(n2143) );
  BUFFD0 U2127 ( .I(n2145), .Z(n2144) );
  BUFFD0 U2128 ( .I(n2146), .Z(n2145) );
  BUFFD0 U2129 ( .I(n2147), .Z(n2146) );
  BUFFD0 U2130 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2131 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2132 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2133 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2134 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2135 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2136 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2137 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2138 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2139 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2140 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2141 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2142 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2143 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2144 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2145 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2146 ( .I(n2164), .Z(n2163) );
  BUFFD0 U2147 ( .I(n2165), .Z(n2164) );
  BUFFD0 U2148 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2149 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2150 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2151 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2152 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2153 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2154 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2155 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2156 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2157 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2158 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2159 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2160 ( .I(n2178), .Z(n2177) );
  BUFFD0 U2161 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2162 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2163 ( .I(n2181), .Z(n2180) );
  BUFFD0 U2164 ( .I(n2182), .Z(n2181) );
  BUFFD0 U2165 ( .I(n2183), .Z(n2182) );
  BUFFD0 U2166 ( .I(N57), .Z(n2183) );
  BUFFD0 U2167 ( .I(n4259), .Z(n2184) );
  BUFFD0 U2168 ( .I(n2186), .Z(n2185) );
  BUFFD0 U2169 ( .I(n2187), .Z(n2186) );
  BUFFD0 U2170 ( .I(n2188), .Z(n2187) );
  BUFFD0 U2171 ( .I(n2189), .Z(n2188) );
  BUFFD0 U2172 ( .I(n2190), .Z(n2189) );
  BUFFD0 U2173 ( .I(n2191), .Z(n2190) );
  BUFFD0 U2174 ( .I(n2192), .Z(n2191) );
  BUFFD0 U2175 ( .I(n2193), .Z(n2192) );
  BUFFD0 U2176 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2177 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2178 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2179 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2180 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2181 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2182 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2183 ( .I(n2201), .Z(n2200) );
  BUFFD0 U2184 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2185 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2186 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2187 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2188 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2189 ( .I(n2207), .Z(n2206) );
  BUFFD0 U2190 ( .I(n2208), .Z(n2207) );
  BUFFD0 U2191 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2192 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2193 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2194 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2195 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2196 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2197 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2198 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2199 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2200 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2201 ( .I(n2219), .Z(n2218) );
  BUFFD0 U2202 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2203 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2204 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2205 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2206 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2207 ( .I(n2225), .Z(n2224) );
  BUFFD0 U2208 ( .I(n2226), .Z(n2225) );
  BUFFD0 U2209 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2210 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2211 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2212 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2213 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2214 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2215 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2216 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2217 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2218 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2219 ( .I(n2237), .Z(n2236) );
  BUFFD0 U2220 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2221 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2222 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2223 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2224 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2225 ( .I(n2243), .Z(n2242) );
  BUFFD0 U2226 ( .I(n2244), .Z(n2243) );
  BUFFD0 U2227 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2228 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2229 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2230 ( .I(n2248), .Z(n2247) );
  BUFFD0 U2231 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2232 ( .I(N58), .Z(n2249) );
  BUFFD0 U2233 ( .I(n4246), .Z(n2250) );
  BUFFD0 U2234 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2235 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2236 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2237 ( .I(n2255), .Z(n2254) );
  BUFFD0 U2238 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2239 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2240 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2241 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2242 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2243 ( .I(n2261), .Z(n2260) );
  BUFFD0 U2244 ( .I(n2262), .Z(n2261) );
  BUFFD0 U2245 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2246 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2247 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2248 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2249 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2250 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2251 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2252 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2253 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2254 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2255 ( .I(n2273), .Z(n2272) );
  BUFFD0 U2256 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2257 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2258 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2259 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2260 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2261 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2262 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2263 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2264 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2265 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2266 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2267 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2268 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2269 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2270 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2271 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2272 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2273 ( .I(n2291), .Z(n2290) );
  BUFFD0 U2274 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2275 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2276 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2277 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2278 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2279 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2280 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2281 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2282 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2283 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2284 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2285 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2286 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2287 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2288 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2289 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2290 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2291 ( .I(n2309), .Z(n2308) );
  BUFFD0 U2292 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2293 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2294 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2295 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2296 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2297 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2298 ( .I(N59), .Z(n2315) );
  BUFFD0 U2299 ( .I(n4233), .Z(n2316) );
  BUFFD0 U2300 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2301 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2302 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2303 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2304 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2305 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2306 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2307 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2308 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2309 ( .I(n2327), .Z(n2326) );
  BUFFD0 U2310 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2311 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2312 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2313 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2314 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2315 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2316 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2317 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2318 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2319 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2320 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2321 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2322 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2323 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2324 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2325 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2326 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2327 ( .I(n2345), .Z(n2344) );
  BUFFD0 U2328 ( .I(n2346), .Z(n2345) );
  BUFFD0 U2329 ( .I(n2347), .Z(n2346) );
  BUFFD0 U2330 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2331 ( .I(n2349), .Z(n2348) );
  BUFFD0 U2332 ( .I(n2350), .Z(n2349) );
  BUFFD0 U2333 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2334 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2335 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2336 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2337 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2338 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2339 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2340 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2341 ( .I(n2359), .Z(n2358) );
  BUFFD0 U2342 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2343 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2344 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2345 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2346 ( .I(n2364), .Z(n2363) );
  BUFFD0 U2347 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2348 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2349 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2350 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2351 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2352 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2353 ( .I(n2371), .Z(n2370) );
  BUFFD0 U2354 ( .I(n2372), .Z(n2371) );
  BUFFD0 U2355 ( .I(n2373), .Z(n2372) );
  BUFFD0 U2356 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2357 ( .I(n2375), .Z(n2374) );
  BUFFD0 U2358 ( .I(n2376), .Z(n2375) );
  BUFFD0 U2359 ( .I(n2377), .Z(n2376) );
  BUFFD0 U2360 ( .I(n2378), .Z(n2377) );
  BUFFD0 U2361 ( .I(n2379), .Z(n2378) );
  BUFFD0 U2362 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2363 ( .I(n2381), .Z(n2380) );
  BUFFD0 U2364 ( .I(N60), .Z(n2381) );
  BUFFD0 U2365 ( .I(n4220), .Z(n2382) );
  BUFFD0 U2366 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2367 ( .I(n2385), .Z(n2384) );
  BUFFD0 U2368 ( .I(n2386), .Z(n2385) );
  BUFFD0 U2369 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2370 ( .I(n2388), .Z(n2387) );
  BUFFD0 U2371 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2372 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2373 ( .I(n2391), .Z(n2390) );
  BUFFD0 U2374 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2375 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2376 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2377 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2378 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2379 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2380 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2381 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2382 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2383 ( .I(n2401), .Z(n2400) );
  BUFFD0 U2384 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2385 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2386 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2387 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2388 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2389 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2390 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2391 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2392 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2393 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2394 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2395 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2396 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2397 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2398 ( .I(n2416), .Z(n2415) );
  BUFFD0 U2399 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2400 ( .I(n2418), .Z(n2417) );
  BUFFD0 U2401 ( .I(n2419), .Z(n2418) );
  BUFFD0 U2402 ( .I(n2420), .Z(n2419) );
  BUFFD0 U2403 ( .I(n2421), .Z(n2420) );
  BUFFD0 U2404 ( .I(n2422), .Z(n2421) );
  BUFFD0 U2405 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2406 ( .I(n2424), .Z(n2423) );
  BUFFD0 U2407 ( .I(n2425), .Z(n2424) );
  BUFFD0 U2408 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2409 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2410 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2411 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2412 ( .I(n2430), .Z(n2429) );
  BUFFD0 U2413 ( .I(n2431), .Z(n2430) );
  BUFFD0 U2414 ( .I(n2432), .Z(n2431) );
  BUFFD0 U2415 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2416 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2417 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2418 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2419 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2420 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2421 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2422 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2423 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2424 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2425 ( .I(n2443), .Z(n2442) );
  BUFFD0 U2426 ( .I(n2444), .Z(n2443) );
  BUFFD0 U2427 ( .I(n2445), .Z(n2444) );
  BUFFD0 U2428 ( .I(n2446), .Z(n2445) );
  BUFFD0 U2429 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2430 ( .I(N61), .Z(n2447) );
  BUFFD0 U2431 ( .I(n4207), .Z(n2448) );
  BUFFD0 U2432 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2433 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2434 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2435 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2436 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2437 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2438 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2439 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2440 ( .I(n2458), .Z(n2457) );
  BUFFD0 U2441 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2442 ( .I(n2460), .Z(n2459) );
  BUFFD0 U2443 ( .I(n2461), .Z(n2460) );
  BUFFD0 U2444 ( .I(n2462), .Z(n2461) );
  BUFFD0 U2445 ( .I(n2463), .Z(n2462) );
  BUFFD0 U2446 ( .I(n2464), .Z(n2463) );
  BUFFD0 U2447 ( .I(n2465), .Z(n2464) );
  BUFFD0 U2448 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2449 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2450 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2451 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2452 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2453 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2454 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2455 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2456 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2457 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2458 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2459 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2460 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2461 ( .I(n2479), .Z(n2478) );
  BUFFD0 U2462 ( .I(n2480), .Z(n2479) );
  BUFFD0 U2463 ( .I(n2481), .Z(n2480) );
  BUFFD0 U2464 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2465 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2466 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2467 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2468 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2469 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2470 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2471 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2472 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2473 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2474 ( .I(n2492), .Z(n2491) );
  BUFFD0 U2475 ( .I(n2493), .Z(n2492) );
  BUFFD0 U2476 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2477 ( .I(n2495), .Z(n2494) );
  BUFFD0 U2478 ( .I(n2496), .Z(n2495) );
  BUFFD0 U2479 ( .I(n2497), .Z(n2496) );
  BUFFD0 U2480 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2481 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2482 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2483 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2484 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2485 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2486 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2487 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2488 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2489 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2490 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2491 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2492 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2493 ( .I(n2511), .Z(n2510) );
  BUFFD0 U2494 ( .I(n2512), .Z(n2511) );
  BUFFD0 U2495 ( .I(n2513), .Z(n2512) );
  BUFFD0 U2496 ( .I(N62), .Z(n2513) );
  BUFFD0 U2497 ( .I(n4194), .Z(n2514) );
  BUFFD0 U2498 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2499 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2500 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2501 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2502 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2503 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2504 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2505 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2506 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2507 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2508 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2509 ( .I(n2527), .Z(n2526) );
  BUFFD0 U2510 ( .I(n2528), .Z(n2527) );
  BUFFD0 U2511 ( .I(n2529), .Z(n2528) );
  BUFFD0 U2512 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2513 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2514 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2515 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2516 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2517 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2518 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2519 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2520 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2521 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2522 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2523 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2524 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2525 ( .I(n2543), .Z(n2542) );
  BUFFD0 U2526 ( .I(n2544), .Z(n2543) );
  BUFFD0 U2527 ( .I(n2545), .Z(n2544) );
  BUFFD0 U2528 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2529 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2530 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2531 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2532 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2533 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2534 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2535 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2536 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2537 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2538 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2539 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2540 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2541 ( .I(n2559), .Z(n2558) );
  BUFFD0 U2542 ( .I(n2560), .Z(n2559) );
  BUFFD0 U2543 ( .I(n2561), .Z(n2560) );
  BUFFD0 U2544 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2545 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2546 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2547 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2548 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2549 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2550 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2551 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2552 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2553 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2554 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2555 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2556 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2557 ( .I(n2575), .Z(n2574) );
  BUFFD0 U2558 ( .I(n2576), .Z(n2575) );
  BUFFD0 U2559 ( .I(n2577), .Z(n2576) );
  BUFFD0 U2560 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2561 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2562 ( .I(N63), .Z(n2579) );
  BUFFD0 U2563 ( .I(n4181), .Z(n2580) );
  BUFFD0 U2564 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2565 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2566 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2567 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2568 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2569 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2570 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2571 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2572 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2573 ( .I(n2591), .Z(n2590) );
  BUFFD0 U2574 ( .I(n2592), .Z(n2591) );
  BUFFD0 U2575 ( .I(n2593), .Z(n2592) );
  BUFFD0 U2576 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2577 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2578 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2579 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2580 ( .I(n2598), .Z(n2597) );
  BUFFD0 U2581 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2582 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2583 ( .I(n2601), .Z(n2600) );
  BUFFD0 U2584 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2585 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2586 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2587 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2588 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2589 ( .I(n2607), .Z(n2606) );
  BUFFD0 U2590 ( .I(n2608), .Z(n2607) );
  BUFFD0 U2591 ( .I(n2609), .Z(n2608) );
  BUFFD0 U2592 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2593 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2594 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2595 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2596 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2597 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2598 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2599 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2600 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2601 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2602 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2603 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2604 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2605 ( .I(n2623), .Z(n2622) );
  BUFFD0 U2606 ( .I(n2624), .Z(n2623) );
  BUFFD0 U2607 ( .I(n2625), .Z(n2624) );
  BUFFD0 U2608 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2609 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2610 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2611 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2612 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2613 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2614 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2615 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2616 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2617 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2618 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2619 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2620 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2621 ( .I(n2639), .Z(n2638) );
  BUFFD0 U2622 ( .I(n2640), .Z(n2639) );
  BUFFD0 U2623 ( .I(n2641), .Z(n2640) );
  BUFFD0 U2624 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2625 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2626 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2627 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2628 ( .I(N64), .Z(n2645) );
  BUFFD0 U2629 ( .I(n4168), .Z(n2646) );
  BUFFD0 U2630 ( .I(n2648), .Z(n2647) );
  BUFFD0 U2631 ( .I(n2649), .Z(n2648) );
  BUFFD0 U2632 ( .I(n2650), .Z(n2649) );
  BUFFD0 U2633 ( .I(n2651), .Z(n2650) );
  BUFFD0 U2634 ( .I(n2652), .Z(n2651) );
  BUFFD0 U2635 ( .I(n2653), .Z(n2652) );
  BUFFD0 U2636 ( .I(n2654), .Z(n2653) );
  BUFFD0 U2637 ( .I(n2655), .Z(n2654) );
  BUFFD0 U2638 ( .I(n2656), .Z(n2655) );
  BUFFD0 U2639 ( .I(n2657), .Z(n2656) );
  BUFFD0 U2640 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2641 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2642 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2643 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2644 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2645 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2646 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2647 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2648 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2649 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2650 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2651 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2652 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2653 ( .I(n2671), .Z(n2670) );
  BUFFD0 U2654 ( .I(n2672), .Z(n2671) );
  BUFFD0 U2655 ( .I(n2673), .Z(n2672) );
  BUFFD0 U2656 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2657 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2658 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2659 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2660 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2661 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2662 ( .I(n2680), .Z(n2679) );
  BUFFD0 U2663 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2664 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2665 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2666 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2667 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2668 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2669 ( .I(n2687), .Z(n2686) );
  BUFFD0 U2670 ( .I(n2688), .Z(n2687) );
  BUFFD0 U2671 ( .I(n2689), .Z(n2688) );
  BUFFD0 U2672 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2673 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2674 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2675 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2676 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2677 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2678 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2679 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2680 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2681 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2682 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2683 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2684 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2685 ( .I(n2703), .Z(n2702) );
  BUFFD0 U2686 ( .I(n2704), .Z(n2703) );
  BUFFD0 U2687 ( .I(n2705), .Z(n2704) );
  BUFFD0 U2688 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2689 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2690 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2691 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2692 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2693 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2694 ( .I(N65), .Z(n2711) );
  BUFFD0 U2695 ( .I(n4155), .Z(n2712) );
  BUFFD0 U2696 ( .I(n2714), .Z(n2713) );
  BUFFD0 U2697 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2698 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2699 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2700 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2701 ( .I(n2719), .Z(n2718) );
  BUFFD0 U2702 ( .I(n2720), .Z(n2719) );
  BUFFD0 U2703 ( .I(n2721), .Z(n2720) );
  BUFFD0 U2704 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2705 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2706 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2707 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2708 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2709 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2710 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2711 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2712 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2713 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2714 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2715 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2716 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2717 ( .I(n2735), .Z(n2734) );
  BUFFD0 U2718 ( .I(n2736), .Z(n2735) );
  BUFFD0 U2719 ( .I(n2737), .Z(n2736) );
  BUFFD0 U2720 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2721 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2722 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2723 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2724 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2725 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2726 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2727 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2728 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2729 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2730 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2731 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2732 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2733 ( .I(n2751), .Z(n2750) );
  BUFFD0 U2734 ( .I(n2752), .Z(n2751) );
  BUFFD0 U2735 ( .I(n2753), .Z(n2752) );
  BUFFD0 U2736 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2737 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2738 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2739 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2740 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2741 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2742 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2743 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2744 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2745 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2746 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2747 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2748 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2749 ( .I(n2767), .Z(n2766) );
  BUFFD0 U2750 ( .I(n2768), .Z(n2767) );
  BUFFD0 U2751 ( .I(n2769), .Z(n2768) );
  BUFFD0 U2752 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2753 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2754 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2755 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2756 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2757 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2758 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2759 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2760 ( .I(N66), .Z(n2777) );
  BUFFD0 U2761 ( .I(n4142), .Z(n2778) );
  BUFFD0 U2762 ( .I(n2780), .Z(n2779) );
  BUFFD0 U2763 ( .I(n2781), .Z(n2780) );
  BUFFD0 U2764 ( .I(n2782), .Z(n2781) );
  BUFFD0 U2765 ( .I(n2783), .Z(n2782) );
  BUFFD0 U2766 ( .I(n2784), .Z(n2783) );
  BUFFD0 U2767 ( .I(n2785), .Z(n2784) );
  BUFFD0 U2768 ( .I(n2786), .Z(n2785) );
  BUFFD0 U2769 ( .I(n2787), .Z(n2786) );
  BUFFD0 U2770 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2771 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2772 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2773 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2774 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2775 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2776 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2777 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2778 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2779 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2780 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2781 ( .I(n2799), .Z(n2798) );
  BUFFD0 U2782 ( .I(n2800), .Z(n2799) );
  BUFFD0 U2783 ( .I(n2801), .Z(n2800) );
  BUFFD0 U2784 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2785 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2786 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2787 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2788 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2789 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2790 ( .I(n2808), .Z(n2807) );
  BUFFD0 U2791 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2792 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2793 ( .I(n2811), .Z(n2810) );
  BUFFD0 U2794 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2795 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2796 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2797 ( .I(n2815), .Z(n2814) );
  BUFFD0 U2798 ( .I(n2816), .Z(n2815) );
  BUFFD0 U2799 ( .I(n2817), .Z(n2816) );
  BUFFD0 U2800 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2801 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2802 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2803 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2804 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2805 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2806 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2807 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2808 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2809 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2810 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2811 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2812 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2813 ( .I(n2831), .Z(n2830) );
  BUFFD0 U2814 ( .I(n2832), .Z(n2831) );
  BUFFD0 U2815 ( .I(n2833), .Z(n2832) );
  BUFFD0 U2816 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2817 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2818 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2819 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2820 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2821 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2822 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2823 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2824 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2825 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2826 ( .I(N67), .Z(n2843) );
  BUFFD0 U2827 ( .I(n4129), .Z(n2844) );
  BUFFD0 U2828 ( .I(n2846), .Z(n2845) );
  BUFFD0 U2829 ( .I(n2847), .Z(n2846) );
  BUFFD0 U2830 ( .I(n2848), .Z(n2847) );
  BUFFD0 U2831 ( .I(n2849), .Z(n2848) );
  BUFFD0 U2832 ( .I(n2850), .Z(n2849) );
  BUFFD0 U2833 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2834 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2835 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2836 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2837 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2838 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2839 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2840 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2841 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2842 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2843 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2844 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2845 ( .I(n2863), .Z(n2862) );
  BUFFD0 U2846 ( .I(n2864), .Z(n2863) );
  BUFFD0 U2847 ( .I(n2865), .Z(n2864) );
  BUFFD0 U2848 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2849 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2850 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2851 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2852 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2853 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2854 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2855 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2856 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2857 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2858 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2859 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2860 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2861 ( .I(n2879), .Z(n2878) );
  BUFFD0 U2862 ( .I(n2880), .Z(n2879) );
  BUFFD0 U2863 ( .I(n2881), .Z(n2880) );
  BUFFD0 U2864 ( .I(n2882), .Z(n2881) );
  BUFFD0 U2865 ( .I(n2883), .Z(n2882) );
  BUFFD0 U2866 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2867 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2868 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2869 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2870 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2871 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2872 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2873 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2874 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2875 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2876 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2877 ( .I(n2895), .Z(n2894) );
  BUFFD0 U2878 ( .I(n2896), .Z(n2895) );
  BUFFD0 U2879 ( .I(n2897), .Z(n2896) );
  BUFFD0 U2880 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2881 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2882 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2883 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2884 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2885 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2886 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2887 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2888 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2889 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2890 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2891 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2892 ( .I(N68), .Z(n2909) );
  BUFFD0 U2893 ( .I(n4116), .Z(n2910) );
  BUFFD0 U2894 ( .I(n2912), .Z(n2911) );
  BUFFD0 U2895 ( .I(n2913), .Z(n2912) );
  BUFFD0 U2896 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2897 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2898 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2899 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2900 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2901 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2902 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2903 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2904 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2905 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2906 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2907 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2908 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2909 ( .I(n2927), .Z(n2926) );
  BUFFD0 U2910 ( .I(n2928), .Z(n2927) );
  BUFFD0 U2911 ( .I(n2929), .Z(n2928) );
  BUFFD0 U2912 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2913 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2914 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2915 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2916 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2917 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2918 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2919 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2920 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2921 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2922 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2923 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2924 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2925 ( .I(n2943), .Z(n2942) );
  BUFFD0 U2926 ( .I(n2944), .Z(n2943) );
  BUFFD0 U2927 ( .I(n2945), .Z(n2944) );
  BUFFD0 U2928 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2929 ( .I(n2947), .Z(n2946) );
  BUFFD0 U2930 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2931 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2932 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2933 ( .I(n2951), .Z(n2950) );
  BUFFD0 U2934 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2935 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2936 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2937 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2938 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2939 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2940 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2941 ( .I(n2959), .Z(n2958) );
  BUFFD0 U2942 ( .I(n2960), .Z(n2959) );
  BUFFD0 U2943 ( .I(n2961), .Z(n2960) );
  BUFFD0 U2944 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2945 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2946 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2947 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2948 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2949 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2950 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2951 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2952 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2953 ( .I(n2971), .Z(n2970) );
  BUFFD0 U2954 ( .I(n2972), .Z(n2971) );
  BUFFD0 U2955 ( .I(n2973), .Z(n2972) );
  BUFFD0 U2956 ( .I(n2974), .Z(n2973) );
  BUFFD0 U2957 ( .I(n2975), .Z(n2974) );
  BUFFD0 U2958 ( .I(N69), .Z(n2975) );
  BUFFD0 U2959 ( .I(n4103), .Z(n2976) );
  BUFFD0 U2960 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2961 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2962 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2963 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2964 ( .I(n2982), .Z(n2981) );
  BUFFD0 U2965 ( .I(n2983), .Z(n2982) );
  BUFFD0 U2966 ( .I(n2984), .Z(n2983) );
  BUFFD0 U2967 ( .I(n2985), .Z(n2984) );
  BUFFD0 U2968 ( .I(n2986), .Z(n2985) );
  BUFFD0 U2969 ( .I(n2987), .Z(n2986) );
  BUFFD0 U2970 ( .I(n2988), .Z(n2987) );
  BUFFD0 U2971 ( .I(n2989), .Z(n2988) );
  BUFFD0 U2972 ( .I(n2990), .Z(n2989) );
  BUFFD0 U2973 ( .I(n2991), .Z(n2990) );
  BUFFD0 U2974 ( .I(n2992), .Z(n2991) );
  BUFFD0 U2975 ( .I(n2993), .Z(n2992) );
  BUFFD0 U2976 ( .I(n2994), .Z(n2993) );
  BUFFD0 U2977 ( .I(n2995), .Z(n2994) );
  BUFFD0 U2978 ( .I(n2996), .Z(n2995) );
  BUFFD0 U2979 ( .I(n2997), .Z(n2996) );
  BUFFD0 U2980 ( .I(n2998), .Z(n2997) );
  BUFFD0 U2981 ( .I(n2999), .Z(n2998) );
  BUFFD0 U2982 ( .I(n3000), .Z(n2999) );
  BUFFD0 U2983 ( .I(n3001), .Z(n3000) );
  BUFFD0 U2984 ( .I(n3002), .Z(n3001) );
  BUFFD0 U2985 ( .I(n3003), .Z(n3002) );
  BUFFD0 U2986 ( .I(n3004), .Z(n3003) );
  BUFFD0 U2987 ( .I(n3005), .Z(n3004) );
  BUFFD0 U2988 ( .I(n3006), .Z(n3005) );
  BUFFD0 U2989 ( .I(n3007), .Z(n3006) );
  BUFFD0 U2990 ( .I(n3008), .Z(n3007) );
  BUFFD0 U2991 ( .I(n3009), .Z(n3008) );
  BUFFD0 U2992 ( .I(n3010), .Z(n3009) );
  BUFFD0 U2993 ( .I(n3011), .Z(n3010) );
  BUFFD0 U2994 ( .I(n3012), .Z(n3011) );
  BUFFD0 U2995 ( .I(n3013), .Z(n3012) );
  BUFFD0 U2996 ( .I(n3014), .Z(n3013) );
  BUFFD0 U2997 ( .I(n3015), .Z(n3014) );
  BUFFD0 U2998 ( .I(n3016), .Z(n3015) );
  BUFFD0 U2999 ( .I(n3017), .Z(n3016) );
  BUFFD0 U3000 ( .I(n3018), .Z(n3017) );
  BUFFD0 U3001 ( .I(n3019), .Z(n3018) );
  BUFFD0 U3002 ( .I(n3020), .Z(n3019) );
  BUFFD0 U3003 ( .I(n3021), .Z(n3020) );
  BUFFD0 U3004 ( .I(n3022), .Z(n3021) );
  BUFFD0 U3005 ( .I(n3023), .Z(n3022) );
  BUFFD0 U3006 ( .I(n3024), .Z(n3023) );
  BUFFD0 U3007 ( .I(n3025), .Z(n3024) );
  BUFFD0 U3008 ( .I(n3026), .Z(n3025) );
  BUFFD0 U3009 ( .I(n3027), .Z(n3026) );
  BUFFD0 U3010 ( .I(n3028), .Z(n3027) );
  BUFFD0 U3011 ( .I(n3029), .Z(n3028) );
  BUFFD0 U3012 ( .I(n3030), .Z(n3029) );
  BUFFD0 U3013 ( .I(n3031), .Z(n3030) );
  BUFFD0 U3014 ( .I(n3032), .Z(n3031) );
  BUFFD0 U3015 ( .I(n3033), .Z(n3032) );
  BUFFD0 U3016 ( .I(n3034), .Z(n3033) );
  BUFFD0 U3017 ( .I(n3035), .Z(n3034) );
  BUFFD0 U3018 ( .I(n3036), .Z(n3035) );
  BUFFD0 U3019 ( .I(n3037), .Z(n3036) );
  BUFFD0 U3020 ( .I(n3038), .Z(n3037) );
  BUFFD0 U3021 ( .I(n3039), .Z(n3038) );
  BUFFD0 U3022 ( .I(n3040), .Z(n3039) );
  BUFFD0 U3023 ( .I(n3041), .Z(n3040) );
  BUFFD0 U3024 ( .I(N70), .Z(n3041) );
  BUFFD0 U3025 ( .I(n4090), .Z(n3042) );
  BUFFD0 U3026 ( .I(n3044), .Z(n3043) );
  BUFFD0 U3027 ( .I(n3045), .Z(n3044) );
  BUFFD0 U3028 ( .I(n3046), .Z(n3045) );
  BUFFD0 U3029 ( .I(n3047), .Z(n3046) );
  BUFFD0 U3030 ( .I(n3048), .Z(n3047) );
  BUFFD0 U3031 ( .I(n3049), .Z(n3048) );
  BUFFD0 U3032 ( .I(n3050), .Z(n3049) );
  BUFFD0 U3033 ( .I(n3051), .Z(n3050) );
  BUFFD0 U3034 ( .I(n3052), .Z(n3051) );
  BUFFD0 U3035 ( .I(n3053), .Z(n3052) );
  BUFFD0 U3036 ( .I(n3054), .Z(n3053) );
  BUFFD0 U3037 ( .I(n3055), .Z(n3054) );
  BUFFD0 U3038 ( .I(n3056), .Z(n3055) );
  BUFFD0 U3039 ( .I(n3057), .Z(n3056) );
  BUFFD0 U3040 ( .I(n3058), .Z(n3057) );
  BUFFD0 U3041 ( .I(n3059), .Z(n3058) );
  BUFFD0 U3042 ( .I(n3060), .Z(n3059) );
  BUFFD0 U3043 ( .I(n3061), .Z(n3060) );
  BUFFD0 U3044 ( .I(n3062), .Z(n3061) );
  BUFFD0 U3045 ( .I(n3063), .Z(n3062) );
  BUFFD0 U3046 ( .I(n3064), .Z(n3063) );
  BUFFD0 U3047 ( .I(n3065), .Z(n3064) );
  BUFFD0 U3048 ( .I(n3066), .Z(n3065) );
  BUFFD0 U3049 ( .I(n3067), .Z(n3066) );
  BUFFD0 U3050 ( .I(n3068), .Z(n3067) );
  BUFFD0 U3051 ( .I(n3069), .Z(n3068) );
  BUFFD0 U3052 ( .I(n3070), .Z(n3069) );
  BUFFD0 U3053 ( .I(n3071), .Z(n3070) );
  BUFFD0 U3054 ( .I(n3072), .Z(n3071) );
  BUFFD0 U3055 ( .I(n3073), .Z(n3072) );
  BUFFD0 U3056 ( .I(n3074), .Z(n3073) );
  BUFFD0 U3057 ( .I(n3075), .Z(n3074) );
  BUFFD0 U3058 ( .I(n3076), .Z(n3075) );
  BUFFD0 U3059 ( .I(n3077), .Z(n3076) );
  BUFFD0 U3060 ( .I(n3078), .Z(n3077) );
  BUFFD0 U3061 ( .I(n3079), .Z(n3078) );
  BUFFD0 U3062 ( .I(n3080), .Z(n3079) );
  BUFFD0 U3063 ( .I(n3081), .Z(n3080) );
  BUFFD0 U3064 ( .I(n3082), .Z(n3081) );
  BUFFD0 U3065 ( .I(n3083), .Z(n3082) );
  BUFFD0 U3066 ( .I(n3084), .Z(n3083) );
  BUFFD0 U3067 ( .I(n3085), .Z(n3084) );
  BUFFD0 U3068 ( .I(n3086), .Z(n3085) );
  BUFFD0 U3069 ( .I(n3087), .Z(n3086) );
  BUFFD0 U3070 ( .I(n3088), .Z(n3087) );
  BUFFD0 U3071 ( .I(n3089), .Z(n3088) );
  BUFFD0 U3072 ( .I(n3090), .Z(n3089) );
  BUFFD0 U3073 ( .I(n3091), .Z(n3090) );
  BUFFD0 U3074 ( .I(n3092), .Z(n3091) );
  BUFFD0 U3075 ( .I(n3093), .Z(n3092) );
  BUFFD0 U3076 ( .I(n3094), .Z(n3093) );
  BUFFD0 U3077 ( .I(n3095), .Z(n3094) );
  BUFFD0 U3078 ( .I(n3096), .Z(n3095) );
  BUFFD0 U3079 ( .I(n3097), .Z(n3096) );
  BUFFD0 U3080 ( .I(n3098), .Z(n3097) );
  BUFFD0 U3081 ( .I(n3099), .Z(n3098) );
  BUFFD0 U3082 ( .I(n3100), .Z(n3099) );
  BUFFD0 U3083 ( .I(n3101), .Z(n3100) );
  BUFFD0 U3084 ( .I(n3102), .Z(n3101) );
  BUFFD0 U3085 ( .I(n3103), .Z(n3102) );
  BUFFD0 U3086 ( .I(n3104), .Z(n3103) );
  BUFFD0 U3087 ( .I(n3105), .Z(n3104) );
  BUFFD0 U3088 ( .I(n3106), .Z(n3105) );
  BUFFD0 U3089 ( .I(n3107), .Z(n3106) );
  BUFFD0 U3090 ( .I(N71), .Z(n3107) );
  BUFFD0 U3091 ( .I(n4077), .Z(n3108) );
  BUFFD0 U3092 ( .I(n3113), .Z(n3109) );
  BUFFD0 U3093 ( .I(n3172), .Z(n3110) );
  BUFFD0 U3094 ( .I(n3110), .Z(n3111) );
  BUFFD0 U3095 ( .I(n3111), .Z(n3112) );
  BUFFD0 U3096 ( .I(n3114), .Z(n3113) );
  BUFFD0 U3097 ( .I(n3115), .Z(n3114) );
  BUFFD0 U3098 ( .I(n3116), .Z(n3115) );
  BUFFD0 U3099 ( .I(n3117), .Z(n3116) );
  BUFFD0 U3100 ( .I(n3118), .Z(n3117) );
  BUFFD0 U3101 ( .I(n3119), .Z(n3118) );
  BUFFD0 U3102 ( .I(n3120), .Z(n3119) );
  BUFFD0 U3103 ( .I(n3121), .Z(n3120) );
  BUFFD0 U3104 ( .I(n3122), .Z(n3121) );
  BUFFD0 U3105 ( .I(n3123), .Z(n3122) );
  BUFFD0 U3106 ( .I(n3124), .Z(n3123) );
  BUFFD0 U3107 ( .I(n3125), .Z(n3124) );
  BUFFD0 U3108 ( .I(n3126), .Z(n3125) );
  BUFFD0 U3109 ( .I(n3127), .Z(n3126) );
  BUFFD0 U3110 ( .I(n3128), .Z(n3127) );
  BUFFD0 U3111 ( .I(n3129), .Z(n3128) );
  BUFFD0 U3112 ( .I(n3130), .Z(n3129) );
  BUFFD0 U3113 ( .I(n3131), .Z(n3130) );
  BUFFD0 U3114 ( .I(n3132), .Z(n3131) );
  BUFFD0 U3115 ( .I(n3133), .Z(n3132) );
  BUFFD0 U3116 ( .I(n3134), .Z(n3133) );
  BUFFD0 U3117 ( .I(n3135), .Z(n3134) );
  BUFFD0 U3118 ( .I(n3136), .Z(n3135) );
  BUFFD0 U3119 ( .I(n3137), .Z(n3136) );
  BUFFD0 U3120 ( .I(n3138), .Z(n3137) );
  BUFFD0 U3121 ( .I(n3139), .Z(n3138) );
  BUFFD0 U3122 ( .I(n3140), .Z(n3139) );
  BUFFD0 U3123 ( .I(n3141), .Z(n3140) );
  BUFFD0 U3124 ( .I(n3142), .Z(n3141) );
  BUFFD0 U3125 ( .I(n3143), .Z(n3142) );
  BUFFD0 U3126 ( .I(n3144), .Z(n3143) );
  BUFFD0 U3127 ( .I(n3145), .Z(n3144) );
  BUFFD0 U3128 ( .I(n3146), .Z(n3145) );
  BUFFD0 U3129 ( .I(n3147), .Z(n3146) );
  BUFFD0 U3130 ( .I(n3148), .Z(n3147) );
  BUFFD0 U3131 ( .I(n3149), .Z(n3148) );
  BUFFD0 U3132 ( .I(n3150), .Z(n3149) );
  BUFFD0 U3133 ( .I(n3151), .Z(n3150) );
  BUFFD0 U3134 ( .I(n3152), .Z(n3151) );
  BUFFD0 U3135 ( .I(n3153), .Z(n3152) );
  BUFFD0 U3136 ( .I(n3154), .Z(n3153) );
  BUFFD0 U3137 ( .I(n3155), .Z(n3154) );
  BUFFD0 U3138 ( .I(n3156), .Z(n3155) );
  BUFFD0 U3139 ( .I(n3157), .Z(n3156) );
  BUFFD0 U3140 ( .I(n3158), .Z(n3157) );
  BUFFD0 U3141 ( .I(n3159), .Z(n3158) );
  BUFFD0 U3142 ( .I(n3160), .Z(n3159) );
  BUFFD0 U3143 ( .I(n3161), .Z(n3160) );
  BUFFD0 U3144 ( .I(n3162), .Z(n3161) );
  BUFFD0 U3145 ( .I(n3163), .Z(n3162) );
  BUFFD0 U3146 ( .I(n3164), .Z(n3163) );
  BUFFD0 U3147 ( .I(n3165), .Z(n3164) );
  BUFFD0 U3148 ( .I(n3166), .Z(n3165) );
  BUFFD0 U3149 ( .I(n3167), .Z(n3166) );
  BUFFD0 U3150 ( .I(n3168), .Z(n3167) );
  BUFFD0 U3151 ( .I(n3169), .Z(n3168) );
  BUFFD0 U3152 ( .I(n3171), .Z(n3169) );
  BUFFD0 U3153 ( .I(N72), .Z(n3170) );
  BUFFD0 U3154 ( .I(n3173), .Z(n3171) );
  BUFFD0 U3155 ( .I(n3170), .Z(n3172) );
  BUFFD0 U3156 ( .I(n3112), .Z(n3173) );
  BUFFD0 U3157 ( .I(n3178), .Z(n3174) );
  BUFFD0 U3158 ( .I(n3862), .Z(n3175) );
  BUFFD0 U3159 ( .I(n3175), .Z(n3176) );
  BUFFD0 U3160 ( .I(n3176), .Z(n3177) );
  BUFFD0 U3161 ( .I(n3179), .Z(n3178) );
  BUFFD0 U3162 ( .I(n3180), .Z(n3179) );
  BUFFD0 U3163 ( .I(n3181), .Z(n3180) );
  BUFFD0 U3164 ( .I(n3182), .Z(n3181) );
  BUFFD0 U3165 ( .I(n3183), .Z(n3182) );
  BUFFD0 U3166 ( .I(n3184), .Z(n3183) );
  BUFFD0 U3167 ( .I(n3185), .Z(n3184) );
  BUFFD0 U3168 ( .I(n3186), .Z(n3185) );
  BUFFD0 U3169 ( .I(n3187), .Z(n3186) );
  BUFFD0 U3170 ( .I(n3188), .Z(n3187) );
  BUFFD0 U3171 ( .I(n3189), .Z(n3188) );
  BUFFD0 U3172 ( .I(n3190), .Z(n3189) );
  BUFFD0 U3173 ( .I(n3191), .Z(n3190) );
  BUFFD0 U3174 ( .I(n3192), .Z(n3191) );
  BUFFD0 U3175 ( .I(n3193), .Z(n3192) );
  BUFFD0 U3176 ( .I(n3194), .Z(n3193) );
  BUFFD0 U3177 ( .I(n3195), .Z(n3194) );
  BUFFD0 U3178 ( .I(n3196), .Z(n3195) );
  BUFFD0 U3179 ( .I(n3197), .Z(n3196) );
  BUFFD0 U3180 ( .I(n3198), .Z(n3197) );
  BUFFD0 U3181 ( .I(n3199), .Z(n3198) );
  BUFFD0 U3182 ( .I(n3200), .Z(n3199) );
  BUFFD0 U3183 ( .I(n3201), .Z(n3200) );
  BUFFD0 U3184 ( .I(n3202), .Z(n3201) );
  BUFFD0 U3185 ( .I(n3203), .Z(n3202) );
  BUFFD0 U3186 ( .I(n3204), .Z(n3203) );
  BUFFD0 U3187 ( .I(n3205), .Z(n3204) );
  BUFFD0 U3188 ( .I(n3206), .Z(n3205) );
  BUFFD0 U3189 ( .I(n3207), .Z(n3206) );
  BUFFD0 U3190 ( .I(n3208), .Z(n3207) );
  BUFFD0 U3191 ( .I(n3209), .Z(n3208) );
  BUFFD0 U3192 ( .I(n3210), .Z(n3209) );
  BUFFD0 U3193 ( .I(n3211), .Z(n3210) );
  BUFFD0 U3194 ( .I(n3212), .Z(n3211) );
  BUFFD0 U3195 ( .I(n3213), .Z(n3212) );
  BUFFD0 U3196 ( .I(n3214), .Z(n3213) );
  BUFFD0 U3197 ( .I(n3215), .Z(n3214) );
  BUFFD0 U3198 ( .I(n3216), .Z(n3215) );
  BUFFD0 U3199 ( .I(n3217), .Z(n3216) );
  BUFFD0 U3200 ( .I(n3218), .Z(n3217) );
  BUFFD0 U3201 ( .I(n3219), .Z(n3218) );
  BUFFD0 U3202 ( .I(n3220), .Z(n3219) );
  BUFFD0 U3203 ( .I(n3221), .Z(n3220) );
  BUFFD0 U3204 ( .I(n3222), .Z(n3221) );
  BUFFD0 U3205 ( .I(n3223), .Z(n3222) );
  BUFFD0 U3206 ( .I(n3224), .Z(n3223) );
  BUFFD0 U3207 ( .I(n3225), .Z(n3224) );
  BUFFD0 U3208 ( .I(n3226), .Z(n3225) );
  BUFFD0 U3209 ( .I(n3227), .Z(n3226) );
  BUFFD0 U3210 ( .I(n3228), .Z(n3227) );
  BUFFD0 U3211 ( .I(n3229), .Z(n3228) );
  BUFFD0 U3212 ( .I(n3230), .Z(n3229) );
  BUFFD0 U3213 ( .I(n3231), .Z(n3230) );
  BUFFD0 U3214 ( .I(n3232), .Z(n3231) );
  BUFFD0 U3215 ( .I(n3233), .Z(n3232) );
  BUFFD0 U3216 ( .I(n3234), .Z(n3233) );
  BUFFD0 U3217 ( .I(n3235), .Z(n3234) );
  BUFFD0 U3218 ( .I(n3177), .Z(n3235) );
  BUFFD0 U3219 ( .I(n3241), .Z(n3236) );
  BUFFD0 U3220 ( .I(n3864), .Z(n3237) );
  BUFFD0 U3221 ( .I(n3237), .Z(n3238) );
  BUFFD0 U3222 ( .I(n3238), .Z(n3239) );
  BUFFD0 U3223 ( .I(n3239), .Z(n3240) );
  BUFFD0 U3224 ( .I(n3242), .Z(n3241) );
  BUFFD0 U3225 ( .I(n3243), .Z(n3242) );
  BUFFD0 U3226 ( .I(n3244), .Z(n3243) );
  BUFFD0 U3227 ( .I(n3245), .Z(n3244) );
  BUFFD0 U3228 ( .I(n3246), .Z(n3245) );
  BUFFD0 U3229 ( .I(n3247), .Z(n3246) );
  BUFFD0 U3230 ( .I(n3248), .Z(n3247) );
  BUFFD0 U3231 ( .I(n3249), .Z(n3248) );
  BUFFD0 U3232 ( .I(n3250), .Z(n3249) );
  BUFFD0 U3233 ( .I(n3251), .Z(n3250) );
  BUFFD0 U3234 ( .I(n3252), .Z(n3251) );
  BUFFD0 U3235 ( .I(n3253), .Z(n3252) );
  BUFFD0 U3236 ( .I(n3254), .Z(n3253) );
  BUFFD0 U3237 ( .I(n3255), .Z(n3254) );
  BUFFD0 U3238 ( .I(n3256), .Z(n3255) );
  BUFFD0 U3239 ( .I(n3257), .Z(n3256) );
  BUFFD0 U3240 ( .I(n3258), .Z(n3257) );
  BUFFD0 U3241 ( .I(n3259), .Z(n3258) );
  BUFFD0 U3242 ( .I(n3260), .Z(n3259) );
  BUFFD0 U3243 ( .I(n3261), .Z(n3260) );
  BUFFD0 U3244 ( .I(n3262), .Z(n3261) );
  BUFFD0 U3245 ( .I(n3263), .Z(n3262) );
  BUFFD0 U3246 ( .I(n3264), .Z(n3263) );
  BUFFD0 U3247 ( .I(n3265), .Z(n3264) );
  BUFFD0 U3248 ( .I(n3266), .Z(n3265) );
  BUFFD0 U3249 ( .I(n3267), .Z(n3266) );
  BUFFD0 U3250 ( .I(n3268), .Z(n3267) );
  BUFFD0 U3251 ( .I(n3269), .Z(n3268) );
  BUFFD0 U3252 ( .I(n3270), .Z(n3269) );
  BUFFD0 U3253 ( .I(n3271), .Z(n3270) );
  BUFFD0 U3254 ( .I(n3272), .Z(n3271) );
  BUFFD0 U3255 ( .I(n3273), .Z(n3272) );
  BUFFD0 U3256 ( .I(n3274), .Z(n3273) );
  BUFFD0 U3257 ( .I(n3275), .Z(n3274) );
  BUFFD0 U3258 ( .I(n3276), .Z(n3275) );
  BUFFD0 U3259 ( .I(n3277), .Z(n3276) );
  BUFFD0 U3260 ( .I(n3278), .Z(n3277) );
  BUFFD0 U3261 ( .I(n3279), .Z(n3278) );
  BUFFD0 U3262 ( .I(n3280), .Z(n3279) );
  BUFFD0 U3263 ( .I(n3281), .Z(n3280) );
  BUFFD0 U3264 ( .I(n3282), .Z(n3281) );
  BUFFD0 U3265 ( .I(n3283), .Z(n3282) );
  BUFFD0 U3266 ( .I(n3284), .Z(n3283) );
  BUFFD0 U3267 ( .I(n3285), .Z(n3284) );
  BUFFD0 U3268 ( .I(n3286), .Z(n3285) );
  BUFFD0 U3269 ( .I(n3287), .Z(n3286) );
  BUFFD0 U3270 ( .I(n3288), .Z(n3287) );
  BUFFD0 U3271 ( .I(n3289), .Z(n3288) );
  BUFFD0 U3272 ( .I(n3290), .Z(n3289) );
  BUFFD0 U3273 ( .I(n3291), .Z(n3290) );
  BUFFD0 U3274 ( .I(n3292), .Z(n3291) );
  BUFFD0 U3275 ( .I(n3293), .Z(n3292) );
  BUFFD0 U3276 ( .I(n3294), .Z(n3293) );
  BUFFD0 U3277 ( .I(n3295), .Z(n3294) );
  BUFFD0 U3278 ( .I(n3296), .Z(n3295) );
  BUFFD0 U3279 ( .I(n3240), .Z(n3296) );
  MUX3ND1 U3280 ( .I0(n4023), .I1(n4024), .I2(n3863), .S0(n4641), .S1(n4352), 
        .ZN(N75) );
  BUFFD0 U3281 ( .I(n3798), .Z(n3297) );
  BUFFD0 U3282 ( .I(n3297), .Z(n3298) );
  BUFFD0 U3283 ( .I(n3298), .Z(n3299) );
  BUFFD0 U3284 ( .I(n3299), .Z(n3300) );
  BUFFD0 U3285 ( .I(n3302), .Z(n3301) );
  BUFFD0 U3286 ( .I(n3303), .Z(n3302) );
  BUFFD0 U3287 ( .I(n3304), .Z(n3303) );
  BUFFD0 U3288 ( .I(n3305), .Z(n3304) );
  BUFFD0 U3289 ( .I(n3306), .Z(n3305) );
  BUFFD0 U3290 ( .I(n3307), .Z(n3306) );
  BUFFD0 U3291 ( .I(n3308), .Z(n3307) );
  BUFFD0 U3292 ( .I(n3309), .Z(n3308) );
  BUFFD0 U3293 ( .I(n3310), .Z(n3309) );
  BUFFD0 U3294 ( .I(n3311), .Z(n3310) );
  BUFFD0 U3295 ( .I(n3312), .Z(n3311) );
  BUFFD0 U3296 ( .I(n3313), .Z(n3312) );
  BUFFD0 U3297 ( .I(n3314), .Z(n3313) );
  BUFFD0 U3298 ( .I(n3315), .Z(n3314) );
  BUFFD0 U3299 ( .I(n3316), .Z(n3315) );
  BUFFD0 U3300 ( .I(n3317), .Z(n3316) );
  BUFFD0 U3301 ( .I(n3318), .Z(n3317) );
  BUFFD0 U3302 ( .I(n3319), .Z(n3318) );
  BUFFD0 U3303 ( .I(n3320), .Z(n3319) );
  BUFFD0 U3304 ( .I(n3321), .Z(n3320) );
  BUFFD0 U3305 ( .I(n3322), .Z(n3321) );
  BUFFD0 U3306 ( .I(n3323), .Z(n3322) );
  BUFFD0 U3307 ( .I(n3324), .Z(n3323) );
  BUFFD0 U3308 ( .I(n3325), .Z(n3324) );
  BUFFD0 U3309 ( .I(n3326), .Z(n3325) );
  BUFFD0 U3310 ( .I(n3327), .Z(n3326) );
  BUFFD0 U3311 ( .I(n3328), .Z(n3327) );
  BUFFD0 U3312 ( .I(n3329), .Z(n3328) );
  BUFFD0 U3313 ( .I(n3330), .Z(n3329) );
  BUFFD0 U3314 ( .I(n3331), .Z(n3330) );
  BUFFD0 U3315 ( .I(n3332), .Z(n3331) );
  BUFFD0 U3316 ( .I(n3333), .Z(n3332) );
  BUFFD0 U3317 ( .I(n3334), .Z(n3333) );
  BUFFD0 U3318 ( .I(n3335), .Z(n3334) );
  BUFFD0 U3319 ( .I(n3336), .Z(n3335) );
  BUFFD0 U3320 ( .I(n3337), .Z(n3336) );
  BUFFD0 U3321 ( .I(n3338), .Z(n3337) );
  BUFFD0 U3322 ( .I(n3339), .Z(n3338) );
  BUFFD0 U3323 ( .I(n3340), .Z(n3339) );
  BUFFD0 U3324 ( .I(n3341), .Z(n3340) );
  BUFFD0 U3325 ( .I(n3342), .Z(n3341) );
  BUFFD0 U3326 ( .I(n3343), .Z(n3342) );
  BUFFD0 U3327 ( .I(n3344), .Z(n3343) );
  BUFFD0 U3328 ( .I(n3345), .Z(n3344) );
  BUFFD0 U3329 ( .I(n3346), .Z(n3345) );
  BUFFD0 U3330 ( .I(n3347), .Z(n3346) );
  BUFFD0 U3331 ( .I(n3348), .Z(n3347) );
  BUFFD0 U3332 ( .I(n3349), .Z(n3348) );
  BUFFD0 U3333 ( .I(n3350), .Z(n3349) );
  BUFFD0 U3334 ( .I(n3351), .Z(n3350) );
  BUFFD0 U3335 ( .I(n3352), .Z(n3351) );
  BUFFD0 U3336 ( .I(n3353), .Z(n3352) );
  BUFFD0 U3337 ( .I(n3354), .Z(n3353) );
  BUFFD0 U3338 ( .I(n3355), .Z(n3354) );
  BUFFD0 U3339 ( .I(n3356), .Z(n3355) );
  BUFFD0 U3340 ( .I(n3357), .Z(n3356) );
  BUFFD0 U3341 ( .I(n3358), .Z(n3357) );
  BUFFD0 U3342 ( .I(n3359), .Z(n3358) );
  BUFFD0 U3343 ( .I(n3300), .Z(n3359) );
  BUFFD0 U3344 ( .I(n3365), .Z(n3360) );
  BUFFD0 U3345 ( .I(n3818), .Z(n3361) );
  BUFFD0 U3346 ( .I(n3361), .Z(n3362) );
  BUFFD0 U3347 ( .I(n3362), .Z(n3363) );
  BUFFD0 U3348 ( .I(n3363), .Z(n3364) );
  BUFFD0 U3349 ( .I(n3366), .Z(n3365) );
  BUFFD0 U3350 ( .I(n3367), .Z(n3366) );
  BUFFD0 U3351 ( .I(n3368), .Z(n3367) );
  BUFFD0 U3352 ( .I(n3369), .Z(n3368) );
  BUFFD0 U3353 ( .I(n3370), .Z(n3369) );
  BUFFD0 U3354 ( .I(n3371), .Z(n3370) );
  BUFFD0 U3355 ( .I(n3372), .Z(n3371) );
  BUFFD0 U3356 ( .I(n3373), .Z(n3372) );
  BUFFD0 U3357 ( .I(n3374), .Z(n3373) );
  BUFFD0 U3358 ( .I(n3375), .Z(n3374) );
  BUFFD0 U3359 ( .I(n3376), .Z(n3375) );
  BUFFD0 U3360 ( .I(n3377), .Z(n3376) );
  BUFFD0 U3361 ( .I(n3378), .Z(n3377) );
  BUFFD0 U3362 ( .I(n3379), .Z(n3378) );
  BUFFD0 U3363 ( .I(n3380), .Z(n3379) );
  BUFFD0 U3364 ( .I(n3381), .Z(n3380) );
  BUFFD0 U3365 ( .I(n3382), .Z(n3381) );
  BUFFD0 U3366 ( .I(n3383), .Z(n3382) );
  BUFFD0 U3367 ( .I(n3384), .Z(n3383) );
  BUFFD0 U3368 ( .I(n3385), .Z(n3384) );
  BUFFD0 U3369 ( .I(n3386), .Z(n3385) );
  BUFFD0 U3370 ( .I(n3387), .Z(n3386) );
  BUFFD0 U3371 ( .I(n3388), .Z(n3387) );
  BUFFD0 U3372 ( .I(n3389), .Z(n3388) );
  BUFFD0 U3373 ( .I(n3390), .Z(n3389) );
  BUFFD0 U3374 ( .I(n3391), .Z(n3390) );
  BUFFD0 U3375 ( .I(n3392), .Z(n3391) );
  BUFFD0 U3376 ( .I(n3393), .Z(n3392) );
  BUFFD0 U3377 ( .I(n3394), .Z(n3393) );
  BUFFD0 U3378 ( .I(n3395), .Z(n3394) );
  BUFFD0 U3379 ( .I(n3396), .Z(n3395) );
  BUFFD0 U3380 ( .I(n3397), .Z(n3396) );
  BUFFD0 U3381 ( .I(n3398), .Z(n3397) );
  BUFFD0 U3382 ( .I(n3399), .Z(n3398) );
  BUFFD0 U3383 ( .I(n3400), .Z(n3399) );
  BUFFD0 U3384 ( .I(n3401), .Z(n3400) );
  BUFFD0 U3385 ( .I(n3402), .Z(n3401) );
  BUFFD0 U3386 ( .I(n3403), .Z(n3402) );
  BUFFD0 U3387 ( .I(n3404), .Z(n3403) );
  BUFFD0 U3388 ( .I(n3405), .Z(n3404) );
  BUFFD0 U3389 ( .I(n3406), .Z(n3405) );
  BUFFD0 U3390 ( .I(n3407), .Z(n3406) );
  BUFFD0 U3391 ( .I(n3408), .Z(n3407) );
  BUFFD0 U3392 ( .I(n3409), .Z(n3408) );
  BUFFD0 U3393 ( .I(n3410), .Z(n3409) );
  BUFFD0 U3394 ( .I(n3411), .Z(n3410) );
  BUFFD0 U3395 ( .I(n3412), .Z(n3411) );
  BUFFD0 U3396 ( .I(n3413), .Z(n3412) );
  BUFFD0 U3397 ( .I(n3414), .Z(n3413) );
  BUFFD0 U3398 ( .I(n3415), .Z(n3414) );
  BUFFD0 U3399 ( .I(n3416), .Z(n3415) );
  BUFFD0 U3400 ( .I(n3417), .Z(n3416) );
  BUFFD0 U3401 ( .I(n3418), .Z(n3417) );
  BUFFD0 U3402 ( .I(n3419), .Z(n3418) );
  BUFFD0 U3403 ( .I(n3420), .Z(n3419) );
  BUFFD0 U3404 ( .I(n3421), .Z(n3420) );
  BUFFD0 U3405 ( .I(n3422), .Z(n3421) );
  BUFFD0 U3406 ( .I(n3364), .Z(n3422) );
  BUFFD0 U3407 ( .I(n3427), .Z(n3423) );
  BUFFD0 U3408 ( .I(n3820), .Z(n3424) );
  BUFFD0 U3409 ( .I(n3424), .Z(n3425) );
  BUFFD0 U3410 ( .I(n3425), .Z(n3426) );
  BUFFD0 U3411 ( .I(n3428), .Z(n3427) );
  BUFFD0 U3412 ( .I(n3429), .Z(n3428) );
  BUFFD0 U3413 ( .I(n3430), .Z(n3429) );
  BUFFD0 U3414 ( .I(n3431), .Z(n3430) );
  BUFFD0 U3415 ( .I(n3432), .Z(n3431) );
  BUFFD0 U3416 ( .I(n3433), .Z(n3432) );
  BUFFD0 U3417 ( .I(n3434), .Z(n3433) );
  BUFFD0 U3418 ( .I(n3435), .Z(n3434) );
  BUFFD0 U3419 ( .I(n3436), .Z(n3435) );
  BUFFD0 U3420 ( .I(n3437), .Z(n3436) );
  BUFFD0 U3421 ( .I(n3438), .Z(n3437) );
  BUFFD0 U3422 ( .I(n3439), .Z(n3438) );
  BUFFD0 U3423 ( .I(n3440), .Z(n3439) );
  BUFFD0 U3424 ( .I(n3441), .Z(n3440) );
  BUFFD0 U3425 ( .I(n3442), .Z(n3441) );
  BUFFD0 U3426 ( .I(n3443), .Z(n3442) );
  BUFFD0 U3427 ( .I(n3444), .Z(n3443) );
  BUFFD0 U3428 ( .I(n3445), .Z(n3444) );
  BUFFD0 U3429 ( .I(n3446), .Z(n3445) );
  BUFFD0 U3430 ( .I(n3447), .Z(n3446) );
  BUFFD0 U3431 ( .I(n3448), .Z(n3447) );
  BUFFD0 U3432 ( .I(n3449), .Z(n3448) );
  BUFFD0 U3433 ( .I(n3450), .Z(n3449) );
  BUFFD0 U3434 ( .I(n3451), .Z(n3450) );
  BUFFD0 U3435 ( .I(n3452), .Z(n3451) );
  BUFFD0 U3436 ( .I(n3453), .Z(n3452) );
  BUFFD0 U3437 ( .I(n3454), .Z(n3453) );
  BUFFD0 U3438 ( .I(n3455), .Z(n3454) );
  BUFFD0 U3439 ( .I(n3456), .Z(n3455) );
  BUFFD0 U3440 ( .I(n3457), .Z(n3456) );
  BUFFD0 U3441 ( .I(n3458), .Z(n3457) );
  BUFFD0 U3442 ( .I(n3459), .Z(n3458) );
  BUFFD0 U3443 ( .I(n3460), .Z(n3459) );
  BUFFD0 U3444 ( .I(n3461), .Z(n3460) );
  BUFFD0 U3445 ( .I(n3462), .Z(n3461) );
  BUFFD0 U3446 ( .I(n3463), .Z(n3462) );
  BUFFD0 U3447 ( .I(n3464), .Z(n3463) );
  BUFFD0 U3448 ( .I(n3465), .Z(n3464) );
  BUFFD0 U3449 ( .I(n3466), .Z(n3465) );
  BUFFD0 U3450 ( .I(n3467), .Z(n3466) );
  BUFFD0 U3451 ( .I(n3468), .Z(n3467) );
  BUFFD0 U3452 ( .I(n3469), .Z(n3468) );
  BUFFD0 U3453 ( .I(n3470), .Z(n3469) );
  BUFFD0 U3454 ( .I(n3471), .Z(n3470) );
  BUFFD0 U3455 ( .I(n3472), .Z(n3471) );
  BUFFD0 U3456 ( .I(n3473), .Z(n3472) );
  BUFFD0 U3457 ( .I(n3474), .Z(n3473) );
  BUFFD0 U3458 ( .I(n3475), .Z(n3474) );
  BUFFD0 U3459 ( .I(n3476), .Z(n3475) );
  BUFFD0 U3460 ( .I(n3477), .Z(n3476) );
  BUFFD0 U3461 ( .I(n3478), .Z(n3477) );
  BUFFD0 U3462 ( .I(n3479), .Z(n3478) );
  BUFFD0 U3463 ( .I(n3480), .Z(n3479) );
  BUFFD0 U3464 ( .I(n3481), .Z(n3480) );
  BUFFD0 U3465 ( .I(n3482), .Z(n3481) );
  BUFFD0 U3466 ( .I(n3483), .Z(n3482) );
  BUFFD0 U3467 ( .I(n3484), .Z(n3483) );
  BUFFD0 U3468 ( .I(n3485), .Z(n3484) );
  BUFFD0 U3469 ( .I(n3426), .Z(n3485) );
  BUFFD0 U3470 ( .I(n3490), .Z(n3486) );
  BUFFD0 U3471 ( .I(n3821), .Z(n3487) );
  BUFFD0 U3472 ( .I(n3487), .Z(n3488) );
  BUFFD0 U3473 ( .I(n3488), .Z(n3489) );
  BUFFD0 U3474 ( .I(n3491), .Z(n3490) );
  BUFFD0 U3475 ( .I(n3492), .Z(n3491) );
  BUFFD0 U3476 ( .I(n3493), .Z(n3492) );
  BUFFD0 U3477 ( .I(n3494), .Z(n3493) );
  BUFFD0 U3478 ( .I(n3495), .Z(n3494) );
  BUFFD0 U3479 ( .I(n3496), .Z(n3495) );
  BUFFD0 U3480 ( .I(n3497), .Z(n3496) );
  BUFFD0 U3481 ( .I(n3498), .Z(n3497) );
  BUFFD0 U3482 ( .I(n3499), .Z(n3498) );
  BUFFD0 U3483 ( .I(n3500), .Z(n3499) );
  BUFFD0 U3484 ( .I(n3501), .Z(n3500) );
  BUFFD0 U3485 ( .I(n3502), .Z(n3501) );
  BUFFD0 U3486 ( .I(n3503), .Z(n3502) );
  BUFFD0 U3487 ( .I(n3504), .Z(n3503) );
  BUFFD0 U3488 ( .I(n3505), .Z(n3504) );
  BUFFD0 U3489 ( .I(n3506), .Z(n3505) );
  BUFFD0 U3490 ( .I(n3507), .Z(n3506) );
  BUFFD0 U3491 ( .I(n3508), .Z(n3507) );
  BUFFD0 U3492 ( .I(n3509), .Z(n3508) );
  BUFFD0 U3493 ( .I(n3510), .Z(n3509) );
  BUFFD0 U3494 ( .I(n3511), .Z(n3510) );
  BUFFD0 U3495 ( .I(n3512), .Z(n3511) );
  BUFFD0 U3496 ( .I(n3513), .Z(n3512) );
  BUFFD0 U3497 ( .I(n3514), .Z(n3513) );
  BUFFD0 U3498 ( .I(n3515), .Z(n3514) );
  BUFFD0 U3499 ( .I(n3516), .Z(n3515) );
  BUFFD0 U3500 ( .I(n3517), .Z(n3516) );
  BUFFD0 U3501 ( .I(n3518), .Z(n3517) );
  BUFFD0 U3502 ( .I(n3519), .Z(n3518) );
  BUFFD0 U3503 ( .I(n3520), .Z(n3519) );
  BUFFD0 U3504 ( .I(n3521), .Z(n3520) );
  BUFFD0 U3505 ( .I(n3522), .Z(n3521) );
  BUFFD0 U3506 ( .I(n3523), .Z(n3522) );
  BUFFD0 U3507 ( .I(n3524), .Z(n3523) );
  BUFFD0 U3508 ( .I(n3525), .Z(n3524) );
  BUFFD0 U3509 ( .I(n3526), .Z(n3525) );
  BUFFD0 U3510 ( .I(n3527), .Z(n3526) );
  BUFFD0 U3511 ( .I(n3528), .Z(n3527) );
  BUFFD0 U3512 ( .I(n3529), .Z(n3528) );
  BUFFD0 U3513 ( .I(n3530), .Z(n3529) );
  BUFFD0 U3514 ( .I(n3531), .Z(n3530) );
  BUFFD0 U3515 ( .I(n3532), .Z(n3531) );
  BUFFD0 U3516 ( .I(n3533), .Z(n3532) );
  BUFFD0 U3517 ( .I(n3534), .Z(n3533) );
  BUFFD0 U3518 ( .I(n3535), .Z(n3534) );
  BUFFD0 U3519 ( .I(n3536), .Z(n3535) );
  BUFFD0 U3520 ( .I(n3537), .Z(n3536) );
  BUFFD0 U3521 ( .I(n3538), .Z(n3537) );
  BUFFD0 U3522 ( .I(n3539), .Z(n3538) );
  BUFFD0 U3523 ( .I(n3540), .Z(n3539) );
  BUFFD0 U3524 ( .I(n3541), .Z(n3540) );
  BUFFD0 U3525 ( .I(n3542), .Z(n3541) );
  BUFFD0 U3526 ( .I(n3543), .Z(n3542) );
  BUFFD0 U3527 ( .I(n3544), .Z(n3543) );
  BUFFD0 U3528 ( .I(n3545), .Z(n3544) );
  BUFFD0 U3529 ( .I(n3546), .Z(n3545) );
  BUFFD0 U3530 ( .I(n3548), .Z(n3546) );
  BUFFD0 U3531 ( .I(N78), .Z(n3547) );
  BUFFD0 U3532 ( .I(n3549), .Z(n3548) );
  BUFFD0 U3533 ( .I(n3489), .Z(n3549) );
  BUFFD0 U3534 ( .I(n3554), .Z(n3550) );
  BUFFD0 U3535 ( .I(n3799), .Z(n3551) );
  BUFFD0 U3536 ( .I(n3551), .Z(n3552) );
  BUFFD0 U3537 ( .I(n3552), .Z(n3553) );
  BUFFD0 U3538 ( .I(n3555), .Z(n3554) );
  BUFFD0 U3539 ( .I(n3556), .Z(n3555) );
  BUFFD0 U3540 ( .I(n3557), .Z(n3556) );
  BUFFD0 U3541 ( .I(n3558), .Z(n3557) );
  BUFFD0 U3542 ( .I(n3559), .Z(n3558) );
  BUFFD0 U3543 ( .I(n3560), .Z(n3559) );
  BUFFD0 U3544 ( .I(n3561), .Z(n3560) );
  BUFFD0 U3545 ( .I(n3562), .Z(n3561) );
  BUFFD0 U3546 ( .I(n3563), .Z(n3562) );
  BUFFD0 U3547 ( .I(n3564), .Z(n3563) );
  BUFFD0 U3548 ( .I(n3565), .Z(n3564) );
  BUFFD0 U3549 ( .I(n3566), .Z(n3565) );
  BUFFD0 U3550 ( .I(n3567), .Z(n3566) );
  BUFFD0 U3551 ( .I(n3568), .Z(n3567) );
  BUFFD0 U3552 ( .I(n3569), .Z(n3568) );
  BUFFD0 U3553 ( .I(n3570), .Z(n3569) );
  BUFFD0 U3554 ( .I(n3571), .Z(n3570) );
  BUFFD0 U3555 ( .I(n3572), .Z(n3571) );
  BUFFD0 U3556 ( .I(n3573), .Z(n3572) );
  BUFFD0 U3557 ( .I(n3574), .Z(n3573) );
  BUFFD0 U3558 ( .I(n3575), .Z(n3574) );
  BUFFD0 U3559 ( .I(n3576), .Z(n3575) );
  BUFFD0 U3560 ( .I(n3577), .Z(n3576) );
  BUFFD0 U3561 ( .I(n3578), .Z(n3577) );
  BUFFD0 U3562 ( .I(n3579), .Z(n3578) );
  BUFFD0 U3563 ( .I(n3580), .Z(n3579) );
  BUFFD0 U3564 ( .I(n3581), .Z(n3580) );
  BUFFD0 U3565 ( .I(n3582), .Z(n3581) );
  BUFFD0 U3566 ( .I(n3583), .Z(n3582) );
  BUFFD0 U3567 ( .I(n3584), .Z(n3583) );
  BUFFD0 U3568 ( .I(n3585), .Z(n3584) );
  BUFFD0 U3569 ( .I(n3586), .Z(n3585) );
  BUFFD0 U3570 ( .I(n3587), .Z(n3586) );
  BUFFD0 U3571 ( .I(n3588), .Z(n3587) );
  BUFFD0 U3572 ( .I(n3589), .Z(n3588) );
  BUFFD0 U3573 ( .I(n3590), .Z(n3589) );
  BUFFD0 U3574 ( .I(n3591), .Z(n3590) );
  BUFFD0 U3575 ( .I(n3592), .Z(n3591) );
  BUFFD0 U3576 ( .I(n3593), .Z(n3592) );
  BUFFD0 U3577 ( .I(n3594), .Z(n3593) );
  BUFFD0 U3578 ( .I(n3595), .Z(n3594) );
  BUFFD0 U3579 ( .I(n3596), .Z(n3595) );
  BUFFD0 U3580 ( .I(n3597), .Z(n3596) );
  BUFFD0 U3581 ( .I(n3598), .Z(n3597) );
  BUFFD0 U3582 ( .I(n3599), .Z(n3598) );
  BUFFD0 U3583 ( .I(n3600), .Z(n3599) );
  BUFFD0 U3584 ( .I(n3601), .Z(n3600) );
  BUFFD0 U3585 ( .I(n3602), .Z(n3601) );
  BUFFD0 U3586 ( .I(n3603), .Z(n3602) );
  BUFFD0 U3587 ( .I(n3604), .Z(n3603) );
  BUFFD0 U3588 ( .I(n3605), .Z(n3604) );
  BUFFD0 U3589 ( .I(n3606), .Z(n3605) );
  BUFFD0 U3590 ( .I(n3607), .Z(n3606) );
  BUFFD0 U3591 ( .I(n3608), .Z(n3607) );
  BUFFD0 U3592 ( .I(n3609), .Z(n3608) );
  BUFFD0 U3593 ( .I(n3553), .Z(n3609) );
  MUX3ND1 U3594 ( .I0(n3958), .I1(n3959), .I2(n3867), .S0(n4641), .S1(n4352), 
        .ZN(N80) );
  BUFFD0 U3595 ( .I(n3800), .Z(n3610) );
  BUFFD0 U3596 ( .I(n3610), .Z(n3611) );
  BUFFD0 U3597 ( .I(n3611), .Z(n3612) );
  BUFFD0 U3598 ( .I(n3612), .Z(n3613) );
  BUFFD0 U3599 ( .I(n3615), .Z(n3614) );
  BUFFD0 U3600 ( .I(n3616), .Z(n3615) );
  BUFFD0 U3601 ( .I(n3617), .Z(n3616) );
  BUFFD0 U3602 ( .I(n3618), .Z(n3617) );
  BUFFD0 U3603 ( .I(n3619), .Z(n3618) );
  BUFFD0 U3604 ( .I(n3620), .Z(n3619) );
  BUFFD0 U3605 ( .I(n3621), .Z(n3620) );
  BUFFD0 U3606 ( .I(n3622), .Z(n3621) );
  BUFFD0 U3607 ( .I(n3623), .Z(n3622) );
  BUFFD0 U3608 ( .I(n3624), .Z(n3623) );
  BUFFD0 U3609 ( .I(n3625), .Z(n3624) );
  BUFFD0 U3610 ( .I(n3626), .Z(n3625) );
  BUFFD0 U3611 ( .I(n3627), .Z(n3626) );
  BUFFD0 U3612 ( .I(n3628), .Z(n3627) );
  BUFFD0 U3613 ( .I(n3629), .Z(n3628) );
  BUFFD0 U3614 ( .I(n3630), .Z(n3629) );
  BUFFD0 U3615 ( .I(n3631), .Z(n3630) );
  BUFFD0 U3616 ( .I(n3632), .Z(n3631) );
  BUFFD0 U3617 ( .I(n3633), .Z(n3632) );
  BUFFD0 U3618 ( .I(n3634), .Z(n3633) );
  BUFFD0 U3619 ( .I(n3635), .Z(n3634) );
  BUFFD0 U3620 ( .I(n3636), .Z(n3635) );
  BUFFD0 U3621 ( .I(n3637), .Z(n3636) );
  BUFFD0 U3622 ( .I(n3638), .Z(n3637) );
  BUFFD0 U3623 ( .I(n3639), .Z(n3638) );
  BUFFD0 U3624 ( .I(n3640), .Z(n3639) );
  BUFFD0 U3625 ( .I(n3641), .Z(n3640) );
  BUFFD0 U3626 ( .I(n3642), .Z(n3641) );
  BUFFD0 U3627 ( .I(n3643), .Z(n3642) );
  BUFFD0 U3628 ( .I(n3644), .Z(n3643) );
  BUFFD0 U3629 ( .I(n3645), .Z(n3644) );
  BUFFD0 U3630 ( .I(n3646), .Z(n3645) );
  BUFFD0 U3631 ( .I(n3647), .Z(n3646) );
  BUFFD0 U3632 ( .I(n3648), .Z(n3647) );
  BUFFD0 U3633 ( .I(n3649), .Z(n3648) );
  BUFFD0 U3634 ( .I(n3650), .Z(n3649) );
  BUFFD0 U3635 ( .I(n3651), .Z(n3650) );
  BUFFD0 U3636 ( .I(n3652), .Z(n3651) );
  BUFFD0 U3637 ( .I(n3653), .Z(n3652) );
  BUFFD0 U3638 ( .I(n3654), .Z(n3653) );
  BUFFD0 U3639 ( .I(n3655), .Z(n3654) );
  BUFFD0 U3640 ( .I(n3656), .Z(n3655) );
  BUFFD0 U3641 ( .I(n3657), .Z(n3656) );
  BUFFD0 U3642 ( .I(n3658), .Z(n3657) );
  BUFFD0 U3643 ( .I(n3659), .Z(n3658) );
  BUFFD0 U3644 ( .I(n3660), .Z(n3659) );
  BUFFD0 U3645 ( .I(n3661), .Z(n3660) );
  BUFFD0 U3646 ( .I(n3662), .Z(n3661) );
  BUFFD0 U3647 ( .I(n3663), .Z(n3662) );
  BUFFD0 U3648 ( .I(n3664), .Z(n3663) );
  BUFFD0 U3649 ( .I(n3665), .Z(n3664) );
  BUFFD0 U3650 ( .I(n3666), .Z(n3665) );
  BUFFD0 U3651 ( .I(n3667), .Z(n3666) );
  BUFFD0 U3652 ( .I(n3668), .Z(n3667) );
  BUFFD0 U3653 ( .I(n3669), .Z(n3668) );
  BUFFD0 U3654 ( .I(n3670), .Z(n3669) );
  BUFFD0 U3655 ( .I(n3671), .Z(n3670) );
  BUFFD0 U3656 ( .I(n3672), .Z(n3671) );
  BUFFD0 U3657 ( .I(n3613), .Z(n3672) );
  MUX3ND1 U3658 ( .I0(n3945), .I1(n3946), .I2(n3868), .S0(n4641), .S1(n4352), 
        .ZN(N81) );
  BUFFD0 U3659 ( .I(n3801), .Z(n3673) );
  BUFFD0 U3660 ( .I(n3673), .Z(n3674) );
  BUFFD0 U3661 ( .I(n3674), .Z(n3675) );
  BUFFD0 U3662 ( .I(n3675), .Z(n3676) );
  BUFFD0 U3663 ( .I(n3678), .Z(n3677) );
  BUFFD0 U3664 ( .I(n3679), .Z(n3678) );
  BUFFD0 U3665 ( .I(n3680), .Z(n3679) );
  BUFFD0 U3666 ( .I(n3681), .Z(n3680) );
  BUFFD0 U3667 ( .I(n3682), .Z(n3681) );
  BUFFD0 U3668 ( .I(n3683), .Z(n3682) );
  BUFFD0 U3669 ( .I(n3684), .Z(n3683) );
  BUFFD0 U3670 ( .I(n3685), .Z(n3684) );
  BUFFD0 U3671 ( .I(n3686), .Z(n3685) );
  BUFFD0 U3672 ( .I(n3687), .Z(n3686) );
  BUFFD0 U3673 ( .I(n3688), .Z(n3687) );
  BUFFD0 U3674 ( .I(n3689), .Z(n3688) );
  BUFFD0 U3675 ( .I(n3690), .Z(n3689) );
  BUFFD0 U3676 ( .I(n3691), .Z(n3690) );
  BUFFD0 U3677 ( .I(n3692), .Z(n3691) );
  BUFFD0 U3678 ( .I(n3693), .Z(n3692) );
  BUFFD0 U3679 ( .I(n3694), .Z(n3693) );
  BUFFD0 U3680 ( .I(n3695), .Z(n3694) );
  BUFFD0 U3681 ( .I(n3696), .Z(n3695) );
  BUFFD0 U3682 ( .I(n3697), .Z(n3696) );
  BUFFD0 U3683 ( .I(n3698), .Z(n3697) );
  BUFFD0 U3684 ( .I(n3699), .Z(n3698) );
  BUFFD0 U3685 ( .I(n3700), .Z(n3699) );
  BUFFD0 U3686 ( .I(n3701), .Z(n3700) );
  BUFFD0 U3687 ( .I(n3702), .Z(n3701) );
  BUFFD0 U3688 ( .I(n3703), .Z(n3702) );
  BUFFD0 U3689 ( .I(n3704), .Z(n3703) );
  BUFFD0 U3690 ( .I(n3705), .Z(n3704) );
  BUFFD0 U3691 ( .I(n3706), .Z(n3705) );
  BUFFD0 U3692 ( .I(n3707), .Z(n3706) );
  BUFFD0 U3693 ( .I(n3708), .Z(n3707) );
  BUFFD0 U3694 ( .I(n3709), .Z(n3708) );
  BUFFD0 U3695 ( .I(n3710), .Z(n3709) );
  BUFFD0 U3696 ( .I(n3711), .Z(n3710) );
  BUFFD0 U3697 ( .I(n3712), .Z(n3711) );
  BUFFD0 U3698 ( .I(n3713), .Z(n3712) );
  BUFFD0 U3699 ( .I(n3714), .Z(n3713) );
  BUFFD0 U3700 ( .I(n3715), .Z(n3714) );
  BUFFD0 U3701 ( .I(n3716), .Z(n3715) );
  BUFFD0 U3702 ( .I(n3717), .Z(n3716) );
  BUFFD0 U3703 ( .I(n3718), .Z(n3717) );
  BUFFD0 U3704 ( .I(n3719), .Z(n3718) );
  BUFFD0 U3705 ( .I(n3720), .Z(n3719) );
  BUFFD0 U3706 ( .I(n3721), .Z(n3720) );
  BUFFD0 U3707 ( .I(n3722), .Z(n3721) );
  BUFFD0 U3708 ( .I(n3723), .Z(n3722) );
  BUFFD0 U3709 ( .I(n3724), .Z(n3723) );
  BUFFD0 U3710 ( .I(n3725), .Z(n3724) );
  BUFFD0 U3711 ( .I(n3726), .Z(n3725) );
  BUFFD0 U3712 ( .I(n3727), .Z(n3726) );
  BUFFD0 U3713 ( .I(n3728), .Z(n3727) );
  BUFFD0 U3714 ( .I(n3729), .Z(n3728) );
  BUFFD0 U3715 ( .I(n3730), .Z(n3729) );
  BUFFD0 U3716 ( .I(n3731), .Z(n3730) );
  BUFFD0 U3717 ( .I(n3732), .Z(n3731) );
  BUFFD0 U3718 ( .I(n3733), .Z(n3732) );
  BUFFD0 U3719 ( .I(n3734), .Z(n3733) );
  BUFFD0 U3720 ( .I(n3676), .Z(n3734) );
  BUFFD0 U3721 ( .I(n3740), .Z(n3735) );
  BUFFD0 U3722 ( .I(n3819), .Z(n3736) );
  BUFFD0 U3723 ( .I(n3736), .Z(n3737) );
  BUFFD0 U3724 ( .I(n3737), .Z(n3738) );
  BUFFD0 U3725 ( .I(n3738), .Z(n3739) );
  BUFFD0 U3726 ( .I(n3741), .Z(n3740) );
  BUFFD0 U3727 ( .I(n3742), .Z(n3741) );
  BUFFD0 U3728 ( .I(n3743), .Z(n3742) );
  BUFFD0 U3729 ( .I(n3744), .Z(n3743) );
  BUFFD0 U3730 ( .I(n3745), .Z(n3744) );
  BUFFD0 U3731 ( .I(n3746), .Z(n3745) );
  BUFFD0 U3732 ( .I(n3747), .Z(n3746) );
  BUFFD0 U3733 ( .I(n3748), .Z(n3747) );
  BUFFD0 U3734 ( .I(n3749), .Z(n3748) );
  BUFFD0 U3735 ( .I(n3750), .Z(n3749) );
  BUFFD0 U3736 ( .I(n3751), .Z(n3750) );
  BUFFD0 U3737 ( .I(n3752), .Z(n3751) );
  BUFFD0 U3738 ( .I(n3753), .Z(n3752) );
  BUFFD0 U3739 ( .I(n3754), .Z(n3753) );
  BUFFD0 U3740 ( .I(n3755), .Z(n3754) );
  BUFFD0 U3741 ( .I(n3756), .Z(n3755) );
  BUFFD0 U3742 ( .I(n3757), .Z(n3756) );
  BUFFD0 U3743 ( .I(n3758), .Z(n3757) );
  BUFFD0 U3744 ( .I(n3759), .Z(n3758) );
  BUFFD0 U3745 ( .I(n3760), .Z(n3759) );
  BUFFD0 U3746 ( .I(n3761), .Z(n3760) );
  BUFFD0 U3747 ( .I(n3762), .Z(n3761) );
  BUFFD0 U3748 ( .I(n3763), .Z(n3762) );
  BUFFD0 U3749 ( .I(n3764), .Z(n3763) );
  BUFFD0 U3750 ( .I(n3765), .Z(n3764) );
  BUFFD0 U3751 ( .I(n3766), .Z(n3765) );
  BUFFD0 U3752 ( .I(n3767), .Z(n3766) );
  BUFFD0 U3753 ( .I(n3768), .Z(n3767) );
  BUFFD0 U3754 ( .I(n3769), .Z(n3768) );
  BUFFD0 U3755 ( .I(n3770), .Z(n3769) );
  BUFFD0 U3756 ( .I(n3771), .Z(n3770) );
  BUFFD0 U3757 ( .I(n3772), .Z(n3771) );
  BUFFD0 U3758 ( .I(n3773), .Z(n3772) );
  BUFFD0 U3759 ( .I(n3774), .Z(n3773) );
  BUFFD0 U3760 ( .I(n3775), .Z(n3774) );
  BUFFD0 U3761 ( .I(n3776), .Z(n3775) );
  BUFFD0 U3762 ( .I(n3777), .Z(n3776) );
  BUFFD0 U3763 ( .I(n3778), .Z(n3777) );
  BUFFD0 U3764 ( .I(n3779), .Z(n3778) );
  BUFFD0 U3765 ( .I(n3780), .Z(n3779) );
  BUFFD0 U3766 ( .I(n3781), .Z(n3780) );
  BUFFD0 U3767 ( .I(n3782), .Z(n3781) );
  BUFFD0 U3768 ( .I(n3783), .Z(n3782) );
  BUFFD0 U3769 ( .I(n3784), .Z(n3783) );
  BUFFD0 U3770 ( .I(n3785), .Z(n3784) );
  BUFFD0 U3771 ( .I(n3786), .Z(n3785) );
  BUFFD0 U3772 ( .I(n3787), .Z(n3786) );
  BUFFD0 U3773 ( .I(n3788), .Z(n3787) );
  BUFFD0 U3774 ( .I(n3789), .Z(n3788) );
  BUFFD0 U3775 ( .I(n3790), .Z(n3789) );
  BUFFD0 U3776 ( .I(n3791), .Z(n3790) );
  BUFFD0 U3777 ( .I(n3792), .Z(n3791) );
  BUFFD0 U3778 ( .I(n3793), .Z(n3792) );
  BUFFD0 U3779 ( .I(n3794), .Z(n3793) );
  BUFFD0 U3780 ( .I(n3796), .Z(n3794) );
  BUFFD0 U3781 ( .I(N82), .Z(n3795) );
  BUFFD0 U3782 ( .I(n3797), .Z(n3796) );
  BUFFD0 U3783 ( .I(n3739), .Z(n3797) );
  BUFFD0 U3784 ( .I(N75), .Z(n3798) );
  BUFFD0 U3785 ( .I(n3869), .Z(n3799) );
  BUFFD0 U3786 ( .I(N80), .Z(n3800) );
  BUFFD0 U3787 ( .I(N81), .Z(n3801) );
  BUFFD0 U3788 ( .I(n3803), .Z(n3802) );
  BUFFD0 U3789 ( .I(n3804), .Z(n3803) );
  BUFFD0 U3790 ( .I(n3805), .Z(n3804) );
  BUFFD0 U3791 ( .I(n3806), .Z(n3805) );
  BUFFD0 U3792 ( .I(n3807), .Z(n3806) );
  BUFFD0 U3793 ( .I(n3808), .Z(n3807) );
  BUFFD0 U3794 ( .I(n3809), .Z(n3808) );
  BUFFD0 U3795 ( .I(n3810), .Z(n3809) );
  BUFFD0 U3796 ( .I(n3811), .Z(n3810) );
  BUFFD0 U3797 ( .I(n3812), .Z(n3811) );
  BUFFD0 U3798 ( .I(n3813), .Z(n3812) );
  BUFFD0 U3799 ( .I(n3814), .Z(n3813) );
  BUFFD0 U3800 ( .I(n3815), .Z(n3814) );
  BUFFD0 U3801 ( .I(n3816), .Z(n3815) );
  BUFFD0 U3802 ( .I(n3817), .Z(n3816) );
  BUFFD0 U3803 ( .I(n3822), .Z(n3817) );
  BUFFD0 U3804 ( .I(n3866), .Z(n3818) );
  BUFFD0 U3805 ( .I(n3795), .Z(n3819) );
  BUFFD0 U3806 ( .I(n3871), .Z(n3820) );
  BUFFD0 U3807 ( .I(n3547), .Z(n3821) );
  BUFFD0 U3808 ( .I(n3823), .Z(n3822) );
  BUFFD0 U3809 ( .I(n3824), .Z(n3823) );
  BUFFD0 U3810 ( .I(n3825), .Z(n3824) );
  BUFFD0 U3811 ( .I(n3826), .Z(n3825) );
  BUFFD0 U3812 ( .I(n3827), .Z(n3826) );
  BUFFD0 U3813 ( .I(n3828), .Z(n3827) );
  BUFFD0 U3814 ( .I(n3829), .Z(n3828) );
  BUFFD0 U3815 ( .I(n3830), .Z(n3829) );
  BUFFD0 U3816 ( .I(n3831), .Z(n3830) );
  BUFFD0 U3817 ( .I(n3832), .Z(n3831) );
  BUFFD0 U3818 ( .I(n3833), .Z(n3832) );
  BUFFD0 U3819 ( .I(n3834), .Z(n3833) );
  BUFFD0 U3820 ( .I(n3835), .Z(n3834) );
  BUFFD0 U3821 ( .I(n3836), .Z(n3835) );
  BUFFD0 U3822 ( .I(n3837), .Z(n3836) );
  BUFFD0 U3823 ( .I(n3838), .Z(n3837) );
  BUFFD0 U3824 ( .I(n3839), .Z(n3838) );
  BUFFD0 U3825 ( .I(n3840), .Z(n3839) );
  BUFFD0 U3826 ( .I(n3841), .Z(n3840) );
  BUFFD0 U3827 ( .I(n3842), .Z(n3841) );
  BUFFD0 U3828 ( .I(n3843), .Z(n3842) );
  BUFFD0 U3829 ( .I(n3844), .Z(n3843) );
  BUFFD0 U3830 ( .I(n3845), .Z(n3844) );
  BUFFD0 U3831 ( .I(n3846), .Z(n3845) );
  BUFFD0 U3832 ( .I(n3847), .Z(n3846) );
  BUFFD0 U3833 ( .I(n3848), .Z(n3847) );
  BUFFD0 U3834 ( .I(n3849), .Z(n3848) );
  BUFFD0 U3835 ( .I(n3850), .Z(n3849) );
  BUFFD0 U3836 ( .I(n3851), .Z(n3850) );
  BUFFD0 U3837 ( .I(n3852), .Z(n3851) );
  BUFFD0 U3838 ( .I(n3853), .Z(n3852) );
  BUFFD0 U3839 ( .I(n3854), .Z(n3853) );
  BUFFD0 U3840 ( .I(n3855), .Z(n3854) );
  BUFFD0 U3841 ( .I(n3856), .Z(n3855) );
  BUFFD0 U3842 ( .I(n3857), .Z(n3856) );
  BUFFD0 U3843 ( .I(n3858), .Z(n3857) );
  BUFFD0 U3844 ( .I(n3859), .Z(n3858) );
  BUFFD0 U3845 ( .I(n3860), .Z(n3859) );
  BUFFD0 U3846 ( .I(n3861), .Z(n3860) );
  BUFFD0 U3847 ( .I(n3876), .Z(n3861) );
  BUFFD0 U3848 ( .I(n3873), .Z(n3862) );
  BUFFD0 U3849 ( .I(n4025), .Z(n3863) );
  BUFFD0 U3850 ( .I(n3875), .Z(n3864) );
  BUFFD0 U3851 ( .I(n4064), .Z(n3865) );
  BUFFD0 U3852 ( .I(N76), .Z(n3866) );
  BUFFD0 U3853 ( .I(n3960), .Z(n3867) );
  BUFFD0 U3854 ( .I(n3947), .Z(n3868) );
  BUFFD0 U3855 ( .I(n3878), .Z(n3869) );
  BUFFD0 U3856 ( .I(n3934), .Z(n3870) );
  BUFFD0 U3857 ( .I(N77), .Z(n3871) );
  BUFFD0 U3858 ( .I(n3986), .Z(n3872) );
  BUFFD0 U3859 ( .I(n3879), .Z(n3873) );
  BUFFD0 U3860 ( .I(n4012), .Z(n3874) );
  BUFFD0 U3861 ( .I(n3880), .Z(n3875) );
  BUFFD0 U3862 ( .I(N83), .Z(n3876) );
  BUFFD0 U3863 ( .I(n3999), .Z(n3877) );
  BUFFD0 U3864 ( .I(n3881), .Z(n3878) );
  BUFFD0 U3865 ( .I(N73), .Z(n3879) );
  BUFFD0 U3866 ( .I(n3883), .Z(n3880) );
  BUFFD0 U3867 ( .I(n3884), .Z(n3881) );
  BUFFD0 U3868 ( .I(n4051), .Z(n3882) );
  BUFFD0 U3869 ( .I(N74), .Z(n3883) );
  BUFFD0 U3870 ( .I(N79), .Z(n3884) );
  BUFFD0 U3871 ( .I(n4038), .Z(n3885) );
  BUFFD0 U3872 ( .I(n3973), .Z(n3886) );
  BUFFD0 U3873 ( .I(n3888), .Z(n3887) );
  BUFFD0 U3874 ( .I(n4636), .Z(n3888) );
  CKAN2D0 U3875 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U3876 ( .I(N48), .ZN(n4351) );
  INVD1 U3877 ( .I(DataI[17]), .ZN(n4687) );
  INVD1 U3878 ( .I(DataI[21]), .ZN(n4697) );
  INVD1 U3879 ( .I(DataI[22]), .ZN(n4699) );
  INVD1 U3880 ( .I(DataI[24]), .ZN(n4705) );
  INVD1 U3881 ( .I(DataI[25]), .ZN(n4707) );
  INVD1 U3882 ( .I(DataI[26]), .ZN(n4709) );
  INVD1 U3883 ( .I(DataI[27]), .ZN(n4712) );
  INVD1 U3884 ( .I(DataI[28]), .ZN(n4715) );
  INVD1 U3885 ( .I(DataI[29]), .ZN(n4717) );
  INVD1 U3886 ( .I(DataI[30]), .ZN(n4719) );
  INVD1 U3887 ( .I(DataI[31]), .ZN(n4722) );
  INVD1 U3888 ( .I(DataI[0]), .ZN(n4643) );
  INVD1 U3889 ( .I(DataI[1]), .ZN(n4646) );
  INVD1 U3890 ( .I(DataI[2]), .ZN(n4648) );
  INVD1 U3891 ( .I(DataI[3]), .ZN(n4651) );
  INVD1 U3892 ( .I(DataI[4]), .ZN(n4654) );
  INVD1 U3893 ( .I(DataI[5]), .ZN(n4656) );
  INVD1 U3894 ( .I(DataI[6]), .ZN(n4659) );
  INVD1 U3895 ( .I(DataI[7]), .ZN(n4661) );
  INVD1 U3896 ( .I(DataI[8]), .ZN(n4663) );
  INVD1 U3897 ( .I(DataI[9]), .ZN(n4666) );
  INVD1 U3898 ( .I(DataI[10]), .ZN(n4669) );
  INVD1 U3899 ( .I(DataI[11]), .ZN(n4672) );
  INVD1 U3900 ( .I(DataI[12]), .ZN(n4674) );
  INVD1 U3901 ( .I(DataI[13]), .ZN(n4677) );
  INVD1 U3902 ( .I(DataI[14]), .ZN(n4679) );
  INVD1 U3903 ( .I(DataI[15]), .ZN(n4681) );
  INVD1 U3904 ( .I(DataI[16]), .ZN(n4684) );
  INVD1 U3905 ( .I(DataI[18]), .ZN(n4690) );
  INVD1 U3906 ( .I(DataI[19]), .ZN(n4692) );
  INVD1 U3907 ( .I(DataI[20]), .ZN(n4695) );
  INVD1 U3908 ( .I(DataI[23]), .ZN(n4702) );
  BUFFD1 U3909 ( .I(n4501), .Z(n4424) );
  BUFFD1 U3910 ( .I(n4501), .Z(n4425) );
  BUFFD1 U3911 ( .I(n4501), .Z(n4426) );
  BUFFD1 U3912 ( .I(n4501), .Z(n4427) );
  BUFFD1 U3913 ( .I(n4500), .Z(n4428) );
  BUFFD1 U3914 ( .I(n4500), .Z(n4429) );
  BUFFD1 U3915 ( .I(n4500), .Z(n4430) );
  BUFFD1 U3916 ( .I(n4500), .Z(n4431) );
  BUFFD1 U3917 ( .I(n4499), .Z(n4432) );
  BUFFD1 U3918 ( .I(n4499), .Z(n4433) );
  BUFFD1 U3919 ( .I(n4499), .Z(n4434) );
  BUFFD1 U3920 ( .I(n4499), .Z(n4435) );
  BUFFD1 U3921 ( .I(n4496), .Z(n4436) );
  BUFFD1 U3922 ( .I(n4511), .Z(n4437) );
  BUFFD1 U3923 ( .I(n4499), .Z(n4438) );
  BUFFD1 U3924 ( .I(n4498), .Z(n4439) );
  BUFFD1 U3925 ( .I(n4498), .Z(n4440) );
  BUFFD1 U3926 ( .I(n4498), .Z(n4441) );
  BUFFD1 U3927 ( .I(n4498), .Z(n4442) );
  BUFFD1 U3928 ( .I(n4494), .Z(n4443) );
  BUFFD1 U3929 ( .I(n4511), .Z(n4444) );
  BUFFD1 U3930 ( .I(n4498), .Z(n4445) );
  BUFFD1 U3931 ( .I(n108), .Z(n4446) );
  BUFFD1 U3932 ( .I(n4497), .Z(n4447) );
  BUFFD1 U3933 ( .I(n4497), .Z(n4448) );
  BUFFD1 U3934 ( .I(n4497), .Z(n4449) );
  BUFFD1 U3935 ( .I(n4497), .Z(n4450) );
  BUFFD1 U3936 ( .I(n4496), .Z(n4451) );
  BUFFD1 U3937 ( .I(n4496), .Z(n4452) );
  BUFFD1 U3938 ( .I(n4496), .Z(n4453) );
  BUFFD1 U3939 ( .I(n4496), .Z(n4454) );
  BUFFD1 U3940 ( .I(n4494), .Z(n4455) );
  BUFFD1 U3941 ( .I(n4494), .Z(n4456) );
  BUFFD1 U3942 ( .I(n4494), .Z(n4457) );
  BUFFD1 U3943 ( .I(n4494), .Z(n4458) );
  BUFFD1 U3944 ( .I(n4495), .Z(n4459) );
  BUFFD1 U3945 ( .I(n4495), .Z(n4460) );
  BUFFD1 U3946 ( .I(n4495), .Z(n4461) );
  BUFFD1 U3947 ( .I(n4495), .Z(n4462) );
  BUFFD1 U3948 ( .I(n4494), .Z(n4463) );
  BUFFD1 U3949 ( .I(n4494), .Z(n4464) );
  BUFFD1 U3950 ( .I(n4494), .Z(n4465) );
  BUFFD1 U3951 ( .I(n4494), .Z(n4466) );
  BUFFD1 U3952 ( .I(n4493), .Z(n4467) );
  BUFFD1 U3953 ( .I(n4492), .Z(n4468) );
  BUFFD1 U3954 ( .I(n4507), .Z(n4469) );
  BUFFD1 U3955 ( .I(n4506), .Z(n4470) );
  BUFFD1 U3956 ( .I(n4493), .Z(n4471) );
  BUFFD1 U3957 ( .I(n4493), .Z(n4472) );
  BUFFD1 U3958 ( .I(n4493), .Z(n4473) );
  BUFFD1 U3959 ( .I(n4493), .Z(n4474) );
  BUFFD1 U3960 ( .I(n4492), .Z(n4475) );
  BUFFD1 U3961 ( .I(n4492), .Z(n4476) );
  BUFFD1 U3962 ( .I(n4492), .Z(n4477) );
  BUFFD1 U3963 ( .I(n4492), .Z(n4478) );
  BUFFD1 U3964 ( .I(n4492), .Z(n4479) );
  BUFFD1 U3965 ( .I(n4493), .Z(n4480) );
  BUFFD1 U3966 ( .I(n4492), .Z(n4481) );
  BUFFD1 U3967 ( .I(n4506), .Z(n4482) );
  BUFFD1 U3968 ( .I(n4506), .Z(n4483) );
  BUFFD1 U3969 ( .I(n4506), .Z(n4484) );
  BUFFD1 U3970 ( .I(n4506), .Z(n4485) );
  BUFFD1 U3971 ( .I(n4506), .Z(n4486) );
  BUFFD1 U3972 ( .I(n4499), .Z(n4487) );
  BUFFD1 U3973 ( .I(n4496), .Z(n4488) );
  BUFFD1 U3974 ( .I(n4496), .Z(n4489) );
  BUFFD1 U3975 ( .I(n4507), .Z(n4400) );
  BUFFD1 U3976 ( .I(n4507), .Z(n4401) );
  BUFFD1 U3977 ( .I(n4507), .Z(n4402) );
  BUFFD1 U3978 ( .I(n4507), .Z(n4403) );
  BUFFD1 U3979 ( .I(n4506), .Z(n4404) );
  BUFFD1 U3980 ( .I(n4506), .Z(n4405) );
  BUFFD1 U3981 ( .I(n4506), .Z(n4406) );
  BUFFD1 U3982 ( .I(n4506), .Z(n4407) );
  BUFFD1 U3983 ( .I(n4505), .Z(n4408) );
  BUFFD1 U3984 ( .I(n4505), .Z(n4409) );
  BUFFD1 U3985 ( .I(n4505), .Z(n4410) );
  BUFFD1 U3986 ( .I(n4505), .Z(n4411) );
  BUFFD1 U3987 ( .I(n4504), .Z(n4412) );
  BUFFD1 U3988 ( .I(n4504), .Z(n4413) );
  BUFFD1 U3989 ( .I(n4504), .Z(n4414) );
  BUFFD1 U3990 ( .I(n4504), .Z(n4415) );
  BUFFD1 U3991 ( .I(n4503), .Z(n4416) );
  BUFFD1 U3992 ( .I(n4503), .Z(n4417) );
  BUFFD1 U3993 ( .I(n4503), .Z(n4418) );
  BUFFD1 U3994 ( .I(n4503), .Z(n4419) );
  BUFFD1 U3995 ( .I(n4502), .Z(n4420) );
  BUFFD1 U3996 ( .I(n4502), .Z(n4421) );
  BUFFD1 U3997 ( .I(n4502), .Z(n4422) );
  BUFFD1 U3998 ( .I(n4502), .Z(n4423) );
  BUFFD1 U3999 ( .I(n4510), .Z(n4501) );
  BUFFD1 U4000 ( .I(n4510), .Z(n4500) );
  BUFFD1 U4001 ( .I(n4511), .Z(n4499) );
  BUFFD1 U4002 ( .I(n4510), .Z(n4498) );
  BUFFD1 U4003 ( .I(n4496), .Z(n4497) );
  BUFFD1 U4004 ( .I(n108), .Z(n4496) );
  BUFFD1 U4005 ( .I(n4509), .Z(n4495) );
  BUFFD1 U4006 ( .I(n4398), .Z(n4494) );
  BUFFD1 U4007 ( .I(n4492), .Z(n4493) );
  BUFFD1 U4008 ( .I(n108), .Z(n4492) );
  BUFFD1 U4009 ( .I(n4629), .Z(n4611) );
  BUFFD1 U4010 ( .I(n4612), .Z(n4610) );
  BUFFD1 U4011 ( .I(n4613), .Z(n4609) );
  BUFFD1 U4012 ( .I(n4613), .Z(n4608) );
  BUFFD1 U4013 ( .I(n4614), .Z(n4607) );
  BUFFD1 U4014 ( .I(n4614), .Z(n4606) );
  BUFFD1 U4015 ( .I(n4615), .Z(n4605) );
  BUFFD1 U4016 ( .I(n4615), .Z(n4604) );
  BUFFD1 U4017 ( .I(n4616), .Z(n4603) );
  BUFFD1 U4018 ( .I(n4616), .Z(n4602) );
  BUFFD1 U4019 ( .I(n4617), .Z(n4601) );
  BUFFD1 U4020 ( .I(n4617), .Z(n4600) );
  BUFFD1 U4021 ( .I(n4618), .Z(n4599) );
  BUFFD1 U4022 ( .I(n4618), .Z(n4598) );
  BUFFD1 U4023 ( .I(n4619), .Z(n4597) );
  BUFFD1 U4024 ( .I(n4619), .Z(n4596) );
  BUFFD1 U4025 ( .I(n4620), .Z(n4595) );
  BUFFD1 U4026 ( .I(n4620), .Z(n4594) );
  BUFFD1 U4027 ( .I(n4621), .Z(n4593) );
  BUFFD1 U4028 ( .I(n4621), .Z(n4592) );
  BUFFD1 U4029 ( .I(n4622), .Z(n4591) );
  BUFFD1 U4030 ( .I(n4622), .Z(n4590) );
  BUFFD1 U4031 ( .I(n4623), .Z(n4589) );
  BUFFD1 U4032 ( .I(n4623), .Z(n4588) );
  BUFFD1 U4033 ( .I(n4624), .Z(n4587) );
  BUFFD1 U4034 ( .I(n4624), .Z(n4586) );
  BUFFD1 U4035 ( .I(n4625), .Z(n4585) );
  BUFFD1 U4036 ( .I(n4625), .Z(n4584) );
  BUFFD1 U4037 ( .I(n4626), .Z(n4583) );
  BUFFD1 U4038 ( .I(n4626), .Z(n4582) );
  BUFFD1 U4039 ( .I(n4627), .Z(n4581) );
  BUFFD1 U4040 ( .I(n4627), .Z(n4580) );
  BUFFD1 U4041 ( .I(n4385), .Z(n4389) );
  BUFFD1 U4042 ( .I(n4365), .Z(n4374) );
  BUFFD1 U4043 ( .I(n4365), .Z(n4375) );
  BUFFD1 U4044 ( .I(n4365), .Z(n4376) );
  BUFFD1 U4045 ( .I(n4385), .Z(n4387) );
  BUFFD1 U4046 ( .I(n4385), .Z(n4388) );
  BUFFD1 U4047 ( .I(N44), .Z(n4390) );
  BUFFD1 U4048 ( .I(n4386), .Z(n4391) );
  BUFFD1 U4049 ( .I(n4385), .Z(n4392) );
  BUFFD1 U4050 ( .I(n4384), .Z(n4393) );
  BUFFD1 U4051 ( .I(n4384), .Z(n4394) );
  BUFFD1 U4052 ( .I(n4384), .Z(n4395) );
  BUFFD1 U4053 ( .I(n4383), .Z(n4396) );
  BUFFD1 U4054 ( .I(n4383), .Z(n4397) );
  BUFFD1 U4055 ( .I(n4364), .Z(n4378) );
  BUFFD1 U4056 ( .I(n4364), .Z(n4379) );
  BUFFD1 U4057 ( .I(n4368), .Z(n4381) );
  BUFFD1 U4058 ( .I(n4368), .Z(n4382) );
  BUFFD1 U4059 ( .I(n4366), .Z(n4380) );
  BUFFD1 U4060 ( .I(n4366), .Z(n4372) );
  BUFFD1 U4061 ( .I(n4366), .Z(n4373) );
  BUFFD1 U4062 ( .I(n4364), .Z(n4377) );
  BUFFD1 U4063 ( .I(n4366), .Z(n4371) );
  BUFFD1 U4064 ( .I(n4491), .Z(n4490) );
  BUFFD1 U4065 ( .I(n4508), .Z(n4506) );
  BUFFD1 U4066 ( .I(n4496), .Z(n4505) );
  BUFFD1 U4067 ( .I(n4496), .Z(n4504) );
  BUFFD1 U4068 ( .I(n4509), .Z(n4503) );
  BUFFD1 U4069 ( .I(n4509), .Z(n4502) );
  BUFFD1 U4070 ( .I(n4508), .Z(n4507) );
  BUFFD1 U4071 ( .I(n4398), .Z(n4510) );
  BUFFD1 U4072 ( .I(n4398), .Z(n4511) );
  BUFFD1 U4073 ( .I(n4614), .Z(n4612) );
  BUFFD1 U4074 ( .I(n4632), .Z(n4613) );
  BUFFD1 U4075 ( .I(n4632), .Z(n4614) );
  BUFFD1 U4076 ( .I(n4632), .Z(n4615) );
  BUFFD1 U4077 ( .I(n4631), .Z(n4616) );
  BUFFD1 U4078 ( .I(n4631), .Z(n4617) );
  BUFFD1 U4079 ( .I(n4631), .Z(n4618) );
  BUFFD1 U4080 ( .I(n4630), .Z(n4619) );
  BUFFD1 U4081 ( .I(n4630), .Z(n4620) );
  BUFFD1 U4082 ( .I(n4630), .Z(n4621) );
  BUFFD1 U4083 ( .I(n4629), .Z(n4622) );
  BUFFD1 U4084 ( .I(n4629), .Z(n4623) );
  BUFFD1 U4085 ( .I(n4629), .Z(n4624) );
  BUFFD1 U4086 ( .I(n4628), .Z(n4625) );
  BUFFD1 U4087 ( .I(n4628), .Z(n4626) );
  BUFFD1 U4088 ( .I(n4628), .Z(n4627) );
  INVD1 U4089 ( .I(n4577), .ZN(n4576) );
  BUFFD1 U4090 ( .I(n4367), .Z(n4369) );
  BUFFD1 U4091 ( .I(n4363), .Z(n4365) );
  BUFFD1 U4092 ( .I(N44), .Z(n4385) );
  BUFFD1 U4093 ( .I(N44), .Z(n4386) );
  BUFFD1 U4094 ( .I(n4355), .Z(n4360) );
  BUFFD1 U4095 ( .I(n4355), .Z(n4361) );
  BUFFD1 U4096 ( .I(n4356), .Z(n4359) );
  BUFFD1 U4097 ( .I(n4355), .Z(n4358) );
  BUFFD1 U4098 ( .I(n4355), .Z(n4357) );
  BUFFD1 U4099 ( .I(n4367), .Z(n4370) );
  BUFFD1 U4100 ( .I(n4354), .Z(n4353) );
  BUFFD1 U4101 ( .I(n4386), .Z(n4384) );
  BUFFD1 U4102 ( .I(n4363), .Z(n4366) );
  BUFFD1 U4103 ( .I(n4363), .Z(n4364) );
  BUFFD1 U4104 ( .I(N44), .Z(n4383) );
  BUFFD1 U4105 ( .I(n4367), .Z(n4368) );
  BUFFD1 U4106 ( .I(n4507), .Z(n4491) );
  BUFFD1 U4107 ( .I(n4508), .Z(n4509) );
  BUFFD1 U4108 ( .I(n108), .Z(n4508) );
  BUFFD1 U4109 ( .I(n4399), .Z(n4398) );
  BUFFD1 U4110 ( .I(n4624), .Z(n4632) );
  BUFFD1 U4111 ( .I(n4579), .Z(n4631) );
  BUFFD1 U4112 ( .I(n4579), .Z(n4630) );
  BUFFD1 U4113 ( .I(n4578), .Z(n4629) );
  BUFFD1 U4114 ( .I(n4578), .Z(n4628) );
  INVD1 U4115 ( .I(N85), .ZN(n4577) );
  BUFFD1 U4116 ( .I(n4362), .Z(n4367) );
  BUFFD1 U4117 ( .I(n4640), .Z(n4362) );
  BUFFD1 U4118 ( .I(n4640), .Z(n4363) );
  BUFFD1 U4119 ( .I(N46), .Z(n4356) );
  BUFFD1 U4120 ( .I(n4641), .Z(n4354) );
  BUFFD1 U4121 ( .I(N46), .Z(n4355) );
  INVD1 U4122 ( .I(n4351), .ZN(n4352) );
  BUFFD1 U4123 ( .I(n108), .Z(n4399) );
  BUFFD1 U4124 ( .I(ClockW), .Z(n4579) );
  BUFFD1 U4125 ( .I(ClockW), .Z(n4578) );
  XOR3D1 U4126 ( .A1(n80), .A2(n4667), .A3(n81), .Z(n79) );
  XOR3D1 U4127 ( .A1(n4691), .A2(n4688), .A3(n82), .Z(n81) );
  XOR3D1 U4128 ( .A1(n83), .A2(n4685), .A3(n84), .Z(n82) );
  XOR3D1 U4129 ( .A1(n4655), .A2(n4652), .A3(n76), .Z(n75) );
  XOR3D1 U4130 ( .A1(n77), .A2(n4649), .A3(n78), .Z(n76) );
  XOR3D1 U4131 ( .A1(n4673), .A2(n4670), .A3(n79), .Z(n78) );
  XOR3D1 U4132 ( .A1(n4642), .A2(n74), .A3(n75), .Z(n73) );
  XOR3D1 U4133 ( .A1(N67), .A2(N66), .A3(n92), .Z(n90) );
  XOR3D1 U4134 ( .A1(N65), .A2(n93), .A3(n94), .Z(n92) );
  XOR3D1 U4135 ( .A1(N60), .A2(N59), .A3(n95), .Z(n94) );
  XOR3D1 U4136 ( .A1(n96), .A2(N58), .A3(n97), .Z(n95) );
  XOR3D1 U4137 ( .A1(n3862), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D1 U4138 ( .A1(n3820), .A2(n3818), .A3(n89), .Z(n88) );
  BUFFD1 U4139 ( .I(N45), .Z(n4640) );
  BUFFD1 U4140 ( .I(N47), .Z(n4641) );
  INVD1 U4141 ( .I(n3893), .ZN(n4537) );
  INVD1 U4142 ( .I(n3893), .ZN(n4536) );
  INVD1 U4143 ( .I(n3894), .ZN(n4535) );
  INVD1 U4144 ( .I(n3894), .ZN(n4534) );
  INVD1 U4145 ( .I(n3895), .ZN(n4533) );
  INVD1 U4146 ( .I(n3895), .ZN(n4532) );
  INVD1 U4147 ( .I(n3896), .ZN(n4531) );
  INVD1 U4148 ( .I(n3896), .ZN(n4530) );
  INVD1 U4149 ( .I(n3897), .ZN(n4529) );
  INVD1 U4150 ( .I(n3897), .ZN(n4528) );
  INVD1 U4151 ( .I(n3898), .ZN(n4527) );
  INVD1 U4152 ( .I(n3898), .ZN(n4526) );
  INVD1 U4153 ( .I(n3899), .ZN(n4525) );
  INVD1 U4154 ( .I(n3899), .ZN(n4524) );
  INVD1 U4155 ( .I(n3900), .ZN(n4523) );
  INVD1 U4156 ( .I(n3900), .ZN(n4522) );
  INVD1 U4157 ( .I(n3901), .ZN(n4521) );
  INVD1 U4158 ( .I(n3901), .ZN(n4520) );
  INVD1 U4159 ( .I(n3902), .ZN(n4519) );
  INVD1 U4160 ( .I(n3902), .ZN(n4518) );
  INVD1 U4161 ( .I(n3903), .ZN(n4517) );
  INVD1 U4162 ( .I(n3903), .ZN(n4516) );
  INVD1 U4163 ( .I(n3904), .ZN(n4515) );
  INVD1 U4164 ( .I(n3904), .ZN(n4514) );
  INVD1 U4165 ( .I(n3905), .ZN(n4513) );
  INVD1 U4166 ( .I(n3905), .ZN(n4512) );
  INVD1 U4167 ( .I(n3906), .ZN(n4575) );
  INVD1 U4168 ( .I(n3906), .ZN(n4574) );
  INVD1 U4169 ( .I(n3907), .ZN(n4573) );
  INVD1 U4170 ( .I(n3907), .ZN(n4572) );
  INVD1 U4171 ( .I(n3908), .ZN(n4571) );
  INVD1 U4172 ( .I(n3908), .ZN(n4570) );
  INVD1 U4173 ( .I(n3909), .ZN(n4569) );
  INVD1 U4174 ( .I(n3909), .ZN(n4568) );
  INVD1 U4175 ( .I(n3910), .ZN(n4567) );
  INVD1 U4176 ( .I(n3910), .ZN(n4566) );
  INVD1 U4177 ( .I(n3911), .ZN(n4565) );
  INVD1 U4178 ( .I(n3911), .ZN(n4564) );
  INVD1 U4179 ( .I(n3912), .ZN(n4563) );
  INVD1 U4180 ( .I(n3912), .ZN(n4562) );
  INVD1 U4181 ( .I(n3913), .ZN(n4561) );
  INVD1 U4182 ( .I(n3913), .ZN(n4560) );
  INVD1 U4183 ( .I(n3914), .ZN(n4559) );
  INVD1 U4184 ( .I(n3914), .ZN(n4558) );
  INVD1 U4185 ( .I(n3915), .ZN(n4557) );
  INVD1 U4186 ( .I(n3915), .ZN(n4556) );
  INVD1 U4187 ( .I(n3916), .ZN(n4555) );
  INVD1 U4188 ( .I(n3916), .ZN(n4554) );
  INVD1 U4189 ( .I(n3917), .ZN(n4553) );
  INVD1 U4190 ( .I(n3917), .ZN(n4552) );
  INVD1 U4191 ( .I(n3918), .ZN(n4551) );
  INVD1 U4192 ( .I(n3918), .ZN(n4550) );
  INVD1 U4193 ( .I(n3919), .ZN(n4549) );
  INVD1 U4194 ( .I(n3919), .ZN(n4548) );
  INVD1 U4195 ( .I(n3920), .ZN(n4547) );
  INVD1 U4196 ( .I(n3920), .ZN(n4546) );
  INVD1 U4197 ( .I(n3921), .ZN(n4545) );
  INVD1 U4198 ( .I(n3921), .ZN(n4544) );
  INVD1 U4199 ( .I(n3890), .ZN(n4543) );
  INVD1 U4200 ( .I(n3890), .ZN(n4542) );
  INVD1 U4201 ( .I(n3891), .ZN(n4541) );
  INVD1 U4202 ( .I(n3891), .ZN(n4540) );
  INVD1 U4203 ( .I(n3892), .ZN(n4539) );
  INVD1 U4204 ( .I(n3892), .ZN(n4538) );
  BUFFD1 U4205 ( .I(n4635), .Z(n4638) );
  BUFFD1 U4206 ( .I(n4635), .Z(n4637) );
  BUFFD1 U4207 ( .I(n4636), .Z(n4639) );
  INVD1 U4208 ( .I(n4634), .ZN(n4633) );
  INVD1 U4209 ( .I(Reset), .ZN(n108) );
  INVD1 U4210 ( .I(n1459), .ZN(n4644) );
  INVD1 U4211 ( .I(n1355), .ZN(n4649) );
  INVD1 U4212 ( .I(n1301), .ZN(n4652) );
  INVD1 U4213 ( .I(n985), .ZN(n4667) );
  INVD1 U4214 ( .I(n931), .ZN(n4670) );
  INVD1 U4215 ( .I(n615), .ZN(n4685) );
  INVD1 U4216 ( .I(n561), .ZN(n4688) );
  INVD1 U4217 ( .I(n1251), .ZN(n4655) );
  INVD1 U4218 ( .I(n881), .ZN(n4673) );
  INVD1 U4219 ( .I(n511), .ZN(n4691) );
  INVD1 U4220 ( .I(n1198), .ZN(n4657) );
  INVD1 U4221 ( .I(n1040), .ZN(n4664) );
  INVD1 U4222 ( .I(n828), .ZN(n4675) );
  INVD1 U4223 ( .I(n670), .ZN(n4682) );
  INVD1 U4224 ( .I(n458), .ZN(n4693) );
  INVD1 U4225 ( .I(n300), .ZN(n4700) );
  INVD1 U4226 ( .I(n246), .ZN(n4703) );
  INVD1 U4227 ( .I(n1566), .ZN(n4710) );
  INVD1 U4228 ( .I(n192), .ZN(n4713) );
  INVD1 U4229 ( .I(n11), .ZN(n4720) );
  INVD1 U4230 ( .I(n1198), .ZN(n4658) );
  INVD1 U4231 ( .I(n1040), .ZN(n4665) );
  INVD1 U4232 ( .I(n828), .ZN(n4676) );
  INVD1 U4233 ( .I(n670), .ZN(n4683) );
  INVD1 U4234 ( .I(n458), .ZN(n4694) );
  INVD1 U4235 ( .I(n300), .ZN(n4701) );
  INVD1 U4236 ( .I(n246), .ZN(n4704) );
  INVD1 U4237 ( .I(n1566), .ZN(n4711) );
  INVD1 U4238 ( .I(n192), .ZN(n4714) );
  INVD1 U4239 ( .I(n11), .ZN(n4721) );
  INVD1 U4240 ( .I(n1147), .ZN(n4660) );
  INVD1 U4241 ( .I(n1095), .ZN(n4662) );
  INVD1 U4242 ( .I(n777), .ZN(n4678) );
  INVD1 U4243 ( .I(n725), .ZN(n4680) );
  INVD1 U4244 ( .I(n407), .ZN(n4696) );
  INVD1 U4245 ( .I(n355), .ZN(n4698) );
  INVD1 U4246 ( .I(n1621), .ZN(n4706) );
  INVD1 U4247 ( .I(n1673), .ZN(n4708) );
  INVD1 U4248 ( .I(n141), .ZN(n4716) );
  INVD1 U4249 ( .I(n47), .ZN(n4718) );
  OR2D1 U4250 ( .A1(n69), .A2(n70), .Z(n3890) );
  OR2D1 U4251 ( .A1(n68), .A2(n70), .Z(n3891) );
  OR2D1 U4252 ( .A1(n67), .A2(n70), .Z(n3892) );
  ND3D1 U4253 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  ND3D1 U4254 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U4255 ( .I(AddrW[1]), .ZN(n106) );
  OR2D1 U4256 ( .A1(n70), .A2(n99), .Z(n3893) );
  OR2D1 U4257 ( .A1(n70), .A2(n98), .Z(n3894) );
  OR2D1 U4258 ( .A1(n70), .A2(n85), .Z(n3895) );
  OR2D1 U4259 ( .A1(n70), .A2(n72), .Z(n3896) );
  OR2D1 U4260 ( .A1(n70), .A2(n71), .Z(n3897) );
  OR2D1 U4261 ( .A1(n66), .A2(n69), .Z(n3898) );
  OR2D1 U4262 ( .A1(n66), .A2(n68), .Z(n3899) );
  OR2D1 U4263 ( .A1(n66), .A2(n67), .Z(n3900) );
  OR2D1 U4264 ( .A1(n66), .A2(n99), .Z(n3901) );
  OR2D1 U4265 ( .A1(n66), .A2(n98), .Z(n3902) );
  OR2D1 U4266 ( .A1(n66), .A2(n85), .Z(n3903) );
  OR2D1 U4267 ( .A1(n66), .A2(n72), .Z(n3904) );
  OR2D1 U4268 ( .A1(n66), .A2(n71), .Z(n3905) );
  OR2D1 U4269 ( .A1(n69), .A2(n103), .Z(n3906) );
  OR2D1 U4270 ( .A1(n68), .A2(n103), .Z(n3907) );
  OR2D1 U4271 ( .A1(n67), .A2(n103), .Z(n3908) );
  OR2D1 U4272 ( .A1(n99), .A2(n103), .Z(n3909) );
  OR2D1 U4273 ( .A1(n98), .A2(n103), .Z(n3910) );
  OR2D1 U4274 ( .A1(n85), .A2(n103), .Z(n3911) );
  OR2D1 U4275 ( .A1(n72), .A2(n103), .Z(n3912) );
  OR2D1 U4276 ( .A1(n71), .A2(n103), .Z(n3913) );
  OR2D1 U4277 ( .A1(n69), .A2(n101), .Z(n3914) );
  OR2D1 U4278 ( .A1(n68), .A2(n101), .Z(n3915) );
  OR2D1 U4279 ( .A1(n67), .A2(n101), .Z(n3916) );
  OR2D1 U4280 ( .A1(n99), .A2(n101), .Z(n3917) );
  OR2D1 U4281 ( .A1(n98), .A2(n101), .Z(n3918) );
  OR2D1 U4282 ( .A1(n85), .A2(n101), .Z(n3919) );
  OR2D1 U4283 ( .A1(n72), .A2(n101), .Z(n3920) );
  OR2D1 U4284 ( .A1(n71), .A2(n101), .Z(n3921) );
  BUFFD1 U4285 ( .I(Read), .Z(n4635) );
  BUFFD1 U4286 ( .I(Read), .Z(n4636) );
  INVD1 U4287 ( .I(ClockR), .ZN(n4634) );
  CKAN2D0 U4288 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  MUX4D0 U4289 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(N44), .S1(n4374), .Z(
        n4251) );
  MUX4D0 U4290 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n4384), .S1(n4375), 
        .Z(n4264) );
  MUX4D0 U4291 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n4385), .S1(n4375), 
        .Z(n4277) );
  MUX4D0 U4292 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n4384), .S1(n4376), 
        .Z(n4290) );
  MUX4D0 U4293 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(N44), .S1(n4376), .Z(
        n4316) );
  MUX4D0 U4294 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n4383), .S1(n4374), .Z(
        n4255) );
  MUX4D0 U4295 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n4383), .S1(n4374), 
        .Z(n4253) );
  MUX4D0 U4296 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n4384), .S1(n4375), 
        .Z(n4266) );
  MUX4D0 U4297 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n4384), .S1(n4375), .Z(
        n4268) );
  MUX4D0 U4298 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(N44), .S1(n4375), .Z(
        n4279) );
  MUX4D0 U4299 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n4383), .S1(n4375), .Z(
        n4281) );
  MUX4D0 U4300 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(N44), .S1(n4376), .Z(
        n4294) );
  MUX4D0 U4301 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n4384), .S1(n4376), 
        .Z(n4292) );
  MUX4D0 U4302 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n4384), .S1(n4376), .Z(
        n4307) );
  MUX4D0 U4303 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n4386), .S1(n4376), 
        .Z(n4305) );
  MUX4D0 U4304 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n4386), .S1(n4377), 
        .Z(n4318) );
  MUX4D0 U4305 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(N44), .S1(n4377), .Z(
        n4320) );
  MUX4D0 U4306 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n4384), .S1(n4377), 
        .Z(n4331) );
  MUX4D0 U4307 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n4384), .S1(n4377), .Z(
        n4333) );
  MUX4D0 U4308 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n4383), .S1(n4374), 
        .Z(n4252) );
  MUX4D0 U4309 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n4384), .S1(n4375), 
        .Z(n4265) );
  MUX4D0 U4310 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n4383), .S1(n4375), 
        .Z(n4278) );
  MUX4D0 U4311 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n4383), .S1(n4376), 
        .Z(n4291) );
  MUX4D0 U4312 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n4386), .S1(n4376), 
        .Z(n4304) );
  MUX4D0 U4313 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(N44), .S1(n4377), .Z(
        n4317) );
  MUX4D0 U4314 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n4383), .S1(n4377), 
        .Z(n4330) );
  MUX4D0 U4315 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n4383), .S1(n4375), .Z(
        n4256) );
  MUX4D0 U4316 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(N44), .S1(n4374), .Z(
        n4254) );
  MUX4D0 U4317 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(N44), .S1(n4375), .Z(
        n4267) );
  MUX4D0 U4318 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n4383), .S1(n4375), .Z(
        n4269) );
  MUX4D0 U4319 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n4384), .S1(n4375), 
        .Z(n4280) );
  MUX4D0 U4320 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n4383), .S1(n4375), .Z(
        n4282) );
  MUX4D0 U4321 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n4383), .S1(n4376), .Z(
        n4295) );
  MUX4D0 U4322 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n4383), .S1(n4376), 
        .Z(n4293) );
  MUX4D0 U4323 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n4383), .S1(n4376), .Z(
        n4308) );
  MUX4D0 U4324 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n4397), .S1(n4376), 
        .Z(n4306) );
  MUX4D0 U4325 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n4383), .S1(n4377), 
        .Z(n4319) );
  MUX4D0 U4326 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n4383), .S1(n4377), .Z(
        n4321) );
  MUX4D0 U4327 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n4385), .S1(n4377), 
        .Z(n4332) );
  MUX4D0 U4328 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n4386), .S1(n4377), .Z(
        n4334) );
  MUX4ND0 U4329 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n4396), .S1(n4368), 
        .ZN(n4341) );
  MUX4ND0 U4330 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n4389), .S1(n4369), 
        .ZN(n4250) );
  MUX4ND0 U4331 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n4389), .S1(n4369), 
        .ZN(n4263) );
  MUX4ND0 U4332 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n4383), .S1(n4369), 
        .ZN(n4276) );
  MUX4ND0 U4333 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n4384), .S1(n4369), 
        .ZN(n4289) );
  MUX4ND0 U4334 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n4385), .S1(n4368), 
        .ZN(n4302) );
  MUX4ND0 U4335 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n4383), .S1(n4368), 
        .ZN(n4315) );
  MUX4ND0 U4336 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n4384), .S1(n4368), 
        .ZN(n4328) );
  MUX4D0 U4337 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(N44), .S1(n4377), .Z(
        n4342) );
  MUX4D0 U4338 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n4391), .S1(n4380), .Z(
        n3926) );
  MUX4D0 U4339 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n4392), .S1(n4378), .Z(
        n3939) );
  MUX4D0 U4340 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n4391), .S1(n4379), .Z(
        n3952) );
  MUX4D0 U4341 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n4391), .S1(n4379), .Z(
        n3965) );
  MUX4D0 U4342 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n4391), .S1(n4378), .Z(
        n3978) );
  MUX4D0 U4343 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n4392), .S1(n4378), .Z(
        n3991) );
  MUX4D0 U4344 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n4390), .S1(n4376), .Z(
        n4004) );
  MUX4D0 U4345 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n4393), .S1(n4378), .Z(
        n4017) );
  MUX4D0 U4346 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n4388), .S1(n4381), .Z(
        n4030) );
  MUX4D0 U4347 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n4390), .S1(n4370), .Z(
        n4043) );
  MUX4D0 U4348 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n4390), .S1(n4379), 
        .Z(n4056) );
  MUX4D0 U4349 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n4391), .S1(n4380), 
        .Z(n4069) );
  MUX4D0 U4350 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n4391), .S1(n4381), 
        .Z(n4082) );
  MUX4D0 U4351 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n4392), .S1(n4381), 
        .Z(n4095) );
  MUX4D0 U4352 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n4392), .S1(n4381), 
        .Z(n4108) );
  MUX4D0 U4353 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n4393), .S1(n4382), 
        .Z(n4121) );
  MUX4D0 U4354 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n4393), .S1(n4382), 
        .Z(n4134) );
  MUX4D0 U4355 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n4394), .S1(n4382), 
        .Z(n4147) );
  MUX4D0 U4356 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n4394), .S1(n4371), 
        .Z(n4160) );
  MUX4D0 U4357 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n4395), .S1(n4371), 
        .Z(n4173) );
  MUX4D0 U4358 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n4395), .S1(n4372), 
        .Z(n4186) );
  MUX4D0 U4359 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n4396), .S1(n4372), 
        .Z(n4199) );
  MUX4D0 U4360 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n4396), .S1(n4373), 
        .Z(n4212) );
  MUX4D0 U4361 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n4397), .S1(n4373), 
        .Z(n4225) );
  MUX4D0 U4362 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n4397), .S1(n4374), 
        .Z(n4238) );
  MUX4D0 U4363 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(N44), .S1(n4376), .Z(
        n4303) );
  MUX4D0 U4364 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n4384), .S1(n4377), 
        .Z(n4329) );
  MUX4D0 U4365 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n4385), .S1(n4378), 
        .Z(n4344) );
  MUX4D0 U4366 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n4385), .S1(n4378), .Z(
        n4346) );
  MUX4D0 U4367 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n4386), .S1(n4378), .Z(
        n3930) );
  MUX4D0 U4368 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n4385), .S1(n4378), .Z(
        n3928) );
  MUX4D0 U4369 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n4396), .S1(n4378), .Z(
        n3941) );
  MUX4D0 U4370 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n4385), .S1(n4379), .Z(
        n3943) );
  MUX4D0 U4371 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n4386), .S1(n4379), .Z(
        n3954) );
  MUX4D0 U4372 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n4386), .S1(n4379), .Z(
        n3956) );
  MUX4D0 U4373 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n4392), .S1(n4379), .Z(
        n3969) );
  MUX4D0 U4374 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n4383), .S1(n4379), .Z(
        n3967) );
  MUX4D0 U4375 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n4390), .S1(n4368), .Z(
        n3982) );
  MUX4D0 U4376 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n4390), .S1(n4366), .Z(
        n3980) );
  MUX4D0 U4377 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n4391), .S1(n4372), .Z(
        n3995) );
  MUX4D0 U4378 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n4392), .S1(n4380), .Z(
        n3993) );
  MUX4D0 U4379 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n4393), .S1(n4370), .Z(
        n4006) );
  MUX4D0 U4380 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n4390), .S1(n4381), .Z(
        n4008) );
  MUX4D0 U4381 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n4390), .S1(n4381), .Z(
        n4019) );
  MUX4D0 U4382 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n4388), .S1(n4366), .Z(
        n4021) );
  MUX4D0 U4383 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n4390), .S1(n4364), .Z(
        n4032) );
  MUX4D0 U4384 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n4393), .S1(N45), .Z(n4034) );
  MUX4D0 U4385 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n4390), .S1(n4379), .Z(
        n4047) );
  MUX4D0 U4386 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n4390), .S1(n4374), .Z(
        n4045) );
  MUX4D0 U4387 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n4390), .S1(n4380), .Z(
        n4060) );
  MUX4D0 U4388 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n4390), .S1(n4380), 
        .Z(n4058) );
  MUX4D0 U4389 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n4391), .S1(n4380), .Z(
        n4073) );
  MUX4D0 U4390 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n4391), .S1(n4380), 
        .Z(n4071) );
  MUX4D0 U4391 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n4391), .S1(n4381), 
        .Z(n4084) );
  MUX4D0 U4392 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n4391), .S1(n4381), .Z(
        n4086) );
  MUX4D0 U4393 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n4392), .S1(n4381), 
        .Z(n4097) );
  MUX4D0 U4394 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n4392), .S1(n4382), .Z(
        n4099) );
  MUX4D0 U4395 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n4392), .S1(n4381), .Z(
        n4112) );
  MUX4D0 U4396 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n4392), .S1(n4381), 
        .Z(n4110) );
  MUX4D0 U4397 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n4393), .S1(n4382), .Z(
        n4125) );
  MUX4D0 U4398 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n4393), .S1(n4382), 
        .Z(n4123) );
  MUX4D0 U4399 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n4393), .S1(n4382), 
        .Z(n4136) );
  MUX4D0 U4400 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n4393), .S1(n4380), .Z(
        n4138) );
  MUX4D0 U4401 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n4394), .S1(n4382), .Z(
        n4151) );
  MUX4D0 U4402 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n4394), .S1(n4382), 
        .Z(n4149) );
  MUX4D0 U4403 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n4394), .S1(n4371), .Z(
        n4164) );
  MUX4D0 U4404 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n4394), .S1(n4371), 
        .Z(n4162) );
  MUX4D0 U4405 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n4395), .S1(n4371), 
        .Z(n4175) );
  MUX4D0 U4406 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n4395), .S1(n4372), .Z(
        n4177) );
  MUX4D0 U4407 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n4395), .S1(n4372), 
        .Z(n4188) );
  MUX4D0 U4408 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n4395), .S1(n4372), .Z(
        n4190) );
  MUX4D0 U4409 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n4396), .S1(n4373), .Z(
        n4203) );
  MUX4D0 U4410 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n4396), .S1(n4372), 
        .Z(n4201) );
  MUX4D0 U4411 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n4396), .S1(n4373), .Z(
        n4216) );
  MUX4D0 U4412 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n4396), .S1(n4373), 
        .Z(n4214) );
  MUX4D0 U4413 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n4397), .S1(n4373), 
        .Z(n4227) );
  MUX4D0 U4414 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n4397), .S1(n4373), .Z(
        n4229) );
  MUX4D0 U4415 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n4397), .S1(n4374), .Z(
        n4242) );
  MUX4D0 U4416 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n4397), .S1(n4374), 
        .Z(n4240) );
  MUX4D0 U4417 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(N44), .S1(n4377), .Z(
        n4343) );
  MUX4D0 U4418 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n4397), .S1(n4378), .Z(
        n3927) );
  MUX4D0 U4419 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n4385), .S1(n4378), .Z(
        n3940) );
  MUX4D0 U4420 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n4386), .S1(n4379), .Z(
        n3953) );
  MUX4D0 U4421 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n4392), .S1(n4379), .Z(
        n3966) );
  MUX4D0 U4422 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n4392), .S1(n4368), .Z(
        n3979) );
  MUX4D0 U4423 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n4388), .S1(n4368), .Z(
        n3992) );
  MUX4D0 U4424 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n4393), .S1(n4379), .Z(
        n4005) );
  MUX4D0 U4425 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n4393), .S1(n4379), .Z(
        n4018) );
  MUX4D0 U4426 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n4396), .S1(n4378), .Z(
        n4031) );
  MUX4D0 U4427 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n4390), .S1(n4366), .Z(
        n4044) );
  MUX4D0 U4428 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n4390), .S1(n4382), 
        .Z(n4057) );
  MUX4D0 U4429 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n4391), .S1(n4380), 
        .Z(n4070) );
  MUX4D0 U4430 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n4391), .S1(n4380), 
        .Z(n4083) );
  MUX4D0 U4431 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n4392), .S1(n4381), 
        .Z(n4096) );
  MUX4D0 U4432 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n4392), .S1(n4380), 
        .Z(n4109) );
  MUX4D0 U4433 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n4393), .S1(n4381), 
        .Z(n4122) );
  MUX4D0 U4434 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n4393), .S1(n4381), 
        .Z(n4135) );
  MUX4D0 U4435 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n4394), .S1(n4370), 
        .Z(n4148) );
  MUX4D0 U4436 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n4394), .S1(n4371), 
        .Z(n4161) );
  MUX4D0 U4437 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n4395), .S1(n4371), 
        .Z(n4174) );
  MUX4D0 U4438 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n4395), .S1(n4372), 
        .Z(n4187) );
  MUX4D0 U4439 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n4396), .S1(n4372), 
        .Z(n4200) );
  MUX4D0 U4440 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n4396), .S1(n4373), 
        .Z(n4213) );
  MUX4D0 U4441 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n4397), .S1(n4373), 
        .Z(n4226) );
  MUX4D0 U4442 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n4397), .S1(n4374), 
        .Z(n4239) );
  MUX4D0 U4443 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n4385), .S1(n4378), 
        .Z(n4345) );
  MUX4D0 U4444 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n4397), .S1(n4378), .Z(
        n4347) );
  MUX4D0 U4445 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n4385), .S1(n4378), .Z(
        n3931) );
  MUX4D0 U4446 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n4392), .S1(n4378), .Z(
        n3929) );
  MUX4D0 U4447 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n4385), .S1(n4378), .Z(
        n3942) );
  MUX4D0 U4448 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n4386), .S1(n4379), .Z(
        n3944) );
  MUX4D0 U4449 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n4394), .S1(n4379), .Z(
        n3955) );
  MUX4D0 U4450 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n4396), .S1(n4379), .Z(
        n3957) );
  MUX4D0 U4451 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n4385), .S1(n4381), .Z(
        n3970) );
  MUX4D0 U4452 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n4391), .S1(n4379), .Z(
        n3968) );
  MUX4D0 U4453 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n4393), .S1(n4366), .Z(
        n3983) );
  MUX4D0 U4454 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n4391), .S1(n4378), .Z(
        n3981) );
  MUX4D0 U4455 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n4388), .S1(n4380), .Z(
        n3996) );
  MUX4D0 U4456 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n4391), .S1(n4381), .Z(
        n3994) );
  MUX4D0 U4457 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n4388), .S1(n4374), .Z(
        n4007) );
  MUX4D0 U4458 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n4393), .S1(n4370), .Z(
        n4009) );
  MUX4D0 U4459 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n4393), .S1(n4370), .Z(
        n4020) );
  MUX4D0 U4460 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n4390), .S1(n4379), .Z(
        n4022) );
  MUX4D0 U4461 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n4390), .S1(n4379), .Z(
        n4033) );
  MUX4D0 U4462 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n4392), .S1(n4379), .Z(
        n4035) );
  MUX4D0 U4463 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n4390), .S1(n4640), .Z(
        n4048) );
  MUX4D0 U4464 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n4390), .S1(n4368), .Z(
        n4046) );
  MUX4D0 U4465 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n4390), .S1(n4380), .Z(
        n4061) );
  MUX4D0 U4466 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n4390), .S1(n4380), 
        .Z(n4059) );
  MUX4D0 U4467 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n4391), .S1(n4380), .Z(
        n4074) );
  MUX4D0 U4468 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n4391), .S1(n4380), 
        .Z(n4072) );
  MUX4D0 U4469 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n4391), .S1(n4381), 
        .Z(n4085) );
  MUX4D0 U4470 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n4392), .S1(n4381), .Z(
        n4087) );
  MUX4D0 U4471 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n4392), .S1(n4382), 
        .Z(n4098) );
  MUX4D0 U4472 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n4392), .S1(n4381), .Z(
        n4100) );
  MUX4D0 U4473 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n4393), .S1(n4382), .Z(
        n4113) );
  MUX4D0 U4474 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n4392), .S1(n4382), 
        .Z(n4111) );
  MUX4D0 U4475 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n4393), .S1(n4382), .Z(
        n4126) );
  MUX4D0 U4476 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n4393), .S1(n4382), 
        .Z(n4124) );
  MUX4D0 U4477 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n4393), .S1(n4382), 
        .Z(n4137) );
  MUX4D0 U4478 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n4394), .S1(n4382), .Z(
        n4139) );
  MUX4D0 U4479 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n4394), .S1(n4371), .Z(
        n4152) );
  MUX4D0 U4480 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n4394), .S1(n4380), 
        .Z(n4150) );
  MUX4D0 U4481 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n4395), .S1(n4371), .Z(
        n4165) );
  MUX4D0 U4482 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n4394), .S1(n4371), 
        .Z(n4163) );
  MUX4D0 U4483 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n4395), .S1(n4372), 
        .Z(n4176) );
  MUX4D0 U4484 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n4395), .S1(n4372), .Z(
        n4178) );
  MUX4D0 U4485 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n4395), .S1(n4372), 
        .Z(n4189) );
  MUX4D0 U4486 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n4396), .S1(n4372), .Z(
        n4191) );
  MUX4D0 U4487 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n4396), .S1(n4373), .Z(
        n4204) );
  MUX4D0 U4488 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n4396), .S1(n4372), 
        .Z(n4202) );
  MUX4D0 U4489 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n4397), .S1(n4373), .Z(
        n4217) );
  MUX4D0 U4490 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n4396), .S1(n4373), 
        .Z(n4215) );
  MUX4D0 U4491 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n4397), .S1(n4373), 
        .Z(n4228) );
  MUX4D0 U4492 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n4397), .S1(n4374), .Z(
        n4230) );
  MUX4D0 U4493 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n4386), .S1(n4374), .Z(
        n4243) );
  MUX4D0 U4494 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n4397), .S1(n4374), 
        .Z(n4241) );
  MUX4ND0 U4495 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n4391), .S1(n4371), .ZN(
        n3925) );
  MUX4ND0 U4496 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n4388), .S1(n4371), .ZN(
        n3938) );
  MUX4ND0 U4497 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n4388), .S1(n4371), .ZN(
        n3951) );
  MUX4ND0 U4498 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n4388), .S1(n4370), .ZN(
        n3964) );
  MUX4ND0 U4499 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n4388), .S1(n4370), .ZN(
        n3977) );
  MUX4ND0 U4500 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n4388), .S1(n4370), .ZN(
        n3990) );
  MUX4ND0 U4501 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n4388), .S1(n4370), .ZN(
        n4003) );
  MUX4ND0 U4502 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n4388), .S1(n4370), .ZN(
        n4016) );
  MUX4ND0 U4503 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n4388), .S1(n4370), .ZN(
        n4029) );
  MUX4ND0 U4504 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n4388), .S1(n4370), .ZN(
        n4042) );
  MUX4ND0 U4505 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n4388), .S1(n4370), 
        .ZN(n4055) );
  MUX4ND0 U4506 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n4388), .S1(n4370), 
        .ZN(n4068) );
  MUX4ND0 U4507 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n4388), .S1(n4370), 
        .ZN(n4081) );
  MUX4ND0 U4508 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n4389), .S1(n4370), 
        .ZN(n4094) );
  MUX4ND0 U4509 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n4389), .S1(n4370), 
        .ZN(n4107) );
  MUX4ND0 U4510 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n4389), .S1(n4370), 
        .ZN(n4120) );
  MUX4ND0 U4511 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n4389), .S1(n4369), 
        .ZN(n4133) );
  MUX4ND0 U4512 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n4389), .S1(n4369), 
        .ZN(n4146) );
  MUX4ND0 U4513 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n4389), .S1(n4369), 
        .ZN(n4159) );
  MUX4ND0 U4514 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n4389), .S1(n4369), 
        .ZN(n4172) );
  MUX4ND0 U4515 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n4389), .S1(n4369), 
        .ZN(n4185) );
  MUX4ND0 U4516 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n4389), .S1(n4369), 
        .ZN(n4198) );
  MUX4ND0 U4517 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n4389), .S1(n4369), 
        .ZN(n4211) );
  MUX4ND0 U4518 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n4389), .S1(n4369), 
        .ZN(n4224) );
  MUX4ND0 U4519 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n4389), .S1(n4369), 
        .ZN(n4237) );
  ND3D1 U4520 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U4521 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U4522 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U4523 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U4524 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U4525 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U4526 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U4527 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U4528 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U4529 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  INVD1 U4530 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U4531 ( .I(AddrW[2]), .ZN(n105) );
  INVD1 U4532 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U4533 ( .I(AddrW[4]), .ZN(n102) );
  CKAN2D0 U4534 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U4535 ( .I0(n3923), .I1(n3924), .I2(n3925), .S0(n4382), .S1(N46), 
        .ZN(n3922) );
  MUX3ND0 U4536 ( .I0(n3932), .I1(n3933), .I2(n3870), .S0(n4641), .S1(n4352), 
        .ZN(N82) );
  MUX3ND0 U4537 ( .I0(n3936), .I1(n3937), .I2(n3938), .S0(n4380), .S1(N46), 
        .ZN(n3935) );
  MUX3ND0 U4538 ( .I0(n3949), .I1(n3950), .I2(n3951), .S0(n4370), .S1(n4355), 
        .ZN(n3948) );
  MUX3ND0 U4539 ( .I0(n3962), .I1(n3963), .I2(n3964), .S0(n4362), .S1(n4355), 
        .ZN(n3961) );
  MUX3ND0 U4540 ( .I0(n3971), .I1(n3972), .I2(n3886), .S0(n4641), .S1(n4352), 
        .ZN(N79) );
  MUX3ND0 U4541 ( .I0(n3975), .I1(n3976), .I2(n3977), .S0(n4382), .S1(n4355), 
        .ZN(n3974) );
  MUX3ND0 U4542 ( .I0(n3984), .I1(n3985), .I2(n3872), .S0(n4641), .S1(n4352), 
        .ZN(N78) );
  MUX3ND0 U4543 ( .I0(n3988), .I1(n3989), .I2(n3990), .S0(n4368), .S1(n4355), 
        .ZN(n3987) );
  MUX3ND0 U4544 ( .I0(n3997), .I1(n3998), .I2(n3877), .S0(n4641), .S1(n4352), 
        .ZN(N77) );
  MUX3ND0 U4545 ( .I0(n4001), .I1(n4002), .I2(n4003), .S0(n4366), .S1(n4355), 
        .ZN(n4000) );
  MUX3ND0 U4546 ( .I0(n4010), .I1(n4011), .I2(n3874), .S0(n4641), .S1(n4352), 
        .ZN(N76) );
  MUX3ND0 U4547 ( .I0(n4014), .I1(n4015), .I2(n4016), .S0(n4368), .S1(n4356), 
        .ZN(n4013) );
  MUX3ND0 U4548 ( .I0(n4027), .I1(n4028), .I2(n4029), .S0(n4368), .S1(n4355), 
        .ZN(n4026) );
  MUX3ND0 U4549 ( .I0(n4036), .I1(n4037), .I2(n3885), .S0(n4641), .S1(n4352), 
        .ZN(N74) );
  MUX3ND0 U4550 ( .I0(n4040), .I1(n4041), .I2(n4042), .S0(n4380), .S1(n4355), 
        .ZN(n4039) );
  MUX3ND0 U4551 ( .I0(n4049), .I1(n4050), .I2(n3882), .S0(n4354), .S1(n4352), 
        .ZN(N73) );
  MUX3ND0 U4552 ( .I0(n4053), .I1(n4054), .I2(n4055), .S0(n4366), .S1(n4356), 
        .ZN(n4052) );
  MUX3ND0 U4553 ( .I0(n4062), .I1(n4063), .I2(n3865), .S0(n4641), .S1(n4352), 
        .ZN(N72) );
  MUX3ND0 U4554 ( .I0(n4066), .I1(n4067), .I2(n4068), .S0(n4368), .S1(n4356), 
        .ZN(n4065) );
  MUX3ND0 U4555 ( .I0(n4075), .I1(n4076), .I2(n3108), .S0(n4641), .S1(n4352), 
        .ZN(N71) );
  MUX3ND0 U4556 ( .I0(n4079), .I1(n4080), .I2(n4081), .S0(n4366), .S1(n4360), 
        .ZN(n4078) );
  MUX3ND0 U4557 ( .I0(n4088), .I1(n4089), .I2(n3042), .S0(N47), .S1(n4352), 
        .ZN(N70) );
  MUX3ND0 U4558 ( .I0(n4092), .I1(n4093), .I2(n4094), .S0(n4380), .S1(n4361), 
        .ZN(n4091) );
  MUX3ND0 U4559 ( .I0(n4101), .I1(n4102), .I2(n2976), .S0(N47), .S1(n4352), 
        .ZN(N69) );
  MUX3ND0 U4560 ( .I0(n4105), .I1(n4106), .I2(n4107), .S0(n4366), .S1(n4356), 
        .ZN(n4104) );
  MUX3ND0 U4561 ( .I0(n4114), .I1(n4115), .I2(n2910), .S0(N47), .S1(n4352), 
        .ZN(N68) );
  MUX3ND0 U4562 ( .I0(n4118), .I1(n4119), .I2(n4120), .S0(n4368), .S1(n4355), 
        .ZN(n4117) );
  MUX3ND0 U4563 ( .I0(n4127), .I1(n4128), .I2(n2844), .S0(N47), .S1(n4352), 
        .ZN(N67) );
  MUX3ND0 U4564 ( .I0(n4131), .I1(n4132), .I2(n4133), .S0(n4381), .S1(n4356), 
        .ZN(n4130) );
  MUX3ND0 U4565 ( .I0(n4140), .I1(n4141), .I2(n2778), .S0(N47), .S1(n4352), 
        .ZN(N66) );
  MUX3ND0 U4566 ( .I0(n4144), .I1(n4145), .I2(n4146), .S0(n4382), .S1(n4357), 
        .ZN(n4143) );
  MUX3ND0 U4567 ( .I0(n4153), .I1(n4154), .I2(n2712), .S0(N47), .S1(n4352), 
        .ZN(N65) );
  MUX3ND0 U4568 ( .I0(n4157), .I1(n4158), .I2(n4159), .S0(n4373), .S1(n4356), 
        .ZN(n4156) );
  MUX3ND0 U4569 ( .I0(n4166), .I1(n4167), .I2(n2646), .S0(N47), .S1(n4352), 
        .ZN(N64) );
  MUX3ND0 U4570 ( .I0(n4170), .I1(n4171), .I2(n4172), .S0(n4371), .S1(n4356), 
        .ZN(n4169) );
  MUX3ND0 U4571 ( .I0(n4179), .I1(n4180), .I2(n2580), .S0(N47), .S1(n4352), 
        .ZN(N63) );
  MUX3ND0 U4572 ( .I0(n4183), .I1(n4184), .I2(n4185), .S0(n4373), .S1(n4356), 
        .ZN(n4182) );
  MUX3ND0 U4573 ( .I0(n4192), .I1(n4193), .I2(n2514), .S0(n4354), .S1(N48), 
        .ZN(N62) );
  MUX3ND0 U4574 ( .I0(n4196), .I1(n4197), .I2(n4198), .S0(n4372), .S1(n4356), 
        .ZN(n4195) );
  MUX3ND0 U4575 ( .I0(n4205), .I1(n4206), .I2(n2448), .S0(n4641), .S1(N48), 
        .ZN(N61) );
  MUX3ND0 U4576 ( .I0(n4209), .I1(n4210), .I2(n4211), .S0(n4370), .S1(n4358), 
        .ZN(n4208) );
  MUX3ND0 U4577 ( .I0(n4218), .I1(n4219), .I2(n2382), .S0(N47), .S1(N48), .ZN(
        N60) );
  MUX3ND0 U4578 ( .I0(n4222), .I1(n4223), .I2(n4224), .S0(n4373), .S1(n4361), 
        .ZN(n4221) );
  MUX3ND0 U4579 ( .I0(n4231), .I1(n4232), .I2(n2316), .S0(N47), .S1(N48), .ZN(
        N59) );
  MUX3ND0 U4580 ( .I0(n4235), .I1(n4236), .I2(n4237), .S0(n4368), .S1(n4356), 
        .ZN(n4234) );
  MUX3ND0 U4581 ( .I0(n4244), .I1(n4245), .I2(n2250), .S0(n4354), .S1(N48), 
        .ZN(N58) );
  MUX3ND0 U4582 ( .I0(n4248), .I1(n4249), .I2(n4250), .S0(n4366), .S1(n4356), 
        .ZN(n4247) );
  MUX3ND0 U4583 ( .I0(n4257), .I1(n4258), .I2(n2184), .S0(n4354), .S1(N48), 
        .ZN(N57) );
  MUX3ND0 U4584 ( .I0(n4261), .I1(n4262), .I2(n4263), .S0(n4366), .S1(n4356), 
        .ZN(n4260) );
  MUX3ND0 U4585 ( .I0(n4270), .I1(n4271), .I2(n2118), .S0(n4354), .S1(N48), 
        .ZN(N56) );
  MUX3ND0 U4586 ( .I0(n4274), .I1(n4275), .I2(n4276), .S0(n4366), .S1(n4356), 
        .ZN(n4273) );
  MUX3ND0 U4587 ( .I0(n4283), .I1(n4284), .I2(n2052), .S0(n4353), .S1(N48), 
        .ZN(N55) );
  MUX3ND0 U4588 ( .I0(n4287), .I1(n4288), .I2(n4289), .S0(n4364), .S1(n4357), 
        .ZN(n4286) );
  MUX3ND0 U4589 ( .I0(n4296), .I1(n4297), .I2(n1986), .S0(n4641), .S1(N48), 
        .ZN(N54) );
  MUX3ND0 U4590 ( .I0(n4300), .I1(n4301), .I2(n4302), .S0(n4364), .S1(n4357), 
        .ZN(n4299) );
  MUX3ND0 U4591 ( .I0(n4309), .I1(n4310), .I2(n1920), .S0(N47), .S1(N48), .ZN(
        N53) );
  MUX3ND0 U4592 ( .I0(n4313), .I1(n4314), .I2(n4315), .S0(n4366), .S1(n4357), 
        .ZN(n4312) );
  MUX3ND0 U4593 ( .I0(n4322), .I1(n4323), .I2(n1854), .S0(N47), .S1(N48), .ZN(
        N52) );
  MUX3ND0 U4594 ( .I0(n4326), .I1(n4327), .I2(n4328), .S0(n4368), .S1(n4357), 
        .ZN(n4325) );
  MUX3ND0 U4595 ( .I0(n4335), .I1(n4336), .I2(n1788), .S0(N47), .S1(N48), .ZN(
        N51) );
  MUX3ND0 U4596 ( .I0(n4339), .I1(n4340), .I2(n4341), .S0(n4364), .S1(n4357), 
        .ZN(n4338) );
  MUX3ND0 U4597 ( .I0(n4348), .I1(n4349), .I2(n4350), .S0(n4353), .S1(N48), 
        .ZN(N50) );
  MUX2ND0 U4598 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n4395), 
        .ZN(n3924) );
  MUX2ND0 U4599 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n4385), 
        .ZN(n3923) );
  MUX3ND0 U4600 ( .I0(n3927), .I1(n3926), .I2(n3922), .S0(n4361), .S1(n4641), 
        .ZN(n3934) );
  MUX2ND0 U4601 ( .I0(n3929), .I1(n3928), .S(N46), .ZN(n3933) );
  MUX2ND0 U4602 ( .I0(n3931), .I1(n3930), .S(N46), .ZN(n3932) );
  MUX2ND0 U4603 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n4395), 
        .ZN(n3937) );
  MUX2ND0 U4604 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n4395), 
        .ZN(n3936) );
  MUX3ND0 U4605 ( .I0(n3940), .I1(n3939), .I2(n3935), .S0(n4361), .S1(n4353), 
        .ZN(n3947) );
  MUX2ND0 U4606 ( .I0(n3942), .I1(n3941), .S(n4359), .ZN(n3946) );
  MUX2ND0 U4607 ( .I0(n3944), .I1(n3943), .S(n4360), .ZN(n3945) );
  MUX2ND0 U4608 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n4394), 
        .ZN(n3950) );
  MUX2ND0 U4609 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n4394), 
        .ZN(n3949) );
  MUX3ND0 U4610 ( .I0(n3953), .I1(n3952), .I2(n3948), .S0(n4361), .S1(n4641), 
        .ZN(n3960) );
  MUX2ND0 U4611 ( .I0(n3955), .I1(n3954), .S(n4361), .ZN(n3959) );
  MUX2ND0 U4612 ( .I0(n3957), .I1(n3956), .S(n4356), .ZN(n3958) );
  MUX2ND0 U4613 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n4395), 
        .ZN(n3963) );
  MUX2ND0 U4614 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n4384), 
        .ZN(n3962) );
  MUX3ND0 U4615 ( .I0(n3966), .I1(n3965), .I2(n3961), .S0(n4361), .S1(n4641), 
        .ZN(n3973) );
  MUX2ND0 U4616 ( .I0(n3968), .I1(n3967), .S(N46), .ZN(n3972) );
  MUX2ND0 U4617 ( .I0(n3970), .I1(n3969), .S(n4356), .ZN(n3971) );
  MUX2ND0 U4618 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n4386), 
        .ZN(n3976) );
  MUX2ND0 U4619 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n4397), 
        .ZN(n3975) );
  MUX3ND0 U4620 ( .I0(n3979), .I1(n3978), .I2(n3974), .S0(n4361), .S1(n4641), 
        .ZN(n3986) );
  MUX2ND0 U4621 ( .I0(n3981), .I1(n3980), .S(n4358), .ZN(n3985) );
  MUX2ND0 U4622 ( .I0(n3983), .I1(n3982), .S(N46), .ZN(n3984) );
  MUX2ND0 U4623 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n4385), 
        .ZN(n3989) );
  MUX2ND0 U4624 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n4387), 
        .ZN(n3988) );
  MUX3ND0 U4625 ( .I0(n3992), .I1(n3991), .I2(n3987), .S0(n4360), .S1(n4353), 
        .ZN(n3999) );
  MUX2ND0 U4626 ( .I0(n3994), .I1(n3993), .S(n4355), .ZN(n3998) );
  MUX2ND0 U4627 ( .I0(n3996), .I1(n3995), .S(n4355), .ZN(n3997) );
  MUX2ND0 U4628 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n4387), 
        .ZN(n4002) );
  MUX2ND0 U4629 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n4387), 
        .ZN(n4001) );
  MUX3ND0 U4630 ( .I0(n4005), .I1(n4004), .I2(n4000), .S0(n4360), .S1(n4353), 
        .ZN(n4012) );
  MUX2ND0 U4631 ( .I0(n4007), .I1(n4006), .S(n4359), .ZN(n4011) );
  MUX2ND0 U4632 ( .I0(n4009), .I1(n4008), .S(n4358), .ZN(n4010) );
  MUX2ND0 U4633 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n4387), 
        .ZN(n4015) );
  MUX2ND0 U4634 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n4387), 
        .ZN(n4014) );
  MUX3ND0 U4635 ( .I0(n4018), .I1(n4017), .I2(n4013), .S0(N46), .S1(n4353), 
        .ZN(n4025) );
  MUX2ND0 U4636 ( .I0(n4020), .I1(n4019), .S(N46), .ZN(n4024) );
  MUX2ND0 U4637 ( .I0(n4022), .I1(n4021), .S(N46), .ZN(n4023) );
  MUX2ND0 U4638 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n4388), 
        .ZN(n4028) );
  MUX2ND0 U4639 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n4387), 
        .ZN(n4027) );
  MUX3ND0 U4640 ( .I0(n4031), .I1(n4030), .I2(n4026), .S0(n4361), .S1(n4353), 
        .ZN(n4038) );
  MUX2ND0 U4641 ( .I0(n4033), .I1(n4032), .S(n4355), .ZN(n4037) );
  MUX2ND0 U4642 ( .I0(n4035), .I1(n4034), .S(N46), .ZN(n4036) );
  MUX2ND0 U4643 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n4387), 
        .ZN(n4041) );
  MUX2ND0 U4644 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n4388), 
        .ZN(n4040) );
  MUX3ND0 U4645 ( .I0(n4044), .I1(n4043), .I2(n4039), .S0(n4360), .S1(n4353), 
        .ZN(n4051) );
  MUX2ND0 U4646 ( .I0(n4046), .I1(n4045), .S(n4359), .ZN(n4050) );
  MUX2ND0 U4647 ( .I0(n4048), .I1(n4047), .S(n4357), .ZN(n4049) );
  MUX2ND0 U4648 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n4388), 
        .ZN(n4054) );
  MUX2ND0 U4649 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n4387), 
        .ZN(n4053) );
  MUX3ND0 U4650 ( .I0(n4057), .I1(n4056), .I2(n4052), .S0(n4359), .S1(n4353), 
        .ZN(n4064) );
  MUX2ND0 U4651 ( .I0(n4059), .I1(n4058), .S(n4355), .ZN(n4063) );
  MUX2ND0 U4652 ( .I0(n4061), .I1(n4060), .S(N46), .ZN(n4062) );
  MUX2ND0 U4653 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n4387), 
        .ZN(n4067) );
  MUX2ND0 U4654 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n4387), 
        .ZN(n4066) );
  MUX3ND0 U4655 ( .I0(n4070), .I1(n4069), .I2(n4065), .S0(n4359), .S1(n4353), 
        .ZN(n4077) );
  MUX2ND0 U4656 ( .I0(n4072), .I1(n4071), .S(n4355), .ZN(n4076) );
  MUX2ND0 U4657 ( .I0(n4074), .I1(n4073), .S(n4356), .ZN(n4075) );
  MUX2ND0 U4658 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n4387), 
        .ZN(n4080) );
  MUX2ND0 U4659 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n4387), 
        .ZN(n4079) );
  MUX3ND0 U4660 ( .I0(n4083), .I1(n4082), .I2(n4078), .S0(n4360), .S1(n4353), 
        .ZN(n4090) );
  MUX2ND0 U4661 ( .I0(n4085), .I1(n4084), .S(n4355), .ZN(n4089) );
  MUX2ND0 U4662 ( .I0(n4087), .I1(n4086), .S(n4357), .ZN(n4088) );
  MUX2ND0 U4663 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n4387), 
        .ZN(n4093) );
  MUX2ND0 U4664 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n4387), 
        .ZN(n4092) );
  MUX3ND0 U4665 ( .I0(n4096), .I1(n4095), .I2(n4091), .S0(n4360), .S1(n4353), 
        .ZN(n4103) );
  MUX2ND0 U4666 ( .I0(n4098), .I1(n4097), .S(n4356), .ZN(n4102) );
  MUX2ND0 U4667 ( .I0(n4100), .I1(n4099), .S(n4358), .ZN(n4101) );
  MUX2ND0 U4668 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n4387), 
        .ZN(n4106) );
  MUX2ND0 U4669 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n4387), 
        .ZN(n4105) );
  MUX3ND0 U4670 ( .I0(n4109), .I1(n4108), .I2(n4104), .S0(n4356), .S1(n4353), 
        .ZN(n4116) );
  MUX2ND0 U4671 ( .I0(n4111), .I1(n4110), .S(n4360), .ZN(n4115) );
  MUX2ND0 U4672 ( .I0(n4113), .I1(n4112), .S(n4355), .ZN(n4114) );
  MUX2ND0 U4673 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n4387), 
        .ZN(n4119) );
  MUX2ND0 U4674 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n4387), 
        .ZN(n4118) );
  MUX3ND0 U4675 ( .I0(n4122), .I1(n4121), .I2(n4117), .S0(N46), .S1(n4353), 
        .ZN(n4129) );
  MUX2ND0 U4676 ( .I0(n4124), .I1(n4123), .S(n4355), .ZN(n4128) );
  MUX2ND0 U4677 ( .I0(n4126), .I1(n4125), .S(n4359), .ZN(n4127) );
  MUX2ND0 U4678 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n4387), 
        .ZN(n4132) );
  MUX2ND0 U4679 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n4385), 
        .ZN(n4131) );
  MUX3ND0 U4680 ( .I0(n4135), .I1(n4134), .I2(n4130), .S0(n4360), .S1(n4353), 
        .ZN(n4142) );
  MUX2ND0 U4681 ( .I0(n4137), .I1(n4136), .S(n4359), .ZN(n4141) );
  MUX2ND0 U4682 ( .I0(n4139), .I1(n4138), .S(n4359), .ZN(n4140) );
  MUX2ND0 U4683 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n4386), 
        .ZN(n4145) );
  MUX2ND0 U4684 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n4394), 
        .ZN(n4144) );
  MUX3ND0 U4685 ( .I0(n4148), .I1(n4147), .I2(n4143), .S0(n4360), .S1(n4353), 
        .ZN(n4155) );
  MUX2ND0 U4686 ( .I0(n4150), .I1(n4149), .S(n4359), .ZN(n4154) );
  MUX2ND0 U4687 ( .I0(n4152), .I1(n4151), .S(n4359), .ZN(n4153) );
  MUX2ND0 U4688 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n4386), 
        .ZN(n4158) );
  MUX2ND0 U4689 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n4396), 
        .ZN(n4157) );
  MUX3ND0 U4690 ( .I0(n4161), .I1(n4160), .I2(n4156), .S0(n4360), .S1(n4353), 
        .ZN(n4168) );
  MUX2ND0 U4691 ( .I0(n4163), .I1(n4162), .S(n4359), .ZN(n4167) );
  MUX2ND0 U4692 ( .I0(n4165), .I1(n4164), .S(n4359), .ZN(n4166) );
  MUX2ND0 U4693 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n4386), 
        .ZN(n4171) );
  MUX2ND0 U4694 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n4396), 
        .ZN(n4170) );
  MUX3ND0 U4695 ( .I0(n4174), .I1(n4173), .I2(n4169), .S0(n4359), .S1(n4354), 
        .ZN(n4181) );
  MUX2ND0 U4696 ( .I0(n4176), .I1(n4175), .S(n4359), .ZN(n4180) );
  MUX2ND0 U4697 ( .I0(n4178), .I1(n4177), .S(n4359), .ZN(n4179) );
  MUX2ND0 U4698 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n4397), 
        .ZN(n4184) );
  MUX2ND0 U4699 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n4397), 
        .ZN(n4183) );
  MUX3ND0 U4700 ( .I0(n4187), .I1(n4186), .I2(n4182), .S0(n4360), .S1(n4354), 
        .ZN(n4194) );
  MUX2ND0 U4701 ( .I0(n4189), .I1(n4188), .S(n4359), .ZN(n4193) );
  MUX2ND0 U4702 ( .I0(n4191), .I1(n4190), .S(n4359), .ZN(n4192) );
  MUX2ND0 U4703 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n4396), 
        .ZN(n4197) );
  MUX2ND0 U4704 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n4395), 
        .ZN(n4196) );
  MUX3ND0 U4705 ( .I0(n4200), .I1(n4199), .I2(n4195), .S0(n4359), .S1(n4354), 
        .ZN(n4207) );
  MUX2ND0 U4706 ( .I0(n4202), .I1(n4201), .S(n4359), .ZN(n4206) );
  MUX2ND0 U4707 ( .I0(n4204), .I1(n4203), .S(n4359), .ZN(n4205) );
  MUX2ND0 U4708 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n4396), 
        .ZN(n4210) );
  MUX2ND0 U4709 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n4397), 
        .ZN(n4209) );
  MUX3ND0 U4710 ( .I0(n4213), .I1(n4212), .I2(n4208), .S0(n4361), .S1(n4354), 
        .ZN(n4220) );
  MUX2ND0 U4711 ( .I0(n4215), .I1(n4214), .S(n4358), .ZN(n4219) );
  MUX2ND0 U4712 ( .I0(n4217), .I1(n4216), .S(n4358), .ZN(n4218) );
  MUX2ND0 U4713 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n4385), 
        .ZN(n4223) );
  MUX2ND0 U4714 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n4389), 
        .ZN(n4222) );
  MUX3ND0 U4715 ( .I0(n4226), .I1(n4225), .I2(n4221), .S0(n4360), .S1(n4354), 
        .ZN(n4233) );
  MUX2ND0 U4716 ( .I0(n4228), .I1(n4227), .S(n4358), .ZN(n4232) );
  MUX2ND0 U4717 ( .I0(n4230), .I1(n4229), .S(n4358), .ZN(n4231) );
  MUX2ND0 U4718 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n4397), 
        .ZN(n4236) );
  MUX2ND0 U4719 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n4394), 
        .ZN(n4235) );
  MUX3ND0 U4720 ( .I0(n4239), .I1(n4238), .I2(n4234), .S0(n4360), .S1(n4354), 
        .ZN(n4246) );
  MUX2ND0 U4721 ( .I0(n4241), .I1(n4240), .S(n4358), .ZN(n4245) );
  MUX2ND0 U4722 ( .I0(n4243), .I1(n4242), .S(n4358), .ZN(n4244) );
  MUX2ND0 U4723 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n4386), 
        .ZN(n4249) );
  MUX2ND0 U4724 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n4389), 
        .ZN(n4248) );
  MUX3ND0 U4725 ( .I0(n4252), .I1(n4251), .I2(n4247), .S0(n4360), .S1(n4641), 
        .ZN(n4259) );
  MUX2ND0 U4726 ( .I0(n4254), .I1(n4253), .S(n4358), .ZN(n4258) );
  MUX2ND0 U4727 ( .I0(n4256), .I1(n4255), .S(n4358), .ZN(n4257) );
  MUX2ND0 U4728 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n4386), 
        .ZN(n4262) );
  MUX2ND0 U4729 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n4386), 
        .ZN(n4261) );
  MUX3ND0 U4730 ( .I0(n4265), .I1(n4264), .I2(n4260), .S0(n4361), .S1(n4354), 
        .ZN(n4272) );
  MUX2ND0 U4731 ( .I0(n4267), .I1(n4266), .S(n4358), .ZN(n4271) );
  MUX2ND0 U4732 ( .I0(n4269), .I1(n4268), .S(n4358), .ZN(n4270) );
  MUX2ND0 U4733 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n4389), 
        .ZN(n4275) );
  MUX2ND0 U4734 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n4389), 
        .ZN(n4274) );
  MUX3ND0 U4735 ( .I0(n4278), .I1(n4277), .I2(n4273), .S0(n4360), .S1(n4641), 
        .ZN(n4285) );
  MUX2ND0 U4736 ( .I0(n4280), .I1(n4279), .S(n4358), .ZN(n4284) );
  MUX2ND0 U4737 ( .I0(n4282), .I1(n4281), .S(n4358), .ZN(n4283) );
  MUX2ND0 U4738 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n4386), 
        .ZN(n4288) );
  MUX2ND0 U4739 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n4384), 
        .ZN(n4287) );
  MUX3ND0 U4740 ( .I0(n4291), .I1(n4290), .I2(n4286), .S0(n4361), .S1(n4354), 
        .ZN(n4298) );
  MUX2ND0 U4741 ( .I0(n4293), .I1(n4292), .S(n4358), .ZN(n4297) );
  MUX2ND0 U4742 ( .I0(n4295), .I1(n4294), .S(n4357), .ZN(n4296) );
  MUX2ND0 U4743 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n4395), 
        .ZN(n4301) );
  MUX2ND0 U4744 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n4384), 
        .ZN(n4300) );
  MUX3ND0 U4745 ( .I0(n4304), .I1(n4303), .I2(n4299), .S0(n4361), .S1(n4354), 
        .ZN(n4311) );
  MUX2ND0 U4746 ( .I0(n4306), .I1(n4305), .S(n4357), .ZN(n4310) );
  MUX2ND0 U4747 ( .I0(n4308), .I1(n4307), .S(n4357), .ZN(n4309) );
  MUX2ND0 U4748 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n4395), 
        .ZN(n4314) );
  MUX2ND0 U4749 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n4389), 
        .ZN(n4313) );
  MUX3ND0 U4750 ( .I0(n4317), .I1(n4316), .I2(n4312), .S0(n4361), .S1(n4354), 
        .ZN(n4324) );
  MUX2ND0 U4751 ( .I0(n4319), .I1(n4318), .S(n4357), .ZN(n4323) );
  MUX2ND0 U4752 ( .I0(n4321), .I1(n4320), .S(n4357), .ZN(n4322) );
  MUX2ND0 U4753 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n4394), 
        .ZN(n4327) );
  MUX2ND0 U4754 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n4384), 
        .ZN(n4326) );
  MUX3ND0 U4755 ( .I0(n4330), .I1(n4329), .I2(n4325), .S0(n4361), .S1(n4354), 
        .ZN(n4337) );
  MUX2ND0 U4756 ( .I0(n4332), .I1(n4331), .S(n4357), .ZN(n4336) );
  MUX2ND0 U4757 ( .I0(n4334), .I1(n4333), .S(n4357), .ZN(n4335) );
  MUX2ND0 U4758 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n4389), 
        .ZN(n4340) );
  MUX2ND0 U4759 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n4387), 
        .ZN(n4339) );
  MUX3ND0 U4760 ( .I0(n4343), .I1(n4342), .I2(n4338), .S0(n4361), .S1(n4353), 
        .ZN(n4350) );
  MUX2ND0 U4761 ( .I0(n4345), .I1(n4344), .S(n4357), .ZN(n4349) );
  MUX2ND0 U4762 ( .I0(n4347), .I1(n4346), .S(n4356), .ZN(n4348) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] , n1;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(n1), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  BUFFD0 U1 ( .I(A[0]), .Z(n1) );
  INVD1 U2 ( .I(n1), .ZN(SUM[0]) );
  CKXOR2D0 U3 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
endmodule

