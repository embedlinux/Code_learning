`ifndef RKV_I2C_CONFIGS_SVH
`define RKV_I2C_CONFIGS_SVH

`include "rkv_i2c_defines.svh"
`include "rkv_i2c_config.sv"

`endif // RKV_I2C_CONFIGS_SVH
