
`ifndef RKV_I2C_ELEMENT_SEQUENCES_SVH
`define RKV_I2C_ELEMENT_SEQUENCES_SVH

`include "rkv_apb_base_sequence.sv"
`include "rkv_apb_config_seq.sv"
`include "rkv_apb_tx_seq.sv"
`include "rkv_apb_rx_seq.sv"
`include "rkv_apb_wait_empty_seq.sv"
`include "rkv_apb_intr_enable_seq.sv"

`include "rkv_i2c_slave_base_sequence.sv"
`include "rkv_i2c_slave_rx_seq.sv"


`endif // RKV_I2C_ELEMENT_SEQUENCES_SVH
