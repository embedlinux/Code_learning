library verilog;
use verilog.vl_types.all;
entity TFT_CTRL_tb is
end TFT_CTRL_tb;
