module chkblk ( ck54, p_rst_x, bt_rst, e_cd_en, bl_v_jpg, v_dec_mod, 
    bl_v_dec_mod, v_pic_all, b_buf_rdt, br_buf_valid, bt_pulse1, bt_pulse2, 
    bt_pulse3, bt_pulse4, bt_pulse5, bt_pulse6, bp_bufval, bp_jpg_enc_sta_adr, 
    bp_jpg_enc_end_adr, bp_jpg_dec_sta_adr, bp_jpg_dec_end_adr, p_out_sta, 
    p_mem_pic, p_dec_sta, s_sd_init, e_stfd_byt, b_dec_en, d_acc_unit, 
    d_seq_end, bd_overflow, s_sd_dat, b_sd_dat, b_sd_adr, b_sd_en, p_bs_req, 
    b_cpu_ack, p_bs_dat, b_cpu_irq, b_cpu_req, bd_dt_ava, bd_au_count, 
    bd_bm_count, b_seq_end, bd_cpu_end, bd_au_state, bd_bm_count_32b, 
    bd_chk_seq_end, bd_cpu_ack_cnt, bd_cpu_ack_dly, bd_cpu_req_lt, 
    bd_gop_hdr_exist, bd_mem_au_count, bd_mem_en, bd_overflow_prev, 
    bd_we_dec_adv, bd_wee_red_adv, bd_seq_hdr_exist, bd_underflow_prev, 
    bd_re_enc_adv, bd_bs_req_lt, bd_underflow, bd_stfd_byt_cnt );
input  [31:0] b_buf_rdt;
input  [7:0] bp_jpg_enc_end_adr;
output [18:0] b_sd_adr;
input  [13:0] bp_bufval;
input  [7:0] bp_jpg_enc_sta_adr;
input  [31:0] s_sd_dat;
output [1:0] b_cpu_irq;
output [13:0] bd_bm_count;
output [1:0] bd_au_state;
output [5:0] bd_cpu_ack_cnt;
input  [31:0] p_bs_dat;
output [5:0] bd_au_count;
output [14:0] bd_bm_count_32b;
input  [7:0] bp_jpg_dec_sta_adr;
input  [7:0] bp_jpg_dec_end_adr;
input  [9:0] e_stfd_byt;
output [6:0] bd_mem_au_count;
output [31:0] b_sd_dat;
output [12:0] bd_stfd_byt_cnt;
input  ck54, p_rst_x, bt_rst, e_cd_en, bl_v_jpg, v_dec_mod, bl_v_dec_mod, 
    v_pic_all, br_buf_valid, bt_pulse1, bt_pulse2, bt_pulse3, bt_pulse4, 
    bt_pulse5, bt_pulse6, p_out_sta, p_mem_pic, p_dec_sta, s_sd_init, 
    d_acc_unit, d_seq_end, p_bs_req;
output b_dec_en, bd_overflow, b_sd_en, b_cpu_ack, b_cpu_req, bd_dt_ava, 
    b_seq_end, bd_cpu_end, bd_chk_seq_end, bd_cpu_ack_dly, bd_cpu_req_lt, 
    bd_gop_hdr_exist, bd_mem_en, bd_overflow_prev, bd_we_dec_adv, 
    bd_wee_red_adv, bd_seq_hdr_exist, bd_underflow_prev, bd_re_enc_adv, 
    bd_bs_req_lt, bd_underflow;
    wire bd_w_adr_c_plus_1_4_, blk_with_stfd_cnt_6_, stfd_byt_cnt11156_6_, 
        bd_r_adr_r_plus_1_10_, bd_w_adr_r_10_, bd_w_adr_r_plus_1_6_, 
        bd_mem_au_count11744_3_, n598_25_, bd_sd_adr_8_, 
        bd_cpu_ack_cnt11656_3_, bd_au_count11668_3_, bd_w_adr_r_plus_1_2_, 
        bd_cpu_endb, n598_28_, bd_sd_adr_5_, stfd_byt_cnt11156_2_, 
        blk_with_stfd_cnt_2_, bd_bm_count_32b11622_12_, bd_seq_hdr_exist11078, 
        bd_bm_count_32b11622_10_, n598_23_, bd_w_adr_r_plus_1_9_, 
        bd_au_count11668_5_, stfd_byt_cnt11156_9_, bd_sd_adr_7_, 
        blk_with_stfd_cnt_9_, stfd_byt_cnt11156_0_, bd_w_adr_c_plus_1_2_, 
        bd_mem_au_count11744_5_, bd_overflow_prev11090, n598_27_, b_sd_en11058, 
        bd_bm_count_32b11622_14_, bd_cpu_ack_cnt11656_1_, bd_sd_adr_3_, 
        bd_w_adr_r_plus_1_4_, stfd_byt_cnt11156_11_, blk_with_stfd_cnt_4_, 
        bd_sd_adr_18_, stfd_byt_cnt11156_4_, bd_r_adr_c_plus_1_1_, 
        stfd_byt_cnt11157_9_, bd_sd_dat11062_3_, bd_sd_dat_30_, bd_sd_dat_29_, 
        bd_r_adr_r_plus_1_3_, bd_r_adr_r_9_, bd_sd_dat_0_, 
        bd_bm_count_32b11631_6_, bd_bs_dat11066_27_, bd_sd_dat11062_18_, 
        bd_bs_dat11066_14_, b_sd_dat11070_9_, bd_w_adr_c_2_, bd_r_adr_r_0_, 
        bd_sd_dat_9_, bd_sd_dat_13_, bd_sd_dat_20_, bd_sd_adr_11_, 
        bd_w_adr_r_3_, b_sd_dat11070_26_, bd_bs_dat11066_5_, b_sd_dat11070_0_, 
        bd_r_adr_c_1_, b_sd_dat11070_15_, bd_sd_dat11062_11_, 
        bd_sd_dat11062_22_, bd_bm_count_32b11622_6_, b_sd_dat11070_18_, 
        bd_bs_dat11066_8_, bd_bs_dat11066_23_, bd_bs_dat11066_10_, 
        bd_sd_dat_4_, bd_bm_count_32b11631_2_, bd_sd_adr_15_, 
        bd_r_adr_r_plus_1_7_, n603_31_, n603_28_, bd_sd_dat11062_7_, 
        bd_bm_count_32b11622_2_, bd_au_count11677_4_, stfd_byt_cnt11157_4_, 
        bd_r_adr_c_5_, bd_bs_dat11066_19_, bd_sd_dat11062_15_, bd_w_adr_r_7_, 
        bd_sd_dat11062_26_, b_sd_dat11070_4_, bd_bs_dat11066_1_, 
        b_sd_dat11070_22_, b_sd_dat11070_11_, bd_sd_dat_17_, 
        bd_bm_count_32b11631_13_, bd_sd_dat_24_, bd_r_adr_r_4_, bd_sd_adr_17_, 
        bd_sd_dat11062_17_, bd_sd_dat11062_24_, bd_w_adr_r_5_, 
        bd_bs_dat11066_31_, bd_bs_dat11066_28_, bd_cpu_ack_dly11086, 
        b_sd_dat11070_20_, bd_bs_dat11066_3_, b_sd_dat11070_6_, bd_w_adr_c_4_, 
        b_sd_dat11070_13_, bd_au_state11074_1_, bd_sd_dat_15_, 
        bd_bm_count_32b11631_11_, bd_sd_dat_26_, bd_r_adr_r_6_, 
        bd_bm_count_32b11631_9_, stfd_byt_cnt11157_6_, bd_bm_count_32b11622_9_, 
        n603_19_, bd_sd_dat11062_5_, b_sd_dat11070_30_, b_sd_dat11070_29_, 
        bd_bs_dat11066_21_, bd_bs_dat11066_12_, bd_sd_dat_6_, 
        bd_cpu_req_lt11152, bd_bm_count_32b11631_0_, bd_r_adr_r_plus_1_5_, 
        bd_sd_dat11062_8_, stfd_byt_cnt11157_2_, bd_au_count11677_2_, 
        bd_bm_count_32b11622_4_, bd_r_adr_r_2_, bd_sd_adr_13_, bd_w_adr_c_0_, 
        blk_with_stfd_cnt_11_, bd_sd_dat_11_, bd_r_adr_r_plus_1_8_, 
        bd_sd_dat_22_, bd_w_adr_r_1_, bd_r_adr_c_3_, b_sd_dat11070_2_, 
        bd_bs_dat11066_7_, b_sd_dat11070_24_, b_sd_dat11070_17_, 
        bd_sd_dat11062_13_, bd_r_adr_r_plus_1_1_, bd_sd_dat11062_20_, 
        bd_sd_dat_18_, bd_sd_dat_2_, bd_bm_count_32b11631_4_, 
        bd_bs_dat11066_25_, bd_sd_dat11062_30_, bd_sd_dat11062_29_, 
        bd_bs_dat11066_16_, bd_w_adr_r_8_, bd_r_adr_c_plus_1_3_, 
        bd_sd_dat11062_1_, bd_w_adr_r_plus_1_10_, bd_au_count11677_3_, 
        bd_sd_dat11062_9_, stfd_byt_cnt11157_3_, bd_active_once, n603_26_, 
        bd_w_adr_c_1_, bd_bm_count_32b11622_5_, bd_sd_dat_10_, 
        bd_bm_count_32b11631_14_, bd_r_adr_r_plus_1_9_, bd_sd_dat_23_, 
        bd_sd_adr_16_, bd_sd_adr_12_, bd_r_adr_r_3_, blk_with_stfd_cnt_10_, 
        bd_r_adr_c_2_, bl_v_jpg_q, bd_sd_dat11062_12_, bd_sd_dat11062_21_, 
        bd_w_adr_r_0_, bd_bs_dat11066_6_, b_sd_dat11070_25_, b_sd_dat11070_3_, 
        b_sd_dat11070_16_, bd_sd_dat_3_, bd_bm_count_32b11631_5_, 
        bd_sd_dat_19_, bd_w_adr_r_9_, bd_sd_dat11062_28_, bd_sd_dat11062_31_, 
        bd_bs_dat11066_24_, bd_bs_dat11066_17_, bd_sd_dat11062_0_, 
        bd_r_adr_c_plus_1_2_, bd_w_adr_r_4_, b_sd_dat11070_7_, 
        b_sd_dat11070_21_, bd_bs_dat11066_2_, b_sd_dat11070_12_, 
        bd_sd_dat11062_16_, bd_bs_dat11066_30_, bd_bs_dat11066_29_, 
        bd_r_adr_r_7_, bd_sd_dat11062_25_, bd_bm_count_32b11631_8_, 
        bd_w_adr_c_5_, bd_au_state11074_0_, bd_bm_count_32b11631_10_, 
        bd_sd_dat_14_, bd_sd_dat_27_, bd_bm_count_32b11622_1_, 
        stfd_byt_cnt11157_7_, bd_bm_count_32b11622_8_, bd_sd_dat11062_4_, 
        bd_bs_dat11066_20_, bd_bs_dat11066_13_, b_sd_dat11070_28_, 
        b_sd_dat11070_31_, bd_r_adr_r_plus_1_4_, bd_sd_dat_7_, 
        bd_bm_count_32b11631_1_, bd_bs_dat11066_22_, bd_bs_dat11066_11_, 
        b_sd_dat11070_19_, bd_bs_dat11066_9_, bd_r_adr_r_plus_1_6_, 
        bd_sd_dat_5_, bd_r_adr_r_10_, bd_bm_count_32b11631_3_, n603_29_, 
        n603_30_, bd_r_adr_c_plus_1_4_, bd_sd_dat11062_6_, b_cpu_req11098, 
        bd_bm_count_32b11622_3_, stfd_byt_cnt11157_5_, bd_au_count11677_5_, 
        bd_sd_adr_14_, bd_w_adr_r_6_, bd_bs_dat11066_0_, b_sd_dat11070_23_, 
        b_sd_dat11070_5_, b_sd_dat11070_10_, bd_r_adr_c_4_, bd_cpu_irq011148, 
        bd_sd_dat11062_14_, bd_bs_dat11066_18_, bd_sd_dat11062_27_, 
        bd_r_adr_r_5_, bd_sd_dat_16_, bd_bm_count_32b11631_12_, bd_sd_dat_25_, 
        stfd_byt_cnt11157_8_, bd_sd_dat11062_2_, bd_r_adr_r_8_, bd_sd_dat_1_, 
        bd_bm_count_32b11631_7_, bd_sd_dat_28_, bd_sd_dat_31_, 
        bd_r_adr_r_plus_1_2_, b_sd_dat11070_8_, bd_bs_dat11066_26_, 
        bd_w_adr_c_3_, bd_bs_dat11066_15_, bd_underflow_prev11094, 
        bd_sd_dat11062_19_, bd_sd_dat_12_, bd_sd_dat_21_, bd_r_adr_r_1_, 
        blk_with_stfd_cnt_12_, bd_sd_adr_10_, bd_r_adr_c_0_, bd_sd_dat_8_, 
        bd_sd_dat11062_10_, bd_w_adr_r_2_, bd_sd_dat11062_23_, 
        b_sd_dat11070_1_, b_sd_dat11070_27_, bd_bs_dat11066_4_, 
        b_sd_dat11070_14_, stfd_byt_cnt11157_1_, bd_bm_count_32b11622_7_, 
        n598_26_, bd_w_adr_r_plus_1_5_, blk_with_stfd_cnt_5_, 
        stfd_byt_cnt11156_10_, stfd_byt_cnt11156_5_, bd_sd_adr_6_, 
        bd_bm_count_32b11622_11_, bd_cpu_ack_cnt11656_4_, 
        bd_gop_hdr_exist11082, n598_22_, bd_w_adr_r_plus_1_8_, 
        stfd_byt_cnt11156_8_, bd_au_count11668_4_, blk_with_stfd_cnt_8_, 
        stfd_byt_cnt11156_1_, blk_with_stfd_cnt_1_, bd_w_adr_c_plus_1_3_, 
        bd_w_adr_r_plus_1_1_, bd_sd_adr_4_, bd_w_adr_r_plus_1_3_, n598_30_, 
        bd_mem_au_count11744_6_, n598_29_, stfd_byt_cnt11156_3_, 
        bd_w_adr_c_plus_1_1_, blk_with_stfd_cnt_3_, bd_bm_count_32b11622_13_, 
        blk_with_stfd_cnt_7_, bd_w_adr_c_plus_1_5_, stfd_byt_cnt11156_12_, 
        stfd_byt_cnt11156_7_, bd_w_adr_r_plus_1_7_, bd_sd_adr_9_, 
        bd_mem_au_count11744_2_, bd_cpu_ack_cnt11656_2_, bd_au_count11668_2_, 
        n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12486, n12487, 
        n12488, n12489, n12490, n12491, n12492, n12494, n12495, n12496, n12498, 
        n12499, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, 
        n12509, n12511, n12513, n12514, n12515, n12516, n12517, n12518, n12519, 
        n12520, n12521, n12523, n12526, n12527, n12528, n12529, n12530, n12532, 
        n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, 
        n12542, n12545, n12546, n12547, n12549, n12550, n12553, n12554, n12555, 
        n12557, n12559, n12561, n12564, n12565, n12566, n12568, n12570, n12575, 
        n12577, n12578, n12579, n12580, n12582, n12583, n12586, n12588, n12591, 
        n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, 
        n12618, n12619, n12621, n12622, n12624, n12625, n12641, n12652, n12655, 
        n12656, n12658, n12659, n12660, n12661, n12662, n12663, n12668, n12669, 
        n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, 
        n12679, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, 
        n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, 
        n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, 
        n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, 
        n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, 
        n12725, n12726, n12727, n12728, n12730, n12762, n12763, n12766, n12771, 
        n12776, n12780, n12797, n12798, n12799, n12800, n12801, n12802, n12803, 
        n12804, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, 
        n12843, n12868, n12869, n12871, n12873, n12875, n12877, n12879, n12881, 
        n12883, n12885, n12888, n12897, n12899, n12904, n12906, n12909, n12912, 
        n12915, n12919, n12920, n12921, n12922, n12923, n12925, n12926, n12927, 
        n12930, n12931, n12936, n12938, n12939, n12940, n12943, n12944, n12945, 
        n12946, n12947, n12948, n12949, n12950, n12952, n12955, n12956, n12957, 
        n12959, n12960, n12965, n12966, n12967, n12971, n12972, n12973, n12975, 
        n12976, n12977, n12978, n12979, n12980, n12981, n12983, n12984, n12985, 
        n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12998, 
        n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, 
        n13008, n13009, n13010, n13011, n13013, n13014, n13015, n13016, n13017, 
        n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, 
        n13028, n13029, n13030, n13032, n13033, n13034, n13035, n13036, n13040, 
        n13042, n13043, n13045, n13046, n13047, n13048, n13049, n13050, n13051, 
        n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13064, n13065, 
        n13066, n13068, n13070, n13071, n13072, n13074, n13075, n13076, n13078, 
        n13079, n13080, n13081, n13082, n13083, n13085, n13086, n13088, n13089, 
        n13090, n13091, n13094, n13095, n13097, n13098, n13099, n13101, n13102, 
        n13103, n13104, n13105, n13106, n13107, n13109, n13112, n13113, n13115, 
        n13116, n13117, n13118, n13120, n13122, n13124, n13125, n13126, n13127, 
        n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, 
        n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, 
        n13146, n13147, n13148, n13151, n13153, n13154, n13156, n13157, n13158, 
        n13159, n13160, n13161, n13162, n13163, n13165, n13166, n13167, n13168, 
        n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, 
        n13178, n13179, n13191, n13192, n13193, n13194, n13195, n13198, n13200, 
        n13201, n13202, n13204, n13205, n13206, n13208, n13209, n13211, n13212, 
        n13217, n13219, n13220, n13223, n13224, n13227, n13229, n13230, n13231, 
        n13232, n13234, n13235, n13236, n13237, n13241, n13243, n13244, n13247, 
        n13249, n13250, n13252, n13256, n13257, n13258, n13261, n13262, n13263, 
        n13264, n13265, n13266, n13268, n13271, n13272, n13274, n13275, n13276, 
        n13277, n13279, n13280, n13281, n13283, n13284, n13285, n13286, n13290, 
        n13292, n13293, n13295, n13299, n13300, n13301, n13302, n13303, n13304, 
        n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, 
        n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, 
        n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, 
        n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, 
        n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, 
        n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, 
        n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, 
        n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, 
        n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, 
        n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, 
        n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, 
        n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, 
        n13413, n13414, n13415, gt_278_n15, gt_278_n16, gt_278_n20, gt_278_n22, 
        gt_278_n24, gt_278_n28, gt_278_n30, gt_278_n32, gt_278_n33, gt_278_n34, 
        gt_278_n35, gt_278_n36, gt_278_n37, gt_278_n38, gt_278_n39, gt_278_n40, 
        gt_278_n41, gt_278_n42, gt_278_n43, gt_278_n44, gt_278_n45, gt_278_n46, 
        gt_278_n47, gt_278_n48, gt_278_n49, gt_278_n50, gt_278_n51, 
        gte_275_2_n65, gte_275_2_n66, add_465_carry_9_, add_465_carry_4_, 
        add_465_carry_2_, add_465_carry_6_, add_465_carry_12_, 
        add_465_carry_11_, add_465_carry_10_, add_465_carry_8_, 
        add_465_carry_7_, add_465_carry_3_, add_465_carry_5_, add_465_carry_1_, 
        add_304_carry_4_, add_304_carry_2_, add_304_carry_3_, add_304_carry_5_, 
        add_510_carry_4_, add_510_carry_2_, add_510_carry_3_, add_510_carry_5_, 
        sub_275_n71, sub_275_n90, sub_275_n94, sub_275_n95, sub_275_n99, 
        sub_275_n100, sub_275_n102, sub_275_n104, sub_275_n105, sub_275_n106, 
        sub_275_n107, sub_275_n108, sub_275_n109, sub_275_n110, sub_513_n73, 
        sub_513_n74, sub_513_n78, sub_513_n80, sub_526_n82, sub_526_n83, 
        sub_526_n84, sub_526_n88, sub_526_n89, sub_526_n116, sub_526_n118, 
        sub_526_n119, sub_526_n120, lt_285_n121, sub_478_n123, sub_478_n124, 
        sub_478_n125, sub_478_n126, sub_478_n127, sub_478_n129, sub_478_n131, 
        sub_478_n133, sub_478_n139, sub_478_n143, sub_478_n145, sub_478_n147, 
        sub_478_n150, gte_275_n152, gte_275_n155, gte_275_n156, 
        add_303_carry_4_, add_303_carry_2_, add_303_carry_3_, add_303_carry_5_, 
        add_277_carry_9_, add_277_carry_4_, add_277_carry_2_, 
        add_277_carry_13_, add_277_carry_6_, add_277_carry_11_, 
        add_277_carry_10_, add_277_carry_12_, add_277_carry_8_, 
        add_277_carry_7_, add_277_carry_3_, add_277_carry_5_, add_301_carry_9_, 
        add_301_carry_4_, add_301_carry_2_, add_301_carry_6_, 
        add_301_carry_10_, add_301_carry_7_, add_301_carry_3_, 
        add_301_carry_8_, add_301_carry_5_, add_491_carry_4_, add_491_carry_2_, 
        add_491_carry_3_, add_491_carry_5_, add_475_carry_9_, add_475_carry_4_, 
        add_475_carry_2_, add_475_carry_6_, add_475_carry_13_, 
        add_475_carry_11_, add_475_carry_10_, add_475_carry_14_, 
        add_475_carry_12_, add_475_carry_7_, add_475_carry_3_, 
        add_475_carry_8_, add_475_carry_5_, sub_275_2_n159, sub_275_2_n180, 
        sub_275_2_n185, sub_275_2_n188, sub_275_2_n191, sub_275_2_n197, 
        sub_275_2_n199, sub_275_2_n200, sub_275_2_n203, gte_274_2_n163, 
        gte_274_2_n165, gte_274_2_n166, gte_274_2_n167, gte_274_n169, 
        gte_274_n173, gte_274_n174, gte_274_n175, add_302_carry_9_, 
        add_302_carry_4_, add_302_carry_2_, add_302_carry_6_, 
        add_302_carry_10_, add_302_carry_7_, add_302_carry_3_, 
        add_302_carry_8_, add_302_carry_5_, n13445, n13446, n13447, n13449, 
        n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, 
        n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13472, n13473, 
        n13474, n13483, n13485, n13486, n13487, n13488, n13490, n13491, n13492, 
        n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, 
        n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, 
        n13511, n13512, n13513, n13514, n13515, n13517, n13518, n13519, n13520, 
        n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, 
        n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, 
        n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, 
        n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, 
        n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, 
        n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, 
        n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, 
        n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, 
        n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, 
        n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, 
        n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, 
        n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, 
        n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, 
        n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, 
        n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13656, 
        n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, 
        n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, 
        n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, 
        n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, 
        n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, 
        n13702, n13703, n13704, n13705;
    dfctnq1 stfd_byt_cnt_reg_6_ ( .d(stfd_byt_cnt11156_6_), .cp(ck54), .cdn(
        n12516), .q(bd_stfd_byt_cnt[6]) );
    dfctnq1 stfd_byt_cnt_reg_8_ ( .d(stfd_byt_cnt11156_8_), .cp(ck54), .cdn(
        n12610), .q(bd_stfd_byt_cnt[8]) );
    dfctnq1 stfd_byt_cnt_reg_4_ ( .d(stfd_byt_cnt11156_4_), .cp(ck54), .cdn(
        n12611), .q(bd_stfd_byt_cnt[4]) );
    dfctnq1 stfd_byt_cnt_reg_0_ ( .d(stfd_byt_cnt11156_0_), .cp(ck54), .cdn(
        n12519), .q(bd_stfd_byt_cnt[0]) );
    dfctnq1 stfd_byt_cnt_reg_3_ ( .d(stfd_byt_cnt11156_3_), .cp(ck54), .cdn(
        n12613), .q(bd_stfd_byt_cnt[3]) );
    dfctnq1 stfd_byt_cnt_reg_1_ ( .d(stfd_byt_cnt11156_1_), .cp(ck54), .cdn(
        n12617), .q(bd_stfd_byt_cnt[1]) );
    dfctnq1 bd_cpu_ack_cnt_reg_2_ ( .d(n13339), .cp(ck54), .cdn(n12516), .q(
        bd_cpu_ack_cnt[2]) );
    nd02e1 U4071 ( .a1(n12478), .b1(n12514), .zn(n13116) );
    // or03d1 U4072 ( .a1(n13023), .a2(n12549), .a3(n13021), .z(n12478) );
    an03d1 U4072 ( .a1(n13023), .a2(n12549), .a3(n13021), .z(n12478) );  // change
    nr02d1 U4077 ( .a1(bd_mem_au_count[4]), .a2(bd_mem_au_count[3]), .zn(
        n13103) );
    mx21d1 U4078 ( .i0(n12480), .i1(n13659), .s(n12915), .z(n13369) );
    an02d1 U4079 ( .a1(bd_dt_ava), .a2(n13660), .z(n12480) );
    mi21d1 U4082 ( .i0(bd_sd_dat_27_), .i1(n12482), .s(n13704), .zn(n12539) );
    in01d1 U4083 ( .i(n13383), .zn(n12482) );
    mi21d1 U4084 ( .i0(n12484), .i1(n12483), .s(n13704), .zn(n12555) );
    nd03d1 U4085 ( .a1(n13389), .a2(n13387), .a3(n13390), .zn(n12483) );
    or03d1 U4086 ( .a1(bd_sd_dat_20_), .a2(bd_sd_dat_21_), .a3(bd_sd_dat_23_), 
        .z(n12484) );
    nd02d1 U4087 ( .a1(bd_seq_hdr_exist), .a2(n13122), .zn(n13231) );
    an02d1 U4090 ( .a1(n12957), .a2(n12565), .z(n12956) );
    mx21d1 U4092 ( .i0(bp_jpg_enc_end_adr[2]), .i1(bp_jpg_dec_end_adr[2]), .s( n13295), .z(n13126) );
    mx21d1 U4093 ( .i0(bp_jpg_enc_end_adr[6]), .i1(bp_jpg_dec_end_adr[6]), .s(
        n13295), .z(n13136) );
    mx21d1 U4094 ( .i0(bp_jpg_enc_end_adr[7]), .i1(bp_jpg_dec_end_adr[7]), .s(
        n13295), .z(n13130) );
    mx21d1 U4095 ( .i0(bp_jpg_enc_end_adr[3]), .i1(bp_jpg_dec_end_adr[3]), .s(
        n13295), .z(n13128) );
    mx21d1 U4096 ( .i0(bp_jpg_enc_end_adr[5]), .i1(bp_jpg_dec_end_adr[5]), .s(
        n13295), .z(n13134) );
    mx21d1 U4097 ( .i0(bp_jpg_enc_end_adr[0]), .i1(bp_jpg_dec_end_adr[0]), .s(
        n13295), .z(n13138) );
    mx21d1 U4098 ( .i0(bp_jpg_enc_end_adr[1]), .i1(bp_jpg_dec_end_adr[1]), .s(
        n13295), .z(n13140) );
    mx21d1 U4099 ( .i0(bp_jpg_enc_end_adr[4]), .i1(bp_jpg_dec_end_adr[4]), .s(
        n13295), .z(n13132) );
    mi21d1 U4100 ( .i0(n12487), .i1(bd_sd_dat_3_), .s(n13286), .zn(n12486) );
    in01d1 U4101 ( .i(n12486), .zn(n13010) );
    in01d1 U4102 ( .i(n13407), .zn(n12487) );
    mi21d1 U4103 ( .i0(n12999), .i1(n13403), .s(n12582), .zn(n12998) );
    mi21d1 U4104 ( .i0(bd_sd_dat_18_), .i1(n12488), .s(n13705), .zn(n12515) );
    in01d1 U4105 ( .i(n13392), .zn(n12488) );
    nr02d1 U4106 ( .a1(n12489), .a2(n13076), .zn(n12537) );
    nd02d1 U4109 ( .a1(n12490), .a2(n13112), .zn(n13172) );
    aon21d1 U4110 ( .a1(n12491), .a2(n12575), .b(n12971), .z(n12490) );
    or02d1 U4111 ( .a1(n12559), .a2(n13004), .z(n13112) );
    in01d1 U4116 ( .i(n13076), .zn(n13078) );
    oan22d1 U4118 ( .a1(n13124), .a2(n12663), .b1(n13542), .b2(n13116), .z(
        n12492) );
    dfctnq1 bd_wee_red_adv_reg ( .d(n13377), .cp(ck54), .cdn(n12612), .q(
        bd_wee_red_adv) );
    oan21d1 U4124 ( .a1(n12494), .a2(n13117), .b(n13244), .z(n12975) );
    oai21d1 U4125 ( .a1(n12541), .a2(n12663), .b(n13085), .zn(n12494) );
    aon211d1 U4127 ( .a1(bd_au_state[0]), .a2(n13117), .b(n13118), .c(n12495), 
        .z(n12977) );
    oan211d1 U4128 ( .a1(n13411), .a2(n13120), .b(bd_gop_hdr_exist), .c(n12965
        ), .z(n12495) );
    nd02d1 U4130 ( .a1(n12496), .a2(n12532), .zn(n12946) );
    nd02d1 U4131 ( .a1(n12945), .a2(n12762), .zn(n12496) );
    nd02d1 U4132 ( .a1(d_acc_unit), .a2(n13091), .zn(n13094) );
    mx21d1 U4135 ( .i0(n12498), .i1(n13258), .s(bl_v_jpg_q), .z(n13050) );
    nd02d1 U4137 ( .a1(n13256), .a2(n13048), .zn(n13047) );
    mx21d1 U4138 ( .i0(n12499), .i1(n13056), .s(bl_v_jpg_q), .z(n13058) );
    oai21d1 U4140 ( .a1(n12762), .a2(n13051), .b(n12502), .zn(n13057) );
    or04d1 U4143 ( .a1(n13539), .a2(bd_cpu_ack_cnt[2]), .a3(n12501), .a4(
        n13105), .z(n13227) );
    nd02d1 U4145 ( .a1(bd_cpu_ack_cnt[1]), .a2(bd_cpu_ack_cnt[3]), .zn(n12501)
         );
    an03d1 U4146 ( .a1(n13045), .a2(n12696), .a3(n13046), .z(n12502) );
    an04d1 U4148 ( .a1(n13102), .a2(n13099), .a3(n13103), .a4(n13104), .z(
        n12503) );
    in01d1 U4149 ( .i(n12503), .zn(n13097) );
    an02d1 U4150 ( .a1(n12946), .a2(n12532), .z(n12504) );
    in01d1 U4152 ( .i(n12946), .zn(n13059) );
    mx21d1 U4153 ( .i0(bd_au_count11668_5_), .i1(bd_au_count11677_5_), .s(
        n13272), .z(n12871) );
    mx21d1 U4154 ( .i0(bd_au_count11668_4_), .i1(bd_au_count11677_4_), .s(
        n13272), .z(n12873) );
    mx21d1 U4156 ( .i0(bd_au_count11668_3_), .i1(bd_au_count11677_3_), .s(
        n13272), .z(n12875) );
    mx21d1 U4157 ( .i0(bd_au_count11668_2_), .i1(bd_au_count11677_2_), .s(
        n13272), .z(n12877) );
    an02d1 U4160 ( .a1(n12959), .a2(n12696), .z(n12506) );
    oai22h1 U4161 ( .a1(n12780), .a2(n12813), .b1(n12507), .b2(
        bd_w_adr_r_plus_1_2_), .zn(n13307) );
    aon22d1 U4162 ( .a1(n13691), .a2(n13257), .b1(n12507), .b2(
        bd_w_adr_r_plus_1_1_), .z(n13308) );
    oai22h1 U4163 ( .a1(n12776), .a2(n12813), .b1(n12507), .b2(n12776), .zn(
        n13309) );
    oai21d1 U4164 ( .a1(n12763), .a2(n13040), .b(n12502), .zn(n12813) );
    an03d1 U4165 ( .a1(n12502), .a2(n12813), .a3(n13050), .z(n12507) );
    an03d1 U4193 ( .a1(n12502), .a2(n13057), .a3(n13058), .z(n12533) );
    in01d1 U4194 ( .i(n13057), .zn(n12944) );
    in01d1 U4196 ( .i(n12883), .zn(n12508) );
    nr02d1 U4197 ( .a1(p_mem_pic), .a2(n13095), .zn(n12509) );
    oai22h1 U4199 ( .a1(n12906), .a2(n13672), .b1(n13671), .b2(n13274), .zn(
        n13358) );
    nd02e1 U4205 ( .a1(n12621), .b1(bt_pulse4), .zn(n12915) );
    nr02d1 U4207 ( .a1(n13101), .a2(n12763), .zn(n12511) );
    nd02d1 U4209 ( .a1(n12763), .a2(n12502), .zn(n12912) );
    oan21d1 U4210 ( .a1(n13048), .a2(n13051), .b(n13256), .z(n12530) );
    an02d1 U4211 ( .a1(n13293), .a2(stfd_byt_cnt11157_7_), .z(
        stfd_byt_cnt11156_7_) );
    an02d1 U4212 ( .a1(n13293), .a2(stfd_byt_cnt11157_5_), .z(
        stfd_byt_cnt11156_5_) );
    an02d1 U4213 ( .a1(n13293), .a2(stfd_byt_cnt11157_2_), .z(
        stfd_byt_cnt11156_2_) );
    nd02d1 U4214 ( .a1(n13293), .a2(b_cpu_ack), .zn(n13106) );
    dfctnq1 bd_mem_en_reg ( .d(n13361), .cp(ck54), .cdn(n12609), .q(bd_mem_en)
         );
    nd02d1 U4217 ( .a1(n12586), .a2(n12663), .zn(n13217) );
    or03d1 U4218 ( .a1(n13390), .a2(n13389), .a3(n13387), .z(n13166) );
    nd03d1 U4219 ( .a1(bd_sd_dat_23_), .a2(bd_sd_dat_20_), .a3(bd_sd_dat_21_), 
        .zn(n13165) );
    or02d1 U4220 ( .a1(bd_sd_dat_29_), .a2(bd_sd_dat_28_), .z(n13160) );
    mi21d1 U4227 ( .i0(n13009), .i1(n13406), .s(n13704), .zn(n13008) );
    mi21d1 U4228 ( .i0(n13007), .i1(n13405), .s(n12582), .zn(n13006) );
    mi21d1 U4229 ( .i0(n13030), .i1(n13398), .s(bl_v_dec_mod), .zn(n13029) );
    an02d1 U4230 ( .a1(n12521), .a2(n12547), .z(n13036) );
    ni01d2 U4231 ( .i(bd_bm_count_32b[8]), .z(bd_bm_count[7]) );
    nd02e1 U4241 ( .a1(n13032), .b1(n13013), .zn(n13086) );
    nd02e1 U4245 ( .a1(n13019), .b1(n12528), .zn(n13277) );
    aon31d1 U4250 ( .a1(n13223), .a2(n13236), .a3(n12542), .b(n12976), .z(
        n13271) );
    an03d1 U4251 ( .a1(n13139), .a2(n13137), .a3(n13178), .z(n13179) );
    xn02d1 U4252 ( .a1(bd_w_adr_r_4_), .a2(n13140), .zn(n13139) );
    xn02d1 U4253 ( .a1(bd_w_adr_r_3_), .a2(n13138), .zn(n13137) );
    an03d1 U4254 ( .a1(bd_w_adr_r_1_), .a2(bd_w_adr_r_0_), .a3(bd_w_adr_r_2_), 
        .z(n13178) );
    an03d1 U4255 ( .a1(n13127), .a2(n13125), .a3(n13129), .z(n13176) );
    xn02d1 U4256 ( .a1(bd_w_adr_r_6_), .a2(n13128), .zn(n13127) );
    xn02d1 U4257 ( .a1(bd_w_adr_r_5_), .a2(n13126), .zn(n13125) );
    xn02d1 U4258 ( .a1(bd_w_adr_r_10_), .a2(n13130), .zn(n13129) );
    an03d1 U4259 ( .a1(n13133), .a2(n13131), .a3(n13135), .z(n13177) );
    xn02d1 U4260 ( .a1(bd_w_adr_r_8_), .a2(n13134), .zn(n13133) );
    xn02d1 U4261 ( .a1(bd_w_adr_r_7_), .a2(n13132), .zn(n13131) );
    xn02d1 U4262 ( .a1(bd_w_adr_r_9_), .a2(n13136), .zn(n13135) );
    nr03d2 U4264 ( .a1(bd_w_adr_r_10_), .a2(bd_w_adr_r_4_), .a3(bd_w_adr_r_3_), 
        .zn(n13153) );
    an03d1 U4267 ( .a1(n13148), .a2(n13147), .a3(n13193), .z(n13194) );
    xn02d1 U4268 ( .a1(bd_r_adr_r_9_), .a2(n13136), .zn(n13148) );
    xn02d1 U4269 ( .a1(bd_r_adr_r_5_), .a2(n13126), .zn(n13147) );
    an03d1 U4270 ( .a1(bd_r_adr_r_0_), .a2(bd_r_adr_r_1_), .a3(bd_r_adr_r_2_), 
        .z(n13193) );
    an03d1 U4271 ( .a1(n13142), .a2(n13141), .a3(n13143), .z(n13191) );
    xn02d1 U4272 ( .a1(bd_r_adr_r_8_), .a2(n13134), .zn(n13142) );
    xn02d1 U4273 ( .a1(bd_r_adr_r_6_), .a2(n13128), .zn(n13141) );
    xn02d1 U4274 ( .a1(bd_r_adr_r_10_), .a2(n13130), .zn(n13143) );
    an03d1 U4275 ( .a1(n13145), .a2(n13144), .a3(n13146), .z(n13192) );
    xn02d1 U4276 ( .a1(bd_r_adr_r_7_), .a2(n13132), .zn(n13145) );
    xn02d1 U4277 ( .a1(bd_r_adr_r_4_), .a2(n13140), .zn(n13144) );
    xn02d1 U4278 ( .a1(bd_r_adr_r_3_), .a2(n13138), .zn(n13146) );
    nr03d2 U4280 ( .a1(bd_r_adr_r_6_), .a2(bd_r_adr_r_4_), .a3(bd_r_adr_r_3_), 
        .zn(n13156) );
    nd02e1 U4282 ( .a1(bd_r_adr_r_10_), .b1(bd_r_adr_r_8_), .zn(n13195) );
    an03d1 U4284 ( .a1(bd_w_adr_c_3_), .a2(bd_w_adr_c_2_), .a3(bd_w_adr_c_4_), 
        .z(n13042) );
    an03d1 U4286 ( .a1(bd_r_adr_c_3_), .a2(bd_r_adr_c_2_), .a3(bd_r_adr_c_4_), 
        .z(n13053) );
    xn02d1 U4288 ( .a1(bl_v_jpg_q), .a2(bl_v_jpg), .zn(n13045) );
    mi21d1 U4289 ( .i0(n13001), .i1(n13409), .s(n12582), .zn(n13000) );
    nd02d1 U4292 ( .a1(n12503), .a2(d_acc_unit), .zn(n12960) );
    nd02d1 U4293 ( .a1(n13081), .a2(n13283), .zn(n12983) );
    nd02e1 U4295 ( .a1(n13247), .b1(n12976), .zn(n13283) );
    nd02e1 U4298 ( .a1(n13542), .b1(n12586), .zn(n13122) );
    in01d1 U4299 ( .i(n13122), .zn(n13124) );
    mi21d1 U4301 ( .i0(n13171), .i1(n13172), .s(n13411), .zn(n13170) );
    aon21d1 U4302 ( .a1(n13237), .a2(n13115), .b(n13074), .z(n13280) );
    nd02e1 U4304 ( .a1(n13411), .b1(bd_au_state[1]), .zn(n13074) );
    nd02d1 U4305 ( .a1(bd_au_state[1]), .a2(n13411), .zn(n12976) );
    in01d1 U4306 ( .i(n12976), .zn(n13244) );
    in01d1 U4309 ( .i(n13281), .zn(n13118) );
    nd02e1 U4310 ( .a1(n12973), .b1(n12575), .zn(n13281) );
    nd03d1 U4316 ( .a1(n13177), .a2(n13176), .a3(n13179), .zn(n13258) );
    nd03d1 U4317 ( .a1(n13192), .a2(n13191), .a3(n13194), .zn(n13056) );
    or02d1 U4320 ( .a1(n12622), .a2(p_mem_pic), .z(n13098) );
    nd02e1 U4321 ( .a1(n13292), .b1(n12883), .zn(n13095) );
    nd02e1 U4324 ( .a1(bl_v_jpg_q), .b1(n12502), .zn(n13048) );
    nr02e1 U4326 ( .a1(bd_active_once), .b1(bd_underflow), .zn(n12985) );
    an02d1 U4327 ( .a1(n13412), .a2(bd_we_dec_adv), .z(n13230) );
    an02d1 U4329 ( .a1(bd_bs_req_lt), .a2(bd_re_enc_adv), .z(n12943) );
    aon31d1 U4331 ( .a1(n13285), .a2(n13284), .a3(n13249), .b(n12659), .z(
        n12656) );
    aon221d1 U4351 ( .a1(bd_bm_count_32b11622_13_), .a2(n12504), .b1(
        bd_bm_count_32b11631_13_), .b2(n12505), .c(n12843), .z(n13322) );
    nd02e1 U4379 ( .a1(n12662), .b1(bd_au_state[1]), .zn(n12660) );
    nd02e1 U4382 ( .a1(n12513), .b1(br_buf_valid), .zn(n12938) );
    oai22d2 U4390 ( .a1(n12661), .a2(n12659), .b1(n12662), .b2(n12663), .zn(
        bd_gop_hdr_exist11082) );
    aoi221d1 U4391 ( .a1(n12977), .a2(n12978), .b1(n12979), .b2(n12980), .c(
        n12975), .zn(n12661) );
    or02d1 U4392 ( .a1(n12621), .a2(n13415), .z(n12659) );
    nd02d1 U4394 ( .a1(bd_bm_count_32b11631_0_), .a2(n12505), .zn(n12868) );
    nd02d1 U4395 ( .a1(bd_bm_count_32b11631_0_), .a2(n12504), .zn(n12869) );
    nd02e1 U4396 ( .a1(n12536), .b1(n13204), .zn(n13268) );
    in01d1 U4401 ( .i(n13094), .zn(n13272) );
    nd02d1 U4403 ( .a1(bd_w_adr_r_plus_1_10_), .a2(n12507), .zn(n12798) );
    nd02d1 U4405 ( .a1(bd_w_adr_r_plus_1_9_), .a2(n12507), .zn(n12800) );
    nd02d1 U4407 ( .a1(bd_w_adr_r_plus_1_8_), .a2(n12507), .zn(n12802) );
    nd02d1 U4409 ( .a1(bd_w_adr_r_plus_1_7_), .a2(n12507), .zn(n12804) );
    nd02d1 U4411 ( .a1(bd_w_adr_r_plus_1_6_), .a2(n12507), .zn(n12806) );
    nd02d1 U4413 ( .a1(bd_w_adr_r_plus_1_5_), .a2(n12507), .zn(n12808) );
    nd02d1 U4415 ( .a1(bd_w_adr_r_plus_1_4_), .a2(n12507), .zn(n12810) );
    nd02d1 U4417 ( .a1(bd_w_adr_r_plus_1_3_), .a2(n12507), .zn(n12812) );
    in01d1 U4418 ( .i(n12813), .zn(n13257) );
    in01d1 U4425 ( .i(n12988), .zn(n13261) );
    in01d1 U4427 ( .i(n12989), .zn(n13262) );
    in01d1 U4429 ( .i(n12990), .zn(n13263) );
    in01d1 U4431 ( .i(n12991), .zn(n13264) );
    in01d1 U4433 ( .i(n12992), .zn(n13265) );
    in01d1 U4436 ( .i(n12993), .zn(n13266) );
    aon31d1 U4442 ( .a1(bd_mem_en), .a2(n13097), .a3(d_acc_unit), .b(n13098), 
        .z(n12883) );
    nd02d1 U4450 ( .a1(p_out_sta), .a2(n12535), .zn(n12904) );
    mx21d1 U4452 ( .i0(bl_v_jpg), .i1(n13674), .s(n12624), .z(n13356) );
    in01d1 U4458 ( .i(n12925), .zn(n13205) );
    aon31d1 U4459 ( .a1(n13275), .a2(n13229), .a3(n13276), .b(n13106), .z(
        n12927) );
    nd02e1 U4461 ( .a1(n12939), .b1(bl_v_dec_mod), .zn(n12925) );
    nd02d1 U4463 ( .a1(n13274), .a2(n13656), .zn(n12930) );
    in01d1 U4464 ( .i(e_cd_en), .zn(n13107) );
    in01d1 U4469 ( .i(n12909), .zn(n13274) );
    aoi21d2 U4471 ( .a1(n12939), .a2(n12940), .b(n13292), .zn(n13378) );
    nd02e1 U4472 ( .a1(n13412), .b1(p_bs_req), .zn(n12939) );
    nd02e1 U4473 ( .a1(bt_pulse4), .b1(n13230), .zn(n12940) );
    in01d1 U4493 ( .i(s_sd_dat[31]), .zn(n12695) );
    in01d1 U4494 ( .i(s_sd_dat[30]), .zn(n12694) );
    in01d1 U4495 ( .i(s_sd_dat[29]), .zn(n12693) );
    in01d1 U4496 ( .i(s_sd_dat[28]), .zn(n12692) );
    in01d1 U4497 ( .i(s_sd_dat[27]), .zn(n12691) );
    in01d1 U4498 ( .i(s_sd_dat[26]), .zn(n12690) );
    in01d1 U4499 ( .i(s_sd_dat[25]), .zn(n12689) );
    in01d1 U4500 ( .i(s_sd_dat[24]), .zn(n12688) );
    in01d1 U4501 ( .i(s_sd_dat[23]), .zn(n12687) );
    in01d1 U4502 ( .i(s_sd_dat[22]), .zn(n12686) );
    in01d1 U4503 ( .i(s_sd_dat[21]), .zn(n12685) );
    in01d1 U4504 ( .i(s_sd_dat[20]), .zn(n12684) );
    in01d1 U4505 ( .i(s_sd_dat[19]), .zn(n12683) );
    in01d1 U4506 ( .i(s_sd_dat[18]), .zn(n12682) );
    in01d1 U4507 ( .i(s_sd_dat[17]), .zn(n12681) );
    in01d1 U4509 ( .i(s_sd_dat[15]), .zn(n12679) );
    in01d1 U4510 ( .i(s_sd_dat[14]), .zn(n12678) );
    in01d1 U4511 ( .i(s_sd_dat[13]), .zn(n12677) );
    in01d1 U4512 ( .i(s_sd_dat[12]), .zn(n12676) );
    in01d1 U4513 ( .i(s_sd_dat[11]), .zn(n12675) );
    in01d1 U4514 ( .i(s_sd_dat[10]), .zn(n12674) );
    in01d1 U4515 ( .i(s_sd_dat[9]), .zn(n12673) );
    in01d1 U4516 ( .i(s_sd_dat[8]), .zn(n12672) );
    in01d1 U4517 ( .i(s_sd_dat[7]), .zn(n12671) );
    in01d1 U4518 ( .i(s_sd_dat[6]), .zn(n12670) );
    in01d1 U4519 ( .i(s_sd_dat[5]), .zn(n12669) );
    in01d1 U4520 ( .i(s_sd_dat[4]), .zn(n12668) );
    in01d1 U4525 ( .i(p_bs_dat[31]), .zn(n12728) );
    in01d1 U4526 ( .i(p_bs_dat[30]), .zn(n12727) );
    in01d1 U4527 ( .i(p_bs_dat[29]), .zn(n12726) );
    in01d1 U4528 ( .i(p_bs_dat[28]), .zn(n12725) );
    in01d1 U4529 ( .i(p_bs_dat[27]), .zn(n12724) );
    in01d1 U4530 ( .i(p_bs_dat[26]), .zn(n12723) );
    in01d1 U4531 ( .i(p_bs_dat[25]), .zn(n12722) );
    in01d1 U4532 ( .i(p_bs_dat[24]), .zn(n12721) );
    in01d1 U4533 ( .i(p_bs_dat[23]), .zn(n12720) );
    in01d1 U4534 ( .i(p_bs_dat[22]), .zn(n12719) );
    in01d1 U4535 ( .i(p_bs_dat[21]), .zn(n12718) );
    in01d1 U4536 ( .i(p_bs_dat[20]), .zn(n12717) );
    in01d1 U4537 ( .i(p_bs_dat[19]), .zn(n12716) );
    in01d1 U4538 ( .i(p_bs_dat[18]), .zn(n12715) );
    in01d1 U4539 ( .i(p_bs_dat[17]), .zn(n12714) );
    in01d1 U4540 ( .i(p_bs_dat[16]), .zn(n12713) );
    in01d1 U4541 ( .i(p_bs_dat[15]), .zn(n12712) );
    in01d1 U4542 ( .i(p_bs_dat[14]), .zn(n12711) );
    in01d1 U4543 ( .i(p_bs_dat[13]), .zn(n12710) );
    in01d1 U4544 ( .i(p_bs_dat[12]), .zn(n12709) );
    in01d1 U4545 ( .i(p_bs_dat[11]), .zn(n12708) );
    in01d1 U4546 ( .i(p_bs_dat[10]), .zn(n12707) );
    in01d1 U4547 ( .i(p_bs_dat[9]), .zn(n12706) );
    in01d1 U4548 ( .i(p_bs_dat[8]), .zn(n12705) );
    in01d1 U4549 ( .i(p_bs_dat[7]), .zn(n12704) );
    in01d1 U4551 ( .i(p_bs_dat[6]), .zn(n12703) );
    in01d1 U4554 ( .i(p_bs_dat[5]), .zn(n12702) );
    in01d1 U4555 ( .i(p_bs_dat[4]), .zn(n12701) );
    in01d1 U4556 ( .i(p_bs_dat[3]), .zn(n12700) );
    in01d1 U4558 ( .i(p_bs_dat[2]), .zn(n12699) );
    in01d1 U4559 ( .i(p_bs_dat[1]), .zn(n12698) );
    in01d1 U4560 ( .i(p_bs_dat[0]), .zn(n12697) );
    ni01d2 U4618 ( .i(n12609), .z(n12612) );
    ni01d2 U4627 ( .i(n12609), .z(n12614) );
    ni01d2 U4633 ( .i(n12610), .z(n12616) );
    ni01d2 U4638 ( .i(n12610), .z(n12615) );
    ni01d2 U4642 ( .i(n12610), .z(n12618) );
    aoi21d2 U4643 ( .a1(n12762), .a2(n12763), .b(n12619), .zn(b_sd_en11058) );
    nd02e1 U4644 ( .a1(n13054), .b1(n13055), .zn(n12762) );
    nd02e1 U4645 ( .a1(n12529), .b1(n13043), .zn(n12763) );
    in01d1 U4647 ( .i(n12763), .zn(n12945) );
    in01d1 U4648 ( .i(n13106), .zn(bd_cpu_ack_dly11086) );
    ni01d2 U4651 ( .i(n12609), .z(n12613) );
    an02d1 U4652 ( .a1(bd_underflow), .a2(n12696), .z(bd_underflow_prev11094)
         );
    in01d1 U4653 ( .i(bt_rst), .zn(n12696) );
    nd03d1 U4657 ( .a1(bd_mem_en), .a2(n12503), .a3(d_acc_unit), .zn(n13175)
         );
    dfctnqn1 bd_au_state_reg_0_ ( .d(bd_au_state11074_0_), .cp(ck54), .cdn(
        n12519), .qn(n13411) );
    in01d1 U4660 ( .i(n13411), .zn(bd_au_state[0]) );
    dfctnq1 bd_bm_count_32b_reg_2_ ( .d(n13333), .cp(ck54), .cdn(n12516), .q(
        bd_bm_count[1]) );
    in01d1 U4669 ( .i(bd_w_adr_r_2_), .zn(n12780) );
    in01d1 U4671 ( .i(bd_w_adr_r_0_), .zn(n12776) );
    in01d1 U4688 ( .i(bd_chk_seq_end), .zn(n12920) );
    in01d1 U4691 ( .i(bd_w_adr_c_4_), .zn(n12771) );
    in01d1 U4693 ( .i(n13654), .zn(n12766) );
    in01d1 U4696 ( .i(bd_sd_dat_31_), .zn(n13020) );
    in01d1 U4698 ( .i(bd_sd_dat_19_), .zn(n13014) );
    in01d1 U4699 ( .i(bd_sd_dat_17_), .zn(n13016) );
    in01d1 U4700 ( .i(bd_sd_dat_16_), .zn(n13033) );
    in01d1 U4701 ( .i(bd_sd_dat_15_), .zn(n13028) );
    in01d1 U4702 ( .i(bd_sd_dat_13_), .zn(n13026) );
    in01d1 U4703 ( .i(bd_sd_dat_10_), .zn(n13022) );
    in01d1 U4704 ( .i(bd_sd_dat_6_), .zn(n13003) );
    in01d1 U4705 ( .i(bd_sd_dat_5_), .zn(n13007) );
    in01d1 U4706 ( .i(bd_sd_dat_4_), .zn(n13009) );
    in01d1 U4707 ( .i(bd_sd_dat_2_), .zn(n13005) );
    in01d1 U4708 ( .i(bd_sd_dat_1_), .zn(n13001) );
    in01d1 U4710 ( .i(n13380), .zn(n13159) );
    in01d1 U4711 ( .i(n13385), .zn(n13071) );
    in01d1 U4712 ( .i(n13388), .zn(n13158) );
    in01d1 U4713 ( .i(n13412), .zn(bd_cpu_req_lt) );
    in01d1 U4714 ( .i(n13413), .zn(bd_overflow_prev) );
    in01d1 U4715 ( .i(n13414), .zn(b_cpu_req) );
    or02d1 U4716 ( .a1(bd_au_state[1]), .a2(n13411), .z(n13082) );
    nr02d1 U4718 ( .a1(bt_pulse6), .a2(bd_wee_red_adv), .zn(n12513) );
    an04d1 U4719 ( .a1(n13029), .a2(n13025), .a3(n13027), .a4(n12545), .z(
        n12514) );
    dfctnq1 bd_bm_count_32b_reg_14_ ( .d(n13321), .cp(ck54), .cdn(n12611), .q(
        bd_bm_count_32b[14]) );
    dfctnq1 bd_bm_count_32b_reg_9_ ( .d(n13326), .cp(ck54), .cdn(n12617), .q(
        bd_bm_count[8]) );
    dfctnq1 bd_bm_count_32b_reg_4_ ( .d(n13331), .cp(ck54), .cdn(n12610), .q(
        bd_bm_count[3]) );
    ni01d2 U4737 ( .i(n12609), .z(n12516) );
    ni01d2 U4738 ( .i(n12609), .z(n12517) );
    ni01d2 U4739 ( .i(p_rst_x), .z(n12609) );
    ni01d2 U4740 ( .i(n12609), .z(n12611) );
    ni01d2 U4741 ( .i(n12610), .z(n12518) );
    ni01d2 U4742 ( .i(n12610), .z(n12519) );
    ni01d2 U4743 ( .i(p_rst_x), .z(n12610) );
    ni01d2 U4744 ( .i(n12610), .z(n12617) );
    ni01d2 U4745 ( .i(v_dec_mod), .z(n13295) );
    mi21d1 U4747 ( .i0(n13580), .i1(bp_jpg_dec_sta_adr[4]), .s(n13295), .zn(
        n12989) );
    mi21d1 U4749 ( .i0(n13581), .i1(bp_jpg_dec_sta_adr[5]), .s(n13295), .zn(
        n12988) );
    mi21d1 U4751 ( .i0(n13579), .i1(bp_jpg_dec_sta_adr[2]), .s(n13295), .zn(
        n12991) );
    mi21d1 U4752 ( .i0(n13577), .i1(bp_jpg_dec_sta_adr[0]), .s(n13295), .zn(
        n12993) );
    mi21d1 U4753 ( .i0(n13578), .i1(bp_jpg_dec_sta_adr[1]), .s(n13295), .zn(
        n12992) );
    xn02d1 U4754 ( .a1(n13705), .a2(v_dec_mod), .zn(n13046) );
    dfctnq1 bd_bm_count_32b_reg_13_ ( .d(n13322), .cp(ck54), .cdn(n12517), .q(
        bd_bm_count[12]) );
    dfctnq1 bd_bm_count_32b_reg_3_ ( .d(n13332), .cp(ck54), .cdn(p_rst_x), .q(
        bd_bm_count[2]) );
    dfctnq1 bd_bm_count_32b_reg_5_ ( .d(n13330), .cp(ck54), .cdn(n12615), .q(
        bd_bm_count[4]) );
    dfctnq1 bd_bm_count_32b_reg_12_ ( .d(n13323), .cp(ck54), .cdn(n12611), .q(
        bd_bm_count[11]) );
    dfctnq1 bd_bm_count_32b_reg_6_ ( .d(n13329), .cp(ck54), .cdn(n12618), .q(
        bd_bm_count[5]) );
    dfctnq1 bd_bm_count_32b_reg_1_ ( .d(n13334), .cp(ck54), .cdn(n12611), .q(
        bd_bm_count_32b[1]) );
    dfctnq1 bd_bm_count_32b_reg_11_ ( .d(n13324), .cp(ck54), .cdn(n12517), .q(
        bd_bm_count_32b[11]) );
    dfctnq1 bd_bm_count_32b_reg_7_ ( .d(n13328), .cp(ck54), .cdn(n12518), .q(
        bd_bm_count[6]) );
    dfctnq1 bd_au_state_reg_1_ ( .d(bd_au_state11074_1_), .cp(ck54), .cdn(
        n12614), .q(bd_au_state[1]) );
    dfctnq1 bd_bm_count_32b_reg_10_ ( .d(n13325), .cp(ck54), .cdn(n12614), .q(
        bd_bm_count[9]) );
    dfctnq1 bd_bm_count_32b_reg_8_ ( .d(n13327), .cp(ck54), .cdn(n12616), .q(
        bd_bm_count_32b[8]) );
    in01d1 U4756 ( .i(bd_wee_red_adv), .zn(n13109) );
    mi21d1 U4757 ( .i0(n12943), .i1(bd_wee_red_adv), .s(bl_v_dec_mod), .zn(
        n13054) );
    dfctnq2 bd_cpu_ack_cnt_reg_1_ ( .d(n13340), .cp(ck54), .cdn(n12618), .q(
        bd_cpu_ack_cnt[1]) );
    nr02d1 U4758 ( .a1(bd_cpu_ack_cnt[0]), .a2(bd_cpu_ack_cnt[3]), .zn(n13201)
         );
    dfctnq2 bd_cpu_ack_cnt_reg_3_ ( .d(n13338), .cp(ck54), .cdn(n12612), .q(
        bd_cpu_ack_cnt[3]) );
    mi21d1 U4759 ( .i0(n13286), .i1(n13105), .s(bd_cpu_ack_cnt[3]), .zn(n13276
        ) );
    dfctnq2 bd_mem_au_count_reg_4_ ( .d(n13350), .cp(ck54), .cdn(n12614), .q(
        bd_mem_au_count[4]) );
    dfctnq2 bd_au_count_reg_5_ ( .d(n13342), .cp(ck54), .cdn(n12614), .q(
        bd_au_count[5]) );
    in01d1 U4772 ( .i(bd_au_count[4]), .zn(n12888) );
    dfctnq2 bd_au_count_reg_4_ ( .d(n13343), .cp(ck54), .cdn(n12615), .q(
        bd_au_count[4]) );
    in01d1 U4774 ( .i(bd_mem_au_count[0]), .zn(n13099) );
    dfctnq2 bd_mem_au_count_reg_0_ ( .d(n13354), .cp(ck54), .cdn(n12613), .q(
        bd_mem_au_count[0]) );
    in01d1 U4777 ( .i(bd_seq_hdr_exist), .zn(n12971) );
    dfctnq2 bd_seq_hdr_exist_reg ( .d(bd_seq_hdr_exist11078), .cp(ck54), .cdn(
        n12615), .q(bd_seq_hdr_exist) );
    in01d1 U4779 ( .i(bd_gop_hdr_exist), .zn(n12663) );
    nr02d1 U4780 ( .a1(bd_gop_hdr_exist), .a2(n13019), .zn(n12957) );
    aoi21d2 U4781 ( .a1(bd_gop_hdr_exist), .a2(n13529), .b(n12538), .zn(n12973
        ) );
    dfctnq2 bd_gop_hdr_exist_reg ( .d(bd_gop_hdr_exist11082), .cp(ck54), .cdn(
        n12517), .q(bd_gop_hdr_exist) );
    dfctnq2 bd_bm_count_32b_reg_0_ ( .d(n13335), .cp(ck54), .cdn(n12617), .q(
        bd_bm_count_32b[0]) );
    in01d1 U4784 ( .i(bd_cpu_ack_cnt[0]), .zn(n13105) );
    mi21d1 U4785 ( .i0(bd_cpu_ack_cnt[0]), .i1(n12582), .s(bd_cpu_ack_cnt[1]), 
        .zn(n13275) );
    dfctnq2 bd_cpu_ack_cnt_reg_0_ ( .d(n13341), .cp(ck54), .cdn(p_rst_x), .q(
        bd_cpu_ack_cnt[0]) );
    dfctnq2 bd_au_count_reg_3_ ( .d(n13344), .cp(ck54), .cdn(n12618), .q(
        bd_au_count[3]) );
    dfctnq2 bd_au_count_reg_2_ ( .d(n13345), .cp(ck54), .cdn(n12518), .q(
        bd_au_count[2]) );
    in01d1 U4791 ( .i(bd_au_count[1]), .zn(n12897) );
    dfctnq2 bd_au_count_reg_1_ ( .d(n13346), .cp(ck54), .cdn(n12519), .q(
        bd_au_count[1]) );
    dfctnq2 bd_au_count_reg_0_ ( .d(n13347), .cp(ck54), .cdn(n12517), .q(
        bd_au_count[0]) );
    mi21d1 U4794 ( .i0(n13026), .i1(n13397), .s(n12582), .zn(n13025) );
    nd02d1 U4797 ( .a1(n13032), .a2(n13015), .zn(n13089) );
    mi21d1 U4801 ( .i0(bd_sd_dat_26_), .i1(n12520), .s(n13705), .zn(n12523) );
    in01d1 U4802 ( .i(n13384), .zn(n12520) );
    mi21d1 U4804 ( .i0(n12526), .i1(bd_sd_dat_24_), .s(n13286), .zn(n12579) );
    in01d1 U4809 ( .i(n13386), .zn(n12526) );
    mx21d1 U4815 ( .i0(n13030), .i1(n13398), .s(n12582), .z(n12527) );
    in01d1 U4816 ( .i(bd_sd_dat_12_), .zn(n13030) );
    or02d1 U4817 ( .a1(n13080), .a2(n12984), .z(n13079) );
    mx21d1 U4819 ( .i0(n13036), .i1(n13035), .s(n13019), .z(n12528) );
    oan32d1 U4826 ( .a1(n13168), .a2(n13080), .a3(n12984), .b1(n13088), .b2(
        n12515), .z(n13167) );
    nd04d1 U4828 ( .a1(n13220), .a3(n13219), .a4(n12553), .a2(n12577), .zn(
        n13083) );
    mi21d1 U4832 ( .i0(n13503), .i1(n13502), .s(bl_v_dec_mod), .zn(bd_dt_ava)
         );
    oan21d1 U4833 ( .a1(n12945), .a2(n12762), .b(n12696), .z(n12532) );
    aoi211d1 U4835 ( .a1(n12502), .a2(n13056), .b(n12944), .c(n13047), .zn(
        n12534) );
    ni01d2 U4836 ( .i(n12730), .z(n13290) );
    ni01d2 U4837 ( .i(n12730), .z(n12625) );
    an04d1 U4839 ( .a1(n13010), .a2(n13078), .a3(n12564), .a4(n13498), .z(
        n12538) );
    oan211d1 U4841 ( .a1(n13494), .a2(n12967), .b(n13232), .c(n13234), .z(
        n12541) );
    oan22d1 U4842 ( .a1(n13021), .a2(n13079), .b1(n12580), .b2(n13090), .z(
        n12542) );
    in01d1 U4843 ( .i(n13027), .zn(n13208) );
    mi21d1 U4844 ( .i0(bd_sd_dat_25_), .i1(n13071), .s(n13705), .zn(n13070) );
    mi21d1 U4845 ( .i0(n13028), .i1(n13395), .s(bl_v_dec_mod), .zn(n13027) );
    nd02e1 U4846 ( .a1(n13088), .b1(n12515), .zn(n13236) );
    in01d1 U4850 ( .i(bd_sd_dat_7_), .zn(n12999) );
    mi21d1 U4851 ( .i0(bd_sd_dat_14_), .i1(n12546), .s(n12582), .zn(n12545) );
    in01d1 U4852 ( .i(n13396), .zn(n12546) );
    in01d1 U4856 ( .i(bd_sd_dat_9_), .zn(n13024) );
    or02d1 U4859 ( .a1(n12591), .a2(n12659), .z(n12922) );
    in01d1 U4862 ( .i(n13399), .zn(n12550) );
    mi21d1 U4864 ( .i0(n13020), .i1(n13379), .s(n12582), .zn(n13019) );
    mi21d1 U4867 ( .i0(n13005), .i1(n13408), .s(n13705), .zn(n13004) );
    mi21d1 U4869 ( .i0(bd_sd_dat_22_), .i1(n13158), .s(n13704), .zn(n13219) );
    nr02e1 U4871 ( .a1(n12566), .b1(n13034), .zn(n12565) );
    an03d1 U4876 ( .a1(n12577), .a2(n12554), .a3(n12583), .z(n13234) );
    mi21d1 U4881 ( .i0(n13160), .i1(n13161), .s(n12582), .zn(n13209) );
    in01d1 U4893 ( .i(n12575), .zn(n12965) );
    in01d1 U4897 ( .i(bd_sd_dat_24_), .zn(n13017) );
    in01d1 U4901 ( .i(n12583), .zn(n13066) );
    aoi22h1 U4908 ( .a1(n12540), .a2(n13250), .b1(n12580), .b2(n13243), .zn(
        n13249) );
    in01d1 U4911 ( .i(n12580), .zn(n13081) );
    in01d1 U4916 ( .i(bd_au_state[1]), .zn(n12978) );
    ni01d2 U4918 ( .i(bd_bm_count[1]), .z(bd_bm_count_32b[2]) );
    ni01d2 U4920 ( .i(bd_bm_count[3]), .z(bd_bm_count_32b[4]) );
    ni01d2 U4921 ( .i(bd_bm_count[4]), .z(bd_bm_count_32b[5]) );
    ni01d2 U4922 ( .i(bd_bm_count[5]), .z(bd_bm_count_32b[6]) );
    ni01d2 U4923 ( .i(bd_bm_count[6]), .z(bd_bm_count_32b[7]) );
    ni01d2 U4925 ( .i(bd_bm_count[8]), .z(bd_bm_count_32b[9]) );
    ni01d2 U4926 ( .i(bd_bm_count[9]), .z(bd_bm_count_32b[10]) );
    ni01d2 U4928 ( .i(bd_bm_count[11]), .z(bd_bm_count_32b[12]) );
    ni01d2 U4929 ( .i(bd_bm_count[12]), .z(bd_bm_count_32b[13]) );
    nr02d1 U4931 ( .a1(n13292), .a2(n12641), .zn(bd_overflow_prev11090) );
    nr02d1 U4932 ( .a1(n12624), .a2(n13499), .zn(stfd_byt_cnt11156_0_) );
    nr02d1 U4939 ( .a1(n12621), .a2(n13541), .zn(stfd_byt_cnt11156_10_) );
    nr02d1 U4940 ( .a1(n13292), .a2(n13540), .zn(stfd_byt_cnt11156_11_) );
    nr02d1 U4941 ( .a1(n12624), .a2(n13501), .zn(stfd_byt_cnt11156_12_) );
    nr02d1 U4944 ( .a1(n13292), .a2(n12655), .zn(bd_seq_hdr_exist11078) );
    oai21d1 U4946 ( .a1(n12658), .a2(n12659), .b(n12660), .zn(
        bd_au_state11074_1_) );
    nr02d1 U4952 ( .a1(n12621), .a2(n12668), .zn(bd_sd_dat11062_4_) );
    nr02d1 U4953 ( .a1(n13292), .a2(n12669), .zn(bd_sd_dat11062_5_) );
    nr02d1 U4954 ( .a1(n12624), .a2(n12670), .zn(bd_sd_dat11062_6_) );
    nr02d1 U4955 ( .a1(n12622), .a2(n12671), .zn(bd_sd_dat11062_7_) );
    nr02d1 U4956 ( .a1(n13292), .a2(n12672), .zn(bd_sd_dat11062_8_) );
    nr02d1 U4957 ( .a1(n12619), .a2(n12673), .zn(bd_sd_dat11062_9_) );
    nr02d1 U4958 ( .a1(n12622), .a2(n12674), .zn(bd_sd_dat11062_10_) );
    nr02d1 U4959 ( .a1(n12624), .a2(n12675), .zn(bd_sd_dat11062_11_) );
    nr02d1 U4960 ( .a1(n12619), .a2(n12676), .zn(bd_sd_dat11062_12_) );
    nr02d1 U4961 ( .a1(n12621), .a2(n12677), .zn(bd_sd_dat11062_13_) );
    nr02d1 U4962 ( .a1(n13292), .a2(n12678), .zn(bd_sd_dat11062_14_) );
    nr02d1 U4963 ( .a1(n13292), .a2(n12679), .zn(bd_sd_dat11062_15_) );
    nr02d1 U4965 ( .a1(n13292), .a2(n12681), .zn(bd_sd_dat11062_17_) );
    nr02d1 U4966 ( .a1(n12619), .a2(n12682), .zn(bd_sd_dat11062_18_) );
    nr02d1 U4967 ( .a1(n12622), .a2(n12683), .zn(bd_sd_dat11062_19_) );
    nr02d1 U4968 ( .a1(n12624), .a2(n12684), .zn(bd_sd_dat11062_20_) );
    nr02d1 U4969 ( .a1(n13292), .a2(n12685), .zn(bd_sd_dat11062_21_) );
    nr02d1 U4970 ( .a1(n12621), .a2(n12686), .zn(bd_sd_dat11062_22_) );
    nr02d1 U4971 ( .a1(n13292), .a2(n12687), .zn(bd_sd_dat11062_23_) );
    nr02d1 U4972 ( .a1(n12624), .a2(n12688), .zn(bd_sd_dat11062_24_) );
    nr02d1 U4973 ( .a1(n12622), .a2(n12689), .zn(bd_sd_dat11062_25_) );
    nr02d1 U4974 ( .a1(n12622), .a2(n12690), .zn(bd_sd_dat11062_26_) );
    nr02d1 U4975 ( .a1(n12619), .a2(n12691), .zn(bd_sd_dat11062_27_) );
    nr02d1 U4976 ( .a1(n13292), .a2(n12692), .zn(bd_sd_dat11062_28_) );
    nr02d1 U4977 ( .a1(n12624), .a2(n12693), .zn(bd_sd_dat11062_29_) );
    nr02d1 U4978 ( .a1(n12621), .a2(n12694), .zn(bd_sd_dat11062_30_) );
    nr02d1 U4979 ( .a1(n12622), .a2(n12695), .zn(bd_sd_dat11062_31_) );
    nr02d1 U4980 ( .a1(n12619), .a2(n12697), .zn(bd_bs_dat11066_0_) );
    nr02d1 U4981 ( .a1(n12619), .a2(n12698), .zn(bd_bs_dat11066_1_) );
    nr02d1 U4982 ( .a1(n12624), .a2(n12699), .zn(bd_bs_dat11066_2_) );
    nr02d1 U4983 ( .a1(n12622), .a2(n12700), .zn(bd_bs_dat11066_3_) );
    nr02d1 U4984 ( .a1(n13292), .a2(n12701), .zn(bd_bs_dat11066_4_) );
    nr02d1 U4985 ( .a1(n12624), .a2(n12702), .zn(bd_bs_dat11066_5_) );
    nr02d1 U4986 ( .a1(n12621), .a2(n12703), .zn(bd_bs_dat11066_6_) );
    nr02d1 U4987 ( .a1(n12619), .a2(n12704), .zn(bd_bs_dat11066_7_) );
    nr02d1 U4988 ( .a1(n12619), .a2(n12705), .zn(bd_bs_dat11066_8_) );
    nr02d1 U4989 ( .a1(n12621), .a2(n12706), .zn(bd_bs_dat11066_9_) );
    nr02d1 U4990 ( .a1(n12624), .a2(n12707), .zn(bd_bs_dat11066_10_) );
    nr02d1 U4991 ( .a1(n12621), .a2(n12708), .zn(bd_bs_dat11066_11_) );
    nr02d1 U4992 ( .a1(n12622), .a2(n12709), .zn(bd_bs_dat11066_12_) );
    nr02d1 U4993 ( .a1(n12619), .a2(n12710), .zn(bd_bs_dat11066_13_) );
    nr02d1 U4994 ( .a1(n12619), .a2(n12711), .zn(bd_bs_dat11066_14_) );
    nr02d1 U4995 ( .a1(n12621), .a2(n12712), .zn(bd_bs_dat11066_15_) );
    nr02d1 U4996 ( .a1(n13292), .a2(n12713), .zn(bd_bs_dat11066_16_) );
    nr02d1 U4997 ( .a1(n12624), .a2(n12714), .zn(bd_bs_dat11066_17_) );
    nr02d1 U4998 ( .a1(n12621), .a2(n12715), .zn(bd_bs_dat11066_18_) );
    nr02d1 U4999 ( .a1(n12619), .a2(n12716), .zn(bd_bs_dat11066_19_) );
    nr02d1 U5000 ( .a1(n12619), .a2(n12717), .zn(bd_bs_dat11066_20_) );
    nr02d1 U5001 ( .a1(n12622), .a2(n12718), .zn(bd_bs_dat11066_21_) );
    nr02d1 U5002 ( .a1(n12619), .a2(n12719), .zn(bd_bs_dat11066_22_) );
    nr02d1 U5003 ( .a1(n12621), .a2(n12720), .zn(bd_bs_dat11066_23_) );
    nr02d1 U5004 ( .a1(n12621), .a2(n12721), .zn(bd_bs_dat11066_24_) );
    nr02d1 U5005 ( .a1(n12624), .a2(n12722), .zn(bd_bs_dat11066_25_) );
    nr02d1 U5006 ( .a1(n13292), .a2(n12723), .zn(bd_bs_dat11066_26_) );
    nr02d1 U5007 ( .a1(n12622), .a2(n12724), .zn(bd_bs_dat11066_27_) );
    nr02d1 U5008 ( .a1(n12624), .a2(n12725), .zn(bd_bs_dat11066_28_) );
    nr02d1 U5009 ( .a1(n12621), .a2(n12726), .zn(bd_bs_dat11066_29_) );
    nr02d1 U5010 ( .a1(n12622), .a2(n12727), .zn(bd_bs_dat11066_30_) );
    nr02d1 U5011 ( .a1(n12619), .a2(n12728), .zn(bd_bs_dat11066_31_) );
    nd02d1 U5012 ( .a1(n12797), .a2(n12798), .zn(n13299) );
    nd02d1 U5013 ( .a1(n12799), .a2(n12800), .zn(n13300) );
    nd02d1 U5014 ( .a1(n12801), .a2(n12802), .zn(n13301) );
    nd02d1 U5015 ( .a1(n12803), .a2(n12804), .zn(n13302) );
    nd02d1 U5017 ( .a1(n12807), .a2(n12808), .zn(n13304) );
    nd02d1 U5018 ( .a1(n12809), .a2(n12810), .zn(n13305) );
    nd02d1 U5019 ( .a1(n12811), .a2(n12812), .zn(n13306) );
    oai21d1 U5031 ( .a1(n12919), .a2(n13665), .b(n12921), .zn(n13365) );
    nd02d1 U5032 ( .a1(n12922), .a2(n12923), .zn(n13366) );
    oai211d1 U5034 ( .a1(n12624), .a2(n12925), .b(n12926), .c(n12927), .zn(
        n13368) );
    oai211d1 U5035 ( .a1(n12906), .a2(n13500), .b(n12930), .c(n12530), .zn(
        n13372) );
    nd02d1 U5036 ( .a1(n12922), .a2(n12931), .zn(n13373) );
    nr02d1 U5039 ( .a1(n12622), .a2(n12936), .zn(n13376) );
    nr02e1 U5041 ( .a1(bd_cpu_ack_cnt11656_4_), .b1(n12947), .zn(n13337) );
    nr02e1 U5042 ( .a1(bd_cpu_ack_cnt11656_3_), .b1(n12947), .zn(n13338) );
    nr02e1 U5043 ( .a1(bd_cpu_ack_cnt11656_2_), .b1(n12947), .zn(n13339) );
    nr02e1 U5044 ( .a1(bd_cpu_ack_cnt11656_1_), .b1(n12947), .zn(n13340) );
    nd02d1 U5053 ( .a1(n13382), .a2(n13381), .zn(n13161) );
    nr02d1 U5060 ( .a1(n13023), .a2(n13021), .zn(n13064) );
    nr02d1 U5062 ( .a1(n13013), .a2(n13015), .zn(n13068) );
    nr02d1 U5071 ( .a1(bd_mem_au_count[6]), .a2(bd_mem_au_count[5]), .zn(
        n13104) );
    nd02d1 U5073 ( .a1(n12502), .a2(n13040), .zn(n13101) );
    nr02d1 U5074 ( .a1(n12621), .a2(d_seq_end), .zn(n12921) );
    nd02d1 U5076 ( .a1(n12535), .a2(n13583), .zn(n12652) );
    nr02d1 U5077 ( .a1(n13032), .a2(n13498), .zn(n13241) );
    nd02d1 U5078 ( .a1(n12491), .a2(n13244), .zn(n13243) );
    nr02d1 U5080 ( .a1(bd_au_state[1]), .a2(n13411), .zn(n13247) );
    in01d1 U5090 ( .i(n13074), .zn(n12979) );
    nd02d1 U5096 ( .a1(b_seq_end), .a2(n12619), .zn(n12923) );
    oai21d1 U5098 ( .a1(n12624), .a2(n13107), .b(bd_cpu_end), .zn(n12931) );
    oai21d1 U5099 ( .a1(n13113), .a2(n13235), .b(n13244), .zn(n13279) );
    mi21d1 U5101 ( .i0(n13109), .i1(n13151), .s(bl_v_dec_mod), .zn(n13043) );
    mi21d1 U5102 ( .i0(n13522), .i1(n12579), .s(n12539), .zn(n13162) );
    oai211d1 U5103 ( .a1(bd_au_state[1]), .a2(n13170), .b(n13279), .c(n13280), 
        .zn(n13173) );
    dfctnq1 b_sd_adr_reg_2_ ( .d(1'b0), .cp(ck54), .cdn(n12617), .q(b_sd_adr
        [2]) );
    dfctnq1 b_sd_adr_reg_1_ ( .d(1'b0), .cp(ck54), .cdn(n12516), .q(b_sd_adr
        [1]) );
    dfctnq1 b_sd_adr_reg_0_ ( .d(1'b0), .cp(ck54), .cdn(n12618), .q(b_sd_adr
        [0]) );
    dfctnq1 bd_w_adr_r_reg_10_ ( .d(n13299), .cp(ck54), .cdn(n12609), .q(
        bd_w_adr_r_10_) );
    dfctnq1 bd_w_adr_r_reg_9_ ( .d(n13300), .cp(ck54), .cdn(n12612), .q(
        bd_w_adr_r_9_) );
    dfctnq1 bd_w_adr_r_reg_8_ ( .d(n13301), .cp(ck54), .cdn(n12618), .q(
        bd_w_adr_r_8_) );
    dfctnq1 bd_w_adr_r_reg_7_ ( .d(n13302), .cp(ck54), .cdn(n12517), .q(
        bd_w_adr_r_7_) );
    dfctnq1 bd_w_adr_r_reg_6_ ( .d(n13303), .cp(ck54), .cdn(n12615), .q(
        bd_w_adr_r_6_) );
    dfctnq1 bd_w_adr_r_reg_5_ ( .d(n13304), .cp(ck54), .cdn(n12609), .q(
        bd_w_adr_r_5_) );
    dfctnq1 bd_w_adr_r_reg_4_ ( .d(n13305), .cp(ck54), .cdn(n12611), .q(
        bd_w_adr_r_4_) );
    dfctnq1 bd_w_adr_r_reg_3_ ( .d(n13306), .cp(ck54), .cdn(n12517), .q(
        bd_w_adr_r_3_) );
    dfctnq1 bd_w_adr_r_reg_2_ ( .d(n13307), .cp(ck54), .cdn(n12517), .q(
        bd_w_adr_r_2_) );
    dfctnq1 bd_w_adr_r_reg_1_ ( .d(n13308), .cp(ck54), .cdn(n12615), .q(
        bd_w_adr_r_1_) );
    dfctnq1 bd_w_adr_r_reg_0_ ( .d(n13309), .cp(ck54), .cdn(n12618), .q(
        bd_w_adr_r_0_) );
    dfctnq1 bd_r_adr_r_reg_10_ ( .d(n13310), .cp(ck54), .cdn(n12517), .q(
        bd_r_adr_r_10_) );
    dfctnq1 bd_r_adr_r_reg_9_ ( .d(n13311), .cp(ck54), .cdn(n12614), .q(
        bd_r_adr_r_9_) );
    dfctnq1 bd_r_adr_r_reg_8_ ( .d(n13312), .cp(ck54), .cdn(n12617), .q(
        bd_r_adr_r_8_) );
    dfctnq1 bd_r_adr_r_reg_7_ ( .d(n13313), .cp(ck54), .cdn(n12611), .q(
        bd_r_adr_r_7_) );
    dfctnq1 bd_r_adr_r_reg_6_ ( .d(n13314), .cp(ck54), .cdn(n12519), .q(
        bd_r_adr_r_6_) );
    dfctnq1 bd_r_adr_r_reg_5_ ( .d(n13315), .cp(ck54), .cdn(n12516), .q(
        bd_r_adr_r_5_) );
    dfctnq1 bd_r_adr_r_reg_4_ ( .d(n13316), .cp(ck54), .cdn(n12617), .q(
        bd_r_adr_r_4_) );
    dfctnq1 bd_r_adr_r_reg_3_ ( .d(n13317), .cp(ck54), .cdn(n12517), .q(
        bd_r_adr_r_3_) );
    dfctnq1 bd_r_adr_r_reg_2_ ( .d(n13318), .cp(ck54), .cdn(n12611), .q(
        bd_r_adr_r_2_) );
    dfctnq1 bd_r_adr_r_reg_1_ ( .d(n13319), .cp(ck54), .cdn(n12612), .q(
        bd_r_adr_r_1_) );
    dfctnq1 bd_r_adr_r_reg_0_ ( .d(n13320), .cp(ck54), .cdn(n12518), .q(
        bd_r_adr_r_0_) );
    dfctnq1 bd_cpu_ack_cnt_reg_5_ ( .d(n13336), .cp(ck54), .cdn(n12609), .q(
        bd_cpu_ack_cnt[5]) );
    dfctnq1 bd_cpu_ack_cnt_reg_4_ ( .d(n13337), .cp(ck54), .cdn(n12612), .q(
        bd_cpu_ack_cnt[4]) );
    dfctnq1 bd_mem_au_count_reg_6_ ( .d(n13348), .cp(ck54), .cdn(n12615), .q(
        bd_mem_au_count[6]) );
    dfctnq1 bd_mem_au_count_reg_5_ ( .d(n13349), .cp(ck54), .cdn(n12616), .q(
        bd_mem_au_count[5]) );
    dfctnq1 bd_mem_au_count_reg_3_ ( .d(n13351), .cp(ck54), .cdn(n12615), .q(
        bd_mem_au_count[3]) );
    dfctnq1 bd_mem_au_count_reg_2_ ( .d(n13352), .cp(ck54), .cdn(n12612), .q(
        bd_mem_au_count[2]) );
    dfctnq1 bd_mem_au_count_reg_1_ ( .d(n13353), .cp(ck54), .cdn(n12519), .q(
        bd_mem_au_count[1]) );
    dfctnq1 bd_active_once_reg ( .d(n13355), .cp(ck54), .cdn(n12617), .q(
        bd_active_once) );
    dfctnq1 bl_v_jpg_q_reg ( .d(n13356), .cp(ck54), .cdn(n12616), .q(
        bl_v_jpg_q) );
    dfptnq1 bd_r_adr_c_reg_2_ ( .d(n13357), .cp(ck54), .sdn(n12618), .q(
        bd_r_adr_c_2_) );
    dfctnq1 bd_r_adr_c_reg_0_ ( .d(n13358), .cp(ck54), .cdn(n12616), .q(
        bd_r_adr_c_0_) );
    dfctnq1 bd_r_adr_c_reg_4_ ( .d(n13359), .cp(ck54), .cdn(n12519), .q(
        bd_r_adr_c_4_) );
    dfptnq1 bd_w_adr_c_reg_5_ ( .d(n13360), .cp(ck54), .sdn(n12611), .q(
        bd_w_adr_c_5_) );
    dfctnq1 bd_bs_req_lt_reg ( .d(n13362), .cp(ck54), .cdn(n12612), .q(
        bd_bs_req_lt) );
    dfptnq1 bd_w_adr_c_reg_1_ ( .d(n13363), .cp(ck54), .sdn(n12615), .q(
        bd_w_adr_c_1_) );
    dfptnq1 bd_w_adr_c_reg_3_ ( .d(n13364), .cp(ck54), .sdn(n12614), .q(
        bd_w_adr_c_3_) );
    dfptnq1 bd_chk_seq_end_reg ( .d(n13365), .cp(ck54), .sdn(n12519), .q(
        bd_chk_seq_end) );
    dfctnq1 b_seq_end_reg ( .d(n13366), .cp(ck54), .cdn(n12611), .q(b_seq_end)
         );
    dfptnq1 bd_w_adr_c_reg_2_ ( .d(n13367), .cp(ck54), .sdn(n12616), .q(
        bd_w_adr_c_2_) );
    dfctnq1 b_cpu_ack_reg ( .d(n13368), .cp(ck54), .cdn(n12516), .q(b_cpu_ack)
         );
    dfctnq1 bd_re_enc_adv_reg ( .d(n13369), .cp(ck54), .cdn(n12616), .q(
        bd_re_enc_adv) );
    dfctnq1 bd_w_adr_c_reg_0_ ( .d(n13370), .cp(ck54), .cdn(n12518), .q(
        bd_w_adr_c_0_) );
    dfctnq1 bd_w_adr_c_reg_4_ ( .d(n13371), .cp(ck54), .cdn(n12610), .q(
        bd_w_adr_c_4_) );
    dfptnq1 bd_r_adr_c_reg_5_ ( .d(n13372), .cp(ck54), .sdn(n12613), .q(
        bd_r_adr_c_5_) );
    dfctnq1 bd_cpu_end_reg ( .d(n13373), .cp(ck54), .cdn(n12519), .q(
        bd_cpu_endb) );
    dfptnq1 bd_r_adr_c_reg_1_ ( .d(n13374), .cp(ck54), .sdn(n12614), .q(
        bd_r_adr_c_1_) );
    dfptnq1 bd_r_adr_c_reg_3_ ( .d(n13375), .cp(ck54), .sdn(n12612), .q(
        bd_r_adr_c_3_) );
    dfctnq1 b_dec_en_reg ( .d(n13376), .cp(ck54), .cdn(n12613), .q(b_dec_en)
         );
    dfctnq1 bd_we_dec_adv_reg ( .d(n13378), .cp(ck54), .cdn(n12609), .q(
        bd_we_dec_adv) );
    dfctnq1 b_sd_adr_reg_18_ ( .d(bd_sd_adr_18_), .cp(ck54), .cdn(n12518), .q(
        b_sd_adr[18]) );
    dfctnq1 b_sd_adr_reg_17_ ( .d(bd_sd_adr_17_), .cp(ck54), .cdn(n12616), .q(
        b_sd_adr[17]) );
    dfctnq1 b_sd_adr_reg_16_ ( .d(bd_sd_adr_16_), .cp(ck54), .cdn(p_rst_x), 
        .q(b_sd_adr[16]) );
    dfctnq1 b_sd_adr_reg_15_ ( .d(bd_sd_adr_15_), .cp(ck54), .cdn(n12519), .q(
        b_sd_adr[15]) );
    dfctnq1 b_sd_adr_reg_14_ ( .d(bd_sd_adr_14_), .cp(ck54), .cdn(n12518), .q(
        b_sd_adr[14]) );
    dfctnq1 b_sd_adr_reg_13_ ( .d(bd_sd_adr_13_), .cp(ck54), .cdn(n12611), .q(
        b_sd_adr[13]) );
    dfctnq1 b_sd_adr_reg_12_ ( .d(bd_sd_adr_12_), .cp(ck54), .cdn(n12613), .q(
        b_sd_adr[12]) );
    dfctnq1 b_sd_adr_reg_11_ ( .d(bd_sd_adr_11_), .cp(ck54), .cdn(p_rst_x), 
        .q(b_sd_adr[11]) );
    dfctnq1 b_sd_adr_reg_10_ ( .d(bd_sd_adr_10_), .cp(ck54), .cdn(n12516), .q(
        b_sd_adr[10]) );
    dfctnq1 b_sd_adr_reg_9_ ( .d(bd_sd_adr_9_), .cp(ck54), .cdn(n12614), .q(
        b_sd_adr[9]) );
    dfctnq1 b_sd_adr_reg_8_ ( .d(bd_sd_adr_8_), .cp(ck54), .cdn(n12615), .q(
        b_sd_adr[8]) );
    dfctnq1 b_sd_adr_reg_7_ ( .d(bd_sd_adr_7_), .cp(ck54), .cdn(n12616), .q(
        b_sd_adr[7]) );
    dfctnq1 b_sd_adr_reg_6_ ( .d(bd_sd_adr_6_), .cp(ck54), .cdn(n12519), .q(
        b_sd_adr[6]) );
    dfctnq1 b_sd_adr_reg_5_ ( .d(bd_sd_adr_5_), .cp(ck54), .cdn(n12618), .q(
        b_sd_adr[5]) );
    dfctnq1 b_sd_adr_reg_4_ ( .d(bd_sd_adr_4_), .cp(ck54), .cdn(n12519), .q(
        b_sd_adr[4]) );
    dfctnq1 b_sd_adr_reg_3_ ( .d(bd_sd_adr_3_), .cp(ck54), .cdn(p_rst_x), .q(
        b_sd_adr[3]) );
    dfctnq1 bd_sd_dat_reg_31_ ( .d(bd_sd_dat11062_31_), .cp(ck54), .cdn(n12613
        ), .q(bd_sd_dat_31_) );
    dfctnq1 bd_sd_dat_reg_30_ ( .d(bd_sd_dat11062_30_), .cp(ck54), .cdn(n12613
        ), .q(bd_sd_dat_30_) );
    dfctnq1 bd_sd_dat_reg_29_ ( .d(bd_sd_dat11062_29_), .cp(ck54), .cdn(n12516
        ), .q(bd_sd_dat_29_) );
    dfctnq1 bd_sd_dat_reg_28_ ( .d(bd_sd_dat11062_28_), .cp(ck54), .cdn(n12614
        ), .q(bd_sd_dat_28_) );
    dfctnq1 bd_sd_dat_reg_27_ ( .d(bd_sd_dat11062_27_), .cp(ck54), .cdn(n12518
        ), .q(bd_sd_dat_27_) );
    dfctnq1 bd_sd_dat_reg_26_ ( .d(bd_sd_dat11062_26_), .cp(ck54), .cdn(n12616
        ), .q(bd_sd_dat_26_) );
    dfctnq1 bd_sd_dat_reg_25_ ( .d(bd_sd_dat11062_25_), .cp(ck54), .cdn(n12615
        ), .q(bd_sd_dat_25_) );
    dfctnq1 bd_sd_dat_reg_24_ ( .d(bd_sd_dat11062_24_), .cp(ck54), .cdn(n12519
        ), .q(bd_sd_dat_24_) );
    dfctnq1 bd_sd_dat_reg_23_ ( .d(bd_sd_dat11062_23_), .cp(ck54), .cdn(n12617
        ), .q(bd_sd_dat_23_) );
    dfctnq1 bd_sd_dat_reg_22_ ( .d(bd_sd_dat11062_22_), .cp(ck54), .cdn(n12611
        ), .q(bd_sd_dat_22_) );
    dfctnq1 bd_sd_dat_reg_21_ ( .d(bd_sd_dat11062_21_), .cp(ck54), .cdn(n12613
        ), .q(bd_sd_dat_21_) );
    dfctnq1 bd_sd_dat_reg_20_ ( .d(bd_sd_dat11062_20_), .cp(ck54), .cdn(n12613
        ), .q(bd_sd_dat_20_) );
    dfctnq1 bd_sd_dat_reg_19_ ( .d(bd_sd_dat11062_19_), .cp(ck54), .cdn(n12516
        ), .q(bd_sd_dat_19_) );
    dfctnq1 bd_sd_dat_reg_18_ ( .d(bd_sd_dat11062_18_), .cp(ck54), .cdn(n12614
        ), .q(bd_sd_dat_18_) );
    dfctnq1 bd_sd_dat_reg_17_ ( .d(bd_sd_dat11062_17_), .cp(ck54), .cdn(n12615
        ), .q(bd_sd_dat_17_) );
    dfctnq1 bd_sd_dat_reg_16_ ( .d(bd_sd_dat11062_16_), .cp(ck54), .cdn(n12616
        ), .q(bd_sd_dat_16_) );
    dfctnq1 bd_sd_dat_reg_15_ ( .d(bd_sd_dat11062_15_), .cp(ck54), .cdn(n12618
        ), .q(bd_sd_dat_15_) );
    dfctnq1 bd_sd_dat_reg_14_ ( .d(bd_sd_dat11062_14_), .cp(ck54), .cdn(n12618
        ), .q(bd_sd_dat_14_) );
    dfctnq1 bd_sd_dat_reg_13_ ( .d(bd_sd_dat11062_13_), .cp(ck54), .cdn(n12609
        ), .q(bd_sd_dat_13_) );
    dfctnq1 bd_sd_dat_reg_12_ ( .d(bd_sd_dat11062_12_), .cp(ck54), .cdn(
        p_rst_x), .q(bd_sd_dat_12_) );
    dfctnq1 bd_sd_dat_reg_11_ ( .d(bd_sd_dat11062_11_), .cp(ck54), .cdn(
        p_rst_x), .q(bd_sd_dat_11_) );
    dfctnq1 bd_sd_dat_reg_10_ ( .d(bd_sd_dat11062_10_), .cp(ck54), .cdn(n12517
        ), .q(bd_sd_dat_10_) );
    dfctnq1 bd_sd_dat_reg_9_ ( .d(bd_sd_dat11062_9_), .cp(ck54), .cdn(n12612), 
        .q(bd_sd_dat_9_) );
    dfctnq1 bd_sd_dat_reg_8_ ( .d(bd_sd_dat11062_8_), .cp(ck54), .cdn(n12614), 
        .q(bd_sd_dat_8_) );
    dfctnq1 bd_sd_dat_reg_7_ ( .d(bd_sd_dat11062_7_), .cp(ck54), .cdn(n12610), 
        .q(bd_sd_dat_7_) );
    dfctnq1 bd_sd_dat_reg_6_ ( .d(bd_sd_dat11062_6_), .cp(ck54), .cdn(n12616), 
        .q(bd_sd_dat_6_) );
    dfctnq1 bd_sd_dat_reg_5_ ( .d(bd_sd_dat11062_5_), .cp(ck54), .cdn(n12610), 
        .q(bd_sd_dat_5_) );
    dfctnq1 bd_sd_dat_reg_4_ ( .d(bd_sd_dat11062_4_), .cp(ck54), .cdn(n12617), 
        .q(bd_sd_dat_4_) );
    dfctnq1 bd_sd_dat_reg_3_ ( .d(bd_sd_dat11062_3_), .cp(ck54), .cdn(n12618), 
        .q(bd_sd_dat_3_) );
    dfctnq1 bd_sd_dat_reg_2_ ( .d(bd_sd_dat11062_2_), .cp(ck54), .cdn(n12516), 
        .q(bd_sd_dat_2_) );
    dfctnq1 bd_sd_dat_reg_1_ ( .d(bd_sd_dat11062_1_), .cp(ck54), .cdn(n12517), 
        .q(bd_sd_dat_1_) );
    dfctnq1 bd_sd_dat_reg_0_ ( .d(bd_sd_dat11062_0_), .cp(ck54), .cdn(n12610), 
        .q(bd_sd_dat_0_) );
    dfctnqn1 bd_bs_dat_reg_31_ ( .d(bd_bs_dat11066_31_), .cp(ck54), .cdn(
        n12517), .qn(n13379) );
    dfctnqn1 bd_bs_dat_reg_30_ ( .d(bd_bs_dat11066_30_), .cp(ck54), .cdn(
        n12517), .qn(n13380) );
    dfctnqn1 bd_bs_dat_reg_29_ ( .d(bd_bs_dat11066_29_), .cp(ck54), .cdn(
        n12618), .qn(n13381) );
    dfctnqn1 bd_bs_dat_reg_28_ ( .d(bd_bs_dat11066_28_), .cp(ck54), .cdn(
        n12518), .qn(n13382) );
    dfctnqn1 bd_bs_dat_reg_27_ ( .d(bd_bs_dat11066_27_), .cp(ck54), .cdn(
        n12617), .qn(n13383) );
    dfctnqn1 bd_bs_dat_reg_26_ ( .d(bd_bs_dat11066_26_), .cp(ck54), .cdn(
        n12518), .qn(n13384) );
    dfctnqn1 bd_bs_dat_reg_25_ ( .d(bd_bs_dat11066_25_), .cp(ck54), .cdn(
        n12609), .qn(n13385) );
    dfctnqn1 bd_bs_dat_reg_24_ ( .d(bd_bs_dat11066_24_), .cp(ck54), .cdn(
        n12516), .qn(n13386) );
    dfctnqn1 bd_bs_dat_reg_23_ ( .d(bd_bs_dat11066_23_), .cp(ck54), .cdn(
        n12611), .qn(n13387) );
    dfctnqn1 bd_bs_dat_reg_22_ ( .d(bd_bs_dat11066_22_), .cp(ck54), .cdn(
        n12611), .qn(n13388) );
    dfctnqn1 bd_bs_dat_reg_21_ ( .d(bd_bs_dat11066_21_), .cp(ck54), .cdn(
        n12612), .qn(n13389) );
    dfctnqn1 bd_bs_dat_reg_20_ ( .d(bd_bs_dat11066_20_), .cp(ck54), .cdn(
        n12610), .qn(n13390) );
    dfctnqn1 bd_bs_dat_reg_19_ ( .d(bd_bs_dat11066_19_), .cp(ck54), .cdn(
        n12617), .qn(n13391) );
    dfctnqn1 bd_bs_dat_reg_18_ ( .d(bd_bs_dat11066_18_), .cp(ck54), .cdn(
        n12519), .qn(n13392) );
    dfctnqn1 bd_bs_dat_reg_17_ ( .d(bd_bs_dat11066_17_), .cp(ck54), .cdn(
        n12615), .qn(n13393) );
    dfctnqn1 bd_bs_dat_reg_16_ ( .d(bd_bs_dat11066_16_), .cp(ck54), .cdn(
        n12618), .qn(n13394) );
    dfctnqn1 bd_bs_dat_reg_15_ ( .d(bd_bs_dat11066_15_), .cp(ck54), .cdn(
        n12610), .qn(n13395) );
    dfctnqn1 bd_bs_dat_reg_14_ ( .d(bd_bs_dat11066_14_), .cp(ck54), .cdn(
        n12612), .qn(n13396) );
    dfctnqn1 bd_bs_dat_reg_13_ ( .d(bd_bs_dat11066_13_), .cp(ck54), .cdn(
        n12612), .qn(n13397) );
    dfctnqn1 bd_bs_dat_reg_12_ ( .d(bd_bs_dat11066_12_), .cp(ck54), .cdn(
        n12517), .qn(n13398) );
    dfctnqn1 bd_bs_dat_reg_11_ ( .d(bd_bs_dat11066_11_), .cp(ck54), .cdn(
        n12609), .qn(n13399) );
    dfctnqn1 bd_bs_dat_reg_10_ ( .d(bd_bs_dat11066_10_), .cp(ck54), .cdn(
        n12613), .qn(n13400) );
    dfctnqn1 bd_bs_dat_reg_9_ ( .d(bd_bs_dat11066_9_), .cp(ck54), .cdn(n12519), 
        .qn(n13401) );
    dfctnqn1 bd_bs_dat_reg_8_ ( .d(bd_bs_dat11066_8_), .cp(ck54), .cdn(n12518), 
        .qn(n13402) );
    dfctnqn1 bd_bs_dat_reg_7_ ( .d(bd_bs_dat11066_7_), .cp(ck54), .cdn(n12610), 
        .qn(n13403) );
    dfctnqn1 bd_bs_dat_reg_6_ ( .d(bd_bs_dat11066_6_), .cp(ck54), .cdn(n12615), 
        .qn(n13404) );
    dfctnqn1 bd_bs_dat_reg_5_ ( .d(bd_bs_dat11066_5_), .cp(ck54), .cdn(n12518), 
        .qn(n13405) );
    dfctnqn1 bd_bs_dat_reg_4_ ( .d(bd_bs_dat11066_4_), .cp(ck54), .cdn(n12613), 
        .qn(n13406) );
    dfctnqn1 bd_bs_dat_reg_3_ ( .d(bd_bs_dat11066_3_), .cp(ck54), .cdn(n12516), 
        .qn(n13407) );
    dfctnqn1 bd_bs_dat_reg_2_ ( .d(bd_bs_dat11066_2_), .cp(ck54), .cdn(n12613), 
        .qn(n13408) );
    dfctnqn1 bd_bs_dat_reg_1_ ( .d(bd_bs_dat11066_1_), .cp(ck54), .cdn(p_rst_x
        ), .qn(n13409) );
    dfctnqn1 bd_bs_dat_reg_0_ ( .d(bd_bs_dat11066_0_), .cp(ck54), .cdn(n12611), 
        .qn(n13410) );
    dfctnq1 b_sd_dat_reg_31_ ( .d(b_sd_dat11070_31_), .cp(ck54), .cdn(n12612), 
        .q(b_sd_dat[31]) );
    dfctnq1 b_sd_dat_reg_30_ ( .d(b_sd_dat11070_30_), .cp(ck54), .cdn(n12614), 
        .q(b_sd_dat[30]) );
    dfctnq1 b_sd_dat_reg_29_ ( .d(b_sd_dat11070_29_), .cp(ck54), .cdn(n12610), 
        .q(b_sd_dat[29]) );
    dfctnq1 b_sd_dat_reg_28_ ( .d(b_sd_dat11070_28_), .cp(ck54), .cdn(n12616), 
        .q(b_sd_dat[28]) );
    dfctnq1 b_sd_dat_reg_27_ ( .d(b_sd_dat11070_27_), .cp(ck54), .cdn(n12617), 
        .q(b_sd_dat[27]) );
    dfctnq1 b_sd_dat_reg_26_ ( .d(b_sd_dat11070_26_), .cp(ck54), .cdn(n12617), 
        .q(b_sd_dat[26]) );
    dfctnq1 b_sd_dat_reg_25_ ( .d(b_sd_dat11070_25_), .cp(ck54), .cdn(n12609), 
        .q(b_sd_dat[25]) );
    dfctnq1 b_sd_dat_reg_24_ ( .d(b_sd_dat11070_24_), .cp(ck54), .cdn(n12516), 
        .q(b_sd_dat[24]) );
    dfctnq1 b_sd_dat_reg_23_ ( .d(b_sd_dat11070_23_), .cp(ck54), .cdn(n12613), 
        .q(b_sd_dat[23]) );
    dfctnq1 b_sd_dat_reg_22_ ( .d(b_sd_dat11070_22_), .cp(ck54), .cdn(n12516), 
        .q(b_sd_dat[22]) );
    dfctnq1 b_sd_dat_reg_21_ ( .d(b_sd_dat11070_21_), .cp(ck54), .cdn(n12612), 
        .q(b_sd_dat[21]) );
    dfctnq1 b_sd_dat_reg_20_ ( .d(b_sd_dat11070_20_), .cp(ck54), .cdn(n12614), 
        .q(b_sd_dat[20]) );
    dfctnq1 b_sd_dat_reg_19_ ( .d(b_sd_dat11070_19_), .cp(ck54), .cdn(n12618), 
        .q(b_sd_dat[19]) );
    dfctnq1 b_sd_dat_reg_18_ ( .d(b_sd_dat11070_18_), .cp(ck54), .cdn(n12616), 
        .q(b_sd_dat[18]) );
    dfctnq1 b_sd_dat_reg_17_ ( .d(b_sd_dat11070_17_), .cp(ck54), .cdn(n12518), 
        .q(b_sd_dat[17]) );
    dfctnq1 b_sd_dat_reg_16_ ( .d(b_sd_dat11070_16_), .cp(ck54), .cdn(n12519), 
        .q(b_sd_dat[16]) );
    dfctnq1 b_sd_dat_reg_15_ ( .d(b_sd_dat11070_15_), .cp(ck54), .cdn(n12615), 
        .q(b_sd_dat[15]) );
    dfctnq1 b_sd_dat_reg_14_ ( .d(b_sd_dat11070_14_), .cp(ck54), .cdn(n12613), 
        .q(b_sd_dat[14]) );
    dfctnq1 b_sd_dat_reg_13_ ( .d(b_sd_dat11070_13_), .cp(ck54), .cdn(p_rst_x), 
        .q(b_sd_dat[13]) );
    dfctnq1 b_sd_dat_reg_12_ ( .d(b_sd_dat11070_12_), .cp(ck54), .cdn(n12612), 
        .q(b_sd_dat[12]) );
    dfctnq1 b_sd_dat_reg_11_ ( .d(b_sd_dat11070_11_), .cp(ck54), .cdn(n12611), 
        .q(b_sd_dat[11]) );
    dfctnq1 b_sd_dat_reg_10_ ( .d(b_sd_dat11070_10_), .cp(ck54), .cdn(n12614), 
        .q(b_sd_dat[10]) );
    dfctnq1 b_sd_dat_reg_9_ ( .d(b_sd_dat11070_9_), .cp(ck54), .cdn(p_rst_x), 
        .q(b_sd_dat[9]) );
    dfctnq1 b_sd_dat_reg_8_ ( .d(b_sd_dat11070_8_), .cp(ck54), .cdn(n12616), 
        .q(b_sd_dat[8]) );
    dfctnq1 b_sd_dat_reg_7_ ( .d(b_sd_dat11070_7_), .cp(ck54), .cdn(n12617), 
        .q(b_sd_dat[7]) );
    dfctnq1 b_sd_dat_reg_6_ ( .d(b_sd_dat11070_6_), .cp(ck54), .cdn(n12617), 
        .q(b_sd_dat[6]) );
    dfctnq1 b_sd_dat_reg_5_ ( .d(b_sd_dat11070_5_), .cp(ck54), .cdn(n12518), 
        .q(b_sd_dat[5]) );
    dfctnq1 b_sd_dat_reg_4_ ( .d(b_sd_dat11070_4_), .cp(ck54), .cdn(n12612), 
        .q(b_sd_dat[4]) );
    dfctnq1 b_sd_dat_reg_3_ ( .d(b_sd_dat11070_3_), .cp(ck54), .cdn(n12613), 
        .q(b_sd_dat[3]) );
    dfctnq1 b_sd_dat_reg_2_ ( .d(b_sd_dat11070_2_), .cp(ck54), .cdn(n12611), 
        .q(b_sd_dat[2]) );
    dfctnq1 b_sd_dat_reg_1_ ( .d(b_sd_dat11070_1_), .cp(ck54), .cdn(n12517), 
        .q(b_sd_dat[1]) );
    dfctnq1 b_sd_dat_reg_0_ ( .d(b_sd_dat11070_0_), .cp(ck54), .cdn(n12614), 
        .q(b_sd_dat[0]) );
    dfctnq1 stfd_byt_cnt_reg_12_ ( .d(stfd_byt_cnt11156_12_), .cp(ck54), .cdn(
        n12518), .q(bd_stfd_byt_cnt[12]) );
    dfctnq1 stfd_byt_cnt_reg_11_ ( .d(stfd_byt_cnt11156_11_), .cp(ck54), .cdn(
        n12616), .q(bd_stfd_byt_cnt[11]) );
    dfctnq1 stfd_byt_cnt_reg_10_ ( .d(stfd_byt_cnt11156_10_), .cp(ck54), .cdn(
        n12518), .q(bd_stfd_byt_cnt[10]) );
    dfctnq1 stfd_byt_cnt_reg_9_ ( .d(stfd_byt_cnt11156_9_), .cp(ck54), .cdn(
        n12617), .q(bd_stfd_byt_cnt[9]) );
    dfctnq1 stfd_byt_cnt_reg_7_ ( .d(stfd_byt_cnt11156_7_), .cp(ck54), .cdn(
        n12516), .q(bd_stfd_byt_cnt[7]) );
    dfctnq1 stfd_byt_cnt_reg_5_ ( .d(stfd_byt_cnt11156_5_), .cp(ck54), .cdn(
        n12516), .q(bd_stfd_byt_cnt[5]) );
    dfctnq1 stfd_byt_cnt_reg_2_ ( .d(stfd_byt_cnt11156_2_), .cp(ck54), .cdn(
        n12615), .q(bd_stfd_byt_cnt[2]) );
    dfctnqn1 bd_cpu_req_lt_reg ( .d(bd_cpu_req_lt11152), .cp(ck54), .cdn(
        n12615), .qn(n13412) );
    dfctnqn1 bd_overflow_prev_reg ( .d(bd_overflow_prev11090), .cp(ck54), 
        .cdn(n12519), .qn(n13413) );
    dfctnqn1 b_cpu_req_reg ( .d(b_cpu_req11098), .cp(ck54), .cdn(n12618), .qn(
        n13414) );
    dfctnq1 b_sd_en_reg ( .d(b_sd_en11058), .cp(ck54), .cdn(n12618), .q(
        b_sd_en) );
    dfctnqn1 bd_cpu_ack_dly_reg ( .d(bd_cpu_ack_dly11086), .cp(ck54), .cdn(
        n12518), .qn(n13415) );
    dfctnq1 bd_cpu_irq0_reg ( .d(bd_cpu_irq011148), .cp(ck54), .cdn(n12517), 
        .q(b_cpu_irq[0]) );
    dfctnq1 bd_underflow_prev_reg ( .d(bd_underflow_prev11094), .cp(ck54), 
        .cdn(n12613), .q(bd_underflow_prev) );
    nd02e1 gt_278_U7 ( .a1(bp_bufval[3]), .b1(blk_with_stfd_cnt_3_), .zn(
        gt_278_n39) );
    nd02e1 gt_278_U12 ( .a1(bp_bufval[2]), .b1(blk_with_stfd_cnt_2_), .zn(
        gt_278_n37) );
    in01d1 gt_278_U19 ( .i(blk_with_stfd_cnt_6_), .zn(gt_278_n33) );
    nd02e1 gt_278_U21 ( .a1(bp_bufval[9]), .b1(blk_with_stfd_cnt_9_), .zn(
        gt_278_n47) );
    aon31d1 gt_278_U23 ( .a1(gt_278_n41), .a2(gt_278_n42), .a3(gt_278_n43), 
        .b(gt_278_n32), .z(gt_278_n40) );
    nd02e1 gt_278_U26 ( .a1(bp_bufval[8]), .b1(blk_with_stfd_cnt_8_), .zn(
        gt_278_n45) );
    in01d1 gt_278_U33 ( .i(blk_with_stfd_cnt_12_), .zn(gt_278_n35) );
    nd02e1 gt_278_U35 ( .a1(bp_bufval[13]), .b1(gt_278_n48), .zn(gt_278_n16)
         );
    aon31d1 gt_278_U36 ( .a1(gt_278_n49), .a2(gt_278_n50), .a3(gt_278_n51), 
        .b(gt_278_n34), .z(gt_278_n48) );
    nr02d1 gt_278_U45 ( .a1(bp_bufval[6]), .a2(gt_278_n33), .zn(gt_278_n32) );
    nr02d1 gt_278_U46 ( .a1(bp_bufval[12]), .a2(gt_278_n35), .zn(gt_278_n34)
         );
    nr03d2 gte_275_2_U8 ( .a1(n603_30_), .a2(bd_bm_count[0]), .a3(n603_26_), 
        .zn(gte_275_2_n66) );
    an02d1 add_465_U5 ( .a1(bd_stfd_byt_cnt[11]), .a2(add_465_carry_11_), .z(
        add_465_carry_12_) );
    an02d1 add_465_U7 ( .a1(bd_stfd_byt_cnt[10]), .a2(add_465_carry_10_), .z(
        add_465_carry_11_) );
    an02d1 add_465_U9 ( .a1(e_stfd_byt[0]), .a2(bd_stfd_byt_cnt[0]), .z(
        add_465_carry_1_) );
    ad01d1 add_465_U1_1 ( .a(bd_stfd_byt_cnt[1]), .b(e_stfd_byt[1]), .ci(
        add_465_carry_1_), .s(stfd_byt_cnt11157_1_), .co(add_465_carry_2_) );
    ad01d1 add_465_U1_6 ( .a(bd_stfd_byt_cnt[6]), .b(e_stfd_byt[6]), .ci(
        add_465_carry_6_), .s(stfd_byt_cnt11157_6_), .co(add_465_carry_7_) );
    ad01d1 add_465_U1_8 ( .a(bd_stfd_byt_cnt[8]), .b(e_stfd_byt[8]), .ci(
        add_465_carry_8_), .s(stfd_byt_cnt11157_8_), .co(add_465_carry_9_) );
    ad01d1 add_465_U1_7 ( .a(bd_stfd_byt_cnt[7]), .b(e_stfd_byt[7]), .ci(
        add_465_carry_7_), .s(stfd_byt_cnt11157_7_), .co(add_465_carry_8_) );
    ad01d1 add_465_U1_2 ( .a(bd_stfd_byt_cnt[2]), .b(e_stfd_byt[2]), .ci(
        add_465_carry_2_), .s(stfd_byt_cnt11157_2_), .co(add_465_carry_3_) );
    ad01d1 add_465_U1_9 ( .a(bd_stfd_byt_cnt[9]), .b(e_stfd_byt[9]), .ci(
        add_465_carry_9_), .s(stfd_byt_cnt11157_9_), .co(add_465_carry_10_) );
    ad01d1 add_465_U1_3 ( .a(bd_stfd_byt_cnt[3]), .b(e_stfd_byt[3]), .ci(
        add_465_carry_3_), .s(stfd_byt_cnt11157_3_), .co(add_465_carry_4_) );
    ad01d1 add_465_U1_4 ( .a(bd_stfd_byt_cnt[4]), .b(e_stfd_byt[4]), .ci(
        add_465_carry_4_), .s(stfd_byt_cnt11157_4_), .co(add_465_carry_5_) );
    ad01d1 add_465_U1_5 ( .a(bd_stfd_byt_cnt[5]), .b(e_stfd_byt[5]), .ci(
        add_465_carry_5_), .s(stfd_byt_cnt11157_5_), .co(add_465_carry_6_) );
    ah01d1 add_304_U1_1 ( .a(bd_r_adr_c_1_), .b(bd_r_adr_c_0_), .s(
        bd_r_adr_c_plus_1_1_), .co(add_304_carry_2_) );
    ah01d1 add_304_U1_2 ( .a(bd_r_adr_c_2_), .b(add_304_carry_2_), .s(
        bd_r_adr_c_plus_1_2_), .co(add_304_carry_3_) );
    ah01d1 add_304_U1_3 ( .a(bd_r_adr_c_3_), .b(add_304_carry_3_), .s(
        bd_r_adr_c_plus_1_3_), .co(add_304_carry_4_) );
    ah01d1 add_304_U1_4 ( .a(bd_r_adr_c_4_), .b(add_304_carry_4_), .s(
        bd_r_adr_c_plus_1_4_), .co(add_304_carry_5_) );
    xo02d1 add_510_U1_5 ( .a1(bd_au_count[5]), .a2(add_510_carry_5_), .z(
        bd_au_count11668_5_) );
    ah01d1 add_510_U1_1 ( .a(bd_au_count[1]), .b(bd_au_count[0]), .co(
        add_510_carry_2_) );
    ah01d1 add_510_U1_2 ( .a(bd_au_count[2]), .b(add_510_carry_2_), .s(
        bd_au_count11668_2_), .co(add_510_carry_3_) );
    ah01d1 add_510_U1_3 ( .a(bd_au_count[3]), .b(add_510_carry_3_), .s(
        bd_au_count11668_3_), .co(add_510_carry_4_) );
    ah01d1 add_510_U1_4 ( .a(bd_au_count[4]), .b(add_510_carry_4_), .s(
        bd_au_count11668_4_), .co(add_510_carry_5_) );
    aon21d1 sub_275_U4 ( .a1(sub_275_n95), .a2(sub_275_n105), .b(sub_275_n104), 
        .z(sub_275_n94) );
    or02d1 sub_275_U5 ( .a1(sub_275_n107), .a2(sub_275_n106), .z(sub_275_n90)
         );
    xo02d1 sub_275_U6 ( .a1(bd_bm_count[9]), .a2(sub_275_n108), .z(n598_23_)
         );
    nd02e1 sub_275_U9 ( .a1(sub_275_n94), .b1(bd_bm_count[6]), .zn(
        sub_275_n106) );
    nd02d1 sub_275_U10 ( .a1(bd_bm_count[3]), .a2(sub_275_n109), .zn(
        sub_275_n95) );
    or03d1 sub_275_U11 ( .a1(bd_bm_count[0]), .a2(bd_bm_count[2]), .a3(
        bd_bm_count[1]), .z(sub_275_n109) );
    xn02d1 sub_275_U15 ( .a1(bd_bm_count[10]), .a2(sub_275_n71), .zn(n598_22_)
         );
    nr02d1 sub_275_U16 ( .a1(bd_bm_count[9]), .a2(sub_275_n108), .zn(
        sub_275_n71) );
    xn02d1 sub_275_U17 ( .a1(bd_bm_count[2]), .a2(sub_275_n99), .zn(n598_30_)
         );
    xn02d1 sub_275_U18 ( .a1(sub_275_n95), .a2(bd_bm_count[4]), .zn(n598_28_)
         );
    nd02e1 sub_275_U22 ( .a1(bd_bm_count[8]), .b1(sub_275_n90), .zn(
        sub_275_n108) );
    in01d1 sub_275_U23 ( .i(bd_bm_count[7]), .zn(sub_275_n107) );
    in01d1 sub_275_U25 ( .i(bd_bm_count[5]), .zn(sub_275_n104) );
    in01d1 sub_275_U32 ( .i(bd_bm_count[12]), .zn(sub_275_n100) );
    in01d1 sub_275_U35 ( .i(bd_bm_count[4]), .zn(sub_275_n105) );
    nr02d1 sub_275_U57 ( .a1(bd_bm_count[1]), .a2(bd_bm_count[0]), .zn(
        sub_275_n99) );
    xn02d1 sub_513_U6 ( .a1(bd_au_count[5]), .a2(sub_513_n80), .zn(
        bd_au_count11677_5_) );
    nr02d1 sub_513_U7 ( .a1(bd_au_count[3]), .a2(sub_513_n78), .zn(sub_513_n73
        ) );
    nr02d1 sub_513_U9 ( .a1(bd_au_count[0]), .a2(bd_au_count[1]), .zn(
        sub_513_n74) );
    xn02d1 sub_513_U13 ( .a1(sub_513_n73), .a2(n12888), .zn(
        bd_au_count11677_4_) );
    nd02d1 sub_513_U14 ( .a1(sub_513_n73), .a2(n12888), .zn(sub_513_n80) );
    nd02e1 sub_513_U17 ( .a1(bd_au_count[2]), .b1(sub_513_n74), .zn(
        sub_513_n78) );
    an02d1 sub_526_U9 ( .a1(bd_mem_au_count[1]), .a2(bd_mem_au_count[0]), .z(
        sub_526_n83) );
    or02d1 sub_526_U10 ( .a1(bd_mem_au_count[0]), .a2(bd_mem_au_count[1]), .z(
        sub_526_n88) );
    xn02d1 sub_526_U11 ( .a1(n13678), .a2(sub_526_n118), .zn(
        bd_mem_au_count11744_6_) );
    in01d1 sub_526_U12 ( .i(sub_526_n84), .zn(sub_526_n119) );
    in01d1 sub_526_U16 ( .i(sub_526_n88), .zn(sub_526_n116) );
    xn02d1 sub_526_U17 ( .a1(sub_526_n119), .a2(sub_526_n120), .zn(
        bd_mem_au_count11744_5_) );
    nd02d1 sub_526_U18 ( .a1(sub_526_n119), .a2(sub_526_n120), .zn(
        sub_526_n118) );
    in01d1 sub_526_U19 ( .i(bd_mem_au_count[5]), .zn(sub_526_n120) );
    nd02e1 sub_526_U21 ( .a1(bd_mem_au_count[4]), .b1(sub_526_n82), .zn(
        sub_526_n84) );
    nd02e1 sub_526_U23 ( .a1(bd_mem_au_count[2]), .b1(sub_526_n116), .zn(
        sub_526_n89) );
    or03d1 lt_285_U7 ( .a1(bd_au_count[1]), .a2(bd_au_count[2]), .a3(
        bd_au_count[5]), .z(lt_285_n121) );
    nr02d1 sub_478_U9 ( .a1(bd_bm_count[2]), .a2(sub_478_n143), .zn(
        sub_478_n123) );
    or02d1 sub_478_U12 ( .a1(bd_bm_count[4]), .a2(sub_478_n133), .z(
        sub_478_n147) );
    nr02d1 sub_478_U15 ( .a1(bd_bm_count[11]), .a2(sub_478_n139), .zn(
        sub_478_n124) );
    nr02d1 sub_478_U18 ( .a1(bd_bm_count_32b[0]), .a2(bd_bm_count[0]), .zn(
        sub_478_n125) );
    or02d1 sub_478_U21 ( .a1(bd_bm_count[5]), .a2(sub_478_n147), .z(
        sub_478_n145) );
    nr02d1 sub_478_U23 ( .a1(bd_bm_count[9]), .a2(sub_478_n127), .zn(
        sub_478_n126) );
    or02d1 sub_478_U25 ( .a1(bd_bm_count[8]), .a2(sub_478_n129), .z(
        sub_478_n127) );
    or02d1 sub_478_U26 ( .a1(bd_bm_count[7]), .a2(sub_478_n131), .z(
        sub_478_n129) );
    or02d1 sub_478_U27 ( .a1(bd_bm_count[6]), .a2(sub_478_n145), .z(
        sub_478_n131) );
    xn02d1 sub_478_U28 ( .a1(bd_bm_count[13]), .a2(sub_478_n150), .zn(
        bd_bm_count_32b11631_14_) );
    nd02e1 sub_478_U30 ( .a1(bd_bm_count[1]), .b1(sub_478_n125), .zn(
        sub_478_n143) );
    nd02d1 sub_478_U31 ( .a1(sub_478_n124), .a2(sub_275_n100), .zn(
        sub_478_n150) );
    nd02e1 sub_478_U33 ( .a1(bd_bm_count[3]), .b1(sub_478_n123), .zn(
        sub_478_n133) );
    nd02e1 sub_478_U37 ( .a1(bd_bm_count[10]), .b1(sub_478_n126), .zn(
        sub_478_n139) );
    xn02d1 sub_478_U39 ( .a1(sub_478_n124), .a2(sub_275_n100), .zn(
        bd_bm_count_32b11631_13_) );
    in01d1 sub_478_U41 ( .i(bd_bm_count_32b[0]), .zn(bd_bm_count_32b11631_0_)
         );
    nr03d2 gte_275_U7 ( .a1(n598_27_), .a2(n598_29_), .a3(n598_25_), .zn(
        gte_275_n155) );
    or03d1 gte_275_U8 ( .a1(n598_28_), .a2(n598_26_), .a3(n598_23_), .z(
        gte_275_n152) );
    xo02d1 add_303_U1_5 ( .a1(bd_w_adr_c_5_), .a2(add_303_carry_5_), .z(
        bd_w_adr_c_plus_1_5_) );
    ah01d1 add_303_U1_1 ( .a(bd_w_adr_c_1_), .b(bd_w_adr_c_0_), .s(
        bd_w_adr_c_plus_1_1_), .co(add_303_carry_2_) );
    ah01d1 add_303_U1_2 ( .a(bd_w_adr_c_2_), .b(add_303_carry_2_), .s(
        bd_w_adr_c_plus_1_2_), .co(add_303_carry_3_) );
    ah01d1 add_303_U1_3 ( .a(bd_w_adr_c_3_), .b(add_303_carry_3_), .s(
        bd_w_adr_c_plus_1_3_), .co(add_303_carry_4_) );
    ah01d1 add_303_U1_4 ( .a(bd_w_adr_c_4_), .b(add_303_carry_4_), .s(
        bd_w_adr_c_plus_1_4_), .co(add_303_carry_5_) );
    an02d1 add_277_U5 ( .a1(bd_stfd_byt_cnt[0]), .a2(bd_bm_count[1]), .z(
        add_277_carry_2_) );
    xo02d1 add_277_U6 ( .a1(bd_stfd_byt_cnt[0]), .a2(bd_bm_count[1]), .z(
        blk_with_stfd_cnt_1_) );
    ad01d1 add_277_U1_6 ( .a(bd_bm_count[6]), .b(bd_stfd_byt_cnt[5]), .ci(
        add_277_carry_6_), .s(blk_with_stfd_cnt_6_), .co(add_277_carry_7_) );
    ad01d1 add_277_U1_8 ( .a(bd_bm_count[8]), .b(bd_stfd_byt_cnt[7]), .ci(
        add_277_carry_8_), .s(blk_with_stfd_cnt_8_), .co(add_277_carry_9_) );
    ad01d1 add_277_U1_11 ( .a(bd_bm_count[11]), .b(bd_stfd_byt_cnt[10]), .ci(
        add_277_carry_11_), .s(blk_with_stfd_cnt_11_), .co(add_277_carry_12_)
         );
    ad01d1 add_277_U1_7 ( .a(bd_bm_count[7]), .b(bd_stfd_byt_cnt[6]), .ci(
        add_277_carry_7_), .s(blk_with_stfd_cnt_7_), .co(add_277_carry_8_) );
    ad01d1 add_277_U1_2 ( .a(bd_bm_count[2]), .b(bd_stfd_byt_cnt[1]), .ci(
        add_277_carry_2_), .s(blk_with_stfd_cnt_2_), .co(add_277_carry_3_) );
    ad01d1 add_277_U1_9 ( .a(bd_bm_count[9]), .b(bd_stfd_byt_cnt[8]), .ci(
        add_277_carry_9_), .s(blk_with_stfd_cnt_9_), .co(add_277_carry_10_) );
    ad01d1 add_277_U1_10 ( .a(bd_bm_count[10]), .b(bd_stfd_byt_cnt[9]), .ci(
        add_277_carry_10_), .s(blk_with_stfd_cnt_10_), .co(add_277_carry_11_)
         );
    ad01d1 add_277_U1_3 ( .a(bd_bm_count[3]), .b(bd_stfd_byt_cnt[2]), .ci(
        add_277_carry_3_), .s(blk_with_stfd_cnt_3_), .co(add_277_carry_4_) );
    ad01d1 add_277_U1_4 ( .a(bd_bm_count[4]), .b(bd_stfd_byt_cnt[3]), .ci(
        add_277_carry_4_), .s(blk_with_stfd_cnt_4_), .co(add_277_carry_5_) );
    ad01d1 add_277_U1_5 ( .a(bd_bm_count[5]), .b(bd_stfd_byt_cnt[4]), .ci(
        add_277_carry_5_), .s(blk_with_stfd_cnt_5_), .co(add_277_carry_6_) );
    ad01d1 add_277_U1_12 ( .a(bd_bm_count[12]), .b(bd_stfd_byt_cnt[11]), .ci(
        add_277_carry_12_), .s(blk_with_stfd_cnt_12_), .co(add_277_carry_13_)
         );
    xo02d1 add_301_U1_10 ( .a1(bd_w_adr_r_10_), .a2(add_301_carry_10_), .z(
        bd_w_adr_r_plus_1_10_) );
    ah01d1 add_301_U1_1 ( .a(bd_w_adr_r_1_), .b(bd_w_adr_r_0_), .s(
        bd_w_adr_r_plus_1_1_), .co(add_301_carry_2_) );
    ah01d1 add_301_U1_8 ( .a(bd_w_adr_r_8_), .b(add_301_carry_8_), .s(
        bd_w_adr_r_plus_1_8_), .co(add_301_carry_9_) );
    ah01d1 add_301_U1_6 ( .a(bd_w_adr_r_6_), .b(add_301_carry_6_), .s(
        bd_w_adr_r_plus_1_6_), .co(add_301_carry_7_) );
    ah01d1 add_301_U1_2 ( .a(bd_w_adr_r_2_), .b(add_301_carry_2_), .s(
        bd_w_adr_r_plus_1_2_), .co(add_301_carry_3_) );
    ah01d1 add_301_U1_7 ( .a(bd_w_adr_r_7_), .b(add_301_carry_7_), .s(
        bd_w_adr_r_plus_1_7_), .co(add_301_carry_8_) );
    ah01d1 add_301_U1_9 ( .a(bd_w_adr_r_9_), .b(add_301_carry_9_), .s(
        bd_w_adr_r_plus_1_9_), .co(add_301_carry_10_) );
    ah01d1 add_301_U1_3 ( .a(bd_w_adr_r_3_), .b(add_301_carry_3_), .s(
        bd_w_adr_r_plus_1_3_), .co(add_301_carry_4_) );
    ah01d1 add_301_U1_4 ( .a(bd_w_adr_r_4_), .b(add_301_carry_4_), .s(
        bd_w_adr_r_plus_1_4_), .co(add_301_carry_5_) );
    ah01d1 add_301_U1_5 ( .a(bd_w_adr_r_5_), .b(add_301_carry_5_), .s(
        bd_w_adr_r_plus_1_5_), .co(add_301_carry_6_) );
    ah01d1 add_491_U1_1 ( .a(bd_cpu_ack_cnt[1]), .b(bd_cpu_ack_cnt[0]), .s(
        bd_cpu_ack_cnt11656_1_), .co(add_491_carry_2_) );
    ah01d1 add_491_U1_2 ( .a(bd_cpu_ack_cnt[2]), .b(add_491_carry_2_), .s(
        bd_cpu_ack_cnt11656_2_), .co(add_491_carry_3_) );
    ah01d1 add_491_U1_3 ( .a(bd_cpu_ack_cnt[3]), .b(add_491_carry_3_), .s(
        bd_cpu_ack_cnt11656_3_), .co(add_491_carry_4_) );
    ah01d1 add_491_U1_4 ( .a(bd_cpu_ack_cnt[4]), .b(add_491_carry_4_), .s(
        bd_cpu_ack_cnt11656_4_), .co(add_491_carry_5_) );
    xo02d1 add_475_U1_14 ( .a1(bd_bm_count[13]), .a2(add_475_carry_14_), .z(
        bd_bm_count_32b11622_14_) );
    ah01d1 add_475_U1_1 ( .a(bd_bm_count[0]), .b(bd_bm_count_32b[0]), .s(
        bd_bm_count_32b11622_1_), .co(add_475_carry_2_) );
    ah01d1 add_475_U1_8 ( .a(bd_bm_count[7]), .b(add_475_carry_8_), .s(
        bd_bm_count_32b11622_8_), .co(add_475_carry_9_) );
    ah01d1 add_475_U1_11 ( .a(bd_bm_count[10]), .b(add_475_carry_11_), .s(
        bd_bm_count_32b11622_11_), .co(add_475_carry_12_) );
    ah01d1 add_475_U1_6 ( .a(bd_bm_count[5]), .b(add_475_carry_6_), .s(
        bd_bm_count_32b11622_6_), .co(add_475_carry_7_) );
    ah01d1 add_475_U1_2 ( .a(bd_bm_count[1]), .b(add_475_carry_2_), .s(
        bd_bm_count_32b11622_2_), .co(add_475_carry_3_) );
    ah01d1 add_475_U1_7 ( .a(bd_bm_count[6]), .b(add_475_carry_7_), .s(
        bd_bm_count_32b11622_7_), .co(add_475_carry_8_) );
    ah01d1 add_475_U1_9 ( .a(bd_bm_count[8]), .b(add_475_carry_9_), .s(
        bd_bm_count_32b11622_9_), .co(add_475_carry_10_) );
    ah01d1 add_475_U1_10 ( .a(bd_bm_count[9]), .b(add_475_carry_10_), .s(
        bd_bm_count_32b11622_10_), .co(add_475_carry_11_) );
    ah01d1 add_475_U1_3 ( .a(bd_bm_count[2]), .b(add_475_carry_3_), .s(
        bd_bm_count_32b11622_3_), .co(add_475_carry_4_) );
    ah01d1 add_475_U1_4 ( .a(bd_bm_count[3]), .b(add_475_carry_4_), .s(
        bd_bm_count_32b11622_4_), .co(add_475_carry_5_) );
    ah01d1 add_475_U1_5 ( .a(bd_bm_count[4]), .b(add_475_carry_5_), .s(
        bd_bm_count_32b11622_5_), .co(add_475_carry_6_) );
    ah01d1 add_475_U1_12 ( .a(bd_bm_count[11]), .b(add_475_carry_12_), .s(
        bd_bm_count_32b11622_12_), .co(add_475_carry_13_) );
    ah01d1 add_475_U1_13 ( .a(bd_bm_count[12]), .b(add_475_carry_13_), .s(
        bd_bm_count_32b11622_13_), .co(add_475_carry_14_) );
    or02d1 sub_275_2_U4 ( .a1(sub_275_2_n200), .a2(bd_bm_count[10]), .z(
        sub_275_2_n191) );
    or02d1 sub_275_2_U5 ( .a1(sub_275_n107), .a2(sub_275_2_n197), .z(
        sub_275_2_n180) );
    xo02d1 sub_275_2_U6 ( .a1(bd_bm_count[2]), .a2(sub_275_2_n188), .z(
        n603_30_) );
    xn02d1 sub_275_2_U10 ( .a1(bd_bm_count[4]), .a2(sub_275_2_n185), .zn(
        n603_28_) );
    oai21d1 sub_275_2_U11 ( .a1(sub_275_2_n188), .a2(bd_bm_count[2]), .b(
        bd_bm_count[3]), .zn(sub_275_2_n185) );
    nd02e1 sub_275_2_U27 ( .a1(bd_bm_count[8]), .b1(sub_275_2_n180), .zn(
        sub_275_2_n199) );
    xo02d1 sub_275_2_U30 ( .a1(bd_bm_count[0]), .a2(bd_bm_count[1]), .z(
        n603_31_) );
    aoi21d2 sub_275_2_U36 ( .a1(sub_275_2_n185), .a2(sub_275_n105), .b(
        sub_275_n104), .zn(sub_275_2_n159) );
    nr02d1 sub_275_2_U60 ( .a1(bd_bm_count[4]), .a2(bd_bm_count[5]), .zn(
        sub_275_2_n203) );
    nr03d2 gte_274_2_U8 ( .a1(bd_bm_count[11]), .a2(bd_bm_count[5]), .a3(
        bd_bm_count[8]), .zn(gte_274_2_n167) );
    nr02d1 gte_274_2_U12 ( .a1(bd_bm_count[2]), .a2(bd_bm_count[6]), .zn(
        gte_274_2_n165) );
    nr02d1 gte_274_2_U13 ( .a1(bd_bm_count[13]), .a2(bd_bm_count[1]), .zn(
        gte_274_2_n166) );
    nr03d2 gte_274_U7 ( .a1(bd_bm_count[12]), .a2(bd_bm_count[10]), .a3(
        bd_bm_count[7]), .zn(gte_274_n175) );
    nr02d1 gte_274_U13 ( .a1(bd_bm_count[0]), .a2(bd_bm_count[11]), .zn(
        gte_274_n173) );
    nr02d1 gte_274_U14 ( .a1(bd_bm_count[5]), .a2(bd_bm_count[3]), .zn(
        gte_274_n174) );
    xo02d1 add_302_U1_10 ( .a1(bd_r_adr_r_10_), .a2(add_302_carry_10_), .z(
        bd_r_adr_r_plus_1_10_) );
    ah01d1 add_302_U1_1 ( .a(bd_r_adr_r_1_), .b(bd_r_adr_r_0_), .s(
        bd_r_adr_r_plus_1_1_), .co(add_302_carry_2_) );
    ah01d1 add_302_U1_8 ( .a(bd_r_adr_r_8_), .b(add_302_carry_8_), .s(
        bd_r_adr_r_plus_1_8_), .co(add_302_carry_9_) );
    ah01d1 add_302_U1_6 ( .a(bd_r_adr_r_6_), .b(add_302_carry_6_), .s(
        bd_r_adr_r_plus_1_6_), .co(add_302_carry_7_) );
    ah01d1 add_302_U1_2 ( .a(bd_r_adr_r_2_), .b(add_302_carry_2_), .s(
        bd_r_adr_r_plus_1_2_), .co(add_302_carry_3_) );
    ah01d1 add_302_U1_7 ( .a(bd_r_adr_r_7_), .b(add_302_carry_7_), .s(
        bd_r_adr_r_plus_1_7_), .co(add_302_carry_8_) );
    ah01d1 add_302_U1_9 ( .a(bd_r_adr_r_9_), .b(add_302_carry_9_), .s(
        bd_r_adr_r_plus_1_9_), .co(add_302_carry_10_) );
    ah01d1 add_302_U1_3 ( .a(bd_r_adr_r_3_), .b(add_302_carry_3_), .s(
        bd_r_adr_r_plus_1_3_), .co(add_302_carry_4_) );
    ah01d1 add_302_U1_4 ( .a(bd_r_adr_r_4_), .b(add_302_carry_4_), .s(
        bd_r_adr_r_plus_1_4_), .co(add_302_carry_5_) );
    ah01d1 add_302_U1_5 ( .a(bd_r_adr_r_5_), .b(add_302_carry_5_), .s(
        bd_r_adr_r_plus_1_5_), .co(add_302_carry_6_) );
    an02d1 U5128 ( .a1(bd_w_adr_r_9_), .a2(bd_w_adr_r_8_), .z(n13445) );
    an02d1 U5129 ( .a1(bd_r_adr_r_9_), .a2(bd_r_adr_r_5_), .z(n13446) );
    oan2111d1 U5130 ( .a1(bp_bufval[13]), .a2(n13528), .b(gt_278_n16), .c(
        gt_278_n15), .d(n13447), .z(n13464) );
    in01d1 U5131 ( .i(bd_active_once), .zn(n13447) );
    xn02d1 U5140 ( .a1(bd_bm_count_32b[8]), .a2(sub_275_2_n197), .zn(n13486)
         );
    nd04d2 U5142 ( .a1(bd_w_adr_c_5_), .a3(bd_w_adr_c_1_), .a4(n13042), .a2(
        bd_w_adr_c_0_), .zn(n13040) );
    nr04d2 U5143 ( .a1(bd_bm_count[9]), .a2(bd_bm_count[4]), .a3(bd_bm_count
        [3]), .a4(n13495), .zn(gte_274_2_n163) );
    an04d1 U5144 ( .a1(gte_274_n174), .a2(gte_274_n173), .a3(gte_274_n175), 
        .a4(gte_274_n169), .z(n13502) );
    an04d1 U5145 ( .a1(gte_274_2_n163), .a2(gte_274_2_n166), .a3(
        gte_274_2_n165), .a4(gte_274_2_n167), .z(n13503) );
    oai31d1 U5147 ( .a1(bd_bm_count[2]), .a2(bd_bm_count[3]), .a3(
        sub_275_2_n188), .b(sub_275_2_n185), .zn(n603_29_) );
    xn02d1 U5148 ( .a1(bd_bm_count[6]), .a2(sub_275_2_n159), .zn(n603_26_) );
    xn02d1 U5149 ( .a1(bd_bm_count[9]), .a2(sub_478_n127), .zn(
        bd_bm_count_32b11631_10_) );
    xn02d1 U5150 ( .a1(bd_bm_count[6]), .a2(sub_478_n145), .zn(
        bd_bm_count_32b11631_7_) );
    xn02d1 U5151 ( .a1(bd_bm_count[8]), .a2(sub_478_n129), .zn(
        bd_bm_count_32b11631_9_) );
    xn02d1 U5152 ( .a1(bd_bm_count[5]), .a2(sub_478_n147), .zn(
        bd_bm_count_32b11631_6_) );
    xn02d1 U5153 ( .a1(bd_bm_count[4]), .a2(sub_478_n133), .zn(
        bd_bm_count_32b11631_5_) );
    xn02d1 U5154 ( .a1(bd_bm_count[2]), .a2(sub_478_n143), .zn(
        bd_bm_count_32b11631_3_) );
    xo02d1 U5155 ( .a1(bd_bm_count[3]), .a2(sub_478_n123), .z(
        bd_bm_count_32b11631_4_) );
    xn02d1 U5156 ( .a1(bd_bm_count[11]), .a2(sub_478_n139), .zn(
        bd_bm_count_32b11631_12_) );
    xn02d1 U5158 ( .a1(bd_mem_au_count[2]), .a2(sub_526_n88), .zn(
        bd_mem_au_count11744_2_) );
    xo02d1 U5160 ( .a1(bd_au_count[2]), .a2(sub_513_n74), .z(
        bd_au_count11677_2_) );
    xn02d1 U5161 ( .a1(bd_au_count[3]), .a2(sub_513_n78), .zn(
        bd_au_count11677_3_) );
    nd02e1 U5162 ( .a1(bd_bm_count_32b[11]), .b1(sub_275_n71), .zn(
        sub_275_n102) );
    in01d1 U5164 ( .i(n13509), .zn(n13449) );
    or03d1 U5165 ( .a1(bd_bm_count_32b[11]), .a2(bd_bm_count[11]), .a3(n13450), 
        .z(sub_275_n110) );
    in01d1 U5166 ( .i(sub_275_n71), .zn(n13450) );
    xo02d1 U5167 ( .a1(bd_bm_count_32b[8]), .a2(sub_275_n106), .z(n598_25_) );
    xn02d1 U5168 ( .a1(bd_bm_count[3]), .a2(sub_275_n109), .zn(n598_29_) );
    aon31d1 U5169 ( .a1(sub_275_n95), .a2(sub_275_n105), .a3(sub_275_n104), 
        .b(n13451), .z(n598_27_) );
    in01d1 U5170 ( .i(sub_275_n94), .zn(n13451) );
    xo02d1 U5171 ( .a1(sub_275_n94), .a2(bd_bm_count[6]), .z(n598_26_) );
    aoi211d1 U5172 ( .a1(sub_275_2_n185), .a2(sub_275_2_n203), .b(n603_31_), 
        .c(sub_275_2_n159), .zn(gte_275_2_n65) );
    oai222d1 U5173 ( .a1(n13452), .a2(bp_bufval[10]), .b1(n13453), .b2(
        bp_bufval[11]), .c1(gt_278_n44), .c2(gt_278_n20), .zn(gt_278_n50) );
    in01d1 U5174 ( .i(blk_with_stfd_cnt_10_), .zn(n13452) );
    in01d1 U5175 ( .i(blk_with_stfd_cnt_11_), .zn(n13453) );
    oai222d1 U5176 ( .a1(n13454), .a2(blk_with_stfd_cnt_7_), .b1(n13455), .b2(
        blk_with_stfd_cnt_8_), .c1(gt_278_n30), .c2(gt_278_n40), .zn(
        gt_278_n46) );
    in01d1 U5177 ( .i(bp_bufval[7]), .zn(n13454) );
    in01d1 U5178 ( .i(bp_bufval[8]), .zn(n13455) );
    oai222d1 U5179 ( .a1(n13456), .a2(bp_bufval[4]), .b1(n13457), .b2(
        bp_bufval[5]), .c1(gt_278_n36), .c2(gt_278_n28), .zn(gt_278_n42) );
    in01d1 U5180 ( .i(blk_with_stfd_cnt_4_), .zn(n13456) );
    in01d1 U5181 ( .i(blk_with_stfd_cnt_5_), .zn(n13457) );
    oai222d1 U5182 ( .a1(n13458), .a2(blk_with_stfd_cnt_1_), .b1(n13459), .b2(
        blk_with_stfd_cnt_2_), .c1(gt_278_n22), .c2(gt_278_n24), .zn(
        gt_278_n38) );
    in01d1 U5183 ( .i(bp_bufval[1]), .zn(n13458) );
    in01d1 U5184 ( .i(bp_bufval[2]), .zn(n13459) );
    nr02e1 U5185 ( .a1(blk_with_stfd_cnt_7_), .b1(bp_bufval[7]), .zn(
        gt_278_n30) );
    nr02e1 U5187 ( .a1(blk_with_stfd_cnt_1_), .b1(bp_bufval[1]), .zn(
        gt_278_n22) );
    aon32d1 U5189 ( .a1(gt_278_n47), .a2(gt_278_n45), .a3(gt_278_n46), .b1(
        bp_bufval[9]), .b2(n13460), .z(gt_278_n44) );
    in01d1 U5190 ( .i(blk_with_stfd_cnt_9_), .zn(n13460) );
    aon32d1 U5191 ( .a1(gt_278_n37), .a2(gt_278_n38), .a3(gt_278_n39), .b1(
        bp_bufval[3]), .b2(n13461), .z(gt_278_n36) );
    in01d1 U5192 ( .i(blk_with_stfd_cnt_3_), .zn(n13461) );
    nd03d1 U5193 ( .a1(n12479), .a2(n13074), .a3(bd_au_state[1]), .zn(n13250)
         );
    an04d1 U5195 ( .a1(bd_r_adr_r_0_), .a2(bd_r_adr_r_1_), .a3(bd_r_adr_r_2_), 
        .a4(n13446), .z(n13157) );
    an04d1 U5196 ( .a1(bd_w_adr_r_1_), .a2(bd_w_adr_r_0_), .a3(bd_w_adr_r_2_), 
        .a4(n13445), .z(n13154) );
    oan211d1 U5197 ( .a1(n12536), .a2(n13206), .b(n13268), .c(n12696), .z(
        n13341) );
    nr02e1 U5198 ( .a1(s_sd_dat[16]), .b1(bt_rst), .zn(bd_sd_dat11062_16_) );
    nr02e1 U5199 ( .a1(stfd_byt_cnt11157_8_), .b1(bt_rst), .zn(
        stfd_byt_cnt11156_8_) );
    nr02e1 U5200 ( .a1(stfd_byt_cnt11157_3_), .b1(bt_rst), .zn(
        stfd_byt_cnt11156_3_) );
    nr02e1 U5201 ( .a1(stfd_byt_cnt11157_1_), .b1(bt_rst), .zn(
        stfd_byt_cnt11156_1_) );
    nr02e1 U5203 ( .a1(bd_dt_ava), .b1(n13198), .zn(n12536) );
    nr04d2 U5204 ( .a1(n12920), .a2(lt_285_n121), .a3(bd_au_count[3]), .a4(
        bd_au_count[4]), .zn(bd_underflow) );
    in01d1 U5206 ( .i(bd_underflow_prev), .zn(n13462) );
    oai22h1 U5208 ( .a1(n13637), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[26]), 
        .zn(b_sd_dat11070_26_) );
    oai22h1 U5209 ( .a1(n13639), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[27]), 
        .zn(b_sd_dat11070_27_) );
    oai22h1 U5210 ( .a1(n13642), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[28]), 
        .zn(b_sd_dat11070_28_) );
    oai22h1 U5211 ( .a1(n13644), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[29]), 
        .zn(b_sd_dat11070_29_) );
    oai22h1 U5212 ( .a1(n13645), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[30]), 
        .zn(b_sd_dat11070_30_) );
    oai22h1 U5213 ( .a1(n13647), .a2(n12730), .b1(n12535), .b2(b_buf_rdt[31]), 
        .zn(b_sd_dat11070_31_) );
    oai221d1 U5218 ( .a1(n13464), .a2(bt_rst), .b1(n13465), .b2(n12730), .c(
        n12904), .zn(n13355) );
    in01d1 U5219 ( .i(p_dec_sta), .zn(n13465) );
    oai21d1 U5220 ( .a1(sub_526_n116), .a2(sub_526_n83), .b(n12509), .zn(
        n12899) );
    or04d1 U5221 ( .a1(n13204), .a2(n12536), .a3(bt_rst), .a4(n13205), .z(
        n12947) );
    aoi22h1 U5222 ( .a1(n13257), .a2(bd_w_adr_r_3_), .b1(n13049), .b2(n12993), 
        .zn(n12811) );
    aoi22h1 U5223 ( .a1(n13257), .a2(bd_w_adr_r_4_), .b1(n13049), .b2(n12992), 
        .zn(n12809) );
    aoi22h1 U5224 ( .a1(n13257), .a2(bd_w_adr_r_5_), .b1(n13049), .b2(n12991), 
        .zn(n12807) );
    aoi22h1 U5226 ( .a1(n13257), .a2(bd_w_adr_r_7_), .b1(n13049), .b2(n12989), 
        .zn(n12803) );
    aoi22h1 U5227 ( .a1(n13257), .a2(bd_w_adr_r_8_), .b1(n13049), .b2(n12988), 
        .zn(n12801) );
    aoi22h1 U5228 ( .a1(n13257), .a2(bd_w_adr_r_9_), .b1(n13049), .b2(n12987), 
        .zn(n12799) );
    aoi22h1 U5229 ( .a1(n13257), .a2(n13692), .b1(n13049), .b2(n12986), .zn(
        n12797) );
    aon22d1 U5230 ( .a1(n12881), .a2(n12506), .b1(n13697), .b2(n13573), .z(
        n13347) );
    aoi32d1 U5242 ( .a1(n13124), .a2(n12491), .a3(n12983), .b1(n12981), .b2(
        n12540), .zn(n12658) );
    nr02e1 U5243 ( .a1(n12939), .b1(bd_we_dec_adv), .zn(n13151) );
    nd04d2 U5244 ( .a1(bd_r_adr_c_5_), .a3(bd_r_adr_c_1_), .a4(n13053), .a2(
        bd_r_adr_c_0_), .zn(n13051) );
    nd04d2 U5245 ( .a1(n13286), .a3(bt_pulse4), .a4(bd_active_once), .a2(
        p_bs_req), .zn(n13198) );
    an04d1 U5246 ( .a1(n13201), .a2(n13200), .a3(n13202), .a4(n12925), .z(
        n13204) );
    oan31d1 U5247 ( .a1(n12491), .a2(n12965), .a3(n12971), .b(n13112), .z(
        n13115) );
    oai211d2 U5248 ( .a1(n13034), .a2(n12565), .b(n12491), .c(n13122), .zn(
        n13284) );
    or04d1 U5249 ( .a1(n13086), .a2(n12570), .a3(n13015), .a4(n13472), .z(
        n13085) );
    in01d1 U5250 ( .i(n12515), .zn(n13472) );
    oai21d1 U5251 ( .a1(n12971), .a2(n12541), .b(n13236), .zn(n13235) );
    aoi22h1 U5252 ( .a1(n13277), .a2(bd_seq_hdr_exist), .b1(n13072), .b2(
        n12521), .zn(n13237) );
    or03d1 U5253 ( .a1(n13004), .a2(n13000), .a3(n13002), .z(n13076) );
    aon211d1 U5254 ( .a1(n13116), .a2(n13217), .b(bd_seq_hdr_exist), .c(n13542
        ), .z(n13090) );
    oai32d1 U5255 ( .a1(n13473), .a2(bt_rst), .a3(n13668), .b1(n13474), .b2(
        n12915), .zn(n13362) );
    in01d1 U5256 ( .i(bd_bs_req_lt), .zn(n13473) );
    in01d1 U5257 ( .i(p_bs_req), .zn(n13474) );
    nd02e1 U5258 ( .a1(n13095), .b1(p_mem_pic), .zn(n12885) );
    nr03d2 U5270 ( .a1(n12945), .a2(n12762), .a3(bt_rst), .zn(n12505) );
    nd04d2 U5271 ( .a1(n13483), .a3(n13156), .a4(n13157), .a2(bd_r_adr_r_7_), 
        .zn(n12499) );
    in01d1 U5272 ( .i(n13195), .zn(n13483) );
    nd04d2 U5273 ( .a1(n13550), .a3(n13153), .a4(n13154), .a2(bd_w_adr_r_7_), 
        .zn(n12498) );
    oai21d1 U5275 ( .a1(n12492), .a2(n12580), .b(n13281), .zn(n13117) );
    oan31d1 U5276 ( .a1(n12948), .a2(bd_seq_hdr_exist), .a3(n12965), .b(n13112
        ), .z(n13224) );
    aon21d1 U5277 ( .a1(n13120), .a2(bd_seq_hdr_exist), .b(n13113), .z(n13171)
         );
    or04d1 U5278 ( .a1(n13008), .a2(n12998), .a3(n13006), .a4(n13010), .z(
        n12489) );
    oan32d1 U5279 ( .a1(n13494), .a2(n12481), .a3(n13066), .b1(n13085), .b2(
        bd_seq_hdr_exist), .z(n13223) );
    an04d1 U5280 ( .a1(n13488), .a2(n13487), .a3(n13486), .a4(n13485), .z(
        n13493) );
    xn02d1 U5281 ( .a1(bd_bm_count[10]), .a2(sub_275_2_n200), .zn(n13485) );
    nr02d1 U5283 ( .a1(n603_28_), .a2(n603_29_), .zn(n13488) );
    oan21d1 U5284 ( .a1(n13549), .a2(bd_bm_count[12]), .b(bd_bm_count[13]), 
        .z(n13511) );
    nd02d1 U5286 ( .a1(gt_278_n33), .a2(bp_bufval[6]), .zn(gt_278_n43) );
    nd02d1 U5287 ( .a1(gt_278_n35), .a2(bp_bufval[12]), .zn(gt_278_n51) );
    or02d1 U5288 ( .a1(bd_bm_count[0]), .a2(bd_bm_count[1]), .z(sub_275_2_n188
        ) );
    nd02d1 U5289 ( .a1(bd_bm_count[6]), .a2(sub_275_2_n159), .zn(
        sub_275_2_n197) );
    an03d1 U5290 ( .a1(n13492), .a2(n13491), .a3(n13490), .z(gte_275_n156) );
    xn02d1 U5291 ( .a1(sub_275_n102), .a2(bd_bm_count[11]), .zn(n13490) );
    xn02d1 U5292 ( .a1(bd_bm_count[0]), .a2(bd_bm_count[1]), .zn(n13491) );
    xo02d1 U5293 ( .a1(sub_275_n90), .a2(bd_bm_count[8]), .z(n13492) );
    xn02d1 U5294 ( .a1(bd_bm_count[12]), .a2(sub_275_n110), .zn(n13510) );
    oan21d1 U5295 ( .a1(sub_275_n110), .a2(bd_bm_count[12]), .b(bd_bm_count
        [13]), .z(n13509) );
    nd02d1 U5296 ( .a1(n12577), .a2(n12553), .zn(n13494) );
    in01d1 U5297 ( .i(n13494), .zn(n12479) );
    or03d1 U5298 ( .a1(bd_bm_count[12]), .a2(bd_bm_count[10]), .a3(bd_bm_count
        [7]), .z(n13495) );
    nr04d1 U5299 ( .a1(n13497), .a2(n13496), .a3(n13511), .a4(n603_19_), .zn(
        n13505) );
    nd04d2 U5300 ( .a1(gte_275_2_n66), .a3(n13507), .a4(n13506), .a2(
        gte_275_2_n65), .zn(n13496) );
    nd02d1 U5301 ( .a1(n13508), .a2(n13493), .zn(n13497) );
    mi21d1 U5302 ( .i0(bd_au_count[0]), .i1(bd_au_count[0]), .s(n13272), .zn(
        n12881) );
    nr02d1 U5303 ( .a1(sub_275_n100), .a2(n12946), .zn(n12843) );
    an02d1 U5304 ( .a1(n13293), .a2(stfd_byt_cnt11157_4_), .z(
        stfd_byt_cnt11156_4_) );
    an02d1 U5306 ( .a1(n13293), .a2(stfd_byt_cnt11157_6_), .z(
        stfd_byt_cnt11156_6_) );
    nd02d1 U5307 ( .a1(n13075), .a2(n12575), .zn(n12559) );
    ni01d2 U5310 ( .i(bd_bm_count_32b[14]), .z(bd_bm_count[13]) );
    mi21d1 U5311 ( .i0(n13505), .i1(n13504), .s(bl_v_dec_mod), .zn(n12641) );
    xn02d1 U5314 ( .a1(e_stfd_byt[0]), .a2(n13703), .zn(n13499) );
    xn02d1 U5315 ( .a1(n13656), .a2(add_304_carry_5_), .zn(n13500) );
    xn02d1 U5321 ( .a1(sub_275_2_n191), .a2(bd_bm_count[11]), .zn(n13506) );
    xo02d1 U5322 ( .a1(sub_275_2_n180), .a2(bd_bm_count[8]), .z(n13507) );
    oai21d1 U5324 ( .a1(n13048), .a2(n13040), .b(n13256), .zn(n13512) );
    aon222d1 U5325 ( .a1(bd_bm_count_32b11631_2_), .a2(n12505), .b1(n12504), 
        .b2(bd_bm_count_32b11622_2_), .c1(bd_bm_count[1]), .c2(n13059), .z(
        n13333) );
    aon21d1 U5326 ( .a1(n12586), .a2(n13542), .b(n12966), .z(n13232) );
    oan211d1 U5327 ( .a1(bd_sd_dat_25_), .a2(n13521), .b(bd_sd_dat_29_), .c(
        bd_sd_dat_28_), .z(n12952) );
    xn02d1 U5328 ( .a1(bd_mem_au_count[3]), .a2(sub_526_n89), .zn(
        bd_mem_au_count11744_3_) );
    aon221d1 U5329 ( .a1(n13277), .a2(bd_gop_hdr_exist), .b1(n12521), .b2(
        n13553), .c(n13118), .z(n12980) );
    oai33d1 U5330 ( .a1(n13513), .a2(n13514), .a3(n12513), .b1(n13109), .b2(
        bt_pulse5), .b3(bt_pulse6), .zn(n13538) );
    in01d1 U5331 ( .i(br_buf_valid), .zn(n13513) );
    in01d1 U5332 ( .i(bd_dt_ava), .zn(n13514) );
    aoi211d1 U5333 ( .a1(n13385), .a2(n12950), .b(n13382), .c(n13381), .zn(
        n12949) );
    an04d1 U5334 ( .a1(n12555), .a2(n12515), .a3(n13219), .a4(n13068), .z(
        n12583) );
    an04d1 U5335 ( .a1(n12586), .a2(n13542), .a3(n12568), .a4(n12967), .z(
        n12575) );
    an04d1 U5336 ( .a1(n13065), .a2(n12545), .a3(n13064), .a4(n13515), .z(
        n12586) );
    in01d1 U5337 ( .i(n13025), .zn(n13515) );
    aon222d1 U5339 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_10_), .b1(n12534), 
        .b2(n13570), .c1(n13690), .c2(n12944), .z(n13310) );
    aon222d1 U5340 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_9_), .b1(n12534), .b2(
        n13569), .c1(n13689), .c2(n12944), .z(n13311) );
    aon222d1 U5341 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_8_), .b1(n12534), .b2(
        n13261), .c1(n13688), .c2(n12944), .z(n13312) );
    aon222d1 U5342 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_7_), .b1(n12534), .b2(
        n13262), .c1(n13687), .c2(n12944), .z(n13313) );
    aon222d1 U5343 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_6_), .b1(n12534), .b2(
        n13263), .c1(n13686), .c2(n12944), .z(n13314) );
    aon222d1 U5344 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_5_), .b1(n12534), .b2(
        n13264), .c1(n13685), .c2(n12944), .z(n13315) );
    aon222d1 U5345 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_4_), .b1(n12534), .b2(
        n13265), .c1(n13684), .c2(n12944), .z(n13316) );
    aon222d1 U5346 ( .a1(n12533), .a2(bd_r_adr_r_plus_1_3_), .b1(n12534), .b2(
        n13266), .c1(n13683), .c2(n12944), .z(n13317) );
    xo02d1 U5348 ( .a1(bd_bm_count_32b[11]), .a2(sub_478_n126), .z(
        bd_bm_count_32b11631_11_) );
    xn02d1 U5349 ( .a1(bd_bm_count_32b[8]), .a2(sub_478_n131), .zn(
        bd_bm_count_32b11631_8_) );
    xn02d1 U5350 ( .a1(bd_bm_count_32b[0]), .a2(bd_bm_count_32b[1]), .zn(
        bd_bm_count_32b11631_1_) );
    xo02d1 U5351 ( .a1(bd_bm_count[1]), .a2(sub_478_n125), .z(
        bd_bm_count_32b11631_2_) );
    nr02e1 U5352 ( .a1(bd_bm_count_32b[1]), .b1(bp_bufval[0]), .zn(gt_278_n24)
         );
    aon221d1 U5354 ( .a1(bd_r_adr_c_plus_1_3_), .a2(n13566), .b1(n13653), .b2(
        n13274), .c(n13517), .z(n13375) );
    aon221d1 U5355 ( .a1(bd_r_adr_c_plus_1_1_), .a2(n13566), .b1(n13654), .b2(
        n13274), .c(n13517), .z(n13374) );
    aon221d1 U5356 ( .a1(n12511), .a2(bd_w_adr_c_plus_1_2_), .b1(n13663), .b2(
        n13520), .c(n13512), .z(n13367) );
    aon221d1 U5357 ( .a1(n12511), .a2(bd_w_adr_c_plus_1_3_), .b1(n13666), .b2(
        n13520), .c(n13512), .z(n13364) );
    aon221d1 U5358 ( .a1(n12511), .a2(bd_w_adr_c_plus_1_1_), .b1(n13667), .b2(
        n13520), .c(n13512), .z(n13363) );
    aon221d1 U5359 ( .a1(n12511), .a2(bd_w_adr_c_plus_1_5_), .b1(n13669), .b2(
        n13520), .c(n13512), .z(n13360) );
    aon221d1 U5360 ( .a1(bd_r_adr_c_plus_1_2_), .a2(n13566), .b1(n13673), .b2(
        n13274), .c(n13517), .z(n13357) );
    in01d1 U5362 ( .i(n12530), .zn(n13517) );
    aon222d1 U5363 ( .a1(n13099), .a2(n12509), .b1(n13697), .b2(n13519), .c1(
        n13696), .c2(n12508), .z(n13354) );
    oai221d1 U5364 ( .a1(n12897), .a2(n12885), .b1(n13518), .b2(n12883), .c(
        n12899), .zn(n13353) );
    in01d1 U5365 ( .i(bd_mem_au_count[1]), .zn(n13518) );
    aon222d1 U5366 ( .a1(n12509), .a2(bd_mem_au_count11744_2_), .b1(n13693), 
        .b2(n13519), .c1(n13675), .c2(n12508), .z(n13352) );
    aon222d1 U5367 ( .a1(bd_mem_au_count11744_3_), .a2(n12509), .b1(n13694), 
        .b2(n13519), .c1(n13676), .c2(n12508), .z(n13351) );
    aon222d1 U5369 ( .a1(n12509), .a2(bd_mem_au_count11744_5_), .b1(n13699), 
        .b2(n13519), .c1(n13677), .c2(n12508), .z(n13349) );
    in01d1 U5370 ( .i(n12885), .zn(n13519) );
    nr02e1 U5371 ( .a1(s_sd_dat[3]), .b1(bt_rst), .zn(bd_sd_dat11062_3_) );
    nr02e1 U5372 ( .a1(s_sd_dat[2]), .b1(bt_rst), .zn(bd_sd_dat11062_2_) );
    nr02e1 U5373 ( .a1(s_sd_dat[1]), .b1(bt_rst), .zn(bd_sd_dat11062_1_) );
    nr02e1 U5374 ( .a1(s_sd_dat[0]), .b1(bt_rst), .zn(bd_sd_dat11062_0_) );
    oai21d1 U5375 ( .a1(n13701), .a2(n12662), .b(n12656), .zn(
        bd_au_state11074_0_) );
    nr03d2 U5376 ( .a1(bd_overflow), .a2(n12915), .a3(s_sd_init), .zn(
        b_cpu_req11098) );
    oai32d1 U5377 ( .a1(n13582), .a2(n12730), .a3(bd_underflow), .b1(n12641), 
        .b2(n12652), .zn(bd_cpu_irq011148) );
    nr02e1 U5378 ( .a1(stfd_byt_cnt11157_9_), .b1(bt_rst), .zn(
        stfd_byt_cnt11156_9_) );
    oai211d2 U5379 ( .a1(n13542), .a2(n13032), .b(n12586), .c(n12568), .zn(
        n13120) );
    an04d1 U5380 ( .a1(n12583), .a2(n12537), .a3(n13241), .a4(n13124), .z(
        n12540) );
    oai211d2 U5382 ( .a1(bd_bm_count_32b11631_0_), .a2(n12946), .b(n12868), 
        .c(n12869), .zn(n13335) );
    aon222d1 U5383 ( .a1(n12504), .a2(bd_bm_count_32b11622_8_), .b1(n12505), 
        .b2(bd_bm_count_32b11631_8_), .c1(bd_bm_count[7]), .c2(n13059), .z(
        n13327) );
    aon222d1 U5384 ( .a1(n12504), .a2(bd_bm_count_32b11622_10_), .b1(
        bd_bm_count_32b11631_10_), .b2(n12505), .c1(bd_bm_count[9]), .c2(
        n13059), .z(n13325) );
    aon222d1 U5385 ( .a1(n12504), .a2(bd_bm_count_32b11622_7_), .b1(
        bd_bm_count_32b11631_7_), .b2(n12505), .c1(bd_bm_count[6]), .c2(n13059
        ), .z(n13328) );
    aon222d1 U5386 ( .a1(n12504), .a2(bd_bm_count_32b11622_1_), .b1(n12505), 
        .b2(bd_bm_count_32b11631_1_), .c1(bd_bm_count[0]), .c2(n13059), .z(
        n13334) );
    aon222d1 U5387 ( .a1(n12504), .a2(bd_bm_count_32b11622_11_), .b1(n12505), 
        .b2(bd_bm_count_32b11631_11_), .c1(bd_bm_count[10]), .c2(n13059), .z(
        n13324) );
    aon222d1 U5388 ( .a1(n12504), .a2(bd_bm_count_32b11622_6_), .b1(
        bd_bm_count_32b11631_6_), .b2(n12505), .c1(bd_bm_count[5]), .c2(n13059
        ), .z(n13329) );
    aon222d1 U5389 ( .a1(n12504), .a2(bd_bm_count_32b11622_12_), .b1(
        bd_bm_count_32b11631_12_), .b2(n12505), .c1(bd_bm_count[11]), .c2(
        n13059), .z(n13323) );
    aon222d1 U5390 ( .a1(n12504), .a2(bd_bm_count_32b11622_5_), .b1(
        bd_bm_count_32b11631_5_), .b2(n12505), .c1(bd_bm_count[4]), .c2(n13059
        ), .z(n13330) );
    aon222d1 U5391 ( .a1(n12504), .a2(bd_bm_count_32b11622_3_), .b1(
        bd_bm_count_32b11631_3_), .b2(n12505), .c1(bd_bm_count[2]), .c2(n13059
        ), .z(n13332) );
    aon222d1 U5392 ( .a1(n12504), .a2(bd_bm_count_32b11622_4_), .b1(
        bd_bm_count_32b11631_4_), .b2(n12505), .c1(bd_bm_count[3]), .c2(n13059
        ), .z(n13331) );
    aon222d1 U5393 ( .a1(n12504), .a2(bd_bm_count_32b11622_9_), .b1(
        bd_bm_count_32b11631_9_), .b2(n12505), .c1(bd_bm_count[8]), .c2(n13059
        ), .z(n13326) );
    aon222d1 U5394 ( .a1(n12504), .a2(bd_bm_count_32b11622_14_), .b1(n12505), 
        .b2(bd_bm_count_32b11631_14_), .c1(bd_bm_count[13]), .c2(n13059), .z(
        n13321) );
    nd03d1 U5396 ( .a1(n12479), .a2(n13074), .a3(bd_au_state[1]), .zn(n12981)
         );
    nd03d1 U5397 ( .a1(n13081), .a2(n12491), .a3(n13247), .zn(n13285) );
    nd03d1 U5398 ( .a1(n12479), .a2(n13220), .a3(n13219), .zn(n12570) );
    oai221d1 U5399 ( .a1(n12580), .a2(n13231), .b1(n13021), .b2(n13079), .c(
        n13115), .zn(n13113) );
    mx21d1 U5400 ( .i0(n12511), .i1(n13520), .s(n13657), .z(n13370) );
    in01d1 U5401 ( .i(n12912), .zn(n13520) );
    xn03d1 U5402 ( .a1(bd_au_count[1]), .a2(bd_au_count[0]), .a3(n13094), .zn(
        n12879) );
    aon211d1 U5403 ( .a1(n12502), .a2(n13258), .b(n13047), .c(n13257), .z(
        n13049) );
    nd04d2 U5404 ( .a1(n12514), .a3(n13542), .a4(n13023), .a2(n12549), .zn(
        n13080) );
    or03d1 U5405 ( .a1(n13032), .a2(bd_seq_hdr_exist), .a3(bd_gop_hdr_exist), 
        .z(n12481) );
    nd02e1 U5407 ( .a1(n13528), .b1(gt_278_n48), .zn(gt_278_n15) );
    an02d1 U5408 ( .a1(bp_bufval[4]), .a2(n13456), .z(gt_278_n28) );
    nd02d1 U5409 ( .a1(n13457), .a2(bp_bufval[5]), .zn(gt_278_n41) );
    or02d1 U5410 ( .a1(bd_bm_count[9]), .a2(sub_275_2_n199), .z(sub_275_2_n200
        ) );
    nd02d1 U5411 ( .a1(n12521), .a2(n12967), .zn(n12966) );
    in01d1 U5412 ( .i(n12950), .zn(n13521) );
    xn02d1 U5413 ( .a1(bd_bm_count[9]), .a2(sub_275_2_n199), .zn(n13487) );
    an02d1 U5414 ( .a1(bp_bufval[10]), .a2(n13452), .z(gt_278_n20) );
    nd02d1 U5415 ( .a1(n13453), .a2(bp_bufval[11]), .zn(gt_278_n49) );
    nd02d1 U5416 ( .a1(n12523), .a2(n13070), .zn(n13522) );
    in01d1 U5417 ( .i(n13522), .zn(n12561) );
    mi21d1 U5418 ( .i0(n13402), .i1(n13523), .s(n13286), .zn(n13542) );
    in01d1 U5419 ( .i(bd_sd_dat_8_), .zn(n13523) );
    nd02d1 U5420 ( .a1(n13032), .a2(n12568), .zn(n12984) );
    nr02d1 U5421 ( .a1(n12523), .a2(n13034), .zn(n12557) );
    an03d1 U5422 ( .a1(n13526), .a2(n13525), .a3(n13524), .z(n13504) );
    oan31d1 U5423 ( .a1(sub_275_n110), .a2(bd_bm_count[12]), .a3(
        bd_bm_count_32b[14]), .b(n13449), .z(n13524) );
    an03d1 U5424 ( .a1(gte_275_n155), .a2(n13510), .a3(gte_275_n156), .z(
        n13525) );
    nr04d2 U5425 ( .a1(gte_275_n152), .a2(n598_30_), .a3(n598_22_), .a4(n13509
        ), .zn(n13526) );
    an02d1 U5426 ( .a1(bd_cpu_ack_cnt[5]), .a2(n13527), .z(n13229) );
    nr02d1 U5427 ( .a1(bd_cpu_ack_cnt[4]), .a2(bd_cpu_ack_cnt[2]), .zn(n13527)
         );
    or02d1 U5428 ( .a1(bl_v_jpg), .a2(n12502), .z(n13256) );
    xn03d1 U5429 ( .a1(bd_bm_count[13]), .a2(bd_stfd_byt_cnt[12]), .a3(
        add_277_carry_13_), .zn(n13528) );
    nr02d1 U5430 ( .a1(bd_mem_au_count[3]), .a2(sub_526_n89), .zn(sub_526_n82)
         );
    nd02d1 U5431 ( .a1(n13498), .a2(n12537), .zn(n13529) );
    in01d1 U5432 ( .i(n13529), .zn(n12491) );
    nd02d1 U5433 ( .a1(n13032), .a2(n12568), .zn(n12580) );
    oan211d1 U5434 ( .a1(n12978), .a2(n13532), .b(n13531), .c(n13530), .z(
        n12591) );
    nd03d1 U5435 ( .a1(n13075), .a2(n12575), .a3(n13004), .zn(n13530) );
    or04d1 U5436 ( .a1(n13168), .a2(n13082), .a3(n13080), .a4(n12984), .z(
        n13531) );
    mx21d1 U5437 ( .i0(n13169), .i1(n13167), .s(n13411), .z(n13532) );
    an02d1 U5438 ( .a1(n12696), .a2(b_cpu_req), .z(bd_cpu_req_lt11152) );
    oai22h1 U5439 ( .a1(n13588), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[0]), 
        .zn(b_sd_dat11070_0_) );
    oai22h1 U5440 ( .a1(n13589), .a2(n12625), .b1(n13534), .b2(b_buf_rdt[1]), 
        .zn(b_sd_dat11070_1_) );
    oai22h1 U5441 ( .a1(n13591), .a2(n12730), .b1(n13534), .b2(b_buf_rdt[2]), 
        .zn(b_sd_dat11070_2_) );
    oai22h1 U5442 ( .a1(n13593), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[3]), 
        .zn(b_sd_dat11070_3_) );
    oai22h1 U5443 ( .a1(n13595), .a2(n12625), .b1(n13534), .b2(b_buf_rdt[4]), 
        .zn(b_sd_dat11070_4_) );
    oai22h1 U5444 ( .a1(n13597), .a2(n12730), .b1(n13533), .b2(b_buf_rdt[5]), 
        .zn(b_sd_dat11070_5_) );
    oai22h1 U5445 ( .a1(n13599), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[6]), 
        .zn(b_sd_dat11070_6_) );
    oai22h1 U5446 ( .a1(n13601), .a2(n12625), .b1(n13533), .b2(b_buf_rdt[7]), 
        .zn(b_sd_dat11070_7_) );
    oai22h1 U5447 ( .a1(n13603), .a2(n12625), .b1(n13533), .b2(b_buf_rdt[8]), 
        .zn(b_sd_dat11070_8_) );
    oai22h1 U5448 ( .a1(n13605), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[9]), 
        .zn(b_sd_dat11070_9_) );
    oai22h1 U5449 ( .a1(n13607), .a2(n12625), .b1(n13534), .b2(b_buf_rdt[10]), 
        .zn(b_sd_dat11070_10_) );
    oai22h1 U5450 ( .a1(n13609), .a2(n12730), .b1(n13533), .b2(b_buf_rdt[11]), 
        .zn(b_sd_dat11070_11_) );
    oai22h1 U5451 ( .a1(n13612), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[12]), 
        .zn(b_sd_dat11070_12_) );
    oai22h1 U5452 ( .a1(n13613), .a2(n12625), .b1(n13533), .b2(b_buf_rdt[13]), 
        .zn(b_sd_dat11070_13_) );
    oai22h1 U5453 ( .a1(n13615), .a2(n12730), .b1(n13533), .b2(b_buf_rdt[14]), 
        .zn(b_sd_dat11070_14_) );
    oai22h1 U5454 ( .a1(n13617), .a2(n13290), .b1(n13533), .b2(b_buf_rdt[15]), 
        .zn(b_sd_dat11070_15_) );
    oai22h1 U5455 ( .a1(n13619), .a2(n12625), .b1(n13533), .b2(b_buf_rdt[16]), 
        .zn(b_sd_dat11070_16_) );
    oai22h1 U5456 ( .a1(n13621), .a2(n13290), .b1(n13533), .b2(b_buf_rdt[17]), 
        .zn(b_sd_dat11070_17_) );
    oai22h1 U5457 ( .a1(n13623), .a2(n13290), .b1(n13533), .b2(b_buf_rdt[18]), 
        .zn(b_sd_dat11070_18_) );
    oai22h1 U5458 ( .a1(n13625), .a2(n12625), .b1(n13533), .b2(b_buf_rdt[19]), 
        .zn(b_sd_dat11070_19_) );
    in01d1 U5459 ( .i(n13576), .zn(n13533) );
    oai22h1 U5460 ( .a1(n13628), .a2(n13290), .b1(n13534), .b2(b_buf_rdt[20]), 
        .zn(b_sd_dat11070_20_) );
    in01d1 U5461 ( .i(n13576), .zn(n13534) );
    oai22h1 U5462 ( .a1(n13630), .a2(n13290), .b1(n12535), .b2(b_buf_rdt[21]), 
        .zn(b_sd_dat11070_21_) );
    oai22h1 U5463 ( .a1(n13631), .a2(n12625), .b1(n12535), .b2(b_buf_rdt[22]), 
        .zn(b_sd_dat11070_22_) );
    oai22h1 U5464 ( .a1(n13634), .a2(n13290), .b1(n12535), .b2(b_buf_rdt[23]), 
        .zn(b_sd_dat11070_23_) );
    oai22h1 U5465 ( .a1(n13635), .a2(n13290), .b1(n12535), .b2(b_buf_rdt[24]), 
        .zn(b_sd_dat11070_24_) );
    oai22h1 U5466 ( .a1(n13636), .a2(n12625), .b1(n12535), .b2(b_buf_rdt[25]), 
        .zn(b_sd_dat11070_25_) );
    oai22h1 U5467 ( .a1(n13535), .a2(n12766), .b1(n13463), .b2(n13649), .zn(
        bd_sd_adr_3_) );
    oai22h1 U5472 ( .a1(n12529), .a2(n12776), .b1(n13055), .b2(n13680), .zn(
        bd_sd_adr_8_) );
    oai22h1 U5474 ( .a1(n12529), .a2(n12780), .b1(n13055), .b2(n13682), .zn(
        bd_sd_adr_10_) );
    mi21d1 U5480 ( .i0(bt_pulse2), .i1(bt_pulse1), .s(bl_v_dec_mod), .zn(
        n13535) );
    mi21d1 U5482 ( .i0(bt_pulse1), .i1(bt_pulse2), .s(n13704), .zn(n12529) );
    nr02d1 U5483 ( .a1(n13415), .a2(n12591), .zn(n12919) );
    nd02d1 U5484 ( .a1(n12502), .a2(n12762), .zn(n12909) );
    nd02d1 U5485 ( .a1(n13293), .a2(bl_v_dec_mod), .zn(n12730) );
    nr02d1 U5486 ( .a1(n13536), .a2(n12947), .zn(n13336) );
    xn02d1 U5487 ( .a1(n13679), .a2(add_491_carry_5_), .zn(n13536) );
    nd02d1 U5488 ( .a1(n12925), .a2(n13695), .zn(n13206) );
    nd02d1 U5489 ( .a1(n13293), .a2(n13415), .zn(n12662) );
    an02d1 U5490 ( .a1(n13293), .a2(n13537), .z(n13361) );
    aon21d1 U5491 ( .a1(n13702), .a2(n12960), .b(p_mem_pic), .z(n13537) );
    oai22h1 U5492 ( .a1(n13576), .a2(n12938), .b1(n13293), .b2(n13538), .zn(
        n13377) );
    aoi21d2 U5493 ( .a1(n12491), .a2(n12663), .b(n12538), .zn(n12948) );
    an03d1 U5494 ( .a1(n13208), .a2(n12527), .a3(n12549), .z(n13065) );
    nr02d1 U5495 ( .a1(n13019), .a2(n12950), .zn(n12972) );
    mi21d1 U5496 ( .i0(n13003), .i1(n13404), .s(n12582), .zn(n13002) );
    mi21d1 U5497 ( .i0(n13165), .i1(n13166), .s(n12582), .zn(n13220) );
    mi21d1 U5498 ( .i0(bd_sd_dat_11_), .i1(n12550), .s(n13705), .zn(n12549) );
    mi21d1 U5499 ( .i0(n13401), .i1(n13024), .s(n13286), .zn(n13023) );
    an03d1 U5500 ( .a1(n13542), .a2(n12554), .a3(n12967), .z(n12955) );
    mi21d1 U5501 ( .i0(n13016), .i1(n13393), .s(n13704), .zn(n13015) );
    an02d1 U5502 ( .a1(n12554), .a2(n12950), .z(n12553) );
    mi21d1 U5503 ( .i0(n13017), .i1(n13386), .s(n12582), .zn(n12950) );
    an02d1 U5504 ( .a1(n12578), .a2(n12561), .z(n12577) );
    an03d1 U5505 ( .a1(n13209), .a2(n13163), .a3(n12539), .z(n12578) );
    an03d1 U5506 ( .a1(n13162), .a2(n13163), .a3(n13543), .z(n13035) );
    an02d1 U5507 ( .a1(n12578), .a2(n12561), .z(n12547) );
    an03d1 U5508 ( .a1(n13000), .a2(n12564), .a3(n13211), .z(n13075) );
    an03d1 U5509 ( .a1(n13006), .a2(n13008), .a3(n12998), .z(n12564) );
    an03d1 U5510 ( .a1(n13212), .a2(n13011), .a3(n12486), .z(n13211) );
    in01d1 U5511 ( .i(n13002), .zn(n13212) );
    or03d1 U5512 ( .a1(n13089), .a2(n13013), .a3(n13083), .z(n13088) );
    nd02d1 U5513 ( .a1(n12566), .a2(n12557), .zn(n13169) );
    nd03d1 U5514 ( .a1(n12583), .a2(n12955), .a3(n12586), .zn(n12566) );
    mi21d1 U5515 ( .i0(n12526), .i1(bd_sd_dat_24_), .s(n13286), .zn(n12521) );
    nr02d1 U5516 ( .a1(bd_cpu_ack_cnt[1]), .a2(bd_cpu_ack_cnt[5]), .zn(n13200)
         );
    nr02d1 U5517 ( .a1(bd_cpu_ack_cnt[4]), .a2(bd_cpu_ack_cnt[2]), .zn(n13202)
         );
    in01d1 U5518 ( .i(n13021), .zn(n13168) );
    nr02d1 U5519 ( .a1(bd_mem_au_count[2]), .a2(bd_mem_au_count[1]), .zn(
        n13102) );
    in01d1 U5520 ( .i(n12641), .zn(bd_overflow) );
    ni01d2 U5521 ( .i(bd_bm_count_32b[11]), .z(bd_bm_count[10]) );
    mi21d1 U5524 ( .i0(n13175), .i1(n13174), .s(n13286), .zn(b_cpu_irq[1]) );
    nd02e1 U5525 ( .a1(n12591), .b1(bd_cpu_ack_dly), .zn(n13174) );
    in01d1 U5526 ( .i(n13415), .zn(bd_cpu_ack_dly) );
    or02d1 U5527 ( .a1(bd_cpu_ack_cnt[5]), .a2(bd_cpu_ack_cnt[4]), .z(n13539)
         );
    xn02d1 U5528 ( .a1(n13585), .a2(add_465_carry_11_), .zn(n13540) );
    xn02d1 U5529 ( .a1(n13584), .a2(add_465_carry_10_), .zn(n13541) );
    an03d1 U5530 ( .a1(n12972), .a2(n12547), .a3(n12583), .z(n12568) );
    mi21d1 U5531 ( .i0(bd_sd_dat_30_), .i1(n13159), .s(n13704), .zn(n13163) );
    mx21d1 U5532 ( .i0(n12952), .i1(n12949), .s(n12582), .z(n13543) );
    in01d1 U5533 ( .i(n13019), .zn(n12554) );
    mi21d1 U5534 ( .i0(n13014), .i1(n13391), .s(n12588), .zn(n13013) );
    mi21d1 U5535 ( .i0(n13036), .i1(n13035), .s(n13019), .zn(n13034) );
    mi21d1 U5536 ( .i0(n13022), .i1(n13400), .s(n13705), .zn(n13021) );
    in01d1 U5537 ( .i(n13032), .zn(n12967) );
    mi21d1 U5538 ( .i0(n13033), .i1(n13394), .s(n12582), .zn(n13032) );
    ni01d2 U5540 ( .i(bd_bm_count_32b[1]), .z(bd_bm_count[0]) );
    ni01d2 U5541 ( .i(n12588), .z(n12582) );
    nr04d2 U5543 ( .a1(bd_bm_count_32b[14]), .a2(bd_bm_count[8]), .a3(n13552), 
        .a4(n13551), .zn(gte_274_n169) );
    mx21d1 U5544 ( .i0(bp_jpg_enc_sta_adr[6]), .i1(bp_jpg_dec_sta_adr[6]), .s(
        v_dec_mod), .z(n13569) );
    mx21d1 U5545 ( .i0(bp_jpg_enc_sta_adr[7]), .i1(bp_jpg_dec_sta_adr[7]), .s(
        v_dec_mod), .z(n13570) );
    oai31d1 U5546 ( .a1(n13549), .a2(bd_bm_count[12]), .a3(bd_bm_count_32b[14]
        ), .b(n13544), .zn(n603_19_) );
    in01d1 U5547 ( .i(n13511), .zn(n13544) );
    oai221d1 U5548 ( .a1(n13571), .a2(n12813), .b1(n12990), .b2(n13049), .c(
        n12806), .zn(n13303) );
    mi21d1 U5549 ( .i0(bp_jpg_enc_sta_adr[3]), .i1(bp_jpg_dec_sta_adr[3]), .s(
        v_dec_mod), .zn(n12990) );
    aoi22h1 U5550 ( .a1(n12511), .a2(bd_w_adr_c_plus_1_4_), .b1(n12771), .b2(
        n12912), .zn(n13545) );
    in01d1 U5551 ( .i(n13545), .zn(n13371) );
    xn02d1 U5552 ( .a1(bd_bm_count[12]), .a2(n13549), .zn(n13508) );
    oai21d1 U5553 ( .a1(n13547), .a2(n13546), .b(n12979), .zn(n13252) );
    oan21d1 U5554 ( .a1(n12956), .a2(n13553), .b(n12971), .z(n13546) );
    nr02d1 U5555 ( .a1(n13072), .a2(n12521), .zn(n13547) );
    or02d1 U5556 ( .a1(n13415), .a2(n13548), .z(n13091) );
    oan2111d1 U5557 ( .a1(n12542), .a2(n13082), .b(n13224), .c(n13252), .d(
        n13271), .z(n13548) );
    aon22d1 U5558 ( .a1(n13681), .a2(n12944), .b1(n12533), .b2(
        bd_r_adr_r_plus_1_1_), .z(n13319) );
    aon22d1 U5559 ( .a1(n13682), .a2(n12944), .b1(n12533), .b2(
        bd_r_adr_r_plus_1_2_), .z(n13318) );
    aon22d1 U5560 ( .a1(n13693), .a2(n13573), .b1(n12877), .b2(n12506), .z(
        n13345) );
    aon22d1 U5561 ( .a1(n13694), .a2(n13573), .b1(n12875), .b2(n12506), .z(
        n13344) );
    mx21d1 U5562 ( .i0(bd_sd_dat_0_), .i1(n13587), .s(n12582), .z(n13011) );
    or03d1 U5563 ( .a1(bd_bm_count_32b[11]), .a2(bd_bm_count[11]), .a3(
        sub_275_2_n200), .z(n13549) );
    an02d1 U5564 ( .a1(n13571), .a2(bd_w_adr_r_5_), .z(n13550) );
    mi21d1 U5565 ( .i0(bd_sd_dat_0_), .i1(n13587), .s(bl_v_dec_mod), .zn(
        n13498) );
    or03d1 U5566 ( .a1(bd_bm_count[9]), .a2(bd_bm_count[4]), .a3(bd_bm_count
        [1]), .z(n13551) );
    or02d1 U5567 ( .a1(bd_bm_count[2]), .a2(bd_bm_count[6]), .z(n13552) );
    an03d1 U5568 ( .a1(n12523), .a2(n13019), .a3(n12565), .z(n13553) );
    in01d1 U5569 ( .i(n13553), .zn(n13072) );
    xo02d1 U5570 ( .a1(n13586), .a2(add_465_carry_12_), .z(n13501) );
    oai22h1 U5571 ( .a1(n13535), .a2(n13554), .b1(n13463), .b2(n13650), .zn(
        bd_sd_adr_4_) );
    in01d1 U5572 ( .i(n13673), .zn(n13554) );
    oai22h1 U5573 ( .a1(n13535), .a2(n13555), .b1(n13463), .b2(n13651), .zn(
        bd_sd_adr_5_) );
    in01d1 U5574 ( .i(n13653), .zn(n13555) );
    oai22d2 U5575 ( .a1(n12529), .a2(n12771), .b1(n13535), .b2(n13670), .zn(
        bd_sd_adr_6_) );
    in01d1 U5576 ( .i(n13535), .zn(n13055) );
    oai22h1 U5577 ( .a1(n13535), .a2(n13556), .b1(n13463), .b2(n13652), .zn(
        bd_sd_adr_7_) );
    in01d1 U5578 ( .i(n13656), .zn(n13556) );
    oai22h1 U5579 ( .a1(n12529), .a2(n13557), .b1(n13055), .b2(n13681), .zn(
        bd_sd_adr_9_) );
    in01d1 U5580 ( .i(n13691), .zn(n13557) );
    oai22h1 U5581 ( .a1(n12529), .a2(n13558), .b1(n13055), .b2(n13683), .zn(
        bd_sd_adr_11_) );
    in01d1 U5582 ( .i(bd_w_adr_r_3_), .zn(n13558) );
    oai22h1 U5583 ( .a1(n12529), .a2(n13559), .b1(n13055), .b2(n13684), .zn(
        bd_sd_adr_12_) );
    in01d1 U5584 ( .i(bd_w_adr_r_4_), .zn(n13559) );
    oai22h1 U5585 ( .a1(n12529), .a2(n13560), .b1(n13055), .b2(n13685), .zn(
        bd_sd_adr_13_) );
    in01d1 U5586 ( .i(bd_w_adr_r_5_), .zn(n13560) );
    oai22h1 U5587 ( .a1(n12529), .a2(n13571), .b1(n13055), .b2(n13686), .zn(
        bd_sd_adr_14_) );
    oai22h1 U5588 ( .a1(n12529), .a2(n13561), .b1(n13055), .b2(n13687), .zn(
        bd_sd_adr_15_) );
    in01d1 U5589 ( .i(bd_w_adr_r_7_), .zn(n13561) );
    oai22h1 U5590 ( .a1(n13562), .a2(n12529), .b1(n13055), .b2(n13688), .zn(
        bd_sd_adr_16_) );
    in01d1 U5591 ( .i(bd_w_adr_r_8_), .zn(n13562) );
    oai22h1 U5592 ( .a1(n13563), .a2(n12529), .b1(n13055), .b2(n13689), .zn(
        bd_sd_adr_17_) );
    in01d1 U5593 ( .i(bd_w_adr_r_9_), .zn(n13563) );
    oai22h1 U5594 ( .a1(n13564), .a2(n12529), .b1(n13055), .b2(n13690), .zn(
        bd_sd_adr_18_) );
    in01d1 U5595 ( .i(n13692), .zn(n13564) );
    in01d1 U5596 ( .i(n12529), .zn(n13463) );
    mi21d1 U5597 ( .i0(n12985), .i1(b_dec_en), .s(n13565), .zn(n12936) );
    in01d1 U5598 ( .i(bt_pulse3), .zn(n13565) );
    or02d1 U5599 ( .a1(n13227), .a2(n13576), .z(n12926) );
    in01d1 U5600 ( .i(n13576), .zn(n12535) );
    oai22h1 U5601 ( .a1(n13670), .a2(n12909), .b1(n13566), .b2(
        bd_r_adr_c_plus_1_4_), .zn(n13359) );
    an03d1 U5602 ( .a1(n12909), .a2(n12502), .a3(n13051), .z(n13566) );
    in01d1 U5603 ( .i(n13566), .zn(n12906) );
    oai22h1 U5604 ( .a1(n12883), .a2(n13567), .b1(n12509), .b2(
        bd_mem_au_count11744_6_), .zn(n13348) );
    in01d1 U5605 ( .i(n13678), .zn(n13567) );
    mx21d1 U5606 ( .i0(n12944), .i1(n12533), .s(n13568), .z(n13320) );
    in01d1 U5607 ( .i(n13680), .zn(n13568) );
    in01d1 U5608 ( .i(n13569), .zn(n12987) );
    in01d1 U5609 ( .i(n13570), .zn(n12986) );
    in01d1 U5610 ( .i(bd_w_adr_r_6_), .zn(n13571) );
    oai22h1 U5611 ( .a1(n12897), .a2(n12959), .b1(n12879), .b2(n12506), .zn(
        n13346) );
    mi21d1 U5612 ( .i0(bd_seq_hdr_exist), .i1(n13173), .s(bd_cpu_ack_dly), 
        .zn(n12655) );
    oai22h1 U5613 ( .a1(n12888), .a2(n12959), .b1(n12873), .b2(n12506), .zn(
        n13343) );
    oai22h1 U5614 ( .a1(n13572), .a2(n12959), .b1(n12871), .b2(n12506), .zn(
        n13342) );
    in01d1 U5615 ( .i(n13699), .zn(n13572) );
    oan211d1 U5616 ( .a1(d_acc_unit), .a2(n13091), .b(n12696), .c(n13094), .z(
        n13573) );
    in01d1 U5617 ( .i(n13573), .zn(n12959) );
    oai222d1 U5618 ( .a1(n13574), .a2(n13575), .b1(n12888), .b2(n12885), .c1(
        n13700), .c2(n12883), .zn(n13350) );
    in01d1 U5619 ( .i(n12509), .zn(n13574) );
    xn02d1 U5620 ( .a1(bd_mem_au_count[4]), .a2(sub_526_n82), .zn(n13575) );
    nd02e1 U5621 ( .a1(bl_v_dec_mod), .b1(n13293), .zn(n13576) );
    in01d3 U5622 ( .i(n13286), .zn(n12588) );
    in01d1 U5623 ( .i(n13286), .zn(n13705) );
    ni01d1 U5624 ( .i(bd_bm_count[2]), .z(bd_bm_count_32b[3]) );
    in01d3 U5625 ( .i(bt_rst), .zn(n13293) );
    ni01d2 U5626 ( .i(bp_jpg_enc_sta_adr[0]), .z(n13577) );
    ni01d2 U5627 ( .i(bp_jpg_enc_sta_adr[1]), .z(n13578) );
    ni01d2 U5628 ( .i(bp_jpg_enc_sta_adr[2]), .z(n13579) );
    ni01d2 U5629 ( .i(bp_jpg_enc_sta_adr[4]), .z(n13580) );
    ni01d2 U5630 ( .i(bp_jpg_enc_sta_adr[5]), .z(n13581) );
    ni01d2 U5631 ( .i(n13462), .z(n13582) );
    ni01d2 U5632 ( .i(n13413), .z(n13583) );
    ni01d2 U5633 ( .i(bd_stfd_byt_cnt[10]), .z(n13584) );
    ni01d2 U5634 ( .i(bd_stfd_byt_cnt[11]), .z(n13585) );
    in01d1 U5635 ( .i(bd_stfd_byt_cnt[12]), .zn(n13586) );
    in01d1 U5636 ( .i(n13410), .zn(n13587) );
    in01d1 U5637 ( .i(n13587), .zn(n13588) );
    ni01d2 U5638 ( .i(n13590), .z(n13589) );
    ni01d1 U5639 ( .i(n13409), .z(n13590) );
    ni01d2 U5640 ( .i(n13592), .z(n13591) );
    ni01d1 U5641 ( .i(n13408), .z(n13592) );
    ni01d2 U5642 ( .i(n13594), .z(n13593) );
    ni01d1 U5643 ( .i(n13407), .z(n13594) );
    ni01d2 U5644 ( .i(n13596), .z(n13595) );
    ni01d1 U5645 ( .i(n13406), .z(n13596) );
    ni01d2 U5646 ( .i(n13598), .z(n13597) );
    ni01d1 U5647 ( .i(n13405), .z(n13598) );
    ni01d2 U5648 ( .i(n13600), .z(n13599) );
    ni01d1 U5649 ( .i(n13404), .z(n13600) );
    ni01d2 U5650 ( .i(n13602), .z(n13601) );
    ni01d1 U5651 ( .i(n13403), .z(n13602) );
    ni01d2 U5652 ( .i(n13604), .z(n13603) );
    ni01d1 U5653 ( .i(n13402), .z(n13604) );
    ni01d2 U5654 ( .i(n13606), .z(n13605) );
    ni01d1 U5655 ( .i(n13401), .z(n13606) );
    ni01d2 U5656 ( .i(n13608), .z(n13607) );
    ni01d1 U5657 ( .i(n13400), .z(n13608) );
    ni01d2 U5658 ( .i(n13610), .z(n13609) );
    ni01d1 U5659 ( .i(n13399), .z(n13610) );
    in01d1 U5660 ( .i(n13398), .zn(n13611) );
    in01d1 U5661 ( .i(n13611), .zn(n13612) );
    ni01d2 U5662 ( .i(n13614), .z(n13613) );
    ni01d1 U5663 ( .i(n13397), .z(n13614) );
    ni01d2 U5664 ( .i(n13616), .z(n13615) );
    ni01d1 U5665 ( .i(n13396), .z(n13616) );
    ni01d2 U5666 ( .i(n13618), .z(n13617) );
    ni01d1 U5667 ( .i(n13395), .z(n13618) );
    ni01d2 U5668 ( .i(n13620), .z(n13619) );
    ni01d1 U5669 ( .i(n13394), .z(n13620) );
    ni01d2 U5670 ( .i(n13622), .z(n13621) );
    ni01d1 U5671 ( .i(n13393), .z(n13622) );
    ni01d2 U5672 ( .i(n13624), .z(n13623) );
    ni01d1 U5673 ( .i(n13392), .z(n13624) );
    ni01d2 U5674 ( .i(n13626), .z(n13625) );
    ni01d1 U5675 ( .i(n13391), .z(n13626) );
    in01d1 U5676 ( .i(n13390), .zn(n13627) );
    in01d1 U5677 ( .i(n13627), .zn(n13628) );
    in01d1 U5678 ( .i(n13389), .zn(n13629) );
    in01d1 U5679 ( .i(n13629), .zn(n13630) );
    ni01d2 U5680 ( .i(n13632), .z(n13631) );
    ni01d1 U5681 ( .i(n13388), .z(n13632) );
    in01d1 U5682 ( .i(n13387), .zn(n13633) );
    in01d1 U5683 ( .i(n13633), .zn(n13634) );
    in01d1 U5684 ( .i(n12526), .zn(n13635) );
    in01d1 U5685 ( .i(n13071), .zn(n13636) );
    ni01d2 U5686 ( .i(n13638), .z(n13637) );
    ni01d1 U5687 ( .i(n13384), .z(n13638) );
    ni01d2 U5688 ( .i(n13640), .z(n13639) );
    ni01d1 U5689 ( .i(n13383), .z(n13640) );
    in01d1 U5690 ( .i(n13382), .zn(n13641) );
    in01d1 U5691 ( .i(n13641), .zn(n13642) );
    in01d1 U5692 ( .i(n13381), .zn(n13643) );
    in01d1 U5693 ( .i(n13643), .zn(n13644) );
    ni01d2 U5694 ( .i(n13646), .z(n13645) );
    ni01d1 U5695 ( .i(n13380), .z(n13646) );
    ni01d2 U5696 ( .i(n13648), .z(n13647) );
    ni01d1 U5697 ( .i(n13379), .z(n13648) );
    ni01d2 U5698 ( .i(n13667), .z(n13649) );
    ni01d2 U5699 ( .i(n13663), .z(n13650) );
    ni01d2 U5700 ( .i(n13666), .z(n13651) );
    ni01d2 U5701 ( .i(n13669), .z(n13652) );
    ni01d1 U5702 ( .i(bd_r_adr_c_5_), .z(n13656) );
    ni01d2 U5703 ( .i(bd_r_adr_c_3_), .z(n13653) );
    ni01d2 U5704 ( .i(bd_r_adr_c_1_), .z(n13654) );
    ni01d1 U5705 ( .i(bd_cpu_endb), .z(bd_cpu_end) );
    ni01d2 U5706 ( .i(n13658), .z(n13657) );
    ni01d1 U5707 ( .i(bd_w_adr_c_0_), .z(n13658) );
    ni01d2 U5708 ( .i(n13662), .z(n13659) );
    ni01d2 U5709 ( .i(bd_active_once), .z(n13660) );
    in01d1 U5710 ( .i(bd_re_enc_adv), .zn(n13661) );
    in01d1 U5711 ( .i(n13661), .zn(n13662) );
    ni01d2 U5712 ( .i(bd_w_adr_c_2_), .z(n13663) );
    in01d1 U5713 ( .i(n12920), .zn(n13664) );
    in01d1 U5714 ( .i(n13664), .zn(n13665) );
    ni01d2 U5715 ( .i(bd_w_adr_c_3_), .z(n13666) );
    ni01d2 U5716 ( .i(bd_w_adr_c_1_), .z(n13667) );
    ni01d2 U5717 ( .i(bt_pulse4), .z(n13668) );
    ni01d2 U5718 ( .i(bd_w_adr_c_5_), .z(n13669) );
    in01d1 U5719 ( .i(bd_r_adr_c_4_), .zn(n13670) );
    ni01d2 U5720 ( .i(n13672), .z(n13671) );
    ni01d2 U5721 ( .i(bd_r_adr_c_0_), .z(n13672) );
    ni01d2 U5722 ( .i(bd_r_adr_c_2_), .z(n13673) );
    ni01d2 U5723 ( .i(bl_v_jpg_q), .z(n13674) );
    ni01d2 U5724 ( .i(bd_mem_au_count[2]), .z(n13675) );
    ni01d2 U5725 ( .i(bd_mem_au_count[3]), .z(n13676) );
    ni01d2 U5726 ( .i(bd_mem_au_count[5]), .z(n13677) );
    ni01d2 U5727 ( .i(bd_mem_au_count[6]), .z(n13678) );
    ni01d2 U5728 ( .i(bd_cpu_ack_cnt[5]), .z(n13679) );
    ni01d2 U5729 ( .i(bd_r_adr_r_0_), .z(n13680) );
    ni01d2 U5730 ( .i(bd_r_adr_r_1_), .z(n13681) );
    ni01d2 U5731 ( .i(bd_r_adr_r_2_), .z(n13682) );
    ni01d2 U5732 ( .i(bd_r_adr_r_3_), .z(n13683) );
    ni01d2 U5733 ( .i(bd_r_adr_r_4_), .z(n13684) );
    ni01d2 U5734 ( .i(bd_r_adr_r_5_), .z(n13685) );
    ni01d2 U5735 ( .i(bd_r_adr_r_6_), .z(n13686) );
    ni01d2 U5736 ( .i(bd_r_adr_r_7_), .z(n13687) );
    ni01d2 U5737 ( .i(bd_r_adr_r_8_), .z(n13688) );
    ni01d2 U5738 ( .i(bd_r_adr_r_9_), .z(n13689) );
    ni01d2 U5739 ( .i(bd_r_adr_r_10_), .z(n13690) );
    ni01d2 U5740 ( .i(bd_w_adr_r_1_), .z(n13691) );
    ni01d2 U5741 ( .i(bd_w_adr_r_10_), .z(n13692) );
    ni01d2 U5742 ( .i(bd_au_count[2]), .z(n13693) );
    ni01d2 U5743 ( .i(bd_au_count[3]), .z(n13694) );
    ni01d2 U5744 ( .i(bd_cpu_ack_cnt[0]), .z(n13695) );
    ni01d2 U5745 ( .i(n13698), .z(n13696) );
    ni01d2 U5746 ( .i(bd_au_count[0]), .z(n13697) );
    in01d1 U5747 ( .i(n13099), .zn(n13698) );
    ni01d2 U5748 ( .i(bd_au_count[5]), .z(n13699) );
    in01d1 U5749 ( .i(bd_mem_au_count[4]), .zn(n13700) );
    ni01d2 U5750 ( .i(n13411), .z(n13701) );
    ni01d2 U5751 ( .i(bd_mem_en), .z(n13702) );
    ni01d2 U5752 ( .i(bd_stfd_byt_cnt[0]), .z(n13703) );
    in01d3 U5753 ( .i(n13293), .zn(n12622) );
    in01d2 U5754 ( .i(n13293), .zn(n13292) );
    in01d2 U5755 ( .i(n13293), .zn(n12621) );
    in01d2 U5756 ( .i(n13293), .zn(n12619) );
    in01d2 U5757 ( .i(n13293), .zn(n12624) );
    in01d2 U5758 ( .i(n13286), .zn(n13704) );
    in01d4 U5759 ( .i(bl_v_dec_mod), .zn(n13286) );
endmodule
