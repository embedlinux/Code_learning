library verilog;
use verilog.vl_types.all;
entity PLL_LED_tb is
end PLL_LED_tb;
