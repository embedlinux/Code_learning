library verilog;
use verilog.vl_types.all;
entity ff_rcv_crv_tb is
    generic(
        test_data       : integer := 51
    );
end ff_rcv_crv_tb;
