
module Deserializer ( ParOut, ParValid, DecoderParClk, FIFOEmpty, FIFOFull, 
        ParOutClk, SerialIn, FIFOReadCmd, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, FIFOReadCmd, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, SerialClk, SerRxToDecode,
         \FIFO_U1/SM_MemWriteCmd , \FIFO_U1/SM_MemReadCmd ,
         \FIFO_U1/FIFO_SM1/N239 , \FIFO_U1/FIFO_SM1/N236 ,
         \FIFO_U1/FIFO_SM1/N233 , \FIFO_U1/FIFO_SM1/N230 ,
         \FIFO_U1/FIFO_SM1/N227 , \FIFO_U1/FIFO_SM1/N224 ,
         \FIFO_U1/FIFO_SM1/N221 , \FIFO_U1/FIFO_SM1/N218 ,
         \FIFO_U1/FIFO_SM1/N215 , \FIFO_U1/FIFO_SM1/N212 ,
         \FIFO_U1/FIFO_SM1/N211 , \FIFO_U1/FIFO_SM1/N210 ,
         \FIFO_U1/FIFO_SM1/N209 , \FIFO_U1/FIFO_SM1/N200 ,
         \FIFO_U1/FIFO_SM1/N199 , \FIFO_U1/FIFO_SM1/N198 ,
         \FIFO_U1/FIFO_SM1/N189 , \FIFO_U1/FIFO_SM1/N188 ,
         \FIFO_U1/FIFO_SM1/N185 , \FIFO_U1/FIFO_SM1/N184 ,
         \FIFO_U1/FIFO_SM1/N182 , \FIFO_U1/FIFO_SM1/N179 ,
         \FIFO_U1/FIFO_SM1/N176 , \FIFO_U1/FIFO_SM1/N173 ,
         \FIFO_U1/FIFO_SM1/N170 , \FIFO_U1/FIFO_SM1/N167 ,
         \FIFO_U1/FIFO_SM1/N165 , \FIFO_U1/FIFO_SM1/N162 ,
         \FIFO_U1/FIFO_SM1/N159 , \FIFO_U1/FIFO_SM1/N156 ,
         \FIFO_U1/FIFO_SM1/N153 , \FIFO_U1/FIFO_SM1/N150 ,
         \FIFO_U1/FIFO_SM1/N148 , \FIFO_U1/FIFO_SM1/N146 ,
         \FIFO_U1/FIFO_SM1/N144 , \FIFO_U1/FIFO_SM1/N142 ,
         \FIFO_U1/FIFO_SM1/N126 , \FIFO_U1/FIFO_SM1/N125 ,
         \FIFO_U1/FIFO_SM1/N124 , \FIFO_U1/FIFO_SM1/N123 ,
         \FIFO_U1/FIFO_SM1/N122 , \FIFO_U1/FIFO_SM1/N109 ,
         \FIFO_U1/FIFO_SM1/N108 , \FIFO_U1/FIFO_SM1/N107 ,
         \FIFO_U1/FIFO_SM1/N106 , \FIFO_U1/FIFO_SM1/N105 ,
         \FIFO_U1/FIFO_SM1/N92 , \FIFO_U1/FIFO_SM1/N91 ,
         \FIFO_U1/FIFO_SM1/N90 , \FIFO_U1/FIFO_SM1/N89 ,
         \FIFO_U1/FIFO_SM1/N88 , \FIFO_U1/FIFO_SM1/N76 ,
         \FIFO_U1/FIFO_SM1/N75 , \FIFO_U1/FIFO_SM1/N74 ,
         \FIFO_U1/FIFO_SM1/N73 , \FIFO_U1/FIFO_SM1/N72 ,
         \FIFO_U1/FIFO_SM1/CurState[1] , \FIFO_U1/FIFO_SM1/N9 ,
         \FIFO_U1/FIFO_SM1/N8 , \FIFO_U1/FIFO_SM1/N7 , \FIFO_U1/FIFO_SM1/N6 ,
         \FIFO_U1/FIFO_SM1/N5 , \FIFO_U1/FIFO_SM1/N4 , \FIFO_U1/FIFO_SM1/N3 ,
         \FIFO_U1/FIFO_SM1/N2 , \FIFO_U1/FIFO_SM1/N1 , \FIFO_U1/FIFO_SM1/N0 ,
         \FIFO_U1/RegFile1/N2423 , \FIFO_U1/RegFile1/N2420 ,
         \FIFO_U1/RegFile1/N2417 , \FIFO_U1/RegFile1/N2414 ,
         \FIFO_U1/RegFile1/N2411 , \FIFO_U1/RegFile1/N2408 ,
         \FIFO_U1/RegFile1/N2405 , \FIFO_U1/RegFile1/N2402 ,
         \FIFO_U1/RegFile1/N2399 , \FIFO_U1/RegFile1/N2396 ,
         \FIFO_U1/RegFile1/N2393 , \FIFO_U1/RegFile1/N2390 ,
         \FIFO_U1/RegFile1/N2387 , \FIFO_U1/RegFile1/N2384 ,
         \FIFO_U1/RegFile1/N2381 , \FIFO_U1/RegFile1/N2378 ,
         \FIFO_U1/RegFile1/N2375 , \FIFO_U1/RegFile1/N2372 ,
         \FIFO_U1/RegFile1/N2369 , \FIFO_U1/RegFile1/N2366 ,
         \FIFO_U1/RegFile1/N2363 , \FIFO_U1/RegFile1/N2360 ,
         \FIFO_U1/RegFile1/N2357 , \FIFO_U1/RegFile1/N2354 ,
         \FIFO_U1/RegFile1/N2351 , \FIFO_U1/RegFile1/N2348 ,
         \FIFO_U1/RegFile1/N2345 , \FIFO_U1/RegFile1/N2342 ,
         \FIFO_U1/RegFile1/N2339 , \FIFO_U1/RegFile1/N2336 ,
         \FIFO_U1/RegFile1/N2333 , \FIFO_U1/RegFile1/N2330 ,
         \FIFO_U1/RegFile1/N2328 , \FIFO_U1/RegFile1/N2327 ,
         \FIFO_U1/RegFile1/N2262 , \FIFO_U1/RegFile1/N2229 ,
         \FIFO_U1/RegFile1/N2196 , \FIFO_U1/RegFile1/N2163 ,
         \FIFO_U1/RegFile1/N2130 , \FIFO_U1/RegFile1/N2097 ,
         \FIFO_U1/RegFile1/N2064 , \FIFO_U1/RegFile1/N2031 ,
         \FIFO_U1/RegFile1/N1998 , \FIFO_U1/RegFile1/N1965 ,
         \FIFO_U1/RegFile1/N1932 , \FIFO_U1/RegFile1/N1899 ,
         \FIFO_U1/RegFile1/N1866 , \FIFO_U1/RegFile1/N1833 ,
         \FIFO_U1/RegFile1/N1800 , \FIFO_U1/RegFile1/N1767 ,
         \FIFO_U1/RegFile1/N1734 , \FIFO_U1/RegFile1/N1701 ,
         \FIFO_U1/RegFile1/N1668 , \FIFO_U1/RegFile1/N1635 ,
         \FIFO_U1/RegFile1/N1602 , \FIFO_U1/RegFile1/N1569 ,
         \FIFO_U1/RegFile1/N1536 , \FIFO_U1/RegFile1/N1503 ,
         \FIFO_U1/RegFile1/N1470 , \FIFO_U1/RegFile1/N1437 ,
         \FIFO_U1/RegFile1/N1404 , \FIFO_U1/RegFile1/N1371 ,
         \FIFO_U1/RegFile1/N1338 , \FIFO_U1/RegFile1/N1305 ,
         \FIFO_U1/RegFile1/N1272 , \FIFO_U1/RegFile1/N1239 ,
         \FIFO_U1/RegFile1/N113 , \FIFO_U1/RegFile1/N112 ,
         \FIFO_U1/RegFile1/N111 , \FIFO_U1/RegFile1/N110 ,
         \FIFO_U1/RegFile1/N109 , \FIFO_U1/RegFile1/N108 ,
         \FIFO_U1/RegFile1/N107 , \FIFO_U1/RegFile1/N106 ,
         \FIFO_U1/RegFile1/N105 , \FIFO_U1/RegFile1/N104 ,
         \FIFO_U1/RegFile1/N103 , \FIFO_U1/RegFile1/N102 ,
         \FIFO_U1/RegFile1/N101 , \FIFO_U1/RegFile1/N100 ,
         \FIFO_U1/RegFile1/N99 , \FIFO_U1/RegFile1/N98 ,
         \FIFO_U1/RegFile1/N97 , \FIFO_U1/RegFile1/N96 ,
         \FIFO_U1/RegFile1/N95 , \FIFO_U1/RegFile1/N94 ,
         \FIFO_U1/RegFile1/N93 , \FIFO_U1/RegFile1/N92 ,
         \FIFO_U1/RegFile1/N91 , \FIFO_U1/RegFile1/N90 ,
         \FIFO_U1/RegFile1/N89 , \FIFO_U1/RegFile1/N88 ,
         \FIFO_U1/RegFile1/N87 , \FIFO_U1/RegFile1/N86 ,
         \FIFO_U1/RegFile1/N85 , \FIFO_U1/RegFile1/N84 ,
         \FIFO_U1/RegFile1/N83 , \FIFO_U1/RegFile1/N82 ,
         \FIFO_U1/RegFile1/Storage[0][0] , \FIFO_U1/RegFile1/Storage[0][1] ,
         \FIFO_U1/RegFile1/Storage[0][2] , \FIFO_U1/RegFile1/Storage[0][3] ,
         \FIFO_U1/RegFile1/Storage[0][4] , \FIFO_U1/RegFile1/Storage[0][5] ,
         \FIFO_U1/RegFile1/Storage[0][6] , \FIFO_U1/RegFile1/Storage[0][7] ,
         \FIFO_U1/RegFile1/Storage[0][8] , \FIFO_U1/RegFile1/Storage[0][9] ,
         \FIFO_U1/RegFile1/Storage[0][10] , \FIFO_U1/RegFile1/Storage[0][11] ,
         \FIFO_U1/RegFile1/Storage[0][12] , \FIFO_U1/RegFile1/Storage[0][13] ,
         \FIFO_U1/RegFile1/Storage[0][14] , \FIFO_U1/RegFile1/Storage[0][15] ,
         \FIFO_U1/RegFile1/Storage[0][16] , \FIFO_U1/RegFile1/Storage[0][17] ,
         \FIFO_U1/RegFile1/Storage[0][18] , \FIFO_U1/RegFile1/Storage[0][19] ,
         \FIFO_U1/RegFile1/Storage[0][20] , \FIFO_U1/RegFile1/Storage[0][21] ,
         \FIFO_U1/RegFile1/Storage[0][22] , \FIFO_U1/RegFile1/Storage[0][23] ,
         \FIFO_U1/RegFile1/Storage[0][24] , \FIFO_U1/RegFile1/Storage[0][25] ,
         \FIFO_U1/RegFile1/Storage[0][26] , \FIFO_U1/RegFile1/Storage[0][27] ,
         \FIFO_U1/RegFile1/Storage[0][28] , \FIFO_U1/RegFile1/Storage[0][29] ,
         \FIFO_U1/RegFile1/Storage[0][30] , \FIFO_U1/RegFile1/Storage[0][31] ,
         \FIFO_U1/RegFile1/Storage[1][0] , \FIFO_U1/RegFile1/Storage[1][1] ,
         \FIFO_U1/RegFile1/Storage[1][2] , \FIFO_U1/RegFile1/Storage[1][3] ,
         \FIFO_U1/RegFile1/Storage[1][4] , \FIFO_U1/RegFile1/Storage[1][5] ,
         \FIFO_U1/RegFile1/Storage[1][6] , \FIFO_U1/RegFile1/Storage[1][7] ,
         \FIFO_U1/RegFile1/Storage[1][8] , \FIFO_U1/RegFile1/Storage[1][9] ,
         \FIFO_U1/RegFile1/Storage[1][10] , \FIFO_U1/RegFile1/Storage[1][11] ,
         \FIFO_U1/RegFile1/Storage[1][12] , \FIFO_U1/RegFile1/Storage[1][13] ,
         \FIFO_U1/RegFile1/Storage[1][14] , \FIFO_U1/RegFile1/Storage[1][15] ,
         \FIFO_U1/RegFile1/Storage[1][16] , \FIFO_U1/RegFile1/Storage[1][17] ,
         \FIFO_U1/RegFile1/Storage[1][18] , \FIFO_U1/RegFile1/Storage[1][19] ,
         \FIFO_U1/RegFile1/Storage[1][20] , \FIFO_U1/RegFile1/Storage[1][21] ,
         \FIFO_U1/RegFile1/Storage[1][22] , \FIFO_U1/RegFile1/Storage[1][23] ,
         \FIFO_U1/RegFile1/Storage[1][24] , \FIFO_U1/RegFile1/Storage[1][25] ,
         \FIFO_U1/RegFile1/Storage[1][26] , \FIFO_U1/RegFile1/Storage[1][27] ,
         \FIFO_U1/RegFile1/Storage[1][28] , \FIFO_U1/RegFile1/Storage[1][29] ,
         \FIFO_U1/RegFile1/Storage[1][30] , \FIFO_U1/RegFile1/Storage[1][31] ,
         \FIFO_U1/RegFile1/Storage[2][0] , \FIFO_U1/RegFile1/Storage[2][1] ,
         \FIFO_U1/RegFile1/Storage[2][2] , \FIFO_U1/RegFile1/Storage[2][3] ,
         \FIFO_U1/RegFile1/Storage[2][4] , \FIFO_U1/RegFile1/Storage[2][5] ,
         \FIFO_U1/RegFile1/Storage[2][6] , \FIFO_U1/RegFile1/Storage[2][7] ,
         \FIFO_U1/RegFile1/Storage[2][8] , \FIFO_U1/RegFile1/Storage[2][9] ,
         \FIFO_U1/RegFile1/Storage[2][10] , \FIFO_U1/RegFile1/Storage[2][11] ,
         \FIFO_U1/RegFile1/Storage[2][12] , \FIFO_U1/RegFile1/Storage[2][13] ,
         \FIFO_U1/RegFile1/Storage[2][14] , \FIFO_U1/RegFile1/Storage[2][15] ,
         \FIFO_U1/RegFile1/Storage[2][16] , \FIFO_U1/RegFile1/Storage[2][17] ,
         \FIFO_U1/RegFile1/Storage[2][18] , \FIFO_U1/RegFile1/Storage[2][19] ,
         \FIFO_U1/RegFile1/Storage[2][20] , \FIFO_U1/RegFile1/Storage[2][21] ,
         \FIFO_U1/RegFile1/Storage[2][22] , \FIFO_U1/RegFile1/Storage[2][23] ,
         \FIFO_U1/RegFile1/Storage[2][24] , \FIFO_U1/RegFile1/Storage[2][25] ,
         \FIFO_U1/RegFile1/Storage[2][26] , \FIFO_U1/RegFile1/Storage[2][27] ,
         \FIFO_U1/RegFile1/Storage[2][28] , \FIFO_U1/RegFile1/Storage[2][29] ,
         \FIFO_U1/RegFile1/Storage[2][30] , \FIFO_U1/RegFile1/Storage[2][31] ,
         \FIFO_U1/RegFile1/Storage[3][0] , \FIFO_U1/RegFile1/Storage[3][1] ,
         \FIFO_U1/RegFile1/Storage[3][2] , \FIFO_U1/RegFile1/Storage[3][3] ,
         \FIFO_U1/RegFile1/Storage[3][4] , \FIFO_U1/RegFile1/Storage[3][5] ,
         \FIFO_U1/RegFile1/Storage[3][6] , \FIFO_U1/RegFile1/Storage[3][7] ,
         \FIFO_U1/RegFile1/Storage[3][8] , \FIFO_U1/RegFile1/Storage[3][9] ,
         \FIFO_U1/RegFile1/Storage[3][10] , \FIFO_U1/RegFile1/Storage[3][11] ,
         \FIFO_U1/RegFile1/Storage[3][12] , \FIFO_U1/RegFile1/Storage[3][13] ,
         \FIFO_U1/RegFile1/Storage[3][14] , \FIFO_U1/RegFile1/Storage[3][15] ,
         \FIFO_U1/RegFile1/Storage[3][16] , \FIFO_U1/RegFile1/Storage[3][17] ,
         \FIFO_U1/RegFile1/Storage[3][18] , \FIFO_U1/RegFile1/Storage[3][19] ,
         \FIFO_U1/RegFile1/Storage[3][20] , \FIFO_U1/RegFile1/Storage[3][21] ,
         \FIFO_U1/RegFile1/Storage[3][22] , \FIFO_U1/RegFile1/Storage[3][23] ,
         \FIFO_U1/RegFile1/Storage[3][24] , \FIFO_U1/RegFile1/Storage[3][25] ,
         \FIFO_U1/RegFile1/Storage[3][26] , \FIFO_U1/RegFile1/Storage[3][27] ,
         \FIFO_U1/RegFile1/Storage[3][28] , \FIFO_U1/RegFile1/Storage[3][29] ,
         \FIFO_U1/RegFile1/Storage[3][30] , \FIFO_U1/RegFile1/Storage[3][31] ,
         \FIFO_U1/RegFile1/Storage[4][0] , \FIFO_U1/RegFile1/Storage[4][1] ,
         \FIFO_U1/RegFile1/Storage[4][2] , \FIFO_U1/RegFile1/Storage[4][3] ,
         \FIFO_U1/RegFile1/Storage[4][4] , \FIFO_U1/RegFile1/Storage[4][5] ,
         \FIFO_U1/RegFile1/Storage[4][6] , \FIFO_U1/RegFile1/Storage[4][7] ,
         \FIFO_U1/RegFile1/Storage[4][8] , \FIFO_U1/RegFile1/Storage[4][9] ,
         \FIFO_U1/RegFile1/Storage[4][10] , \FIFO_U1/RegFile1/Storage[4][11] ,
         \FIFO_U1/RegFile1/Storage[4][12] , \FIFO_U1/RegFile1/Storage[4][13] ,
         \FIFO_U1/RegFile1/Storage[4][14] , \FIFO_U1/RegFile1/Storage[4][15] ,
         \FIFO_U1/RegFile1/Storage[4][16] , \FIFO_U1/RegFile1/Storage[4][17] ,
         \FIFO_U1/RegFile1/Storage[4][18] , \FIFO_U1/RegFile1/Storage[4][19] ,
         \FIFO_U1/RegFile1/Storage[4][20] , \FIFO_U1/RegFile1/Storage[4][21] ,
         \FIFO_U1/RegFile1/Storage[4][22] , \FIFO_U1/RegFile1/Storage[4][23] ,
         \FIFO_U1/RegFile1/Storage[4][24] , \FIFO_U1/RegFile1/Storage[4][25] ,
         \FIFO_U1/RegFile1/Storage[4][26] , \FIFO_U1/RegFile1/Storage[4][27] ,
         \FIFO_U1/RegFile1/Storage[4][28] , \FIFO_U1/RegFile1/Storage[4][29] ,
         \FIFO_U1/RegFile1/Storage[4][30] , \FIFO_U1/RegFile1/Storage[4][31] ,
         \FIFO_U1/RegFile1/Storage[5][0] , \FIFO_U1/RegFile1/Storage[5][1] ,
         \FIFO_U1/RegFile1/Storage[5][2] , \FIFO_U1/RegFile1/Storage[5][3] ,
         \FIFO_U1/RegFile1/Storage[5][4] , \FIFO_U1/RegFile1/Storage[5][5] ,
         \FIFO_U1/RegFile1/Storage[5][6] , \FIFO_U1/RegFile1/Storage[5][7] ,
         \FIFO_U1/RegFile1/Storage[5][8] , \FIFO_U1/RegFile1/Storage[5][9] ,
         \FIFO_U1/RegFile1/Storage[5][10] , \FIFO_U1/RegFile1/Storage[5][11] ,
         \FIFO_U1/RegFile1/Storage[5][12] , \FIFO_U1/RegFile1/Storage[5][13] ,
         \FIFO_U1/RegFile1/Storage[5][14] , \FIFO_U1/RegFile1/Storage[5][15] ,
         \FIFO_U1/RegFile1/Storage[5][16] , \FIFO_U1/RegFile1/Storage[5][17] ,
         \FIFO_U1/RegFile1/Storage[5][18] , \FIFO_U1/RegFile1/Storage[5][19] ,
         \FIFO_U1/RegFile1/Storage[5][20] , \FIFO_U1/RegFile1/Storage[5][21] ,
         \FIFO_U1/RegFile1/Storage[5][22] , \FIFO_U1/RegFile1/Storage[5][23] ,
         \FIFO_U1/RegFile1/Storage[5][24] , \FIFO_U1/RegFile1/Storage[5][25] ,
         \FIFO_U1/RegFile1/Storage[5][26] , \FIFO_U1/RegFile1/Storage[5][27] ,
         \FIFO_U1/RegFile1/Storage[5][28] , \FIFO_U1/RegFile1/Storage[5][29] ,
         \FIFO_U1/RegFile1/Storage[5][30] , \FIFO_U1/RegFile1/Storage[5][31] ,
         \FIFO_U1/RegFile1/Storage[6][0] , \FIFO_U1/RegFile1/Storage[6][1] ,
         \FIFO_U1/RegFile1/Storage[6][2] , \FIFO_U1/RegFile1/Storage[6][3] ,
         \FIFO_U1/RegFile1/Storage[6][4] , \FIFO_U1/RegFile1/Storage[6][5] ,
         \FIFO_U1/RegFile1/Storage[6][6] , \FIFO_U1/RegFile1/Storage[6][7] ,
         \FIFO_U1/RegFile1/Storage[6][8] , \FIFO_U1/RegFile1/Storage[6][9] ,
         \FIFO_U1/RegFile1/Storage[6][10] , \FIFO_U1/RegFile1/Storage[6][11] ,
         \FIFO_U1/RegFile1/Storage[6][12] , \FIFO_U1/RegFile1/Storage[6][13] ,
         \FIFO_U1/RegFile1/Storage[6][14] , \FIFO_U1/RegFile1/Storage[6][15] ,
         \FIFO_U1/RegFile1/Storage[6][16] , \FIFO_U1/RegFile1/Storage[6][17] ,
         \FIFO_U1/RegFile1/Storage[6][18] , \FIFO_U1/RegFile1/Storage[6][19] ,
         \FIFO_U1/RegFile1/Storage[6][20] , \FIFO_U1/RegFile1/Storage[6][21] ,
         \FIFO_U1/RegFile1/Storage[6][22] , \FIFO_U1/RegFile1/Storage[6][23] ,
         \FIFO_U1/RegFile1/Storage[6][24] , \FIFO_U1/RegFile1/Storage[6][25] ,
         \FIFO_U1/RegFile1/Storage[6][26] , \FIFO_U1/RegFile1/Storage[6][27] ,
         \FIFO_U1/RegFile1/Storage[6][28] , \FIFO_U1/RegFile1/Storage[6][29] ,
         \FIFO_U1/RegFile1/Storage[6][30] , \FIFO_U1/RegFile1/Storage[6][31] ,
         \FIFO_U1/RegFile1/Storage[7][0] , \FIFO_U1/RegFile1/Storage[7][1] ,
         \FIFO_U1/RegFile1/Storage[7][2] , \FIFO_U1/RegFile1/Storage[7][3] ,
         \FIFO_U1/RegFile1/Storage[7][4] , \FIFO_U1/RegFile1/Storage[7][5] ,
         \FIFO_U1/RegFile1/Storage[7][6] , \FIFO_U1/RegFile1/Storage[7][7] ,
         \FIFO_U1/RegFile1/Storage[7][8] , \FIFO_U1/RegFile1/Storage[7][9] ,
         \FIFO_U1/RegFile1/Storage[7][10] , \FIFO_U1/RegFile1/Storage[7][11] ,
         \FIFO_U1/RegFile1/Storage[7][12] , \FIFO_U1/RegFile1/Storage[7][13] ,
         \FIFO_U1/RegFile1/Storage[7][14] , \FIFO_U1/RegFile1/Storage[7][15] ,
         \FIFO_U1/RegFile1/Storage[7][16] , \FIFO_U1/RegFile1/Storage[7][17] ,
         \FIFO_U1/RegFile1/Storage[7][18] , \FIFO_U1/RegFile1/Storage[7][19] ,
         \FIFO_U1/RegFile1/Storage[7][20] , \FIFO_U1/RegFile1/Storage[7][21] ,
         \FIFO_U1/RegFile1/Storage[7][22] , \FIFO_U1/RegFile1/Storage[7][23] ,
         \FIFO_U1/RegFile1/Storage[7][24] , \FIFO_U1/RegFile1/Storage[7][25] ,
         \FIFO_U1/RegFile1/Storage[7][26] , \FIFO_U1/RegFile1/Storage[7][27] ,
         \FIFO_U1/RegFile1/Storage[7][28] , \FIFO_U1/RegFile1/Storage[7][29] ,
         \FIFO_U1/RegFile1/Storage[7][30] , \FIFO_U1/RegFile1/Storage[7][31] ,
         \FIFO_U1/RegFile1/Storage[8][0] , \FIFO_U1/RegFile1/Storage[8][1] ,
         \FIFO_U1/RegFile1/Storage[8][2] , \FIFO_U1/RegFile1/Storage[8][3] ,
         \FIFO_U1/RegFile1/Storage[8][4] , \FIFO_U1/RegFile1/Storage[8][5] ,
         \FIFO_U1/RegFile1/Storage[8][6] , \FIFO_U1/RegFile1/Storage[8][7] ,
         \FIFO_U1/RegFile1/Storage[8][8] , \FIFO_U1/RegFile1/Storage[8][9] ,
         \FIFO_U1/RegFile1/Storage[8][10] , \FIFO_U1/RegFile1/Storage[8][11] ,
         \FIFO_U1/RegFile1/Storage[8][12] , \FIFO_U1/RegFile1/Storage[8][13] ,
         \FIFO_U1/RegFile1/Storage[8][14] , \FIFO_U1/RegFile1/Storage[8][15] ,
         \FIFO_U1/RegFile1/Storage[8][16] , \FIFO_U1/RegFile1/Storage[8][17] ,
         \FIFO_U1/RegFile1/Storage[8][18] , \FIFO_U1/RegFile1/Storage[8][19] ,
         \FIFO_U1/RegFile1/Storage[8][20] , \FIFO_U1/RegFile1/Storage[8][21] ,
         \FIFO_U1/RegFile1/Storage[8][22] , \FIFO_U1/RegFile1/Storage[8][23] ,
         \FIFO_U1/RegFile1/Storage[8][24] , \FIFO_U1/RegFile1/Storage[8][25] ,
         \FIFO_U1/RegFile1/Storage[8][26] , \FIFO_U1/RegFile1/Storage[8][27] ,
         \FIFO_U1/RegFile1/Storage[8][28] , \FIFO_U1/RegFile1/Storage[8][29] ,
         \FIFO_U1/RegFile1/Storage[8][30] , \FIFO_U1/RegFile1/Storage[8][31] ,
         \FIFO_U1/RegFile1/Storage[9][0] , \FIFO_U1/RegFile1/Storage[9][1] ,
         \FIFO_U1/RegFile1/Storage[9][2] , \FIFO_U1/RegFile1/Storage[9][3] ,
         \FIFO_U1/RegFile1/Storage[9][4] , \FIFO_U1/RegFile1/Storage[9][5] ,
         \FIFO_U1/RegFile1/Storage[9][6] , \FIFO_U1/RegFile1/Storage[9][7] ,
         \FIFO_U1/RegFile1/Storage[9][8] , \FIFO_U1/RegFile1/Storage[9][9] ,
         \FIFO_U1/RegFile1/Storage[9][10] , \FIFO_U1/RegFile1/Storage[9][11] ,
         \FIFO_U1/RegFile1/Storage[9][12] , \FIFO_U1/RegFile1/Storage[9][13] ,
         \FIFO_U1/RegFile1/Storage[9][14] , \FIFO_U1/RegFile1/Storage[9][15] ,
         \FIFO_U1/RegFile1/Storage[9][16] , \FIFO_U1/RegFile1/Storage[9][17] ,
         \FIFO_U1/RegFile1/Storage[9][18] , \FIFO_U1/RegFile1/Storage[9][19] ,
         \FIFO_U1/RegFile1/Storage[9][20] , \FIFO_U1/RegFile1/Storage[9][21] ,
         \FIFO_U1/RegFile1/Storage[9][22] , \FIFO_U1/RegFile1/Storage[9][23] ,
         \FIFO_U1/RegFile1/Storage[9][24] , \FIFO_U1/RegFile1/Storage[9][25] ,
         \FIFO_U1/RegFile1/Storage[9][26] , \FIFO_U1/RegFile1/Storage[9][27] ,
         \FIFO_U1/RegFile1/Storage[9][28] , \FIFO_U1/RegFile1/Storage[9][29] ,
         \FIFO_U1/RegFile1/Storage[9][30] , \FIFO_U1/RegFile1/Storage[9][31] ,
         \FIFO_U1/RegFile1/Storage[10][0] , \FIFO_U1/RegFile1/Storage[10][1] ,
         \FIFO_U1/RegFile1/Storage[10][2] , \FIFO_U1/RegFile1/Storage[10][3] ,
         \FIFO_U1/RegFile1/Storage[10][4] , \FIFO_U1/RegFile1/Storage[10][5] ,
         \FIFO_U1/RegFile1/Storage[10][6] , \FIFO_U1/RegFile1/Storage[10][7] ,
         \FIFO_U1/RegFile1/Storage[10][8] , \FIFO_U1/RegFile1/Storage[10][9] ,
         \FIFO_U1/RegFile1/Storage[10][10] ,
         \FIFO_U1/RegFile1/Storage[10][11] ,
         \FIFO_U1/RegFile1/Storage[10][12] ,
         \FIFO_U1/RegFile1/Storage[10][13] ,
         \FIFO_U1/RegFile1/Storage[10][14] ,
         \FIFO_U1/RegFile1/Storage[10][15] ,
         \FIFO_U1/RegFile1/Storage[10][16] ,
         \FIFO_U1/RegFile1/Storage[10][17] ,
         \FIFO_U1/RegFile1/Storage[10][18] ,
         \FIFO_U1/RegFile1/Storage[10][19] ,
         \FIFO_U1/RegFile1/Storage[10][20] ,
         \FIFO_U1/RegFile1/Storage[10][21] ,
         \FIFO_U1/RegFile1/Storage[10][22] ,
         \FIFO_U1/RegFile1/Storage[10][23] ,
         \FIFO_U1/RegFile1/Storage[10][24] ,
         \FIFO_U1/RegFile1/Storage[10][25] ,
         \FIFO_U1/RegFile1/Storage[10][26] ,
         \FIFO_U1/RegFile1/Storage[10][27] ,
         \FIFO_U1/RegFile1/Storage[10][28] ,
         \FIFO_U1/RegFile1/Storage[10][29] ,
         \FIFO_U1/RegFile1/Storage[10][30] ,
         \FIFO_U1/RegFile1/Storage[10][31] , \FIFO_U1/RegFile1/Storage[11][0] ,
         \FIFO_U1/RegFile1/Storage[11][1] , \FIFO_U1/RegFile1/Storage[11][2] ,
         \FIFO_U1/RegFile1/Storage[11][3] , \FIFO_U1/RegFile1/Storage[11][4] ,
         \FIFO_U1/RegFile1/Storage[11][5] , \FIFO_U1/RegFile1/Storage[11][6] ,
         \FIFO_U1/RegFile1/Storage[11][7] , \FIFO_U1/RegFile1/Storage[11][8] ,
         \FIFO_U1/RegFile1/Storage[11][9] , \FIFO_U1/RegFile1/Storage[11][10] ,
         \FIFO_U1/RegFile1/Storage[11][11] ,
         \FIFO_U1/RegFile1/Storage[11][12] ,
         \FIFO_U1/RegFile1/Storage[11][13] ,
         \FIFO_U1/RegFile1/Storage[11][14] ,
         \FIFO_U1/RegFile1/Storage[11][15] ,
         \FIFO_U1/RegFile1/Storage[11][16] ,
         \FIFO_U1/RegFile1/Storage[11][17] ,
         \FIFO_U1/RegFile1/Storage[11][18] ,
         \FIFO_U1/RegFile1/Storage[11][19] ,
         \FIFO_U1/RegFile1/Storage[11][20] ,
         \FIFO_U1/RegFile1/Storage[11][21] ,
         \FIFO_U1/RegFile1/Storage[11][22] ,
         \FIFO_U1/RegFile1/Storage[11][23] ,
         \FIFO_U1/RegFile1/Storage[11][24] ,
         \FIFO_U1/RegFile1/Storage[11][25] ,
         \FIFO_U1/RegFile1/Storage[11][26] ,
         \FIFO_U1/RegFile1/Storage[11][27] ,
         \FIFO_U1/RegFile1/Storage[11][28] ,
         \FIFO_U1/RegFile1/Storage[11][29] ,
         \FIFO_U1/RegFile1/Storage[11][30] ,
         \FIFO_U1/RegFile1/Storage[11][31] , \FIFO_U1/RegFile1/Storage[12][0] ,
         \FIFO_U1/RegFile1/Storage[12][1] , \FIFO_U1/RegFile1/Storage[12][2] ,
         \FIFO_U1/RegFile1/Storage[12][3] , \FIFO_U1/RegFile1/Storage[12][4] ,
         \FIFO_U1/RegFile1/Storage[12][5] , \FIFO_U1/RegFile1/Storage[12][6] ,
         \FIFO_U1/RegFile1/Storage[12][7] , \FIFO_U1/RegFile1/Storage[12][8] ,
         \FIFO_U1/RegFile1/Storage[12][9] , \FIFO_U1/RegFile1/Storage[12][10] ,
         \FIFO_U1/RegFile1/Storage[12][11] ,
         \FIFO_U1/RegFile1/Storage[12][12] ,
         \FIFO_U1/RegFile1/Storage[12][13] ,
         \FIFO_U1/RegFile1/Storage[12][14] ,
         \FIFO_U1/RegFile1/Storage[12][15] ,
         \FIFO_U1/RegFile1/Storage[12][16] ,
         \FIFO_U1/RegFile1/Storage[12][17] ,
         \FIFO_U1/RegFile1/Storage[12][18] ,
         \FIFO_U1/RegFile1/Storage[12][19] ,
         \FIFO_U1/RegFile1/Storage[12][20] ,
         \FIFO_U1/RegFile1/Storage[12][21] ,
         \FIFO_U1/RegFile1/Storage[12][22] ,
         \FIFO_U1/RegFile1/Storage[12][23] ,
         \FIFO_U1/RegFile1/Storage[12][24] ,
         \FIFO_U1/RegFile1/Storage[12][25] ,
         \FIFO_U1/RegFile1/Storage[12][26] ,
         \FIFO_U1/RegFile1/Storage[12][27] ,
         \FIFO_U1/RegFile1/Storage[12][28] ,
         \FIFO_U1/RegFile1/Storage[12][29] ,
         \FIFO_U1/RegFile1/Storage[12][30] ,
         \FIFO_U1/RegFile1/Storage[12][31] , \FIFO_U1/RegFile1/Storage[13][0] ,
         \FIFO_U1/RegFile1/Storage[13][1] , \FIFO_U1/RegFile1/Storage[13][2] ,
         \FIFO_U1/RegFile1/Storage[13][3] , \FIFO_U1/RegFile1/Storage[13][4] ,
         \FIFO_U1/RegFile1/Storage[13][5] , \FIFO_U1/RegFile1/Storage[13][6] ,
         \FIFO_U1/RegFile1/Storage[13][7] , \FIFO_U1/RegFile1/Storage[13][8] ,
         \FIFO_U1/RegFile1/Storage[13][9] , \FIFO_U1/RegFile1/Storage[13][10] ,
         \FIFO_U1/RegFile1/Storage[13][11] ,
         \FIFO_U1/RegFile1/Storage[13][12] ,
         \FIFO_U1/RegFile1/Storage[13][13] ,
         \FIFO_U1/RegFile1/Storage[13][14] ,
         \FIFO_U1/RegFile1/Storage[13][15] ,
         \FIFO_U1/RegFile1/Storage[13][16] ,
         \FIFO_U1/RegFile1/Storage[13][17] ,
         \FIFO_U1/RegFile1/Storage[13][18] ,
         \FIFO_U1/RegFile1/Storage[13][19] ,
         \FIFO_U1/RegFile1/Storage[13][20] ,
         \FIFO_U1/RegFile1/Storage[13][21] ,
         \FIFO_U1/RegFile1/Storage[13][22] ,
         \FIFO_U1/RegFile1/Storage[13][23] ,
         \FIFO_U1/RegFile1/Storage[13][24] ,
         \FIFO_U1/RegFile1/Storage[13][25] ,
         \FIFO_U1/RegFile1/Storage[13][26] ,
         \FIFO_U1/RegFile1/Storage[13][27] ,
         \FIFO_U1/RegFile1/Storage[13][28] ,
         \FIFO_U1/RegFile1/Storage[13][29] ,
         \FIFO_U1/RegFile1/Storage[13][30] ,
         \FIFO_U1/RegFile1/Storage[13][31] , \FIFO_U1/RegFile1/Storage[14][0] ,
         \FIFO_U1/RegFile1/Storage[14][1] , \FIFO_U1/RegFile1/Storage[14][2] ,
         \FIFO_U1/RegFile1/Storage[14][3] , \FIFO_U1/RegFile1/Storage[14][4] ,
         \FIFO_U1/RegFile1/Storage[14][5] , \FIFO_U1/RegFile1/Storage[14][6] ,
         \FIFO_U1/RegFile1/Storage[14][7] , \FIFO_U1/RegFile1/Storage[14][8] ,
         \FIFO_U1/RegFile1/Storage[14][9] , \FIFO_U1/RegFile1/Storage[14][10] ,
         \FIFO_U1/RegFile1/Storage[14][11] ,
         \FIFO_U1/RegFile1/Storage[14][12] ,
         \FIFO_U1/RegFile1/Storage[14][13] ,
         \FIFO_U1/RegFile1/Storage[14][14] ,
         \FIFO_U1/RegFile1/Storage[14][15] ,
         \FIFO_U1/RegFile1/Storage[14][16] ,
         \FIFO_U1/RegFile1/Storage[14][17] ,
         \FIFO_U1/RegFile1/Storage[14][18] ,
         \FIFO_U1/RegFile1/Storage[14][19] ,
         \FIFO_U1/RegFile1/Storage[14][20] ,
         \FIFO_U1/RegFile1/Storage[14][21] ,
         \FIFO_U1/RegFile1/Storage[14][22] ,
         \FIFO_U1/RegFile1/Storage[14][23] ,
         \FIFO_U1/RegFile1/Storage[14][24] ,
         \FIFO_U1/RegFile1/Storage[14][25] ,
         \FIFO_U1/RegFile1/Storage[14][26] ,
         \FIFO_U1/RegFile1/Storage[14][27] ,
         \FIFO_U1/RegFile1/Storage[14][28] ,
         \FIFO_U1/RegFile1/Storage[14][29] ,
         \FIFO_U1/RegFile1/Storage[14][30] ,
         \FIFO_U1/RegFile1/Storage[14][31] , \FIFO_U1/RegFile1/Storage[15][0] ,
         \FIFO_U1/RegFile1/Storage[15][1] , \FIFO_U1/RegFile1/Storage[15][2] ,
         \FIFO_U1/RegFile1/Storage[15][3] , \FIFO_U1/RegFile1/Storage[15][4] ,
         \FIFO_U1/RegFile1/Storage[15][5] , \FIFO_U1/RegFile1/Storage[15][6] ,
         \FIFO_U1/RegFile1/Storage[15][7] , \FIFO_U1/RegFile1/Storage[15][8] ,
         \FIFO_U1/RegFile1/Storage[15][9] , \FIFO_U1/RegFile1/Storage[15][10] ,
         \FIFO_U1/RegFile1/Storage[15][11] ,
         \FIFO_U1/RegFile1/Storage[15][12] ,
         \FIFO_U1/RegFile1/Storage[15][13] ,
         \FIFO_U1/RegFile1/Storage[15][14] ,
         \FIFO_U1/RegFile1/Storage[15][15] ,
         \FIFO_U1/RegFile1/Storage[15][16] ,
         \FIFO_U1/RegFile1/Storage[15][17] ,
         \FIFO_U1/RegFile1/Storage[15][18] ,
         \FIFO_U1/RegFile1/Storage[15][19] ,
         \FIFO_U1/RegFile1/Storage[15][20] ,
         \FIFO_U1/RegFile1/Storage[15][21] ,
         \FIFO_U1/RegFile1/Storage[15][22] ,
         \FIFO_U1/RegFile1/Storage[15][23] ,
         \FIFO_U1/RegFile1/Storage[15][24] ,
         \FIFO_U1/RegFile1/Storage[15][25] ,
         \FIFO_U1/RegFile1/Storage[15][26] ,
         \FIFO_U1/RegFile1/Storage[15][27] ,
         \FIFO_U1/RegFile1/Storage[15][28] ,
         \FIFO_U1/RegFile1/Storage[15][29] ,
         \FIFO_U1/RegFile1/Storage[15][30] ,
         \FIFO_U1/RegFile1/Storage[15][31] , \FIFO_U1/RegFile1/Storage[16][0] ,
         \FIFO_U1/RegFile1/Storage[16][1] , \FIFO_U1/RegFile1/Storage[16][2] ,
         \FIFO_U1/RegFile1/Storage[16][3] , \FIFO_U1/RegFile1/Storage[16][4] ,
         \FIFO_U1/RegFile1/Storage[16][5] , \FIFO_U1/RegFile1/Storage[16][6] ,
         \FIFO_U1/RegFile1/Storage[16][7] , \FIFO_U1/RegFile1/Storage[16][8] ,
         \FIFO_U1/RegFile1/Storage[16][9] , \FIFO_U1/RegFile1/Storage[16][10] ,
         \FIFO_U1/RegFile1/Storage[16][11] ,
         \FIFO_U1/RegFile1/Storage[16][12] ,
         \FIFO_U1/RegFile1/Storage[16][13] ,
         \FIFO_U1/RegFile1/Storage[16][14] ,
         \FIFO_U1/RegFile1/Storage[16][15] ,
         \FIFO_U1/RegFile1/Storage[16][16] ,
         \FIFO_U1/RegFile1/Storage[16][17] ,
         \FIFO_U1/RegFile1/Storage[16][18] ,
         \FIFO_U1/RegFile1/Storage[16][19] ,
         \FIFO_U1/RegFile1/Storage[16][20] ,
         \FIFO_U1/RegFile1/Storage[16][21] ,
         \FIFO_U1/RegFile1/Storage[16][22] ,
         \FIFO_U1/RegFile1/Storage[16][23] ,
         \FIFO_U1/RegFile1/Storage[16][24] ,
         \FIFO_U1/RegFile1/Storage[16][25] ,
         \FIFO_U1/RegFile1/Storage[16][26] ,
         \FIFO_U1/RegFile1/Storage[16][27] ,
         \FIFO_U1/RegFile1/Storage[16][28] ,
         \FIFO_U1/RegFile1/Storage[16][29] ,
         \FIFO_U1/RegFile1/Storage[16][30] ,
         \FIFO_U1/RegFile1/Storage[16][31] , \FIFO_U1/RegFile1/Storage[17][0] ,
         \FIFO_U1/RegFile1/Storage[17][1] , \FIFO_U1/RegFile1/Storage[17][2] ,
         \FIFO_U1/RegFile1/Storage[17][3] , \FIFO_U1/RegFile1/Storage[17][4] ,
         \FIFO_U1/RegFile1/Storage[17][5] , \FIFO_U1/RegFile1/Storage[17][6] ,
         \FIFO_U1/RegFile1/Storage[17][7] , \FIFO_U1/RegFile1/Storage[17][8] ,
         \FIFO_U1/RegFile1/Storage[17][9] , \FIFO_U1/RegFile1/Storage[17][10] ,
         \FIFO_U1/RegFile1/Storage[17][11] ,
         \FIFO_U1/RegFile1/Storage[17][12] ,
         \FIFO_U1/RegFile1/Storage[17][13] ,
         \FIFO_U1/RegFile1/Storage[17][14] ,
         \FIFO_U1/RegFile1/Storage[17][15] ,
         \FIFO_U1/RegFile1/Storage[17][16] ,
         \FIFO_U1/RegFile1/Storage[17][17] ,
         \FIFO_U1/RegFile1/Storage[17][18] ,
         \FIFO_U1/RegFile1/Storage[17][19] ,
         \FIFO_U1/RegFile1/Storage[17][20] ,
         \FIFO_U1/RegFile1/Storage[17][21] ,
         \FIFO_U1/RegFile1/Storage[17][22] ,
         \FIFO_U1/RegFile1/Storage[17][23] ,
         \FIFO_U1/RegFile1/Storage[17][24] ,
         \FIFO_U1/RegFile1/Storage[17][25] ,
         \FIFO_U1/RegFile1/Storage[17][26] ,
         \FIFO_U1/RegFile1/Storage[17][27] ,
         \FIFO_U1/RegFile1/Storage[17][28] ,
         \FIFO_U1/RegFile1/Storage[17][29] ,
         \FIFO_U1/RegFile1/Storage[17][30] ,
         \FIFO_U1/RegFile1/Storage[17][31] , \FIFO_U1/RegFile1/Storage[18][0] ,
         \FIFO_U1/RegFile1/Storage[18][1] , \FIFO_U1/RegFile1/Storage[18][2] ,
         \FIFO_U1/RegFile1/Storage[18][3] , \FIFO_U1/RegFile1/Storage[18][4] ,
         \FIFO_U1/RegFile1/Storage[18][5] , \FIFO_U1/RegFile1/Storage[18][6] ,
         \FIFO_U1/RegFile1/Storage[18][7] , \FIFO_U1/RegFile1/Storage[18][8] ,
         \FIFO_U1/RegFile1/Storage[18][9] , \FIFO_U1/RegFile1/Storage[18][10] ,
         \FIFO_U1/RegFile1/Storage[18][11] ,
         \FIFO_U1/RegFile1/Storage[18][12] ,
         \FIFO_U1/RegFile1/Storage[18][13] ,
         \FIFO_U1/RegFile1/Storage[18][14] ,
         \FIFO_U1/RegFile1/Storage[18][15] ,
         \FIFO_U1/RegFile1/Storage[18][16] ,
         \FIFO_U1/RegFile1/Storage[18][17] ,
         \FIFO_U1/RegFile1/Storage[18][18] ,
         \FIFO_U1/RegFile1/Storage[18][19] ,
         \FIFO_U1/RegFile1/Storage[18][20] ,
         \FIFO_U1/RegFile1/Storage[18][21] ,
         \FIFO_U1/RegFile1/Storage[18][22] ,
         \FIFO_U1/RegFile1/Storage[18][23] ,
         \FIFO_U1/RegFile1/Storage[18][24] ,
         \FIFO_U1/RegFile1/Storage[18][25] ,
         \FIFO_U1/RegFile1/Storage[18][26] ,
         \FIFO_U1/RegFile1/Storage[18][27] ,
         \FIFO_U1/RegFile1/Storage[18][28] ,
         \FIFO_U1/RegFile1/Storage[18][29] ,
         \FIFO_U1/RegFile1/Storage[18][30] ,
         \FIFO_U1/RegFile1/Storage[18][31] , \FIFO_U1/RegFile1/Storage[19][0] ,
         \FIFO_U1/RegFile1/Storage[19][1] , \FIFO_U1/RegFile1/Storage[19][2] ,
         \FIFO_U1/RegFile1/Storage[19][3] , \FIFO_U1/RegFile1/Storage[19][4] ,
         \FIFO_U1/RegFile1/Storage[19][5] , \FIFO_U1/RegFile1/Storage[19][6] ,
         \FIFO_U1/RegFile1/Storage[19][7] , \FIFO_U1/RegFile1/Storage[19][8] ,
         \FIFO_U1/RegFile1/Storage[19][9] , \FIFO_U1/RegFile1/Storage[19][10] ,
         \FIFO_U1/RegFile1/Storage[19][11] ,
         \FIFO_U1/RegFile1/Storage[19][12] ,
         \FIFO_U1/RegFile1/Storage[19][13] ,
         \FIFO_U1/RegFile1/Storage[19][14] ,
         \FIFO_U1/RegFile1/Storage[19][15] ,
         \FIFO_U1/RegFile1/Storage[19][16] ,
         \FIFO_U1/RegFile1/Storage[19][17] ,
         \FIFO_U1/RegFile1/Storage[19][18] ,
         \FIFO_U1/RegFile1/Storage[19][19] ,
         \FIFO_U1/RegFile1/Storage[19][20] ,
         \FIFO_U1/RegFile1/Storage[19][21] ,
         \FIFO_U1/RegFile1/Storage[19][22] ,
         \FIFO_U1/RegFile1/Storage[19][23] ,
         \FIFO_U1/RegFile1/Storage[19][24] ,
         \FIFO_U1/RegFile1/Storage[19][25] ,
         \FIFO_U1/RegFile1/Storage[19][26] ,
         \FIFO_U1/RegFile1/Storage[19][27] ,
         \FIFO_U1/RegFile1/Storage[19][28] ,
         \FIFO_U1/RegFile1/Storage[19][29] ,
         \FIFO_U1/RegFile1/Storage[19][30] ,
         \FIFO_U1/RegFile1/Storage[19][31] , \FIFO_U1/RegFile1/Storage[20][0] ,
         \FIFO_U1/RegFile1/Storage[20][1] , \FIFO_U1/RegFile1/Storage[20][2] ,
         \FIFO_U1/RegFile1/Storage[20][3] , \FIFO_U1/RegFile1/Storage[20][4] ,
         \FIFO_U1/RegFile1/Storage[20][5] , \FIFO_U1/RegFile1/Storage[20][6] ,
         \FIFO_U1/RegFile1/Storage[20][7] , \FIFO_U1/RegFile1/Storage[20][8] ,
         \FIFO_U1/RegFile1/Storage[20][9] , \FIFO_U1/RegFile1/Storage[20][10] ,
         \FIFO_U1/RegFile1/Storage[20][11] ,
         \FIFO_U1/RegFile1/Storage[20][12] ,
         \FIFO_U1/RegFile1/Storage[20][13] ,
         \FIFO_U1/RegFile1/Storage[20][14] ,
         \FIFO_U1/RegFile1/Storage[20][15] ,
         \FIFO_U1/RegFile1/Storage[20][16] ,
         \FIFO_U1/RegFile1/Storage[20][17] ,
         \FIFO_U1/RegFile1/Storage[20][18] ,
         \FIFO_U1/RegFile1/Storage[20][19] ,
         \FIFO_U1/RegFile1/Storage[20][20] ,
         \FIFO_U1/RegFile1/Storage[20][21] ,
         \FIFO_U1/RegFile1/Storage[20][22] ,
         \FIFO_U1/RegFile1/Storage[20][23] ,
         \FIFO_U1/RegFile1/Storage[20][24] ,
         \FIFO_U1/RegFile1/Storage[20][25] ,
         \FIFO_U1/RegFile1/Storage[20][26] ,
         \FIFO_U1/RegFile1/Storage[20][27] ,
         \FIFO_U1/RegFile1/Storage[20][28] ,
         \FIFO_U1/RegFile1/Storage[20][29] ,
         \FIFO_U1/RegFile1/Storage[20][30] ,
         \FIFO_U1/RegFile1/Storage[20][31] , \FIFO_U1/RegFile1/Storage[21][0] ,
         \FIFO_U1/RegFile1/Storage[21][1] , \FIFO_U1/RegFile1/Storage[21][2] ,
         \FIFO_U1/RegFile1/Storage[21][3] , \FIFO_U1/RegFile1/Storage[21][4] ,
         \FIFO_U1/RegFile1/Storage[21][5] , \FIFO_U1/RegFile1/Storage[21][6] ,
         \FIFO_U1/RegFile1/Storage[21][7] , \FIFO_U1/RegFile1/Storage[21][8] ,
         \FIFO_U1/RegFile1/Storage[21][9] , \FIFO_U1/RegFile1/Storage[21][10] ,
         \FIFO_U1/RegFile1/Storage[21][11] ,
         \FIFO_U1/RegFile1/Storage[21][12] ,
         \FIFO_U1/RegFile1/Storage[21][13] ,
         \FIFO_U1/RegFile1/Storage[21][14] ,
         \FIFO_U1/RegFile1/Storage[21][15] ,
         \FIFO_U1/RegFile1/Storage[21][16] ,
         \FIFO_U1/RegFile1/Storage[21][17] ,
         \FIFO_U1/RegFile1/Storage[21][18] ,
         \FIFO_U1/RegFile1/Storage[21][19] ,
         \FIFO_U1/RegFile1/Storage[21][20] ,
         \FIFO_U1/RegFile1/Storage[21][21] ,
         \FIFO_U1/RegFile1/Storage[21][22] ,
         \FIFO_U1/RegFile1/Storage[21][23] ,
         \FIFO_U1/RegFile1/Storage[21][24] ,
         \FIFO_U1/RegFile1/Storage[21][25] ,
         \FIFO_U1/RegFile1/Storage[21][26] ,
         \FIFO_U1/RegFile1/Storage[21][27] ,
         \FIFO_U1/RegFile1/Storage[21][28] ,
         \FIFO_U1/RegFile1/Storage[21][29] ,
         \FIFO_U1/RegFile1/Storage[21][30] ,
         \FIFO_U1/RegFile1/Storage[21][31] , \FIFO_U1/RegFile1/Storage[22][0] ,
         \FIFO_U1/RegFile1/Storage[22][1] , \FIFO_U1/RegFile1/Storage[22][2] ,
         \FIFO_U1/RegFile1/Storage[22][3] , \FIFO_U1/RegFile1/Storage[22][4] ,
         \FIFO_U1/RegFile1/Storage[22][5] , \FIFO_U1/RegFile1/Storage[22][6] ,
         \FIFO_U1/RegFile1/Storage[22][7] , \FIFO_U1/RegFile1/Storage[22][8] ,
         \FIFO_U1/RegFile1/Storage[22][9] , \FIFO_U1/RegFile1/Storage[22][10] ,
         \FIFO_U1/RegFile1/Storage[22][11] ,
         \FIFO_U1/RegFile1/Storage[22][12] ,
         \FIFO_U1/RegFile1/Storage[22][13] ,
         \FIFO_U1/RegFile1/Storage[22][14] ,
         \FIFO_U1/RegFile1/Storage[22][15] ,
         \FIFO_U1/RegFile1/Storage[22][16] ,
         \FIFO_U1/RegFile1/Storage[22][17] ,
         \FIFO_U1/RegFile1/Storage[22][18] ,
         \FIFO_U1/RegFile1/Storage[22][19] ,
         \FIFO_U1/RegFile1/Storage[22][20] ,
         \FIFO_U1/RegFile1/Storage[22][21] ,
         \FIFO_U1/RegFile1/Storage[22][22] ,
         \FIFO_U1/RegFile1/Storage[22][23] ,
         \FIFO_U1/RegFile1/Storage[22][24] ,
         \FIFO_U1/RegFile1/Storage[22][25] ,
         \FIFO_U1/RegFile1/Storage[22][26] ,
         \FIFO_U1/RegFile1/Storage[22][27] ,
         \FIFO_U1/RegFile1/Storage[22][28] ,
         \FIFO_U1/RegFile1/Storage[22][29] ,
         \FIFO_U1/RegFile1/Storage[22][30] ,
         \FIFO_U1/RegFile1/Storage[22][31] , \FIFO_U1/RegFile1/Storage[23][0] ,
         \FIFO_U1/RegFile1/Storage[23][1] , \FIFO_U1/RegFile1/Storage[23][2] ,
         \FIFO_U1/RegFile1/Storage[23][3] , \FIFO_U1/RegFile1/Storage[23][4] ,
         \FIFO_U1/RegFile1/Storage[23][5] , \FIFO_U1/RegFile1/Storage[23][6] ,
         \FIFO_U1/RegFile1/Storage[23][7] , \FIFO_U1/RegFile1/Storage[23][8] ,
         \FIFO_U1/RegFile1/Storage[23][9] , \FIFO_U1/RegFile1/Storage[23][10] ,
         \FIFO_U1/RegFile1/Storage[23][11] ,
         \FIFO_U1/RegFile1/Storage[23][12] ,
         \FIFO_U1/RegFile1/Storage[23][13] ,
         \FIFO_U1/RegFile1/Storage[23][14] ,
         \FIFO_U1/RegFile1/Storage[23][15] ,
         \FIFO_U1/RegFile1/Storage[23][16] ,
         \FIFO_U1/RegFile1/Storage[23][17] ,
         \FIFO_U1/RegFile1/Storage[23][18] ,
         \FIFO_U1/RegFile1/Storage[23][19] ,
         \FIFO_U1/RegFile1/Storage[23][20] ,
         \FIFO_U1/RegFile1/Storage[23][21] ,
         \FIFO_U1/RegFile1/Storage[23][22] ,
         \FIFO_U1/RegFile1/Storage[23][23] ,
         \FIFO_U1/RegFile1/Storage[23][24] ,
         \FIFO_U1/RegFile1/Storage[23][25] ,
         \FIFO_U1/RegFile1/Storage[23][26] ,
         \FIFO_U1/RegFile1/Storage[23][27] ,
         \FIFO_U1/RegFile1/Storage[23][28] ,
         \FIFO_U1/RegFile1/Storage[23][29] ,
         \FIFO_U1/RegFile1/Storage[23][30] ,
         \FIFO_U1/RegFile1/Storage[23][31] , \FIFO_U1/RegFile1/Storage[24][0] ,
         \FIFO_U1/RegFile1/Storage[24][1] , \FIFO_U1/RegFile1/Storage[24][2] ,
         \FIFO_U1/RegFile1/Storage[24][3] , \FIFO_U1/RegFile1/Storage[24][4] ,
         \FIFO_U1/RegFile1/Storage[24][5] , \FIFO_U1/RegFile1/Storage[24][6] ,
         \FIFO_U1/RegFile1/Storage[24][7] , \FIFO_U1/RegFile1/Storage[24][8] ,
         \FIFO_U1/RegFile1/Storage[24][9] , \FIFO_U1/RegFile1/Storage[24][10] ,
         \FIFO_U1/RegFile1/Storage[24][11] ,
         \FIFO_U1/RegFile1/Storage[24][12] ,
         \FIFO_U1/RegFile1/Storage[24][13] ,
         \FIFO_U1/RegFile1/Storage[24][14] ,
         \FIFO_U1/RegFile1/Storage[24][15] ,
         \FIFO_U1/RegFile1/Storage[24][16] ,
         \FIFO_U1/RegFile1/Storage[24][17] ,
         \FIFO_U1/RegFile1/Storage[24][18] ,
         \FIFO_U1/RegFile1/Storage[24][19] ,
         \FIFO_U1/RegFile1/Storage[24][20] ,
         \FIFO_U1/RegFile1/Storage[24][21] ,
         \FIFO_U1/RegFile1/Storage[24][22] ,
         \FIFO_U1/RegFile1/Storage[24][23] ,
         \FIFO_U1/RegFile1/Storage[24][24] ,
         \FIFO_U1/RegFile1/Storage[24][25] ,
         \FIFO_U1/RegFile1/Storage[24][26] ,
         \FIFO_U1/RegFile1/Storage[24][27] ,
         \FIFO_U1/RegFile1/Storage[24][28] ,
         \FIFO_U1/RegFile1/Storage[24][29] ,
         \FIFO_U1/RegFile1/Storage[24][30] ,
         \FIFO_U1/RegFile1/Storage[24][31] , \FIFO_U1/RegFile1/Storage[25][0] ,
         \FIFO_U1/RegFile1/Storage[25][1] , \FIFO_U1/RegFile1/Storage[25][2] ,
         \FIFO_U1/RegFile1/Storage[25][3] , \FIFO_U1/RegFile1/Storage[25][4] ,
         \FIFO_U1/RegFile1/Storage[25][5] , \FIFO_U1/RegFile1/Storage[25][6] ,
         \FIFO_U1/RegFile1/Storage[25][7] , \FIFO_U1/RegFile1/Storage[25][8] ,
         \FIFO_U1/RegFile1/Storage[25][9] , \FIFO_U1/RegFile1/Storage[25][10] ,
         \FIFO_U1/RegFile1/Storage[25][11] ,
         \FIFO_U1/RegFile1/Storage[25][12] ,
         \FIFO_U1/RegFile1/Storage[25][13] ,
         \FIFO_U1/RegFile1/Storage[25][14] ,
         \FIFO_U1/RegFile1/Storage[25][15] ,
         \FIFO_U1/RegFile1/Storage[25][16] ,
         \FIFO_U1/RegFile1/Storage[25][17] ,
         \FIFO_U1/RegFile1/Storage[25][18] ,
         \FIFO_U1/RegFile1/Storage[25][19] ,
         \FIFO_U1/RegFile1/Storage[25][20] ,
         \FIFO_U1/RegFile1/Storage[25][21] ,
         \FIFO_U1/RegFile1/Storage[25][22] ,
         \FIFO_U1/RegFile1/Storage[25][23] ,
         \FIFO_U1/RegFile1/Storage[25][24] ,
         \FIFO_U1/RegFile1/Storage[25][25] ,
         \FIFO_U1/RegFile1/Storage[25][26] ,
         \FIFO_U1/RegFile1/Storage[25][27] ,
         \FIFO_U1/RegFile1/Storage[25][28] ,
         \FIFO_U1/RegFile1/Storage[25][29] ,
         \FIFO_U1/RegFile1/Storage[25][30] ,
         \FIFO_U1/RegFile1/Storage[25][31] , \FIFO_U1/RegFile1/Storage[26][0] ,
         \FIFO_U1/RegFile1/Storage[26][1] , \FIFO_U1/RegFile1/Storage[26][2] ,
         \FIFO_U1/RegFile1/Storage[26][3] , \FIFO_U1/RegFile1/Storage[26][4] ,
         \FIFO_U1/RegFile1/Storage[26][5] , \FIFO_U1/RegFile1/Storage[26][6] ,
         \FIFO_U1/RegFile1/Storage[26][7] , \FIFO_U1/RegFile1/Storage[26][8] ,
         \FIFO_U1/RegFile1/Storage[26][9] , \FIFO_U1/RegFile1/Storage[26][10] ,
         \FIFO_U1/RegFile1/Storage[26][11] ,
         \FIFO_U1/RegFile1/Storage[26][12] ,
         \FIFO_U1/RegFile1/Storage[26][13] ,
         \FIFO_U1/RegFile1/Storage[26][14] ,
         \FIFO_U1/RegFile1/Storage[26][15] ,
         \FIFO_U1/RegFile1/Storage[26][16] ,
         \FIFO_U1/RegFile1/Storage[26][17] ,
         \FIFO_U1/RegFile1/Storage[26][18] ,
         \FIFO_U1/RegFile1/Storage[26][19] ,
         \FIFO_U1/RegFile1/Storage[26][20] ,
         \FIFO_U1/RegFile1/Storage[26][21] ,
         \FIFO_U1/RegFile1/Storage[26][22] ,
         \FIFO_U1/RegFile1/Storage[26][23] ,
         \FIFO_U1/RegFile1/Storage[26][24] ,
         \FIFO_U1/RegFile1/Storage[26][25] ,
         \FIFO_U1/RegFile1/Storage[26][26] ,
         \FIFO_U1/RegFile1/Storage[26][27] ,
         \FIFO_U1/RegFile1/Storage[26][28] ,
         \FIFO_U1/RegFile1/Storage[26][29] ,
         \FIFO_U1/RegFile1/Storage[26][30] ,
         \FIFO_U1/RegFile1/Storage[26][31] , \FIFO_U1/RegFile1/Storage[27][0] ,
         \FIFO_U1/RegFile1/Storage[27][1] , \FIFO_U1/RegFile1/Storage[27][2] ,
         \FIFO_U1/RegFile1/Storage[27][3] , \FIFO_U1/RegFile1/Storage[27][4] ,
         \FIFO_U1/RegFile1/Storage[27][5] , \FIFO_U1/RegFile1/Storage[27][6] ,
         \FIFO_U1/RegFile1/Storage[27][7] , \FIFO_U1/RegFile1/Storage[27][8] ,
         \FIFO_U1/RegFile1/Storage[27][9] , \FIFO_U1/RegFile1/Storage[27][10] ,
         \FIFO_U1/RegFile1/Storage[27][11] ,
         \FIFO_U1/RegFile1/Storage[27][12] ,
         \FIFO_U1/RegFile1/Storage[27][13] ,
         \FIFO_U1/RegFile1/Storage[27][14] ,
         \FIFO_U1/RegFile1/Storage[27][15] ,
         \FIFO_U1/RegFile1/Storage[27][16] ,
         \FIFO_U1/RegFile1/Storage[27][17] ,
         \FIFO_U1/RegFile1/Storage[27][18] ,
         \FIFO_U1/RegFile1/Storage[27][19] ,
         \FIFO_U1/RegFile1/Storage[27][20] ,
         \FIFO_U1/RegFile1/Storage[27][21] ,
         \FIFO_U1/RegFile1/Storage[27][22] ,
         \FIFO_U1/RegFile1/Storage[27][23] ,
         \FIFO_U1/RegFile1/Storage[27][24] ,
         \FIFO_U1/RegFile1/Storage[27][25] ,
         \FIFO_U1/RegFile1/Storage[27][26] ,
         \FIFO_U1/RegFile1/Storage[27][27] ,
         \FIFO_U1/RegFile1/Storage[27][28] ,
         \FIFO_U1/RegFile1/Storage[27][29] ,
         \FIFO_U1/RegFile1/Storage[27][30] ,
         \FIFO_U1/RegFile1/Storage[27][31] , \FIFO_U1/RegFile1/Storage[28][0] ,
         \FIFO_U1/RegFile1/Storage[28][1] , \FIFO_U1/RegFile1/Storage[28][2] ,
         \FIFO_U1/RegFile1/Storage[28][3] , \FIFO_U1/RegFile1/Storage[28][4] ,
         \FIFO_U1/RegFile1/Storage[28][5] , \FIFO_U1/RegFile1/Storage[28][6] ,
         \FIFO_U1/RegFile1/Storage[28][7] , \FIFO_U1/RegFile1/Storage[28][8] ,
         \FIFO_U1/RegFile1/Storage[28][9] , \FIFO_U1/RegFile1/Storage[28][10] ,
         \FIFO_U1/RegFile1/Storage[28][11] ,
         \FIFO_U1/RegFile1/Storage[28][12] ,
         \FIFO_U1/RegFile1/Storage[28][13] ,
         \FIFO_U1/RegFile1/Storage[28][14] ,
         \FIFO_U1/RegFile1/Storage[28][15] ,
         \FIFO_U1/RegFile1/Storage[28][16] ,
         \FIFO_U1/RegFile1/Storage[28][17] ,
         \FIFO_U1/RegFile1/Storage[28][18] ,
         \FIFO_U1/RegFile1/Storage[28][19] ,
         \FIFO_U1/RegFile1/Storage[28][20] ,
         \FIFO_U1/RegFile1/Storage[28][21] ,
         \FIFO_U1/RegFile1/Storage[28][22] ,
         \FIFO_U1/RegFile1/Storage[28][23] ,
         \FIFO_U1/RegFile1/Storage[28][24] ,
         \FIFO_U1/RegFile1/Storage[28][25] ,
         \FIFO_U1/RegFile1/Storage[28][26] ,
         \FIFO_U1/RegFile1/Storage[28][27] ,
         \FIFO_U1/RegFile1/Storage[28][28] ,
         \FIFO_U1/RegFile1/Storage[28][29] ,
         \FIFO_U1/RegFile1/Storage[28][30] ,
         \FIFO_U1/RegFile1/Storage[28][31] , \FIFO_U1/RegFile1/Storage[29][0] ,
         \FIFO_U1/RegFile1/Storage[29][1] , \FIFO_U1/RegFile1/Storage[29][2] ,
         \FIFO_U1/RegFile1/Storage[29][3] , \FIFO_U1/RegFile1/Storage[29][4] ,
         \FIFO_U1/RegFile1/Storage[29][5] , \FIFO_U1/RegFile1/Storage[29][6] ,
         \FIFO_U1/RegFile1/Storage[29][7] , \FIFO_U1/RegFile1/Storage[29][8] ,
         \FIFO_U1/RegFile1/Storage[29][9] , \FIFO_U1/RegFile1/Storage[29][10] ,
         \FIFO_U1/RegFile1/Storage[29][11] ,
         \FIFO_U1/RegFile1/Storage[29][12] ,
         \FIFO_U1/RegFile1/Storage[29][13] ,
         \FIFO_U1/RegFile1/Storage[29][14] ,
         \FIFO_U1/RegFile1/Storage[29][15] ,
         \FIFO_U1/RegFile1/Storage[29][16] ,
         \FIFO_U1/RegFile1/Storage[29][17] ,
         \FIFO_U1/RegFile1/Storage[29][18] ,
         \FIFO_U1/RegFile1/Storage[29][19] ,
         \FIFO_U1/RegFile1/Storage[29][20] ,
         \FIFO_U1/RegFile1/Storage[29][21] ,
         \FIFO_U1/RegFile1/Storage[29][22] ,
         \FIFO_U1/RegFile1/Storage[29][23] ,
         \FIFO_U1/RegFile1/Storage[29][24] ,
         \FIFO_U1/RegFile1/Storage[29][25] ,
         \FIFO_U1/RegFile1/Storage[29][26] ,
         \FIFO_U1/RegFile1/Storage[29][27] ,
         \FIFO_U1/RegFile1/Storage[29][28] ,
         \FIFO_U1/RegFile1/Storage[29][29] ,
         \FIFO_U1/RegFile1/Storage[29][30] ,
         \FIFO_U1/RegFile1/Storage[29][31] , \FIFO_U1/RegFile1/Storage[30][0] ,
         \FIFO_U1/RegFile1/Storage[30][1] , \FIFO_U1/RegFile1/Storage[30][2] ,
         \FIFO_U1/RegFile1/Storage[30][3] , \FIFO_U1/RegFile1/Storage[30][4] ,
         \FIFO_U1/RegFile1/Storage[30][5] , \FIFO_U1/RegFile1/Storage[30][6] ,
         \FIFO_U1/RegFile1/Storage[30][7] , \FIFO_U1/RegFile1/Storage[30][8] ,
         \FIFO_U1/RegFile1/Storage[30][9] , \FIFO_U1/RegFile1/Storage[30][10] ,
         \FIFO_U1/RegFile1/Storage[30][11] ,
         \FIFO_U1/RegFile1/Storage[30][12] ,
         \FIFO_U1/RegFile1/Storage[30][13] ,
         \FIFO_U1/RegFile1/Storage[30][14] ,
         \FIFO_U1/RegFile1/Storage[30][15] ,
         \FIFO_U1/RegFile1/Storage[30][16] ,
         \FIFO_U1/RegFile1/Storage[30][17] ,
         \FIFO_U1/RegFile1/Storage[30][18] ,
         \FIFO_U1/RegFile1/Storage[30][19] ,
         \FIFO_U1/RegFile1/Storage[30][20] ,
         \FIFO_U1/RegFile1/Storage[30][21] ,
         \FIFO_U1/RegFile1/Storage[30][22] ,
         \FIFO_U1/RegFile1/Storage[30][23] ,
         \FIFO_U1/RegFile1/Storage[30][24] ,
         \FIFO_U1/RegFile1/Storage[30][25] ,
         \FIFO_U1/RegFile1/Storage[30][26] ,
         \FIFO_U1/RegFile1/Storage[30][27] ,
         \FIFO_U1/RegFile1/Storage[30][28] ,
         \FIFO_U1/RegFile1/Storage[30][29] ,
         \FIFO_U1/RegFile1/Storage[30][30] ,
         \FIFO_U1/RegFile1/Storage[30][31] , \FIFO_U1/RegFile1/Storage[31][0] ,
         \FIFO_U1/RegFile1/Storage[31][1] , \FIFO_U1/RegFile1/Storage[31][2] ,
         \FIFO_U1/RegFile1/Storage[31][3] , \FIFO_U1/RegFile1/Storage[31][4] ,
         \FIFO_U1/RegFile1/Storage[31][5] , \FIFO_U1/RegFile1/Storage[31][6] ,
         \FIFO_U1/RegFile1/Storage[31][7] , \FIFO_U1/RegFile1/Storage[31][8] ,
         \FIFO_U1/RegFile1/Storage[31][9] , \FIFO_U1/RegFile1/Storage[31][10] ,
         \FIFO_U1/RegFile1/Storage[31][11] ,
         \FIFO_U1/RegFile1/Storage[31][12] ,
         \FIFO_U1/RegFile1/Storage[31][13] ,
         \FIFO_U1/RegFile1/Storage[31][14] ,
         \FIFO_U1/RegFile1/Storage[31][15] ,
         \FIFO_U1/RegFile1/Storage[31][16] ,
         \FIFO_U1/RegFile1/Storage[31][17] ,
         \FIFO_U1/RegFile1/Storage[31][18] ,
         \FIFO_U1/RegFile1/Storage[31][19] ,
         \FIFO_U1/RegFile1/Storage[31][20] ,
         \FIFO_U1/RegFile1/Storage[31][21] ,
         \FIFO_U1/RegFile1/Storage[31][22] ,
         \FIFO_U1/RegFile1/Storage[31][23] ,
         \FIFO_U1/RegFile1/Storage[31][24] ,
         \FIFO_U1/RegFile1/Storage[31][25] ,
         \FIFO_U1/RegFile1/Storage[31][26] ,
         \FIFO_U1/RegFile1/Storage[31][27] ,
         \FIFO_U1/RegFile1/Storage[31][28] ,
         \FIFO_U1/RegFile1/Storage[31][29] ,
         \FIFO_U1/RegFile1/Storage[31][30] ,
         \FIFO_U1/RegFile1/Storage[31][31] , \FIFO_U1/RegFile1/ChipClock ,
         \FIFO_U1/RegFile1/N79 , \FIFO_U1/RegFile1/N78 ,
         \FIFO_U1/RegFile1/N76 , \FIFO_U1/RegFile1/N75 ,
         \FIFO_U1/RegFile1/N63 , \FIFO_U1/RegFile1/N62 ,
         \FIFO_U1/RegFile1/N61 , \FIFO_U1/RegFile1/N60 ,
         \FIFO_U1/RegFile1/N59 , \FIFO_U1/RegFile1/N58 ,
         \FIFO_U1/RegFile1/N57 , \FIFO_U1/RegFile1/N56 ,
         \FIFO_U1/RegFile1/N55 , \FIFO_U1/RegFile1/N54 ,
         \FIFO_U1/RegFile1/N53 , \FIFO_U1/RegFile1/N52 ,
         \FIFO_U1/RegFile1/N51 , \FIFO_U1/RegFile1/N50 ,
         \FIFO_U1/RegFile1/N49 , \FIFO_U1/RegFile1/N48 ,
         \FIFO_U1/RegFile1/N47 , \FIFO_U1/RegFile1/N46 ,
         \FIFO_U1/RegFile1/N45 , \FIFO_U1/RegFile1/N44 ,
         \FIFO_U1/RegFile1/N43 , \FIFO_U1/RegFile1/N42 ,
         \FIFO_U1/RegFile1/N41 , \FIFO_U1/RegFile1/N40 ,
         \FIFO_U1/RegFile1/N39 , \FIFO_U1/RegFile1/N38 ,
         \FIFO_U1/RegFile1/N37 , \FIFO_U1/RegFile1/N36 ,
         \FIFO_U1/RegFile1/N35 , \FIFO_U1/RegFile1/N34 ,
         \FIFO_U1/RegFile1/N33 , \FIFO_U1/RegFile1/N32 , \DesDecoder_U1/N70 ,
         \DesDecoder_U1/N69 , \DesDecoder_U1/N68 , \DesDecoder_U1/N67 ,
         \DesDecoder_U1/N66 , \DesDecoder_U1/N65 , \DesDecoder_U1/N63 ,
         \DesDecoder_U1/N62 , \DesDecoder_U1/N53 , \DesDecoder_U1/N52 ,
         \DesDecoder_U1/N51 , \DesDecoder_U1/N50 , \DesDecoder_U1/N49 ,
         \DesDecoder_U1/N44 , \DesDecoder_U1/N12 , \DesDecoder_U1/FrameSR[0] ,
         \DesDecoder_U1/FrameSR[1] , \DesDecoder_U1/FrameSR[2] ,
         \DesDecoder_U1/FrameSR[3] , \DesDecoder_U1/FrameSR[4] ,
         \DesDecoder_U1/FrameSR[5] , \DesDecoder_U1/FrameSR[6] ,
         \DesDecoder_U1/FrameSR[7] , \DesDecoder_U1/FrameSR[8] ,
         \DesDecoder_U1/FrameSR[9] , \DesDecoder_U1/FrameSR[10] ,
         \DesDecoder_U1/FrameSR[11] , \DesDecoder_U1/FrameSR[12] ,
         \DesDecoder_U1/FrameSR[13] , \DesDecoder_U1/FrameSR[14] ,
         \DesDecoder_U1/FrameSR[15] , \DesDecoder_U1/FrameSR[16] ,
         \DesDecoder_U1/FrameSR[17] , \DesDecoder_U1/FrameSR[18] ,
         \DesDecoder_U1/FrameSR[19] , \DesDecoder_U1/FrameSR[20] ,
         \DesDecoder_U1/FrameSR[21] , \DesDecoder_U1/FrameSR[22] ,
         \DesDecoder_U1/FrameSR[23] , \DesDecoder_U1/FrameSR[24] ,
         \DesDecoder_U1/FrameSR[25] , \DesDecoder_U1/FrameSR[26] ,
         \DesDecoder_U1/FrameSR[27] , \DesDecoder_U1/FrameSR[28] ,
         \DesDecoder_U1/FrameSR[29] , \DesDecoder_U1/FrameSR[30] ,
         \DesDecoder_U1/FrameSR[31] , \DesDecoder_U1/FrameSR[32] ,
         \DesDecoder_U1/FrameSR[33] , \DesDecoder_U1/FrameSR[34] ,
         \DesDecoder_U1/FrameSR[35] , \DesDecoder_U1/FrameSR[36] ,
         \DesDecoder_U1/FrameSR[37] , \DesDecoder_U1/FrameSR[38] ,
         \DesDecoder_U1/FrameSR[39] , \DesDecoder_U1/FrameSR[40] ,
         \DesDecoder_U1/FrameSR[41] , \DesDecoder_U1/FrameSR[42] ,
         \DesDecoder_U1/FrameSR[43] , \DesDecoder_U1/FrameSR[44] ,
         \DesDecoder_U1/FrameSR[45] , \DesDecoder_U1/FrameSR[46] ,
         \DesDecoder_U1/FrameSR[47] , \DesDecoder_U1/FrameSR[48] ,
         \DesDecoder_U1/FrameSR[49] , \DesDecoder_U1/FrameSR[50] ,
         \DesDecoder_U1/FrameSR[51] , \DesDecoder_U1/FrameSR[52] ,
         \DesDecoder_U1/FrameSR[53] , \DesDecoder_U1/FrameSR[54] ,
         \DesDecoder_U1/FrameSR[55] , \DesDecoder_U1/FrameSR[56] ,
         \DesDecoder_U1/FrameSR[57] , \DesDecoder_U1/FrameSR[58] ,
         \DesDecoder_U1/FrameSR[59] , \DesDecoder_U1/FrameSR[60] ,
         \DesDecoder_U1/FrameSR[61] , \DesDecoder_U1/FrameSR[62] ,
         \SerialRx_U1/PLL_RxU1/CtrCarry , \SerialRx_U1/PLL_RxU1/SampleWire ,
         \SerialRx_U1/PLL_RxU1/Comp1/N20 , \SerialRx_U1/PLL_RxU1/Comp1/N19 ,
         \SerialRx_U1/PLL_RxU1/Comp1/N9 , \SerialRx_U1/PLL_RxU1/Comp1/N8 ,
         \SerialRx_U1/PLL_RxU1/Comp1/N7 , \SerialRx_U1/PLL_RxU1/Comp1/N6 ,
         \SerialRx_U1/PLL_RxU1/Comp1/N5 ,
         \SerialRx_U1/PLL_RxU1/Comp1/ClockInN[0] ,
         \SerialRx_U1/PLL_RxU1/Comp1/ClockInN[1] ,
         \SerialRx_U1/PLL_RxU1/VFO1/N55 , \SerialRx_U1/PLL_RxU1/VFO1/N54 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N53 , \SerialRx_U1/PLL_RxU1/VFO1/N51 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N49 , \SerialRx_U1/PLL_RxU1/VFO1/N47 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N45 , \SerialRx_U1/PLL_RxU1/VFO1/N21 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N20 , \SerialRx_U1/PLL_RxU1/VFO1/N19 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N18 , \SerialRx_U1/PLL_RxU1/VFO1/N17 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N16 , \SerialRx_U1/PLL_RxU1/VFO1/N14 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N13 , \SerialRx_U1/PLL_RxU1/VFO1/N12 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N11 , \SerialRx_U1/PLL_RxU1/VFO1/N10 ,
         \SerialRx_U1/PLL_RxU1/VFO1/N9 ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[0] ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[2] ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[4] ,
         \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[5] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[0] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[1] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[2] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[3] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[4] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[5] ,
         \SerialRx_U1/PLL_RxU1/VFO1/FastClock ,
         \SerialRx_U1/PLL_RxU1/MCntr1/N5 , \SerialRx_U1/PLL_RxU1/MCntr1/N4 ,
         \SerialRx_U1/PLL_RxU1/MCntr1/N3 , \SerialRx_U1/PLL_RxU1/MCntr1/N2 ,
         \SerialRx_U1/PLL_RxU1/MCntr1/N1 , \U3/U1/Z_0 , \U3/U1/Z_1 ,
         \U3/U1/Z_2 , \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U2/Z_0 ,
         \FIFO_U1/RegFile1/DataOreg[9] , \FIFO_U1/RegFile1/DataOreg[8] ,
         \FIFO_U1/RegFile1/DataOreg[7] , \FIFO_U1/RegFile1/DataOreg[6] ,
         \FIFO_U1/RegFile1/DataOreg[5] , \FIFO_U1/RegFile1/DataOreg[4] ,
         \FIFO_U1/RegFile1/DataOreg[3] , \FIFO_U1/RegFile1/DataOreg[31] ,
         \FIFO_U1/RegFile1/DataOreg[30] , \FIFO_U1/RegFile1/DataOreg[2] ,
         \FIFO_U1/RegFile1/DataOreg[29] , \FIFO_U1/RegFile1/DataOreg[28] ,
         \FIFO_U1/RegFile1/DataOreg[27] , \FIFO_U1/RegFile1/DataOreg[26] ,
         \FIFO_U1/RegFile1/DataOreg[25] , \FIFO_U1/RegFile1/DataOreg[24] ,
         \FIFO_U1/RegFile1/DataOreg[23] , \FIFO_U1/RegFile1/DataOreg[22] ,
         \FIFO_U1/RegFile1/DataOreg[21] , \FIFO_U1/RegFile1/DataOreg[20] ,
         \FIFO_U1/RegFile1/DataOreg[1] , \FIFO_U1/RegFile1/DataOreg[19] ,
         \FIFO_U1/RegFile1/DataOreg[18] , \FIFO_U1/RegFile1/DataOreg[17] ,
         \FIFO_U1/RegFile1/DataOreg[16] , \FIFO_U1/RegFile1/DataOreg[15] ,
         \FIFO_U1/RegFile1/DataOreg[14] , \FIFO_U1/RegFile1/DataOreg[13] ,
         \FIFO_U1/RegFile1/DataOreg[12] , \FIFO_U1/RegFile1/DataOreg[11] ,
         \FIFO_U1/RegFile1/DataOreg[10] , \FIFO_U1/RegFile1/DataOreg[0] , n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n281, n283,
         n285, n287, n289, n291, n293, n295, n297, n299, n301, n303, n305,
         n307, n309, n311, n313, n315, n317, n319, n321, n323, n325, n327,
         n329, n331, n333, n335, n337, n339, n341, n356, n360, n361, n368,
         n374, n375, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n564, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;
  wire   [4:0] \FIFO_U1/SM_WriteAddr ;
  wire   [4:0] \FIFO_U1/SM_ReadAddr ;
  wire   [2:0] \FIFO_U1/FIFO_SM1/NextState ;
  wire   [4:0] \DesDecoder_U1/Count32 ;
  wire   [1:0] \SerialRx_U1/PLL_RxU1/AdjFreq ;
  wire   [5:0] \SerialRx_U1/PLL_RxU1/VFO1/WireD ;
  wire   [3:0] \SerialRx_U1/PLL_RxU1/MCntr1/Ctr ;
  assign SerRxToDecode = SerialIn;

  DEL005 \SerialRx_U1/PLL_RxU1/SampleDelay1  ( .I(DecoderParClk), .Z(
        \SerialRx_U1/PLL_RxU1/SampleWire ) );
  DEL005 \SerialRx_U1/PLL_RxU1/VFO1/DelayLine[4].Delay83ps  ( .I(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [4]), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [5]) );
  DEL005 \SerialRx_U1/PLL_RxU1/VFO1/DelayLine[3].Delay83ps  ( .I(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [3]), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [4]) );
  DEL005 \SerialRx_U1/PLL_RxU1/VFO1/DelayLine[2].Delay83ps  ( .I(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [2]), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [3]) );
  DEL005 \SerialRx_U1/PLL_RxU1/VFO1/DelayLine[1].Delay83ps  ( .I(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [1]), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [2]) );
  DEL005 \SerialRx_U1/PLL_RxU1/VFO1/DelayLine[0].Delay83ps  ( .I(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [0]), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [1]) );
  CKND1 \SerialRx_U1/PLL_RxU1/VFO1/I_2  ( .CLK(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CN(
        \SerialRx_U1/PLL_RxU1/VFO1/WireD [0]) );
  LHQD1 \DesDecoder_U1/Count32_reg[0]  ( .E(\DesDecoder_U1/N69 ), .D(
        \DesDecoder_U1/N65 ), .Q(\DesDecoder_U1/Count32 [0]) );
  LHQD1 \DesDecoder_U1/Count32_reg[1]  ( .E(\DesDecoder_U1/N69 ), .D(
        \DesDecoder_U1/N66 ), .Q(\DesDecoder_U1/Count32 [1]) );
  LHQD1 \DesDecoder_U1/Count32_reg[2]  ( .E(\DesDecoder_U1/N69 ), .D(
        \DesDecoder_U1/N67 ), .Q(\DesDecoder_U1/Count32 [2]) );
  LHQD1 \DesDecoder_U1/Count32_reg[3]  ( .E(\DesDecoder_U1/N69 ), .D(
        \DesDecoder_U1/N68 ), .Q(\DesDecoder_U1/Count32 [3]) );
  LHQD1 \DesDecoder_U1/Count32_reg[4]  ( .E(\DesDecoder_U1/N69 ), .D(
        \DesDecoder_U1/N70 ), .Q(\DesDecoder_U1/Count32 [4]) );
  LHQD1 \DesDecoder_U1/ParClkReg_reg  ( .E(\DesDecoder_U1/N62 ), .D(
        \DesDecoder_U1/N63 ), .Q(DecoderParClk) );
  DFNCND2 \DesDecoder_U1/UnLoad_reg  ( .D(\DesDecoder_U1/N44 ), .CPN(n637), 
        .CDN(n594), .Q(n1242) );
  LHQD1 \FIFO_U1/FIFO_SM1/NextState_reg[0]  ( .E(\FIFO_U1/FIFO_SM1/N188 ), .D(
        \FIFO_U1/FIFO_SM1/N142 ), .Q(\FIFO_U1/FIFO_SM1/NextState [0]) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_reg[0]  ( .E(\FIFO_U1/FIFO_SM1/N198 ), 
        .D(\FIFO_U1/FIFO_SM1/N150 ), .Q(\FIFO_U1/FIFO_SM1/N239 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_reg[0]  ( .E(\FIFO_U1/FIFO_SM1/N209 ), .D(
        \FIFO_U1/FIFO_SM1/N167 ), .Q(\FIFO_U1/FIFO_SM1/N224 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_reg[4]  ( .E(\FIFO_U1/FIFO_SM1/N198 ), 
        .D(\FIFO_U1/FIFO_SM1/N162 ), .Q(\FIFO_U1/FIFO_SM1/N227 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_reg[4]  ( .E(\FIFO_U1/FIFO_SM1/N209 ), .D(
        \FIFO_U1/FIFO_SM1/N179 ), .Q(\FIFO_U1/FIFO_SM1/N212 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/NextState_reg[1]  ( .E(\FIFO_U1/FIFO_SM1/N188 ), .D(
        \FIFO_U1/FIFO_SM1/N144 ), .Q(\FIFO_U1/FIFO_SM1/NextState [1]) );
  LHQD1 \FIFO_U1/FIFO_SM1/NextState_reg[2]  ( .E(\FIFO_U1/FIFO_SM1/N188 ), .D(
        \FIFO_U1/FIFO_SM1/N146 ), .Q(\FIFO_U1/FIFO_SM1/NextState [2]) );
  LHQD1 \FIFO_U1/FIFO_SM1/EmptyFIFOReg_reg  ( .E(\FIFO_U1/FIFO_SM1/N211 ), .D(
        \FIFO_U1/FIFO_SM1/N182 ), .Q(FIFOEmpty) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_tri_enable_reg[4]  ( .E(
        \FIFO_U1/FIFO_SM1/N209 ), .D(\FIFO_U1/FIFO_SM1/N210 ), .Q(
        \FIFO_U1/FIFO_SM1/N0 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_tri_enable_reg[2]  ( .E(
        \FIFO_U1/FIFO_SM1/N209 ), .D(\FIFO_U1/FIFO_SM1/N210 ), .Q(
        \FIFO_U1/FIFO_SM1/N2 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_tri_enable_reg[0]  ( .E(
        \FIFO_U1/FIFO_SM1/N209 ), .D(\FIFO_U1/FIFO_SM1/N210 ), .Q(
        \FIFO_U1/FIFO_SM1/N4 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_tri_enable_reg[1]  ( .E(
        \FIFO_U1/FIFO_SM1/N209 ), .D(\FIFO_U1/FIFO_SM1/N210 ), .Q(
        \FIFO_U1/FIFO_SM1/N3 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_tri_enable_reg[3]  ( .E(
        \FIFO_U1/FIFO_SM1/N209 ), .D(\FIFO_U1/FIFO_SM1/N210 ), .Q(
        \FIFO_U1/FIFO_SM1/N1 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_tri_enable_reg[4]  ( .E(
        \FIFO_U1/FIFO_SM1/N198 ), .D(\FIFO_U1/FIFO_SM1/N199 ), .Q(
        \FIFO_U1/FIFO_SM1/N5 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_tri_enable_reg[2]  ( .E(
        \FIFO_U1/FIFO_SM1/N198 ), .D(\FIFO_U1/FIFO_SM1/N199 ), .Q(
        \FIFO_U1/FIFO_SM1/N7 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_tri_enable_reg[0]  ( .E(
        \FIFO_U1/FIFO_SM1/N198 ), .D(\FIFO_U1/FIFO_SM1/N199 ), .Q(
        \FIFO_U1/FIFO_SM1/N9 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_tri_enable_reg[1]  ( .E(
        \FIFO_U1/FIFO_SM1/N198 ), .D(\FIFO_U1/FIFO_SM1/N199 ), .Q(
        \FIFO_U1/FIFO_SM1/N8 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_tri_enable_reg[3]  ( .E(
        \FIFO_U1/FIFO_SM1/N198 ), .D(\FIFO_U1/FIFO_SM1/N199 ), .Q(
        \FIFO_U1/FIFO_SM1/N6 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/FullFIFOReg_reg  ( .E(\FIFO_U1/FIFO_SM1/N189 ), .D(
        \FIFO_U1/FIFO_SM1/N148 ), .Q(FIFOFull) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_reg[1]  ( .E(\FIFO_U1/FIFO_SM1/N209 ), .D(
        \FIFO_U1/FIFO_SM1/N170 ), .Q(\FIFO_U1/FIFO_SM1/N221 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_reg[1]  ( .E(\FIFO_U1/FIFO_SM1/N198 ), 
        .D(\FIFO_U1/FIFO_SM1/N153 ), .Q(\FIFO_U1/FIFO_SM1/N236 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_reg[2]  ( .E(\FIFO_U1/FIFO_SM1/N198 ), 
        .D(\FIFO_U1/FIFO_SM1/N156 ), .Q(\FIFO_U1/FIFO_SM1/N233 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_reg[2]  ( .E(\FIFO_U1/FIFO_SM1/N209 ), .D(
        \FIFO_U1/FIFO_SM1/N173 ), .Q(\FIFO_U1/FIFO_SM1/N218 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCount_reg[3]  ( .E(\FIFO_U1/FIFO_SM1/N198 ), 
        .D(\FIFO_U1/FIFO_SM1/N159 ), .Q(\FIFO_U1/FIFO_SM1/N230 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCount_reg[3]  ( .E(\FIFO_U1/FIFO_SM1/N209 ), .D(
        \FIFO_U1/FIFO_SM1/N176 ), .Q(\FIFO_U1/FIFO_SM1/N215 ) );
  LHQD1 \FIFO_U1/FIFO_SM1/ReadCmdReg_reg  ( .E(\FIFO_U1/FIFO_SM1/N185 ), .D(
        \FIFO_U1/FIFO_SM1/N184 ), .Q(\FIFO_U1/SM_MemReadCmd ) );
  LHQD1 \FIFO_U1/FIFO_SM1/WriteCmdReg_reg  ( .E(\FIFO_U1/FIFO_SM1/N200 ), .D(
        \FIFO_U1/FIFO_SM1/N165 ), .Q(\FIFO_U1/SM_MemWriteCmd ) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[31]  ( .I(\FIFO_U1/RegFile1/DataOreg[31] ), .OE(n419), .Z(FIFO_Out[31]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[30]  ( .I(\FIFO_U1/RegFile1/DataOreg[30] ), .OE(n419), .Z(FIFO_Out[30]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[29]  ( .I(\FIFO_U1/RegFile1/DataOreg[29] ), .OE(n419), .Z(FIFO_Out[29]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[28]  ( .I(\FIFO_U1/RegFile1/DataOreg[28] ), .OE(n419), .Z(FIFO_Out[28]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[27]  ( .I(\FIFO_U1/RegFile1/DataOreg[27] ), .OE(n419), .Z(FIFO_Out[27]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[26]  ( .I(\FIFO_U1/RegFile1/DataOreg[26] ), .OE(n419), .Z(FIFO_Out[26]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[25]  ( .I(\FIFO_U1/RegFile1/DataOreg[25] ), .OE(n419), .Z(FIFO_Out[25]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[24]  ( .I(\FIFO_U1/RegFile1/DataOreg[24] ), .OE(n419), .Z(FIFO_Out[24]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[23]  ( .I(\FIFO_U1/RegFile1/DataOreg[23] ), .OE(n419), .Z(FIFO_Out[23]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[22]  ( .I(\FIFO_U1/RegFile1/DataOreg[22] ), .OE(n419), .Z(FIFO_Out[22]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[21]  ( .I(\FIFO_U1/RegFile1/DataOreg[21] ), .OE(n419), .Z(FIFO_Out[21]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[20]  ( .I(\FIFO_U1/RegFile1/DataOreg[20] ), .OE(n419), .Z(FIFO_Out[20]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[19]  ( .I(\FIFO_U1/RegFile1/DataOreg[19] ), .OE(n419), .Z(FIFO_Out[19]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[18]  ( .I(\FIFO_U1/RegFile1/DataOreg[18] ), .OE(n419), .Z(FIFO_Out[18]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[17]  ( .I(\FIFO_U1/RegFile1/DataOreg[17] ), .OE(n419), .Z(FIFO_Out[17]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[16]  ( .I(\FIFO_U1/RegFile1/DataOreg[16] ), .OE(n419), .Z(FIFO_Out[16]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[15]  ( .I(\FIFO_U1/RegFile1/DataOreg[15] ), .OE(n419), .Z(FIFO_Out[15]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[14]  ( .I(\FIFO_U1/RegFile1/DataOreg[14] ), .OE(n419), .Z(FIFO_Out[14]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[13]  ( .I(\FIFO_U1/RegFile1/DataOreg[13] ), .OE(n419), .Z(FIFO_Out[13]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[12]  ( .I(\FIFO_U1/RegFile1/DataOreg[12] ), .OE(n419), .Z(FIFO_Out[12]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[11]  ( .I(\FIFO_U1/RegFile1/DataOreg[11] ), .OE(n419), .Z(FIFO_Out[11]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[10]  ( .I(\FIFO_U1/RegFile1/DataOreg[10] ), .OE(n419), .Z(FIFO_Out[10]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[9]  ( .I(\FIFO_U1/RegFile1/DataOreg[9] ), 
        .OE(n419), .Z(FIFO_Out[9]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[8]  ( .I(\FIFO_U1/RegFile1/DataOreg[8] ), 
        .OE(n419), .Z(FIFO_Out[8]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[7]  ( .I(\FIFO_U1/RegFile1/DataOreg[7] ), 
        .OE(n419), .Z(FIFO_Out[7]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[6]  ( .I(\FIFO_U1/RegFile1/DataOreg[6] ), 
        .OE(n419), .Z(FIFO_Out[6]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[5]  ( .I(\FIFO_U1/RegFile1/DataOreg[5] ), 
        .OE(n419), .Z(FIFO_Out[5]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[4]  ( .I(\FIFO_U1/RegFile1/DataOreg[4] ), 
        .OE(n419), .Z(FIFO_Out[4]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[3]  ( .I(\FIFO_U1/RegFile1/DataOreg[3] ), 
        .OE(n419), .Z(FIFO_Out[3]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[2]  ( .I(\FIFO_U1/RegFile1/DataOreg[2] ), 
        .OE(n419), .Z(FIFO_Out[2]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[1]  ( .I(\FIFO_U1/RegFile1/DataOreg[1] ), 
        .OE(n419), .Z(FIFO_Out[1]) );
  BUFTD1 \FIFO_U1/RegFile1/DataO_tri[0]  ( .I(\FIFO_U1/RegFile1/DataOreg[0] ), 
        .OE(n419), .Z(FIFO_Out[0]) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[31]  ( .I(\FIFO_U1/RegFile1/N2330 ), 
        .OE(n418), .Z(\FIFO_U1/RegFile1/DataOreg[31] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[30]  ( .I(\FIFO_U1/RegFile1/N2333 ), 
        .OE(n417), .Z(\FIFO_U1/RegFile1/DataOreg[30] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[29]  ( .I(\FIFO_U1/RegFile1/N2336 ), 
        .OE(n416), .Z(\FIFO_U1/RegFile1/DataOreg[29] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[28]  ( .I(\FIFO_U1/RegFile1/N2339 ), 
        .OE(n415), .Z(\FIFO_U1/RegFile1/DataOreg[28] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[27]  ( .I(\FIFO_U1/RegFile1/N2342 ), 
        .OE(n414), .Z(\FIFO_U1/RegFile1/DataOreg[27] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[26]  ( .I(\FIFO_U1/RegFile1/N2345 ), 
        .OE(n413), .Z(\FIFO_U1/RegFile1/DataOreg[26] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[25]  ( .I(\FIFO_U1/RegFile1/N2348 ), 
        .OE(n412), .Z(\FIFO_U1/RegFile1/DataOreg[25] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[24]  ( .I(\FIFO_U1/RegFile1/N2351 ), 
        .OE(n411), .Z(\FIFO_U1/RegFile1/DataOreg[24] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[23]  ( .I(\FIFO_U1/RegFile1/N2354 ), 
        .OE(n410), .Z(\FIFO_U1/RegFile1/DataOreg[23] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[22]  ( .I(\FIFO_U1/RegFile1/N2357 ), 
        .OE(n409), .Z(\FIFO_U1/RegFile1/DataOreg[22] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[21]  ( .I(\FIFO_U1/RegFile1/N2360 ), 
        .OE(n408), .Z(\FIFO_U1/RegFile1/DataOreg[21] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[20]  ( .I(\FIFO_U1/RegFile1/N2363 ), 
        .OE(n407), .Z(\FIFO_U1/RegFile1/DataOreg[20] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[19]  ( .I(\FIFO_U1/RegFile1/N2366 ), 
        .OE(n406), .Z(\FIFO_U1/RegFile1/DataOreg[19] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[18]  ( .I(\FIFO_U1/RegFile1/N2369 ), 
        .OE(n405), .Z(\FIFO_U1/RegFile1/DataOreg[18] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[17]  ( .I(\FIFO_U1/RegFile1/N2372 ), 
        .OE(n404), .Z(\FIFO_U1/RegFile1/DataOreg[17] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[16]  ( .I(\FIFO_U1/RegFile1/N2375 ), 
        .OE(n403), .Z(\FIFO_U1/RegFile1/DataOreg[16] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[15]  ( .I(\FIFO_U1/RegFile1/N2378 ), 
        .OE(n402), .Z(\FIFO_U1/RegFile1/DataOreg[15] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[14]  ( .I(\FIFO_U1/RegFile1/N2381 ), 
        .OE(n401), .Z(\FIFO_U1/RegFile1/DataOreg[14] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[13]  ( .I(\FIFO_U1/RegFile1/N2384 ), 
        .OE(n400), .Z(\FIFO_U1/RegFile1/DataOreg[13] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[12]  ( .I(\FIFO_U1/RegFile1/N2387 ), 
        .OE(n399), .Z(\FIFO_U1/RegFile1/DataOreg[12] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[11]  ( .I(\FIFO_U1/RegFile1/N2390 ), 
        .OE(n398), .Z(\FIFO_U1/RegFile1/DataOreg[11] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[10]  ( .I(\FIFO_U1/RegFile1/N2393 ), 
        .OE(n397), .Z(\FIFO_U1/RegFile1/DataOreg[10] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[9]  ( .I(\FIFO_U1/RegFile1/N2396 ), 
        .OE(n396), .Z(\FIFO_U1/RegFile1/DataOreg[9] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[8]  ( .I(\FIFO_U1/RegFile1/N2399 ), 
        .OE(n395), .Z(\FIFO_U1/RegFile1/DataOreg[8] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[7]  ( .I(\FIFO_U1/RegFile1/N2402 ), 
        .OE(n394), .Z(\FIFO_U1/RegFile1/DataOreg[7] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[6]  ( .I(\FIFO_U1/RegFile1/N2405 ), 
        .OE(n393), .Z(\FIFO_U1/RegFile1/DataOreg[6] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[5]  ( .I(\FIFO_U1/RegFile1/N2408 ), 
        .OE(n392), .Z(\FIFO_U1/RegFile1/DataOreg[5] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[4]  ( .I(\FIFO_U1/RegFile1/N2411 ), 
        .OE(n391), .Z(\FIFO_U1/RegFile1/DataOreg[4] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[3]  ( .I(\FIFO_U1/RegFile1/N2414 ), 
        .OE(n390), .Z(\FIFO_U1/RegFile1/DataOreg[3] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[2]  ( .I(\FIFO_U1/RegFile1/N2417 ), 
        .OE(n389), .Z(\FIFO_U1/RegFile1/DataOreg[2] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[1]  ( .I(\FIFO_U1/RegFile1/N2420 ), 
        .OE(n388), .Z(\FIFO_U1/RegFile1/DataOreg[1] ) );
  BUFTD1 \FIFO_U1/RegFile1/DataOreg_tri[0]  ( .I(\FIFO_U1/RegFile1/N2423 ), 
        .OE(n387), .Z(\FIFO_U1/RegFile1/DataOreg[0] ) );
  BUFTD1 \FIFO_U1/FIFO_SM1/ReadCount_tri[4]  ( .I(\FIFO_U1/FIFO_SM1/N212 ), 
        .OE(n386), .Z(\FIFO_U1/SM_ReadAddr [4]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/ReadCount_tri[3]  ( .I(\FIFO_U1/FIFO_SM1/N215 ), 
        .OE(n385), .Z(\FIFO_U1/SM_ReadAddr [3]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/ReadCount_tri[2]  ( .I(\FIFO_U1/FIFO_SM1/N218 ), 
        .OE(n384), .Z(\FIFO_U1/SM_ReadAddr [2]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/ReadCount_tri[1]  ( .I(\FIFO_U1/FIFO_SM1/N221 ), 
        .OE(n383), .Z(\FIFO_U1/SM_ReadAddr [1]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/ReadCount_tri[0]  ( .I(\FIFO_U1/FIFO_SM1/N224 ), 
        .OE(n382), .Z(\FIFO_U1/SM_ReadAddr [0]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/WriteCount_tri[4]  ( .I(\FIFO_U1/FIFO_SM1/N227 ), 
        .OE(n381), .Z(\FIFO_U1/SM_WriteAddr [4]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/WriteCount_tri[3]  ( .I(\FIFO_U1/FIFO_SM1/N230 ), 
        .OE(n380), .Z(\FIFO_U1/SM_WriteAddr [3]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/WriteCount_tri[2]  ( .I(\FIFO_U1/FIFO_SM1/N233 ), 
        .OE(n379), .Z(\FIFO_U1/SM_WriteAddr [2]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/WriteCount_tri[1]  ( .I(\FIFO_U1/FIFO_SM1/N236 ), 
        .OE(n378), .Z(\FIFO_U1/SM_WriteAddr [1]) );
  BUFTD1 \FIFO_U1/FIFO_SM1/WriteCount_tri[0]  ( .I(\FIFO_U1/FIFO_SM1/N239 ), 
        .OE(n377), .Z(\FIFO_U1/SM_WriteAddr [0]) );
  Deserializer_DW01_incdec_0 r255 ( .A({
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[5] , 
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[4] , 
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] , 
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[2] , 
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] , 
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[0] }), .INC_DEC(\U3/U2/Z_0 ), 
        .SUM({\SerialRx_U1/PLL_RxU1/VFO1/N55 , \SerialRx_U1/PLL_RxU1/VFO1/N53 , 
        \SerialRx_U1/PLL_RxU1/VFO1/N51 , \SerialRx_U1/PLL_RxU1/VFO1/N49 , 
        \SerialRx_U1/PLL_RxU1/VFO1/N47 , \SerialRx_U1/PLL_RxU1/VFO1/N45 }) );
  Deserializer_DW01_inc_0 \SerialRx_U1/PLL_RxU1/MCntr1/add_16  ( .A({
        \SerialRx_U1/PLL_RxU1/CtrCarry , \SerialRx_U1/PLL_RxU1/MCntr1/Ctr }), 
        .SUM({\SerialRx_U1/PLL_RxU1/MCntr1/N5 , 
        \SerialRx_U1/PLL_RxU1/MCntr1/N4 , \SerialRx_U1/PLL_RxU1/MCntr1/N3 , 
        \SerialRx_U1/PLL_RxU1/MCntr1/N2 , \SerialRx_U1/PLL_RxU1/MCntr1/N1 })
         );
  Deserializer_DW01_inc_1 \DesDecoder_U1/SerClockGen/add_170_C252_S2  ( .A(
        \DesDecoder_U1/Count32 ), .SUM({\DesDecoder_U1/N53 , 
        \DesDecoder_U1/N52 , \DesDecoder_U1/N51 , \DesDecoder_U1/N50 , 
        \DesDecoder_U1/N49 }) );
  Deserializer_DW01_inc_2 \SerialRx_U1/PLL_RxU1/VFO1/ClockOutGen/add_161  ( 
        .A({\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[5] , 
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[4] , 
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[3] , 
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[2] , 
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[1] , 
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[0] }), .SUM({
        \SerialRx_U1/PLL_RxU1/VFO1/N14 , \SerialRx_U1/PLL_RxU1/VFO1/N13 , 
        \SerialRx_U1/PLL_RxU1/VFO1/N12 , \SerialRx_U1/PLL_RxU1/VFO1/N11 , 
        \SerialRx_U1/PLL_RxU1/VFO1/N10 , \SerialRx_U1/PLL_RxU1/VFO1/N9 }) );
  Deserializer_DW01_inc_3 \FIFO_U1/FIFO_SM1/add_183  ( .A({
        \FIFO_U1/FIFO_SM1/N76 , \FIFO_U1/FIFO_SM1/N75 , \FIFO_U1/FIFO_SM1/N74 , 
        \FIFO_U1/FIFO_SM1/N73 , \FIFO_U1/FIFO_SM1/N72 }), .SUM({
        \FIFO_U1/FIFO_SM1/N92 , \FIFO_U1/FIFO_SM1/N91 , \FIFO_U1/FIFO_SM1/N90 , 
        \FIFO_U1/FIFO_SM1/N89 , \FIFO_U1/FIFO_SM1/N88 }) );
  Deserializer_DW01_inc_4 r231 ( .A(\FIFO_U1/SM_WriteAddr ), .SUM({
        \FIFO_U1/FIFO_SM1/N76 , \FIFO_U1/FIFO_SM1/N75 , \FIFO_U1/FIFO_SM1/N74 , 
        \FIFO_U1/FIFO_SM1/N73 , \FIFO_U1/FIFO_SM1/N72 }) );
  Deserializer_DW01_inc_5 \FIFO_U1/FIFO_SM1/add_196  ( .A({
        \FIFO_U1/FIFO_SM1/N126 , \FIFO_U1/FIFO_SM1/N125 , 
        \FIFO_U1/FIFO_SM1/N124 , \FIFO_U1/FIFO_SM1/N123 , 
        \FIFO_U1/FIFO_SM1/N122 }), .SUM({\FIFO_U1/FIFO_SM1/N109 , 
        \FIFO_U1/FIFO_SM1/N108 , \FIFO_U1/FIFO_SM1/N107 , 
        \FIFO_U1/FIFO_SM1/N106 , \FIFO_U1/FIFO_SM1/N105 }) );
  Deserializer_DW01_inc_6 r197 ( .A({\U3/U1/Z_4 , \U3/U1/Z_3 , \U3/U1/Z_2 , 
        \U3/U1/Z_1 , \U3/U1/Z_0 }), .SUM({\FIFO_U1/FIFO_SM1/N126 , 
        \FIFO_U1/FIFO_SM1/N125 , \FIFO_U1/FIFO_SM1/N124 , 
        \FIFO_U1/FIFO_SM1/N123 , \FIFO_U1/FIFO_SM1/N122 }) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[63]  ( .D(\DesDecoder_U1/FrameSR[62] ), 
        .CPN(n636), .CDN(n596), .QN(n375) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n679), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[26][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n687), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[26][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n686), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[26][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n690), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[26][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n670), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[26][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n682), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[26][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n687), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[26][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n687), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[26][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n667), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[26][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n696), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[26][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n683), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[26][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n686), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[26][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n688), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[26][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n694), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[26][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n682), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[26][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n695), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[26][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n677), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[26][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n694), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[26][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n670), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[26][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n670), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[26][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n677), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[26][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n684), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[26][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n685), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[26][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n692), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[26][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n683), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[26][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n687), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[26][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n693), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[26][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n675), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[26][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n696), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[26][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n684), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[26][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n627), .Q(\FIFO_U1/RegFile1/Storage[26][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[26][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2097 ), .CP(n689), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[26][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n688), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[24][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n671), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[24][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n679), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[24][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n681), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[24][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n683), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[24][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n667), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[24][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n696), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[24][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n683), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[24][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n691), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[24][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n689), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[24][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n594), .Q(\FIFO_U1/RegFile1/Storage[24][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n686), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[24][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n685), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[24][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n670), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[24][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n676), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[24][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n686), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[24][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n683), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[24][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n672), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[24][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n685), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[24][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n688), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[24][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n696), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[24][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n687), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[24][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n687), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[24][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n693), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[24][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n691), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[24][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n671), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[24][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n696), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[24][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n679), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[24][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n689), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[24][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n666), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[24][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n669), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[24][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[24][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2031 ), .CP(n687), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[24][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n668), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[30][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n674), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[30][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n684), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[30][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n672), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[30][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n679), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[30][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n667), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[30][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n679), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[30][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n690), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[30][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n618), .Q(\FIFO_U1/RegFile1/Storage[30][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n692), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[30][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n679), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[30][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n677), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[30][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n685), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[30][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n667), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[30][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n696), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[30][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n687), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[30][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n695), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[30][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n681), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[30][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n689), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[30][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n674), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[30][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n689), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[30][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n678), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[30][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n674), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[30][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n695), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[30][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n696), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[30][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n692), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[30][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n693), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[30][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n694), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[30][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n671), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[30][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n679), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[30][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n694), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[30][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[30][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2229 ), .CP(n684), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[30][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[31]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n685), 
        .CDN(n622), .Q(\FIFO_U1/RegFile1/N32 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[30]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n692), 
        .CDN(n633), .Q(\FIFO_U1/RegFile1/N33 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[29]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n679), 
        .CDN(n604), .Q(\FIFO_U1/RegFile1/N34 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[28]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n686), 
        .CDN(n606), .Q(\FIFO_U1/RegFile1/N35 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[27]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n688), 
        .CDN(n605), .Q(\FIFO_U1/RegFile1/N36 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[26]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n687), 
        .CDN(n630), .Q(\FIFO_U1/RegFile1/N37 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[25]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n671), 
        .CDN(n594), .Q(\FIFO_U1/RegFile1/N38 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[24]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n684), 
        .CDN(n606), .Q(\FIFO_U1/RegFile1/N39 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[23]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n675), 
        .CDN(n625), .Q(\FIFO_U1/RegFile1/N40 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[22]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n690), 
        .CDN(n627), .Q(\FIFO_U1/RegFile1/N41 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[21]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n668), 
        .CDN(n602), .Q(\FIFO_U1/RegFile1/N42 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[20]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n681), 
        .CDN(n615), .Q(\FIFO_U1/RegFile1/N43 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[19]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n688), 
        .CDN(n633), .Q(\FIFO_U1/RegFile1/N44 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[18]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n694), 
        .CDN(n620), .Q(\FIFO_U1/RegFile1/N45 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[17]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n695), 
        .CDN(n613), .Q(\FIFO_U1/RegFile1/N46 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[16]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n684), 
        .CDN(n612), .Q(\FIFO_U1/RegFile1/N47 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[15]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n671), 
        .CDN(n614), .Q(\FIFO_U1/RegFile1/N48 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[14]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n692), 
        .CDN(n593), .Q(\FIFO_U1/RegFile1/N49 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[13]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n693), 
        .CDN(n610), .Q(\FIFO_U1/RegFile1/N50 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[12]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n670), 
        .CDN(n635), .Q(\FIFO_U1/RegFile1/N51 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[11]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n676), 
        .CDN(n631), .Q(\FIFO_U1/RegFile1/N52 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[10]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n680), 
        .CDN(n596), .Q(\FIFO_U1/RegFile1/N53 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[9]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n688), 
        .CDN(n604), .Q(\FIFO_U1/RegFile1/N54 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[8]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n695), 
        .CDN(n629), .Q(\FIFO_U1/RegFile1/N55 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[7]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n688), 
        .CDN(n602), .Q(\FIFO_U1/RegFile1/N56 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[6]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n689), 
        .CDN(n593), .Q(\FIFO_U1/RegFile1/N57 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[5]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n685), 
        .CDN(n605), .Q(\FIFO_U1/RegFile1/N58 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[4]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n678), 
        .CDN(n592), .Q(\FIFO_U1/RegFile1/N59 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[3]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n686), 
        .CDN(n615), .Q(\FIFO_U1/RegFile1/N60 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[2]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n680), 
        .CDN(n626), .Q(\FIFO_U1/RegFile1/N61 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[1]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n690), 
        .CDN(n623), .Q(\FIFO_U1/RegFile1/N62 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_tri_enable_reg[0]  ( .D(
        \FIFO_U1/RegFile1/N2328 ), .E(\FIFO_U1/RegFile1/N2327 ), .CP(n683), 
        .CDN(n601), .Q(\FIFO_U1/RegFile1/N63 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n691), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[28][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n671), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[28][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n680), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[28][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n676), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[28][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n673), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[28][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n696), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[28][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n696), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[28][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n695), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[28][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n678), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[28][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n694), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[28][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n675), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[28][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n687), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[28][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n691), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[28][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n680), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[28][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n683), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[28][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n683), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[28][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n692), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[28][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n678), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[28][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n685), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[28][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n670), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[28][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n675), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[28][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n692), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[28][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n667), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[28][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n673), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[28][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n690), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[28][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n673), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[28][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n666), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[28][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n681), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[28][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n685), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[28][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n679), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[28][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n695), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[28][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[28][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2163 ), .CP(n686), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[28][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n687), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[29][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n688), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[29][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n689), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[29][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n690), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[29][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n691), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[29][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n684), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[29][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n669), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[29][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n686), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[29][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n690), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[29][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n689), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[29][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n687), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[29][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n688), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[29][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n681), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[29][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n680), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[29][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n669), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[29][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n696), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[29][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n670), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[29][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n673), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[29][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n688), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[29][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n689), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[29][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n686), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[29][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n684), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[29][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n685), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[29][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n693), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[29][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n679), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[29][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n690), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[29][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n674), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[29][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n694), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[29][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n687), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[29][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n688), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[29][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n666), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[29][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[29][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2196 ), .CP(n668), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[29][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n678), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[27][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n688), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[27][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n668), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[27][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n684), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[27][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n673), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[27][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n695), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[27][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n691), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[27][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n692), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[27][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n696), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[27][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n687), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[27][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n680), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[27][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n684), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[27][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n682), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[27][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n675), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[27][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n695), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[27][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n688), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[27][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n692), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[27][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n670), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[27][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n691), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[27][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n667), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[27][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n694), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[27][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n694), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[27][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n694), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[27][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n676), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[27][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n676), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[27][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n695), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[27][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n696), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[27][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n675), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[27][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n671), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[27][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n670), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[27][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n694), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[27][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[27][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2130 ), .CP(n677), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[27][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n672), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[25][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n677), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[25][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n695), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[25][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n681), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[25][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n669), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[25][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n692), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[25][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n691), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[25][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n674), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[25][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n681), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[25][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n674), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[25][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n685), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[25][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n691), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[25][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n685), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[25][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n696), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[25][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n671), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[25][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n680), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[25][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n684), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[25][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n677), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[25][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n666), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[25][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n691), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[25][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n695), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[25][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n668), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[25][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n689), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[25][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n684), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[25][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n680), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[25][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n690), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[25][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n668), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[25][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n671), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[25][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n620), .Q(\FIFO_U1/RegFile1/Storage[25][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n696), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[25][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n677), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[25][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[25][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2064 ), .CP(n689), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[25][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n674), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[22][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n673), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[22][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n684), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[22][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n681), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[22][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n690), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[22][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n685), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[22][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n680), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[22][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n682), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[22][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n695), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[22][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n690), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[22][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n674), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[22][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n674), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[22][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n672), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[22][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n691), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[22][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n667), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[22][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n667), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[22][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n672), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[22][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n669), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[22][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n684), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[22][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n682), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[22][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n685), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[22][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n695), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[22][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n669), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[22][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n694), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[22][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n690), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[22][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n685), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[22][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n695), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[22][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n691), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[22][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n685), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[22][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n669), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[22][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n675), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[22][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[22][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1965 ), .CP(n668), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[22][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[14][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[14][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[14][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[14][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n673), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n682), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[14][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n691), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[14][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n673), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[14][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n690), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[14][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n679), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[14][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n675), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[14][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n670), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[14][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n669), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[14][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[14][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[14][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[14][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[14][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[14][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[14][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[14][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[14][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1701 ), .CP(n668), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[14][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[6][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[6][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[6][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[6][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[6][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[6][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[6][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n683), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[6][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[6][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[6][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[6][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[6][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n676), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[6][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n695), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[6][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n695), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[6][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n679), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[6][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n696), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[6][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n694), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[6][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n674), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[6][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n696), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[6][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[6][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[6][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[6][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[6][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[6][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n682), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[6][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[6][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[6][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[6][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[6][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[6][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[6][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1437 ), .CP(n681), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[6][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n691), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[18][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n687), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[18][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n668), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[18][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n686), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[18][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n696), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[18][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n682), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[18][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n674), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[18][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n690), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[18][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n696), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[18][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n669), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[18][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n683), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[18][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n694), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[18][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n688), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[18][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n689), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[18][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n672), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[18][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n689), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[18][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n668), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[18][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n670), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[18][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n678), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[18][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n692), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[18][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n675), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[18][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n694), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[18][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n688), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[18][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n672), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[18][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n681), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[18][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n687), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[18][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n672), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[18][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n666), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[18][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n693), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[18][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n668), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[18][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n689), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[18][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[18][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1833 ), .CP(n682), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[18][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n676), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[10][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n677), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n678), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[10][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n686), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n671), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n682), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n680), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n681), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n668), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n667), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n666), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n670), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n685), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[10][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n687), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[10][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n693), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[10][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n692), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[10][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n668), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[10][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n672), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[10][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n684), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n693), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[10][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n679), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[10][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n679), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n673), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n677), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n673), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n669), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n674), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n672), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n675), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n683), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n677), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[10][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[10][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1569 ), .CP(n677), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[10][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n670), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[2][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n677), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[2][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n691), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[2][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n671), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[2][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n692), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[2][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n694), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[2][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n684), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[2][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n691), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[2][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n690), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[2][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n693), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[2][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n689), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[2][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n672), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[2][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n667), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[2][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n679), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[2][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n685), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[2][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n693), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[2][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n669), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[2][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n685), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[2][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n684), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[2][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n686), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[2][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n695), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[2][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n688), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[2][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n676), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[2][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n676), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[2][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n678), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[2][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n688), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[2][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n677), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[2][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n677), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[2][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n676), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[2][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n668), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[2][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n669), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[2][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[2][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1305 ), .CP(n666), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[2][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n692), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[21][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n696), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[21][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n669), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[21][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n690), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[21][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n681), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[21][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n692), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[21][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n667), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[21][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n666), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[21][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n666), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[21][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n681), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[21][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n667), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[21][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n689), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[21][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n693), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[21][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n688), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[21][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n668), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[21][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n681), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[21][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n669), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[21][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n685), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[21][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n692), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[21][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n687), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[21][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n684), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[21][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n689), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[21][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n686), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[21][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n689), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[21][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n678), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[21][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n680), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[21][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n675), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[21][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n689), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[21][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n671), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[21][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n689), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[21][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n687), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[21][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[21][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1932 ), .CP(n688), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[21][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[13][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[13][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[13][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[13][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[13][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[13][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[13][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[13][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n672), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[13][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[13][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[13][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n690), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[13][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n692), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[13][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n669), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[13][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n675), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[13][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n693), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[13][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n680), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[13][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n694), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[13][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n675), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[13][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[13][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[13][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[13][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[13][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[13][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n671), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[13][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1668 ), .CP(n670), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[13][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n686), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[5][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n671), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[5][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n666), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[5][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n667), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[5][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n666), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[5][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n670), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[5][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n693), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[5][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n687), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[5][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n675), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[5][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n674), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[5][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n677), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[5][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n676), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[5][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n696), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[5][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n693), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[5][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n696), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[5][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n692), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[5][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n680), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[5][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n696), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[5][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n684), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[5][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n696), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[5][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n666), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[5][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n691), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[5][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n674), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[5][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n675), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[5][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n674), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[5][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n673), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[5][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n672), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[5][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n677), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[5][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n676), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[5][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n668), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[5][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n683), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[5][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[5][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1404 ), .CP(n683), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[5][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n686), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[17][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n674), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[17][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n689), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[17][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n676), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[17][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n684), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[17][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n685), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[17][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n680), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[17][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n674), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[17][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n689), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[17][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n666), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[17][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n688), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[17][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n679), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[17][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n685), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[17][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n680), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[17][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n677), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[17][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n693), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[17][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n673), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[17][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n673), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[17][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n671), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[17][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n681), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[17][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n694), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[17][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n671), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[17][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n676), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[17][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n676), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[17][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n673), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[17][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n670), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[17][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n693), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[17][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n695), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[17][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n683), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[17][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n684), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[17][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n686), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[17][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[17][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1800 ), .CP(n679), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[17][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n673), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[9][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n667), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[9][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n667), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n693), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[9][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n692), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[9][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n686), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n673), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n668), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n675), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n683), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n672), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n674), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n690), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[9][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n676), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[9][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n691), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[9][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n694), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[9][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n694), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[9][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n693), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[9][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n690), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[9][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n682), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[9][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n669), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n685), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n684), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n690), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[9][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n679), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n673), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n680), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n693), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n692), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n686), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n691), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[9][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1536 ), .CP(n689), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[9][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n671), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[1][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n679), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[1][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n667), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[1][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n666), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[1][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n694), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[1][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n692), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[1][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n693), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[1][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n692), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[1][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n678), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[1][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n672), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[1][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n683), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[1][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n682), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[1][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n675), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[1][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n689), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[1][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n695), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[1][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n687), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[1][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n682), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[1][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n678), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[1][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n694), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[1][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n693), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[1][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n681), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[1][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n680), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[1][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n679), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[1][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n678), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[1][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n685), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[1][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n686), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[1][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n682), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[1][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n682), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[1][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n689), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[1][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n677), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[1][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n676), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[1][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[1][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1272 ), .CP(n670), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[1][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n691), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n694), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n689), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n696), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n683), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n693), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n674), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n680), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n668), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n609), .Q(\FIFO_U1/RegFile1/Storage[20][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n673), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n685), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n683), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[20][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n687), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[20][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n676), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[20][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n695), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[20][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n667), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[20][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n687), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[20][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n695), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[20][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n682), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[20][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n688), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n688), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n693), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n666), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n608), .Q(\FIFO_U1/RegFile1/Storage[20][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n691), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[20][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n684), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[20][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n674), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n696), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n686), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[20][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n695), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[20][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[20][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1899 ), .CP(n668), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[20][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[12][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[12][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[12][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[12][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n684), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n688), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[12][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n668), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[12][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n693), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[12][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n666), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[12][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n694), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[12][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n696), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[12][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n686), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[12][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[12][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n674), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[12][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[12][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[12][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[12][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[12][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[12][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[12][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[12][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[12][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[12][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[12][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1635 ), .CP(n673), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[12][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n670), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[4][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n685), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[4][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n673), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[4][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n672), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[4][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n682), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[4][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n673), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[4][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n666), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[4][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n670), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[4][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n671), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[4][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n678), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[4][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n668), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[4][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n666), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[4][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n695), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[4][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n686), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[4][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n687), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[4][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n692), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[4][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n670), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[4][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n671), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[4][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n677), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[4][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n666), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[4][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n667), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[4][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n675), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[4][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n674), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[4][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n677), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[4][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n675), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[4][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n690), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[4][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n687), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[4][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n686), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[4][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n689), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[4][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n691), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[4][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n672), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[4][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[4][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1371 ), .CP(n669), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[4][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n685), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[23][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n684), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[23][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n627), .Q(\FIFO_U1/RegFile1/Storage[23][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n691), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[23][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n695), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[23][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n682), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[23][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n677), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[23][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n671), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[23][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n682), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[23][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n678), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[23][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n675), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[23][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n685), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[23][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n672), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[23][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n669), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[23][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n681), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[23][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n681), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[23][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n681), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[23][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n695), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[23][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n690), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[23][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n692), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[23][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n686), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[23][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n691), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[23][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n680), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[23][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n671), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[23][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n692), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[23][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n678), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[23][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n681), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[23][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n673), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[23][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n693), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[23][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n690), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[23][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n668), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[23][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[23][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1998 ), .CP(n669), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[23][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n668), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[15][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n667), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[15][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n667), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[15][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n667), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[15][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n667), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[15][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n667), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[15][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[15][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[15][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[15][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[15][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[15][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n686), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[15][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n679), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[15][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n686), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[15][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n666), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[15][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n690), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[15][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n678), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[15][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n669), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[15][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n675), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[15][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n683), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[15][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n684), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[15][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n691), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[15][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n668), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[15][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n694), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[15][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n685), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[15][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n672), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[15][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n696), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[15][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n675), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[15][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n678), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[15][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n677), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[15][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n682), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[15][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[15][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1734 ), .CP(n683), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[15][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n681), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[7][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n681), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[7][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n681), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[7][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n681), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[7][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[7][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[7][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[7][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[7][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[7][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[7][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[7][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[7][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n694), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[7][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n676), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[7][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n678), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[7][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n667), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[7][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[7][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n672), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[7][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n695), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[7][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[7][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[7][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n680), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[7][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[7][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[7][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[7][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[7][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[7][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[7][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[7][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[7][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[7][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[7][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1470 ), .CP(n679), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[7][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n688), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[19][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n691), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[19][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n683), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[19][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n668), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[19][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n681), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[19][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n685), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[19][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n684), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[19][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n669), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[19][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n691), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[19][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n668), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[19][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n695), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n690), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n693), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[19][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n690), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[19][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n694), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[19][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n666), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[19][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n688), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[19][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n693), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[19][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n690), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[19][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n674), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[19][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n689), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n696), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n692), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n694), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[19][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n673), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n690), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n691), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n671), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n684), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n682), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n666), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[19][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1866 ), .CP(n692), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[19][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[11][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[11][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[11][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[11][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[11][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[11][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[11][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[11][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[11][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[11][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n616), .Q(
        \FIFO_U1/RegFile1/Storage[11][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n672), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[11][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n677), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[11][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n673), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[11][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n683), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[11][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n682), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[11][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n687), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[11][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n691), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[11][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n678), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[11][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n676), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[11][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[11][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[11][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1602 ), .CP(n675), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[11][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n693), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[3][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n681), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[3][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n676), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[3][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n691), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[3][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n695), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[3][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n676), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[3][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n667), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[3][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n685), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[3][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n669), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[3][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n687), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[3][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n681), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[3][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n680), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[3][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n668), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[3][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n685), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[3][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n686), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[3][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n669), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[3][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n673), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[3][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n678), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[3][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n689), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[3][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n676), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[3][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n667), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[3][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n666), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[3][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n670), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[3][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n671), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[3][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n675), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[3][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n674), .CDN(n605), .Q(
        \FIFO_U1/RegFile1/Storage[3][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n677), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[3][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n676), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[3][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n673), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[3][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n669), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[3][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n672), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[3][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[3][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1338 ), .CP(n683), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[3][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n672), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[16][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n675), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[16][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n695), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[16][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n669), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[16][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n674), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[16][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n696), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[16][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n670), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[16][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n695), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[16][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n687), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[16][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n683), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[16][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n678), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[16][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n678), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[16][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n690), .CDN(n601), .Q(
        \FIFO_U1/RegFile1/Storage[16][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n677), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[16][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n683), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[16][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n696), .CDN(n635), .Q(
        \FIFO_U1/RegFile1/Storage[16][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n678), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[16][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n681), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[16][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n694), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[16][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n686), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[16][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n667), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[16][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n693), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[16][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n682), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[16][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n684), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[16][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n688), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[16][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n687), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[16][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n689), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[16][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n690), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/Storage[16][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n696), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[16][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n679), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[16][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n691), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[16][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[16][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1767 ), .CP(n684), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[16][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[8][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[8][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[8][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[8][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[8][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/Storage[8][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[8][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n591), .Q(
        \FIFO_U1/RegFile1/Storage[8][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[8][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[8][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n678), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/Storage[8][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n672), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[8][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n687), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[8][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n684), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[8][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n680), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[8][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n688), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/Storage[8][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n687), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[8][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n670), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[8][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n672), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/Storage[8][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n687), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[8][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n679), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/Storage[8][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n683), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/Storage[8][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n692), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[8][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n693), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[8][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n686), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[8][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n684), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[8][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n694), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[8][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n690), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[8][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n676), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[8][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n688), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[8][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n695), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[8][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[8][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1503 ), .CP(n694), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/Storage[8][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n696), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[0][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n667), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[0][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n686), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[0][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n680), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[0][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n684), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[0][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n681), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[0][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n667), .CDN(n600), .Q(
        \FIFO_U1/RegFile1/Storage[0][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n694), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[0][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n668), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[0][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n670), .CDN(n491), .Q(
        \FIFO_U1/RegFile1/Storage[0][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n687), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/Storage[0][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n688), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[0][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n675), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[0][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n683), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[0][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n686), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[0][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n667), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[0][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n676), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[0][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n686), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[0][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n689), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[0][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n689), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[0][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n696), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[0][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n686), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/Storage[0][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n689), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[0][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(\FIFO_U1/RegFile1/ChipClock ), .CDN(
        n624), .Q(\FIFO_U1/RegFile1/Storage[0][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n688), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[0][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n682), .CDN(n594), .Q(
        \FIFO_U1/RegFile1/Storage[0][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n669), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/Storage[0][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n692), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[0][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n694), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[0][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n670), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[0][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n666), .CDN(n619), .Q(
        \FIFO_U1/RegFile1/Storage[0][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[0][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N1239 ), .CP(n684), .CDN(n614), .Q(
        \FIFO_U1/RegFile1/Storage[0][30] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][31]  ( .D(DecodeToFIFO[31]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n685), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[31][31] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][29]  ( .D(DecodeToFIFO[29]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n690), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[31][29] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][27]  ( .D(DecodeToFIFO[27]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n691), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[31][27] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][25]  ( .D(DecodeToFIFO[25]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n692), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/Storage[31][25] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][23]  ( .D(DecodeToFIFO[23]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n680), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[31][23] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][21]  ( .D(DecodeToFIFO[21]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n682), .CDN(n628), .Q(
        \FIFO_U1/RegFile1/Storage[31][21] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][19]  ( .D(DecodeToFIFO[19]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n695), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/Storage[31][19] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][17]  ( .D(DecodeToFIFO[17]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n676), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/Storage[31][17] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][15]  ( .D(DecodeToFIFO[15]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n687), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[31][15] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][13]  ( .D(DecodeToFIFO[13]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n679), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/Storage[31][13] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][11]  ( .D(DecodeToFIFO[11]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n671), .CDN(n618), .Q(
        \FIFO_U1/RegFile1/Storage[31][11] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][9]  ( .D(DecodeToFIFO[9]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n693), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[31][9] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][7]  ( .D(DecodeToFIFO[7]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n692), .CDN(n617), .Q(
        \FIFO_U1/RegFile1/Storage[31][7] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][5]  ( .D(DecodeToFIFO[5]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n681), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/Storage[31][5] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][3]  ( .D(DecodeToFIFO[3]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n692), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/Storage[31][3] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][1]  ( .D(DecodeToFIFO[1]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n696), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/Storage[31][1] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][0]  ( .D(DecodeToFIFO[0]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n671), .CDN(n623), .Q(
        \FIFO_U1/RegFile1/Storage[31][0] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][2]  ( .D(DecodeToFIFO[2]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n685), .CDN(n629), .Q(
        \FIFO_U1/RegFile1/Storage[31][2] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][4]  ( .D(DecodeToFIFO[4]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n688), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[31][4] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][6]  ( .D(DecodeToFIFO[6]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n692), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/Storage[31][6] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][8]  ( .D(DecodeToFIFO[8]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n688), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/Storage[31][8] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][10]  ( .D(DecodeToFIFO[10]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n666), .CDN(n622), .Q(
        \FIFO_U1/RegFile1/Storage[31][10] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][12]  ( .D(DecodeToFIFO[12]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n696), .CDN(n613), .Q(
        \FIFO_U1/RegFile1/Storage[31][12] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][14]  ( .D(DecodeToFIFO[14]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n677), .CDN(n626), .Q(
        \FIFO_U1/RegFile1/Storage[31][14] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][16]  ( .D(DecodeToFIFO[16]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n670), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/Storage[31][16] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][18]  ( .D(DecodeToFIFO[18]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n677), .CDN(n633), .Q(
        \FIFO_U1/RegFile1/Storage[31][18] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][20]  ( .D(DecodeToFIFO[20]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n693), .CDN(n632), .Q(
        \FIFO_U1/RegFile1/Storage[31][20] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][22]  ( .D(DecodeToFIFO[22]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n683), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/Storage[31][22] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][24]  ( .D(DecodeToFIFO[24]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n672), .CDN(n634), .Q(
        \FIFO_U1/RegFile1/Storage[31][24] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][26]  ( .D(DecodeToFIFO[26]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n690), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/Storage[31][26] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][28]  ( .D(DecodeToFIFO[28]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n688), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/Storage[31][28] ) );
  EDFCNQD1 \FIFO_U1/RegFile1/Storage_reg[31][30]  ( .D(DecodeToFIFO[30]), .E(
        \FIFO_U1/RegFile1/N2262 ), .CP(n691), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/Storage[31][30] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[8]  ( .D(\DesDecoder_U1/FrameSR[7] ), 
        .CPN(n637), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[8] ), .QN(n281) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[9]  ( .D(\DesDecoder_U1/FrameSR[8] ), 
        .CPN(n487), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[9] ), .QN(n283) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[10]  ( .D(\DesDecoder_U1/FrameSR[9] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[10] ), .QN(n285) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[11]  ( .D(\DesDecoder_U1/FrameSR[10] ), 
        .CPN(n638), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[11] ), .QN(n287) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[12]  ( .D(\DesDecoder_U1/FrameSR[11] ), 
        .CPN(n638), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[12] ), .QN(n289) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[13]  ( .D(\DesDecoder_U1/FrameSR[12] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[13] ), .QN(n291) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[14]  ( .D(\DesDecoder_U1/FrameSR[13] ), 
        .CPN(n638), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[14] ), .QN(n293) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[15]  ( .D(\DesDecoder_U1/FrameSR[14] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[15] ), .QN(n295) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[18]  ( .D(\DesDecoder_U1/FrameSR[17] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[18] ), .QN(n368) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[19]  ( .D(\DesDecoder_U1/FrameSR[18] ), 
        .CPN(n638), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[19] ), .QN(n374) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[22]  ( .D(\DesDecoder_U1/FrameSR[21] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[22] ), .QN(n1250) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[24]  ( .D(\DesDecoder_U1/FrameSR[23] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[24] ), .QN(n297) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[25]  ( .D(\DesDecoder_U1/FrameSR[24] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[25] ), .QN(n299) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[26]  ( .D(\DesDecoder_U1/FrameSR[25] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[26] ), .QN(n301) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[27]  ( .D(\DesDecoder_U1/FrameSR[26] ), 
        .CPN(n637), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[27] ), .QN(n303) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[28]  ( .D(\DesDecoder_U1/FrameSR[27] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[28] ), .QN(n305) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[29]  ( .D(\DesDecoder_U1/FrameSR[28] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[29] ), .QN(n307) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[30]  ( .D(\DesDecoder_U1/FrameSR[29] ), 
        .CPN(n637), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[30] ), .QN(n309) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[31]  ( .D(\DesDecoder_U1/FrameSR[30] ), 
        .CPN(n636), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[31] ), .QN(n311) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[32]  ( .D(\DesDecoder_U1/FrameSR[31] ), 
        .CPN(n636), .CDN(n600), .Q(\DesDecoder_U1/FrameSR[32] ), .QN(n1249) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[34]  ( .D(\DesDecoder_U1/FrameSR[33] ), 
        .CPN(n636), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[34] ), .QN(n360) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[35]  ( .D(\DesDecoder_U1/FrameSR[34] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[35] ), .QN(n361) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[38]  ( .D(\DesDecoder_U1/FrameSR[37] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[38] ), .QN(n1251) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[40]  ( .D(\DesDecoder_U1/FrameSR[39] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[40] ), .QN(n313) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[41]  ( .D(\DesDecoder_U1/FrameSR[40] ), 
        .CPN(n487), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[41] ), .QN(n315) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[42]  ( .D(\DesDecoder_U1/FrameSR[41] ), 
        .CPN(n638), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[42] ), .QN(n317) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[43]  ( .D(\DesDecoder_U1/FrameSR[42] ), 
        .CPN(n637), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[43] ), .QN(n319) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[44]  ( .D(\DesDecoder_U1/FrameSR[43] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[44] ), .QN(n321) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[45]  ( .D(\DesDecoder_U1/FrameSR[44] ), 
        .CPN(n637), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[45] ), .QN(n323) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[46]  ( .D(\DesDecoder_U1/FrameSR[45] ), 
        .CPN(n487), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[46] ), .QN(n325) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[47]  ( .D(\DesDecoder_U1/FrameSR[46] ), 
        .CPN(n487), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[47] ), .QN(n327) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[48]  ( .D(\DesDecoder_U1/FrameSR[47] ), 
        .CPN(n638), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[48] ), .QN(n356) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[53]  ( .D(\DesDecoder_U1/FrameSR[52] ), 
        .CPN(n638), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[53] ), .QN(n1253) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[55]  ( .D(\DesDecoder_U1/FrameSR[54] ), 
        .CPN(n636), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[55] ), .QN(n1252) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[56]  ( .D(\DesDecoder_U1/FrameSR[55] ), 
        .CPN(n636), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[56] ), .QN(n329) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[57]  ( .D(\DesDecoder_U1/FrameSR[56] ), 
        .CPN(n487), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[57] ), .QN(n331) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[58]  ( .D(\DesDecoder_U1/FrameSR[57] ), 
        .CPN(n637), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[58] ), .QN(n333) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[59]  ( .D(\DesDecoder_U1/FrameSR[58] ), 
        .CPN(n636), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[59] ), .QN(n335) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[60]  ( .D(\DesDecoder_U1/FrameSR[59] ), 
        .CPN(n637), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[60] ), .QN(n337) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[61]  ( .D(\DesDecoder_U1/FrameSR[60] ), 
        .CPN(n487), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[61] ), .QN(n339) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[62]  ( .D(\DesDecoder_U1/FrameSR[61] ), 
        .CPN(n636), .CDN(n596), .Q(\DesDecoder_U1/FrameSR[62] ), .QN(n341) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[31]  ( .D(n486), .CPN(n637), .CDN(n596), 
        .QN(n561) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[30]  ( .D(n485), .CPN(n638), .CDN(n596), 
        .QN(n560) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[29]  ( .D(n484), .CPN(n487), .CDN(n596), 
        .QN(n559) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[28]  ( .D(n483), .CPN(n487), .CDN(n596), 
        .QN(n558) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[27]  ( .D(n482), .CPN(n487), .CDN(n596), 
        .QN(n557) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[26]  ( .D(n481), .CPN(n638), .CDN(n596), 
        .QN(n556) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[25]  ( .D(n480), .CPN(n487), .CDN(n596), 
        .QN(n555) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[24]  ( .D(n479), .CPN(n487), .CDN(n596), 
        .QN(n554) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[23]  ( .D(n478), .CPN(n637), .CDN(n595), 
        .QN(n553) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[22]  ( .D(n477), .CPN(n636), .CDN(n595), 
        .QN(n552) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[21]  ( .D(n476), .CPN(n638), .CDN(n595), 
        .QN(n551) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[20]  ( .D(n475), .CPN(n636), .CDN(n595), 
        .QN(n550) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[19]  ( .D(n474), .CPN(n636), .CDN(n595), 
        .QN(n549) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[18]  ( .D(n473), .CPN(n637), .CDN(n595), 
        .QN(n548) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[17]  ( .D(n472), .CPN(n638), .CDN(n595), 
        .QN(n547) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[16]  ( .D(n471), .CPN(n636), .CDN(n595), 
        .QN(n546) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[15]  ( .D(n470), .CPN(n636), .CDN(n595), 
        .QN(n545) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[14]  ( .D(n469), .CPN(n487), .CDN(n594), 
        .QN(n544) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[13]  ( .D(n468), .CPN(n638), .CDN(n594), 
        .QN(n543) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[12]  ( .D(n467), .CPN(n637), .CDN(n594), 
        .QN(n542) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[11]  ( .D(n466), .CPN(n487), .CDN(n594), 
        .QN(n541) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[10]  ( .D(n465), .CPN(n487), .CDN(n594), 
        .QN(n540) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[9]  ( .D(n464), .CPN(n487), .CDN(n594), 
        .QN(n539) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[8]  ( .D(n463), .CPN(n638), .CDN(n594), 
        .QN(n538) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[7]  ( .D(n462), .CPN(n487), .CDN(n591), 
        .QN(n537) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[6]  ( .D(n461), .CPN(n487), .CDN(n591), 
        .QN(n536) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[5]  ( .D(n460), .CPN(n638), .CDN(n591), 
        .QN(n535) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[4]  ( .D(n459), .CPN(n487), .CDN(n591), 
        .QN(n534) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[3]  ( .D(n458), .CPN(n638), .CDN(n597), 
        .QN(n533) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[2]  ( .D(n457), .CPN(n638), .CDN(n595), 
        .QN(n532) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[1]  ( .D(n456), .CPN(n637), .CDN(n598), 
        .QN(n531) );
  DFNCND1 \DesDecoder_U1/DecodeReg_reg[0]  ( .D(n455), .CPN(n638), .CDN(n601), 
        .QN(n530) );
  DFSNQD1 \SerialRx_U1/PLL_RxU1/Comp1/AdjustFreq_reg[0]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N19 ), .CP(\SerialRx_U1/PLL_RxU1/CtrCarry ), .SDN(n620), .Q(\SerialRx_U1/PLL_RxU1/AdjFreq [0]) );
  DFSNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[4]  ( .D(n489), .CP(
        \SerialRx_U1/PLL_RxU1/SampleWire ), .SDN(n620), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[4] ) );
  DFSNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[0]  ( .D(n454), .CP(
        \SerialRx_U1/PLL_RxU1/SampleWire ), .SDN(n620), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[0] ) );
  DFNCND1 \DesDecoder_U1/doParSync_reg  ( .D(\DesDecoder_U1/N12 ), .CPN(n637), 
        .CDN(n596), .Q(n1248) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[36]  ( .D(\DesDecoder_U1/FrameSR[35] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[36] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[51]  ( .D(\DesDecoder_U1/FrameSR[50] ), 
        .CPN(n636), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[51] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[52]  ( .D(\DesDecoder_U1/FrameSR[51] ), 
        .CPN(n637), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[52] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[0]  ( .D(SerRxToDecode), .CPN(n638), 
        .CDN(n603), .Q(\DesDecoder_U1/FrameSR[0] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[1]  ( .D(\DesDecoder_U1/FrameSR[0] ), 
        .CPN(n637), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[1] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[2]  ( .D(\DesDecoder_U1/FrameSR[1] ), 
        .CPN(n636), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[2] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[4]  ( .D(\DesDecoder_U1/FrameSR[3] ), 
        .CPN(n487), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[4] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[5]  ( .D(\DesDecoder_U1/FrameSR[4] ), 
        .CPN(n638), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[5] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[6]  ( .D(\DesDecoder_U1/FrameSR[5] ), 
        .CPN(n637), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[6] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[16]  ( .D(\DesDecoder_U1/FrameSR[15] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[16] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[17]  ( .D(\DesDecoder_U1/FrameSR[16] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[17] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[20]  ( .D(\DesDecoder_U1/FrameSR[19] ), 
        .CPN(n638), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[20] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[21]  ( .D(\DesDecoder_U1/FrameSR[20] ), 
        .CPN(n637), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[21] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[23]  ( .D(\DesDecoder_U1/FrameSR[22] ), 
        .CPN(n637), .CDN(n601), .Q(\DesDecoder_U1/FrameSR[23] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[33]  ( .D(\DesDecoder_U1/FrameSR[32] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[33] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[37]  ( .D(\DesDecoder_U1/FrameSR[36] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[37] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[39]  ( .D(\DesDecoder_U1/FrameSR[38] ), 
        .CPN(n636), .CDN(n599), .Q(\DesDecoder_U1/FrameSR[39] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[49]  ( .D(\DesDecoder_U1/FrameSR[48] ), 
        .CPN(n487), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[49] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[50]  ( .D(\DesDecoder_U1/FrameSR[49] ), 
        .CPN(n636), .CDN(n598), .Q(\DesDecoder_U1/FrameSR[50] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[54]  ( .D(\DesDecoder_U1/FrameSR[53] ), 
        .CPN(n636), .CDN(n597), .Q(\DesDecoder_U1/FrameSR[54] ) );
  DFCND1 \FIFO_U1/FIFO_SM1/CurState_reg[0]  ( .D(
        \FIFO_U1/FIFO_SM1/NextState [0]), .CP(DecoderParClk), .CDN(n591), .Q(
        n1245), .QN(n528) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[3]  ( .D(\DesDecoder_U1/FrameSR[2] ), 
        .CPN(n636), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[3] ) );
  DFNCND1 \DesDecoder_U1/FrameSR_reg[7]  ( .D(\DesDecoder_U1/FrameSR[6] ), 
        .CPN(n487), .CDN(n602), .Q(\DesDecoder_U1/FrameSR[7] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/MCntr1/Ctr_reg[1]  ( .D(
        \SerialRx_U1/PLL_RxU1/MCntr1/N2 ), .CP(SerialClk), .CDN(n606), .Q(
        \SerialRx_U1/PLL_RxU1/MCntr1/Ctr [1]) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/MCntr1/Ctr_reg[2]  ( .D(
        \SerialRx_U1/PLL_RxU1/MCntr1/N3 ), .CP(SerialClk), .CDN(n607), .Q(
        \SerialRx_U1/PLL_RxU1/MCntr1/Ctr [2]) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/MCntr1/Ctr_reg[3]  ( .D(
        \SerialRx_U1/PLL_RxU1/MCntr1/N4 ), .CP(SerialClk), .CDN(n606), .Q(
        \SerialRx_U1/PLL_RxU1/MCntr1/Ctr [3]) );
  DFSNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[1]  ( .D(n453), .CP(
        \SerialRx_U1/PLL_RxU1/SampleWire ), .SDN(n620), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/MCntr1/Ctr_reg[0]  ( .D(
        \SerialRx_U1/PLL_RxU1/MCntr1/N1 ), .CP(SerialClk), .CDN(n607), .Q(
        \SerialRx_U1/PLL_RxU1/MCntr1/Ctr [0]) );
  EDFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[5]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N55 ), .E(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .CP(\SerialRx_U1/PLL_RxU1/SampleWire ), .CDN(n609), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[5] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/Comp1/AdjustFreq_reg[1]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N20 ), .CP(\SerialRx_U1/PLL_RxU1/CtrCarry ), .CDN(n606), .Q(\SerialRx_U1/PLL_RxU1/AdjFreq [1]) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[5]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N21 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n606), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[5] ) );
  DFNCND1 \DesDecoder_U1/ParValidReg_reg  ( .D(n420), .CPN(n638), .CDN(n591), 
        .Q(n1247) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/Comp1/ClockInN_reg[1]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N6 ), .CP(DecoderParClk), .CDN(n490), .Q(
        \SerialRx_U1/PLL_RxU1/Comp1/ClockInN[1] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/Comp1/ClockInN_reg[0]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N5 ), .CP(DecoderParClk), .CDN(n490), .Q(
        \SerialRx_U1/PLL_RxU1/Comp1/ClockInN[0] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[2]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N18 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n605), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[2] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[3]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N19 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n606), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[3] ) );
  DFCND1 \FIFO_U1/FIFO_SM1/CurState_reg[2]  ( .D(
        \FIFO_U1/FIFO_SM1/NextState [2]), .CP(DecoderParClk), .CDN(n591), .Q(
        n1246), .QN(n529) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[0]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N16 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n605), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[0] ) );
  EDFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[2]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N49 ), .E(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .CP(\SerialRx_U1/PLL_RxU1/SampleWire ), .CDN(n608), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[2] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[1]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N17 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n605), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[1] ) );
  DFCND1 \SerialRx_U1/PLL_RxU1/Comp1/CounterClockN_reg[1]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N8 ), .CP(\SerialRx_U1/PLL_RxU1/CtrCarry ), 
        .CDN(n490), .Q(n1244) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy_reg[4]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N20 ), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n607), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[4] ) );
  EDFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor_reg[3]  ( .D(
        \SerialRx_U1/PLL_RxU1/VFO1/N51 ), .E(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .CP(\SerialRx_U1/PLL_RxU1/SampleWire ), .CDN(n599), .Q(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] ) );
  DFCND1 \SerialRx_U1/PLL_RxU1/Comp1/CounterClockN_reg[0]  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N7 ), .CP(\SerialRx_U1/PLL_RxU1/CtrCarry ), 
        .CDN(n490), .Q(n1243), .QN(\SerialRx_U1/PLL_RxU1/Comp1/N7 ) );
  DFCNQD1 \FIFO_U1/FIFO_SM1/CurState_reg[1]  ( .D(
        \FIFO_U1/FIFO_SM1/NextState [1]), .CP(DecoderParClk), .CDN(n607), .Q(
        \FIFO_U1/FIFO_SM1/CurState[1] ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/MCntr1/Ctr_reg[4]  ( .D(
        \SerialRx_U1/PLL_RxU1/MCntr1/N5 ), .CP(SerialClk), .CDN(n604), .Q(
        \SerialRx_U1/PLL_RxU1/CtrCarry ) );
  DFCNQD1 \SerialRx_U1/PLL_RxU1/VFO1/ClockOutReg_reg  ( .D(n488), .CP(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ), .CDN(n606), .Q(SerialClk) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[0]  ( .D(n452), .CPN(n637), .CDN(n601), 
        .Q(DecodeToFIFO[0]), .QN(n279) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[1]  ( .D(n451), .CPN(n636), .CDN(n598), 
        .Q(DecodeToFIFO[1]), .QN(n278) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[2]  ( .D(n450), .CPN(n487), .CDN(n595), 
        .Q(DecodeToFIFO[2]), .QN(n277) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[3]  ( .D(n449), .CPN(n487), .CDN(n592), 
        .Q(DecodeToFIFO[3]), .QN(n276) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[4]  ( .D(n448), .CPN(n638), .CDN(n591), 
        .Q(DecodeToFIFO[4]), .QN(n275) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[5]  ( .D(n447), .CPN(n637), .CDN(n591), 
        .Q(DecodeToFIFO[5]), .QN(n274) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[6]  ( .D(n446), .CPN(n636), .CDN(n591), 
        .Q(DecodeToFIFO[6]), .QN(n273) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[7]  ( .D(n445), .CPN(n638), .CDN(n591), 
        .Q(DecodeToFIFO[7]), .QN(n272) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[8]  ( .D(n444), .CPN(n637), .CDN(n594), 
        .Q(DecodeToFIFO[8]), .QN(n271) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[9]  ( .D(n443), .CPN(n487), .CDN(n594), 
        .Q(DecodeToFIFO[9]), .QN(n270) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[10]  ( .D(n442), .CPN(n636), .CDN(n594), 
        .Q(DecodeToFIFO[10]), .QN(n269) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[11]  ( .D(n441), .CPN(n638), .CDN(n593), 
        .Q(DecodeToFIFO[11]), .QN(n268) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[12]  ( .D(n440), .CPN(n637), .CDN(n593), 
        .Q(DecodeToFIFO[12]), .QN(n267) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[13]  ( .D(n439), .CPN(n636), .CDN(n593), 
        .Q(DecodeToFIFO[13]), .QN(n266) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[14]  ( .D(n438), .CPN(n487), .CDN(n593), 
        .Q(DecodeToFIFO[14]), .QN(n265) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[15]  ( .D(n437), .CPN(n487), .CDN(n593), 
        .Q(DecodeToFIFO[15]), .QN(n264) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[16]  ( .D(n436), .CPN(n637), .CDN(n593), 
        .Q(DecodeToFIFO[16]), .QN(n263) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[17]  ( .D(n435), .CPN(n638), .CDN(n593), 
        .Q(DecodeToFIFO[17]), .QN(n262) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[18]  ( .D(n434), .CPN(n637), .CDN(n593), 
        .Q(DecodeToFIFO[18]), .QN(n261) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[19]  ( .D(n433), .CPN(n636), .CDN(n593), 
        .Q(DecodeToFIFO[19]), .QN(n260) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[20]  ( .D(n432), .CPN(n637), .CDN(n593), 
        .Q(DecodeToFIFO[20]), .QN(n259) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[21]  ( .D(n431), .CPN(n487), .CDN(n593), 
        .Q(DecodeToFIFO[21]), .QN(n258) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[22]  ( .D(n430), .CPN(n487), .CDN(n592), 
        .Q(DecodeToFIFO[22]), .QN(n257) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[23]  ( .D(n429), .CPN(n638), .CDN(n592), 
        .Q(DecodeToFIFO[23]), .QN(n256) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[24]  ( .D(n428), .CPN(n636), .CDN(n592), 
        .Q(DecodeToFIFO[24]), .QN(n255) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[25]  ( .D(n427), .CPN(n637), .CDN(n592), 
        .Q(DecodeToFIFO[25]), .QN(n254) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[26]  ( .D(n426), .CPN(n638), .CDN(n592), 
        .Q(DecodeToFIFO[26]), .QN(n253) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[27]  ( .D(n425), .CPN(n487), .CDN(n592), 
        .Q(DecodeToFIFO[27]), .QN(n252) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[28]  ( .D(n424), .CPN(n638), .CDN(n592), 
        .Q(DecodeToFIFO[28]), .QN(n251) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[29]  ( .D(n423), .CPN(n637), .CDN(n592), 
        .Q(DecodeToFIFO[29]), .QN(n250) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[30]  ( .D(n422), .CPN(n636), .CDN(n592), 
        .Q(DecodeToFIFO[30]), .QN(n249) );
  DFNCND1 \DesDecoder_U1/ParOutReg_reg[31]  ( .D(n421), .CPN(n487), .CDN(n592), 
        .Q(DecodeToFIFO[31]), .QN(n248) );
  DFCNQD1 ParValidReg_reg ( .D(N35), .CP(ParOutClk), .CDN(n606), .Q(ParValid)
         );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[31]) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[30]) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[29]) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[28]) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[27]) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[26]) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[25]) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[24]) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[23]) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[22]) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n605), .Q(
        ParOut[21]) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[20]) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[19]) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[18]) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[17]) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n603), .Q(
        ParOut[16]) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[15]) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n606), .Q(
        ParOut[14]) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[13]) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[12]) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[11]) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n604), .Q(
        ParOut[10]) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n604), .Q(ParOut[9])
         );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n604), .Q(ParOut[8])
         );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n604), .Q(ParOut[7])
         );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n605), .Q(ParOut[6])
         );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n605), .Q(ParOut[5])
         );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n606), .Q(ParOut[4])
         );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n606), .Q(ParOut[3])
         );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n603), .Q(ParOut[2])
         );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n606), .Q(ParOut[1])
         );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n603), .Q(ParOut[0])
         );
  DFSND1 \SerialRx_U1/PLL_RxU1/Comp1/ZeroCounters_reg  ( .D(
        \SerialRx_U1/PLL_RxU1/Comp1/N9 ), .CP(DecoderParClk), .SDN(n619), .QN(
        n490) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[31]  ( .D(\FIFO_U1/RegFile1/N82 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n668), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/N2330 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[30]  ( .D(\FIFO_U1/RegFile1/N83 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n682), .CDN(n598), .Q(
        \FIFO_U1/RegFile1/N2333 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[29]  ( .D(\FIFO_U1/RegFile1/N84 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n597), .Q(
        \FIFO_U1/RegFile1/N2336 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[28]  ( .D(\FIFO_U1/RegFile1/N85 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n681), .CDN(n599), .Q(
        \FIFO_U1/RegFile1/N2339 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[27]  ( .D(\FIFO_U1/RegFile1/N86 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/N2342 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[26]  ( .D(\FIFO_U1/RegFile1/N87 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n680), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/N2345 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[25]  ( .D(\FIFO_U1/RegFile1/N88 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n621), .Q(
        \FIFO_U1/RegFile1/N2348 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[24]  ( .D(\FIFO_U1/RegFile1/N89 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n695), .CDN(n592), .Q(
        \FIFO_U1/RegFile1/N2351 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[23]  ( .D(\FIFO_U1/RegFile1/N90 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n620), .Q(
        \FIFO_U1/RegFile1/N2354 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[22]  ( .D(\FIFO_U1/RegFile1/N91 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n670), .CDN(n595), .Q(
        \FIFO_U1/RegFile1/N2357 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[21]  ( .D(\FIFO_U1/RegFile1/N92 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n596), .Q(
        \FIFO_U1/RegFile1/N2360 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[20]  ( .D(\FIFO_U1/RegFile1/N93 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n671), .CDN(n625), .Q(
        \FIFO_U1/RegFile1/N2363 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[19]  ( .D(\FIFO_U1/RegFile1/N94 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n630), .Q(
        \FIFO_U1/RegFile1/N2366 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[18]  ( .D(\FIFO_U1/RegFile1/N95 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n667), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/N2369 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[17]  ( .D(\FIFO_U1/RegFile1/N96 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n624), .Q(
        \FIFO_U1/RegFile1/N2372 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[16]  ( .D(\FIFO_U1/RegFile1/N97 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/N2375 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[15]  ( .D(\FIFO_U1/RegFile1/N98 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n602), .Q(
        \FIFO_U1/RegFile1/N2378 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[14]  ( .D(\FIFO_U1/RegFile1/N99 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n677), .CDN(n603), .Q(
        \FIFO_U1/RegFile1/N2381 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[13]  ( .D(\FIFO_U1/RegFile1/N100 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n609), .Q(
        \FIFO_U1/RegFile1/N2384 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[12]  ( .D(\FIFO_U1/RegFile1/N101 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n688), .CDN(n604), .Q(
        \FIFO_U1/RegFile1/N2387 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[11]  ( .D(\FIFO_U1/RegFile1/N102 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n666), .CDN(n608), .Q(
        \FIFO_U1/RegFile1/N2390 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[10]  ( .D(\FIFO_U1/RegFile1/N103 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n678), .CDN(n606), .Q(
        \FIFO_U1/RegFile1/N2393 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[9]  ( .D(\FIFO_U1/RegFile1/N104 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n674), .CDN(n611), .Q(
        \FIFO_U1/RegFile1/N2396 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[8]  ( .D(\FIFO_U1/RegFile1/N105 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n673), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/N2399 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[7]  ( .D(\FIFO_U1/RegFile1/N106 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n689), .CDN(n615), .Q(
        \FIFO_U1/RegFile1/N2402 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[6]  ( .D(\FIFO_U1/RegFile1/N107 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n691), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/N2405 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[5]  ( .D(\FIFO_U1/RegFile1/N108 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n694), .CDN(n593), .Q(
        \FIFO_U1/RegFile1/N2408 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[4]  ( .D(\FIFO_U1/RegFile1/N109 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n693), .CDN(n612), .Q(
        \FIFO_U1/RegFile1/N2411 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[3]  ( .D(\FIFO_U1/RegFile1/N110 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n675), .CDN(n610), .Q(
        \FIFO_U1/RegFile1/N2414 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[2]  ( .D(\FIFO_U1/RegFile1/N111 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n671), .CDN(n631), .Q(
        \FIFO_U1/RegFile1/N2417 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[1]  ( .D(\FIFO_U1/RegFile1/N112 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n685), .CDN(n627), .Q(
        \FIFO_U1/RegFile1/N2420 ) );
  EDFCNQD1 \FIFO_U1/RegFile1/DataOreg_reg[0]  ( .D(\FIFO_U1/RegFile1/N113 ), 
        .E(\FIFO_U1/RegFile1/N2327 ), .CP(n690), .CDN(n607), .Q(
        \FIFO_U1/RegFile1/N2423 ) );
  LHCND1 \DesDecoder_U1/SerClock_reg  ( .E(SerValid), .D(SerialClk), .CDN(n620), .Q(n487) );
  INVD3 U403 ( .I(n527), .ZN(\FIFO_U1/RegFile1/N2327 ) );
  OA21D1 U404 ( .A1(n1148), .A2(n1149), .B(n1150), .Z(n527) );
  INVD1 U405 ( .I(n1150), .ZN(\FIFO_U1/RegFile1/N2328 ) );
  NR2D2P5 U406 ( .A1(n1152), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1734 ) );
  ND3D1 U407 ( .A1(n1163), .A2(\FIFO_U1/RegFile1/N78 ), .A3(
        \FIFO_U1/RegFile1/N2328 ), .ZN(n1162) );
  NR2D2P5 U408 ( .A1(n1159), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1767 ) );
  ND3D1 U409 ( .A1(n1161), .A2(\FIFO_U1/RegFile1/N79 ), .A3(
        \FIFO_U1/RegFile1/N2328 ), .ZN(n1160) );
  NR2D2P5 U410 ( .A1(n1153), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1701 ) );
  NR2D2P5 U411 ( .A1(n1158), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1800 ) );
  NR2D2P5 U412 ( .A1(n1154), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1668 ) );
  NR2D2P5 U413 ( .A1(n1157), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1833 ) );
  NR2D2P5 U414 ( .A1(n1155), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1635 ) );
  NR2D2P5 U415 ( .A1(n1156), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1866 ) );
  NR2D2P5 U416 ( .A1(n1156), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1602 ) );
  NR2D2P5 U417 ( .A1(n1155), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1899 ) );
  NR2D2P5 U418 ( .A1(n1157), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1569 ) );
  NR2D2P5 U419 ( .A1(n1154), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1932 ) );
  NR2D2P5 U420 ( .A1(n1158), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1536 ) );
  NR2D2P5 U421 ( .A1(n1153), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1965 ) );
  NR2D2P5 U422 ( .A1(n1159), .A2(n1162), .ZN(\FIFO_U1/RegFile1/N1503 ) );
  NR2D2P5 U423 ( .A1(n1152), .A2(n1160), .ZN(\FIFO_U1/RegFile1/N1998 ) );
  NR2D2P5 U424 ( .A1(n1152), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1470 ) );
  ND3D1 U425 ( .A1(n1161), .A2(n1163), .A3(\FIFO_U1/RegFile1/N2328 ), .ZN(
        n1164) );
  NR2D2P5 U426 ( .A1(n1151), .A2(n1159), .ZN(\FIFO_U1/RegFile1/N2031 ) );
  ND3D1 U427 ( .A1(\FIFO_U1/RegFile1/N78 ), .A2(\FIFO_U1/RegFile1/N79 ), .A3(
        \FIFO_U1/RegFile1/N2328 ), .ZN(n1151) );
  NR2D2P5 U428 ( .A1(n1153), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1437 ) );
  NR2D2P5 U429 ( .A1(n1151), .A2(n1158), .ZN(\FIFO_U1/RegFile1/N2064 ) );
  NR2D2P5 U430 ( .A1(n1154), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1404 ) );
  NR2D2P5 U431 ( .A1(n1151), .A2(n1157), .ZN(\FIFO_U1/RegFile1/N2097 ) );
  NR2D2P5 U432 ( .A1(n1155), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1371 ) );
  NR2D2P5 U433 ( .A1(n1151), .A2(n1156), .ZN(\FIFO_U1/RegFile1/N2130 ) );
  NR2D2P5 U434 ( .A1(n1156), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1338 ) );
  NR2D2P5 U435 ( .A1(n1151), .A2(n1155), .ZN(\FIFO_U1/RegFile1/N2163 ) );
  NR2D2P5 U436 ( .A1(n1157), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1305 ) );
  NR2D2P5 U437 ( .A1(n1151), .A2(n1154), .ZN(\FIFO_U1/RegFile1/N2196 ) );
  NR2D2P5 U438 ( .A1(n1158), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1272 ) );
  ND3D1 U439 ( .A1(n1166), .A2(n564), .A3(n649), .ZN(n1158) );
  NR2D2P5 U440 ( .A1(n1151), .A2(n1153), .ZN(\FIFO_U1/RegFile1/N2229 ) );
  NR2D2P5 U441 ( .A1(n1159), .A2(n1164), .ZN(\FIFO_U1/RegFile1/N1239 ) );
  NR2D2P5 U442 ( .A1(n1151), .A2(n1152), .ZN(\FIFO_U1/RegFile1/N2262 ) );
  AOI211XD4 U443 ( .A1(\FIFO_U1/SM_MemWriteCmd ), .A2(\FIFO_U1/SM_MemReadCmd ), 
        .B(FIFOFull), .C(FIFOEmpty), .ZN(n419) );
  INVD3 U444 ( .I(n1161), .ZN(\FIFO_U1/RegFile1/N78 ) );
  INVD0 U445 ( .I(n419), .ZN(n1149) );
  IAO21D1 U446 ( .A1(n1174), .A2(n1175), .B(DecoderParClk), .ZN(
        \FIFO_U1/FIFO_SM1/N198 ) );
  IND3D1 U447 ( .A1(n1181), .B1(n1177), .B2(n1182), .ZN(n1174) );
  INVD1 U448 ( .I(FIFOReadCmd), .ZN(n1147) );
  AOI21D1 U449 ( .A1(n1170), .A2(n1115), .B(DecoderParClk), .ZN(
        \FIFO_U1/FIFO_SM1/N209 ) );
  MUX2ND2 U450 ( .I0(n1118), .I1(n1116), .S(n1167), .ZN(\FIFO_U1/RegFile1/N79 ) );
  INR2XD2 U451 ( .A1(n1230), .B1(n1231), .ZN(\DesDecoder_U1/N44 ) );
  AN4D1 U452 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .Z(n1230) );
  BUFFD1 U453 ( .I(n674), .Z(n678) );
  BUFFD1 U454 ( .I(n686), .Z(n676) );
  BUFFD1 U455 ( .I(n689), .Z(n671) );
  BUFFD1 U456 ( .I(n688), .Z(n672) );
  BUFFD1 U457 ( .I(n686), .Z(n679) );
  BUFFD1 U458 ( .I(n685), .Z(n680) );
  BUFFD1 U459 ( .I(n686), .Z(n677) );
  BUFFD1 U460 ( .I(n688), .Z(n673) );
  BUFFD1 U461 ( .I(n687), .Z(n674) );
  BUFFD1 U462 ( .I(n687), .Z(n675) );
  BUFFD1 U463 ( .I(n685), .Z(n681) );
  BUFFD1 U464 ( .I(n684), .Z(n682) );
  BUFFD1 U465 ( .I(n684), .Z(n683) );
  BUFFD1 U466 ( .I(n690), .Z(n669) );
  BUFFD1 U467 ( .I(n689), .Z(n670) );
  BUFFD1 U468 ( .I(n691), .Z(n666) );
  BUFFD1 U469 ( .I(n691), .Z(n667) );
  BUFFD1 U470 ( .I(n690), .Z(n668) );
  BUFFD1 U471 ( .I(n693), .Z(n686) );
  BUFFD1 U472 ( .I(n693), .Z(n688) );
  BUFFD1 U473 ( .I(n693), .Z(n687) );
  BUFFD1 U474 ( .I(n694), .Z(n685) );
  BUFFD1 U475 ( .I(n694), .Z(n684) );
  BUFFD1 U476 ( .I(n692), .Z(n689) );
  BUFFD1 U477 ( .I(n692), .Z(n691) );
  BUFFD1 U478 ( .I(n692), .Z(n690) );
  BUFFD1 U479 ( .I(n695), .Z(n693) );
  BUFFD1 U480 ( .I(n669), .Z(n694) );
  BUFFD1 U481 ( .I(n695), .Z(n692) );
  INVD1 U482 ( .I(n564), .ZN(n661) );
  BUFFD1 U483 ( .I(n629), .Z(n593) );
  BUFFD1 U484 ( .I(n629), .Z(n592) );
  BUFFD1 U485 ( .I(n629), .Z(n594) );
  BUFFD1 U486 ( .I(n629), .Z(n595) );
  BUFFD1 U487 ( .I(n628), .Z(n596) );
  BUFFD1 U488 ( .I(n628), .Z(n597) );
  BUFFD1 U489 ( .I(n628), .Z(n598) );
  BUFFD1 U490 ( .I(n628), .Z(n599) );
  BUFFD1 U491 ( .I(n627), .Z(n600) );
  BUFFD1 U492 ( .I(n627), .Z(n601) );
  BUFFD1 U493 ( .I(n627), .Z(n602) );
  BUFFD1 U494 ( .I(n627), .Z(n603) );
  BUFFD1 U495 ( .I(n626), .Z(n605) );
  BUFFD1 U496 ( .I(n626), .Z(n606) );
  BUFFD1 U497 ( .I(n626), .Z(n604) );
  BUFFD1 U498 ( .I(n626), .Z(n607) );
  BUFFD1 U499 ( .I(n622), .Z(n620) );
  BUFFD1 U500 ( .I(n622), .Z(n619) );
  BUFFD1 U501 ( .I(n623), .Z(n615) );
  BUFFD1 U502 ( .I(n625), .Z(n610) );
  BUFFD1 U503 ( .I(n625), .Z(n611) );
  BUFFD1 U504 ( .I(n623), .Z(n616) );
  BUFFD1 U505 ( .I(n623), .Z(n617) );
  BUFFD1 U506 ( .I(n622), .Z(n618) );
  BUFFD1 U507 ( .I(n615), .Z(n614) );
  BUFFD1 U508 ( .I(n625), .Z(n608) );
  BUFFD1 U509 ( .I(n625), .Z(n609) );
  BUFFD1 U510 ( .I(n624), .Z(n612) );
  BUFFD1 U511 ( .I(n624), .Z(n613) );
  BUFFD1 U512 ( .I(n649), .Z(n646) );
  BUFFD1 U513 ( .I(n647), .Z(n645) );
  BUFFD1 U514 ( .I(n648), .Z(n644) );
  BUFFD1 U515 ( .I(n648), .Z(n643) );
  BUFFD1 U516 ( .I(n649), .Z(n642) );
  BUFFD1 U517 ( .I(n649), .Z(n641) );
  BUFFD1 U518 ( .I(n650), .Z(n640) );
  BUFFD1 U519 ( .I(n650), .Z(n639) );
  BUFFD1 U520 ( .I(n657), .Z(n656) );
  BUFFD1 U521 ( .I(n659), .Z(n653) );
  BUFFD1 U522 ( .I(n658), .Z(n654) );
  BUFFD1 U523 ( .I(n659), .Z(n652) );
  BUFFD1 U524 ( .I(n658), .Z(n655) );
  BUFFD1 U525 ( .I(n622), .Z(n621) );
  BUFFD1 U526 ( .I(n696), .Z(n695) );
  INVD1 U527 ( .I(n564), .ZN(n663) );
  INVD1 U528 ( .I(n564), .ZN(n662) );
  INVD1 U529 ( .I(n564), .ZN(n664) );
  INVD1 U530 ( .I(n564), .ZN(n665) );
  BUFFD1 U531 ( .I(n630), .Z(n591) );
  BUFFD1 U532 ( .I(n631), .Z(n630) );
  BUFFD1 U533 ( .I(n649), .Z(n647) );
  BUFFD1 U534 ( .I(n651), .Z(n648) );
  BUFFD1 U535 ( .I(n651), .Z(n649) );
  BUFFD1 U536 ( .I(n660), .Z(n659) );
  BUFFD1 U537 ( .I(n660), .Z(n658) );
  BUFFD1 U538 ( .I(n651), .Z(n650) );
  BUFFD1 U539 ( .I(n660), .Z(n657) );
  BUFFD1 U540 ( .I(n634), .Z(n623) );
  BUFFD1 U541 ( .I(n633), .Z(n625) );
  BUFFD1 U542 ( .I(n602), .Z(n624) );
  BUFFD1 U543 ( .I(n631), .Z(n629) );
  BUFFD1 U544 ( .I(n632), .Z(n628) );
  BUFFD1 U545 ( .I(n632), .Z(n627) );
  BUFFD1 U546 ( .I(n634), .Z(n622) );
  BUFFD1 U547 ( .I(n633), .Z(n626) );
  BUFFD1 U548 ( .I(\FIFO_U1/RegFile1/ChipClock ), .Z(n696) );
  BUFFD1 U549 ( .I(\FIFO_U1/RegFile1/N75 ), .Z(n651) );
  BUFFD1 U550 ( .I(\FIFO_U1/RegFile1/N76 ), .Z(n660) );
  BUFFD1 U551 ( .I(n635), .Z(n631) );
  BUFFD1 U552 ( .I(n635), .Z(n632) );
  BUFFD1 U553 ( .I(n626), .Z(n634) );
  BUFFD1 U554 ( .I(n635), .Z(n633) );
  MUX2D0 U555 ( .I0(n1122), .I1(n1121), .S(n1167), .Z(n564) );
  BUFFD1 U556 ( .I(n491), .Z(n635) );
  MUX4ND0 U557 ( .I0(\FIFO_U1/RegFile1/Storage[28][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][0] ), .S0(n646), .S1(n658), .ZN(n700) );
  MUX4ND0 U558 ( .I0(\FIFO_U1/RegFile1/Storage[28][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][1] ), .S0(n651), .S1(n657), .ZN(n713) );
  MUX4ND0 U559 ( .I0(\FIFO_U1/RegFile1/Storage[28][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][2] ), .S0(n650), .S1(n656), .ZN(n726) );
  MUX4ND0 U560 ( .I0(\FIFO_U1/RegFile1/Storage[28][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][3] ), .S0(n641), .S1(n659), .ZN(n739) );
  MUX4ND0 U561 ( .I0(\FIFO_U1/RegFile1/Storage[28][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][4] ), .S0(n648), .S1(n653), .ZN(n752) );
  MUX4ND0 U562 ( .I0(\FIFO_U1/RegFile1/Storage[28][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][5] ), .S0(n649), .S1(n660), .ZN(n765) );
  MUX4ND0 U563 ( .I0(\FIFO_U1/RegFile1/Storage[28][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][6] ), .S0(n651), .S1(n652), .ZN(n778) );
  MUX4ND0 U564 ( .I0(\FIFO_U1/RegFile1/Storage[28][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][7] ), .S0(n651), .S1(n653), .ZN(n791) );
  MUX4ND0 U565 ( .I0(\FIFO_U1/RegFile1/Storage[28][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][8] ), .S0(n644), .S1(n660), .ZN(n804) );
  MUX4ND0 U566 ( .I0(\FIFO_U1/RegFile1/Storage[28][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][9] ), .S0(n647), .S1(n652), .ZN(n817) );
  MUX4ND0 U567 ( .I0(\FIFO_U1/RegFile1/Storage[28][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][10] ), .S0(n645), .S1(n657), .ZN(n830)
         );
  MUX4ND0 U568 ( .I0(\FIFO_U1/RegFile1/Storage[28][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][11] ), .S0(n650), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n843) );
  MUX4ND0 U569 ( .I0(\FIFO_U1/RegFile1/Storage[28][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][12] ), .S0(n641), .S1(n653), .ZN(n856)
         );
  MUX4ND0 U570 ( .I0(\FIFO_U1/RegFile1/Storage[28][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][13] ), .S0(n644), .S1(n657), .ZN(n869)
         );
  MUX4ND0 U571 ( .I0(\FIFO_U1/RegFile1/Storage[28][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][14] ), .S0(n644), .S1(n658), .ZN(n882)
         );
  MUX4ND0 U572 ( .I0(\FIFO_U1/RegFile1/Storage[28][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][15] ), .S0(n647), .S1(n659), .ZN(n895)
         );
  MUX4ND0 U573 ( .I0(\FIFO_U1/RegFile1/Storage[28][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][16] ), .S0(n648), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n908) );
  MUX4ND0 U574 ( .I0(\FIFO_U1/RegFile1/Storage[28][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][17] ), .S0(n646), .S1(n657), .ZN(n921)
         );
  MUX4ND0 U575 ( .I0(\FIFO_U1/RegFile1/Storage[28][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][18] ), .S0(n650), .S1(n654), .ZN(n934)
         );
  MUX4ND0 U576 ( .I0(\FIFO_U1/RegFile1/Storage[28][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][19] ), .S0(n648), .S1(n660), .ZN(n947)
         );
  MUX4ND0 U577 ( .I0(\FIFO_U1/RegFile1/Storage[28][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][20] ), .S0(n650), .S1(n654), .ZN(n960)
         );
  MUX4ND0 U578 ( .I0(\FIFO_U1/RegFile1/Storage[28][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][21] ), .S0(\FIFO_U1/RegFile1/N75 ), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n973) );
  MUX4ND0 U579 ( .I0(\FIFO_U1/RegFile1/Storage[28][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][22] ), .S0(n651), .S1(n655), .ZN(n986)
         );
  MUX4ND0 U580 ( .I0(\FIFO_U1/RegFile1/Storage[28][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][23] ), .S0(n649), .S1(n655), .ZN(n999)
         );
  MUX4ND0 U581 ( .I0(\FIFO_U1/RegFile1/Storage[28][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][24] ), .S0(n648), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n1012) );
  MUX4ND0 U582 ( .I0(\FIFO_U1/RegFile1/Storage[28][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][25] ), .S0(n645), .S1(n657), .ZN(n1025)
         );
  MUX4ND0 U583 ( .I0(\FIFO_U1/RegFile1/Storage[28][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][26] ), .S0(n646), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n1038) );
  MUX4ND0 U584 ( .I0(\FIFO_U1/RegFile1/Storage[28][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][27] ), .S0(n649), .S1(
        \FIFO_U1/RegFile1/N76 ), .ZN(n1051) );
  MUX4ND0 U585 ( .I0(\FIFO_U1/RegFile1/Storage[28][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][28] ), .S0(n645), .S1(n660), .ZN(n1064)
         );
  MUX4ND0 U586 ( .I0(\FIFO_U1/RegFile1/Storage[28][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][29] ), .S0(n648), .S1(n660), .ZN(n1077)
         );
  MUX4ND0 U587 ( .I0(\FIFO_U1/RegFile1/Storage[28][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][30] ), .S0(n649), .S1(n652), .ZN(n1090)
         );
  MUX4ND0 U588 ( .I0(\FIFO_U1/RegFile1/Storage[28][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[29][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[30][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[31][31] ), .S0(n644), .S1(n655), .ZN(n1103)
         );
  MUX4D0 U589 ( .I0(\FIFO_U1/RegFile1/Storage[20][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][0] ), .S0(n644), .S1(n660), .Z(n701) );
  MUX4D0 U590 ( .I0(\FIFO_U1/RegFile1/Storage[20][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][1] ), .S0(n646), .S1(n656), .Z(n714) );
  MUX4D0 U591 ( .I0(\FIFO_U1/RegFile1/Storage[20][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][2] ), .S0(n646), .S1(n657), .Z(n727) );
  MUX4D0 U592 ( .I0(\FIFO_U1/RegFile1/Storage[20][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][3] ), .S0(n650), .S1(n652), .Z(n740) );
  MUX4D0 U593 ( .I0(\FIFO_U1/RegFile1/Storage[20][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][4] ), .S0(n639), .S1(n656), .Z(n753) );
  MUX4D0 U594 ( .I0(\FIFO_U1/RegFile1/Storage[20][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][5] ), .S0(n649), .S1(n659), .Z(n766) );
  MUX4D0 U595 ( .I0(\FIFO_U1/RegFile1/Storage[20][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][6] ), .S0(n648), .S1(n658), .Z(n779) );
  MUX4D0 U596 ( .I0(\FIFO_U1/RegFile1/Storage[20][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][7] ), .S0(\FIFO_U1/RegFile1/N75 ), .S1(
        n656), .Z(n792) );
  MUX4D0 U597 ( .I0(\FIFO_U1/RegFile1/Storage[20][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][8] ), .S0(n648), .S1(n660), .Z(n805) );
  MUX4D0 U598 ( .I0(\FIFO_U1/RegFile1/Storage[20][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][9] ), .S0(n648), .S1(n658), .Z(n818) );
  MUX4D0 U599 ( .I0(\FIFO_U1/RegFile1/Storage[20][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][10] ), .S0(n645), .S1(n653), .Z(n831) );
  MUX4D0 U600 ( .I0(\FIFO_U1/RegFile1/Storage[20][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][11] ), .S0(n645), .S1(n659), .Z(n844) );
  MUX4D0 U601 ( .I0(\FIFO_U1/RegFile1/Storage[20][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][12] ), .S0(n646), .S1(n657), .Z(n857) );
  MUX4D0 U602 ( .I0(\FIFO_U1/RegFile1/Storage[20][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][13] ), .S0(n640), .S1(n659), .Z(n870) );
  MUX4D0 U603 ( .I0(\FIFO_U1/RegFile1/Storage[20][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][14] ), .S0(n651), .S1(n658), .Z(n883) );
  MUX4D0 U604 ( .I0(\FIFO_U1/RegFile1/Storage[20][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][15] ), .S0(n647), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n896) );
  MUX4D0 U605 ( .I0(\FIFO_U1/RegFile1/Storage[20][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][16] ), .S0(n639), .S1(n659), .Z(n909) );
  MUX4D0 U606 ( .I0(\FIFO_U1/RegFile1/Storage[20][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][17] ), .S0(n648), .S1(n654), .Z(n922) );
  MUX4D0 U607 ( .I0(\FIFO_U1/RegFile1/Storage[20][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][18] ), .S0(n645), .S1(n653), .Z(n935) );
  MUX4D0 U608 ( .I0(\FIFO_U1/RegFile1/Storage[20][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][19] ), .S0(n645), .S1(n657), .Z(n948) );
  MUX4D0 U609 ( .I0(\FIFO_U1/RegFile1/Storage[20][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][20] ), .S0(n646), .S1(n659), .Z(n961) );
  MUX4D0 U610 ( .I0(\FIFO_U1/RegFile1/Storage[20][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][21] ), .S0(n644), .S1(n659), .Z(n974) );
  MUX4D0 U611 ( .I0(\FIFO_U1/RegFile1/Storage[20][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][22] ), .S0(n644), .S1(n653), .Z(n987) );
  MUX4D0 U612 ( .I0(\FIFO_U1/RegFile1/Storage[20][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][23] ), .S0(n643), .S1(n652), .Z(n1000)
         );
  MUX4D0 U613 ( .I0(\FIFO_U1/RegFile1/Storage[20][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][24] ), .S0(n643), .S1(n652), .Z(n1013)
         );
  MUX4D0 U614 ( .I0(\FIFO_U1/RegFile1/Storage[20][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][25] ), .S0(n642), .S1(n653), .Z(n1026)
         );
  MUX4D0 U615 ( .I0(\FIFO_U1/RegFile1/Storage[20][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][26] ), .S0(n642), .S1(n653), .Z(n1039)
         );
  MUX4D0 U616 ( .I0(\FIFO_U1/RegFile1/Storage[20][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][27] ), .S0(n641), .S1(n654), .Z(n1052)
         );
  MUX4D0 U617 ( .I0(\FIFO_U1/RegFile1/Storage[20][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][28] ), .S0(n641), .S1(n654), .Z(n1065)
         );
  MUX4D0 U618 ( .I0(\FIFO_U1/RegFile1/Storage[20][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][29] ), .S0(n640), .S1(n655), .Z(n1078)
         );
  MUX4D0 U619 ( .I0(\FIFO_U1/RegFile1/Storage[20][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][30] ), .S0(n640), .S1(n655), .Z(n1091)
         );
  MUX4D0 U620 ( .I0(\FIFO_U1/RegFile1/Storage[20][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[21][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[22][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[23][31] ), .S0(n639), .S1(n658), .Z(n1104)
         );
  MUX4D0 U621 ( .I0(\FIFO_U1/RegFile1/Storage[12][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][0] ), .S0(n647), .S1(n656), .Z(n703) );
  MUX4D0 U622 ( .I0(\FIFO_U1/RegFile1/Storage[4][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][0] ), .S0(n646), .S1(n656), .Z(n705) );
  MUX4D0 U623 ( .I0(\FIFO_U1/RegFile1/Storage[12][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][1] ), .S0(n646), .S1(n656), .Z(n716) );
  MUX4D0 U624 ( .I0(\FIFO_U1/RegFile1/Storage[4][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][1] ), .S0(n646), .S1(n656), .Z(n718) );
  MUX4D0 U625 ( .I0(\FIFO_U1/RegFile1/Storage[12][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][2] ), .S0(n646), .S1(n660), .Z(n729) );
  MUX4D0 U626 ( .I0(\FIFO_U1/RegFile1/Storage[4][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][2] ), .S0(n640), .S1(n654), .Z(n731) );
  MUX4D0 U627 ( .I0(\FIFO_U1/RegFile1/Storage[12][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][3] ), .S0(n641), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n742) );
  MUX4D0 U628 ( .I0(\FIFO_U1/RegFile1/Storage[4][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][3] ), .S0(n642), .S1(n653), .Z(n744) );
  MUX4D0 U629 ( .I0(\FIFO_U1/RegFile1/Storage[12][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][4] ), .S0(n647), .S1(n657), .Z(n755) );
  MUX4D0 U630 ( .I0(\FIFO_U1/RegFile1/Storage[4][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][4] ), .S0(n649), .S1(n659), .Z(n757) );
  MUX4D0 U631 ( .I0(\FIFO_U1/RegFile1/Storage[12][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][5] ), .S0(n651), .S1(n660), .Z(n768) );
  MUX4D0 U632 ( .I0(\FIFO_U1/RegFile1/Storage[4][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][5] ), .S0(n639), .S1(n653), .Z(n770) );
  MUX4D0 U633 ( .I0(\FIFO_U1/RegFile1/Storage[12][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][6] ), .S0(n640), .S1(n657), .Z(n781) );
  MUX4D0 U634 ( .I0(\FIFO_U1/RegFile1/Storage[4][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][6] ), .S0(n651), .S1(n659), .Z(n783) );
  MUX4D0 U635 ( .I0(\FIFO_U1/RegFile1/Storage[12][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][7] ), .S0(n649), .S1(n658), .Z(n794) );
  MUX4D0 U636 ( .I0(\FIFO_U1/RegFile1/Storage[4][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][7] ), .S0(n650), .S1(n660), .Z(n796) );
  MUX4D0 U637 ( .I0(\FIFO_U1/RegFile1/Storage[12][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][8] ), .S0(n648), .S1(n653), .Z(n807) );
  MUX4D0 U638 ( .I0(\FIFO_U1/RegFile1/Storage[4][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][8] ), .S0(n649), .S1(n653), .Z(n809) );
  MUX4D0 U639 ( .I0(\FIFO_U1/RegFile1/Storage[12][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][9] ), .S0(n642), .S1(n660), .Z(n820) );
  MUX4D0 U640 ( .I0(\FIFO_U1/RegFile1/Storage[4][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][9] ), .S0(n650), .S1(n659), .Z(n822) );
  MUX4D0 U641 ( .I0(\FIFO_U1/RegFile1/Storage[12][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][10] ), .S0(n643), .S1(n655), .Z(n833) );
  MUX4D0 U642 ( .I0(\FIFO_U1/RegFile1/Storage[4][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][10] ), .S0(n647), .S1(n658), .Z(n835) );
  MUX4D0 U643 ( .I0(\FIFO_U1/RegFile1/Storage[12][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][11] ), .S0(n649), .S1(n654), .Z(n846) );
  MUX4D0 U644 ( .I0(\FIFO_U1/RegFile1/Storage[4][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][11] ), .S0(n645), .S1(n658), .Z(n848) );
  MUX4D0 U645 ( .I0(\FIFO_U1/RegFile1/Storage[12][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][12] ), .S0(n644), .S1(n660), .Z(n859) );
  MUX4D0 U646 ( .I0(\FIFO_U1/RegFile1/Storage[4][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][12] ), .S0(n643), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n861) );
  MUX4D0 U647 ( .I0(\FIFO_U1/RegFile1/Storage[12][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][13] ), .S0(n642), .S1(n657), .Z(n872) );
  MUX4D0 U648 ( .I0(\FIFO_U1/RegFile1/Storage[4][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][13] ), .S0(n639), .S1(n656), .Z(n874) );
  MUX4D0 U649 ( .I0(\FIFO_U1/RegFile1/Storage[12][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][14] ), .S0(n641), .S1(n654), .Z(n885) );
  MUX4D0 U650 ( .I0(\FIFO_U1/RegFile1/Storage[4][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][14] ), .S0(n642), .S1(n656), .Z(n887) );
  MUX4D0 U651 ( .I0(\FIFO_U1/RegFile1/Storage[12][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][15] ), .S0(n643), .S1(n658), .Z(n898) );
  MUX4D0 U652 ( .I0(\FIFO_U1/RegFile1/Storage[4][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][15] ), .S0(n650), .S1(n657), .Z(n900) );
  MUX4D0 U653 ( .I0(\FIFO_U1/RegFile1/Storage[12][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][16] ), .S0(n646), .S1(n656), .Z(n911) );
  MUX4D0 U654 ( .I0(\FIFO_U1/RegFile1/Storage[4][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][16] ), .S0(n643), .S1(n660), .Z(n913) );
  MUX4D0 U655 ( .I0(\FIFO_U1/RegFile1/Storage[12][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][17] ), .S0(n645), .S1(n655), .Z(n924) );
  MUX4D0 U656 ( .I0(\FIFO_U1/RegFile1/Storage[4][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][17] ), .S0(n645), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n926) );
  MUX4D0 U657 ( .I0(\FIFO_U1/RegFile1/Storage[12][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][18] ), .S0(n645), .S1(n660), .Z(n937) );
  MUX4D0 U658 ( .I0(\FIFO_U1/RegFile1/Storage[4][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][18] ), .S0(n645), .S1(n652), .Z(n939) );
  MUX4D0 U659 ( .I0(\FIFO_U1/RegFile1/Storage[12][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][19] ), .S0(n649), .S1(n652), .Z(n950) );
  MUX4D0 U660 ( .I0(\FIFO_U1/RegFile1/Storage[4][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][19] ), .S0(n641), .S1(n656), .Z(n952) );
  MUX4D0 U661 ( .I0(\FIFO_U1/RegFile1/Storage[12][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][20] ), .S0(n642), .S1(n659), .Z(n963) );
  MUX4D0 U662 ( .I0(\FIFO_U1/RegFile1/Storage[4][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][20] ), .S0(n639), .S1(n658), .Z(n965) );
  MUX4D0 U663 ( .I0(\FIFO_U1/RegFile1/Storage[12][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][21] ), .S0(n644), .S1(n654), .Z(n976) );
  MUX4D0 U664 ( .I0(\FIFO_U1/RegFile1/Storage[4][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][21] ), .S0(n644), .S1(n658), .Z(n978) );
  MUX4D0 U665 ( .I0(\FIFO_U1/RegFile1/Storage[12][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][22] ), .S0(n644), .S1(n656), .Z(n989) );
  MUX4D0 U666 ( .I0(\FIFO_U1/RegFile1/Storage[4][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][22] ), .S0(n644), .S1(n654), .Z(n991) );
  MUX4D0 U667 ( .I0(\FIFO_U1/RegFile1/Storage[12][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][23] ), .S0(n643), .S1(n652), .Z(n1002)
         );
  MUX4D0 U668 ( .I0(\FIFO_U1/RegFile1/Storage[4][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][23] ), .S0(n643), .S1(n652), .Z(n1004) );
  MUX4D0 U669 ( .I0(\FIFO_U1/RegFile1/Storage[12][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][24] ), .S0(n643), .S1(n652), .Z(n1015)
         );
  MUX4D0 U670 ( .I0(\FIFO_U1/RegFile1/Storage[4][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][24] ), .S0(n642), .S1(n653), .Z(n1017) );
  MUX4D0 U671 ( .I0(\FIFO_U1/RegFile1/Storage[12][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][25] ), .S0(n642), .S1(n653), .Z(n1028)
         );
  MUX4D0 U672 ( .I0(\FIFO_U1/RegFile1/Storage[4][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][25] ), .S0(n642), .S1(n653), .Z(n1030) );
  MUX4D0 U673 ( .I0(\FIFO_U1/RegFile1/Storage[12][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][26] ), .S0(n642), .S1(n653), .Z(n1041)
         );
  MUX4D0 U674 ( .I0(\FIFO_U1/RegFile1/Storage[4][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][26] ), .S0(n641), .S1(n654), .Z(n1043) );
  MUX4D0 U675 ( .I0(\FIFO_U1/RegFile1/Storage[12][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][27] ), .S0(n641), .S1(n654), .Z(n1054)
         );
  MUX4D0 U676 ( .I0(\FIFO_U1/RegFile1/Storage[4][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][27] ), .S0(n641), .S1(n654), .Z(n1056) );
  MUX4D0 U677 ( .I0(\FIFO_U1/RegFile1/Storage[12][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][28] ), .S0(n640), .S1(n652), .Z(n1067)
         );
  MUX4D0 U678 ( .I0(\FIFO_U1/RegFile1/Storage[4][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][28] ), .S0(n640), .S1(n655), .Z(n1069) );
  MUX4D0 U679 ( .I0(\FIFO_U1/RegFile1/Storage[12][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][29] ), .S0(n640), .S1(n655), .Z(n1080)
         );
  MUX4D0 U680 ( .I0(\FIFO_U1/RegFile1/Storage[4][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][29] ), .S0(n640), .S1(n655), .Z(n1082) );
  MUX4D0 U681 ( .I0(\FIFO_U1/RegFile1/Storage[12][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][30] ), .S0(n639), .S1(n659), .Z(n1093)
         );
  MUX4D0 U682 ( .I0(\FIFO_U1/RegFile1/Storage[4][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][30] ), .S0(n639), .S1(n655), .Z(n1095) );
  MUX4D0 U683 ( .I0(\FIFO_U1/RegFile1/Storage[12][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[13][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[14][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[15][31] ), .S0(n639), .S1(n654), .Z(n1106)
         );
  MUX4D0 U684 ( .I0(\FIFO_U1/RegFile1/Storage[4][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[5][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[6][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[7][31] ), .S0(n639), .S1(n660), .Z(n1108) );
  MUX4D0 U685 ( .I0(\FIFO_U1/RegFile1/Storage[16][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][0] ), .S0(n650), .S1(n656), .Z(n702) );
  MUX4D0 U686 ( .I0(\FIFO_U1/RegFile1/Storage[16][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][1] ), .S0(n646), .S1(n656), .Z(n715) );
  MUX4D0 U687 ( .I0(\FIFO_U1/RegFile1/Storage[16][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][2] ), .S0(n646), .S1(n655), .Z(n728) );
  MUX4D0 U688 ( .I0(\FIFO_U1/RegFile1/Storage[16][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][3] ), .S0(n643), .S1(n658), .Z(n741) );
  MUX4D0 U689 ( .I0(\FIFO_U1/RegFile1/Storage[16][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][4] ), .S0(n644), .S1(n652), .Z(n754) );
  MUX4D0 U690 ( .I0(\FIFO_U1/RegFile1/Storage[16][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][5] ), .S0(n650), .S1(n660), .Z(n767) );
  MUX4D0 U691 ( .I0(\FIFO_U1/RegFile1/Storage[16][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][6] ), .S0(n651), .S1(n660), .Z(n780) );
  MUX4D0 U692 ( .I0(\FIFO_U1/RegFile1/Storage[16][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][7] ), .S0(\FIFO_U1/RegFile1/N75 ), .S1(
        n656), .Z(n793) );
  MUX4D0 U693 ( .I0(\FIFO_U1/RegFile1/Storage[16][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][8] ), .S0(n650), .S1(n654), .Z(n806) );
  MUX4D0 U694 ( .I0(\FIFO_U1/RegFile1/Storage[16][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][9] ), .S0(n651), .S1(n659), .Z(n819) );
  MUX4D0 U695 ( .I0(\FIFO_U1/RegFile1/Storage[16][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][10] ), .S0(n648), .S1(n657), .Z(n832) );
  MUX4D0 U696 ( .I0(\FIFO_U1/RegFile1/Storage[16][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][11] ), .S0(n644), .S1(n654), .Z(n845) );
  MUX4D0 U697 ( .I0(\FIFO_U1/RegFile1/Storage[16][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][12] ), .S0(n642), .S1(n652), .Z(n858) );
  MUX4D0 U698 ( .I0(\FIFO_U1/RegFile1/Storage[16][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][13] ), .S0(n641), .S1(n660), .Z(n871) );
  MUX4D0 U699 ( .I0(\FIFO_U1/RegFile1/Storage[16][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][14] ), .S0(n640), .S1(n660), .Z(n884) );
  MUX4D0 U700 ( .I0(\FIFO_U1/RegFile1/Storage[16][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][15] ), .S0(n643), .S1(n659), .Z(n897) );
  MUX4D0 U701 ( .I0(\FIFO_U1/RegFile1/Storage[16][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][16] ), .S0(n647), .S1(n658), .Z(n910) );
  MUX4D0 U702 ( .I0(\FIFO_U1/RegFile1/Storage[16][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][17] ), .S0(n651), .S1(n659), .Z(n923) );
  MUX4D0 U703 ( .I0(\FIFO_U1/RegFile1/Storage[16][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][18] ), .S0(n645), .S1(n659), .Z(n936) );
  MUX4D0 U704 ( .I0(\FIFO_U1/RegFile1/Storage[16][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][19] ), .S0(n640), .S1(n656), .Z(n949) );
  MUX4D0 U705 ( .I0(\FIFO_U1/RegFile1/Storage[16][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][20] ), .S0(n644), .S1(n652), .Z(n962) );
  MUX4D0 U706 ( .I0(\FIFO_U1/RegFile1/Storage[16][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][21] ), .S0(n644), .S1(n658), .Z(n975) );
  MUX4D0 U707 ( .I0(\FIFO_U1/RegFile1/Storage[16][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][22] ), .S0(n644), .S1(n659), .Z(n988) );
  MUX4D0 U708 ( .I0(\FIFO_U1/RegFile1/Storage[16][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][23] ), .S0(n643), .S1(n657), .Z(n1001)
         );
  MUX4D0 U709 ( .I0(\FIFO_U1/RegFile1/Storage[16][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][24] ), .S0(n643), .S1(n652), .Z(n1014)
         );
  MUX4D0 U710 ( .I0(\FIFO_U1/RegFile1/Storage[16][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][25] ), .S0(n642), .S1(n653), .Z(n1027)
         );
  MUX4D0 U711 ( .I0(\FIFO_U1/RegFile1/Storage[16][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][26] ), .S0(n642), .S1(n653), .Z(n1040)
         );
  MUX4D0 U712 ( .I0(\FIFO_U1/RegFile1/Storage[16][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][27] ), .S0(n641), .S1(n654), .Z(n1053)
         );
  MUX4D0 U713 ( .I0(\FIFO_U1/RegFile1/Storage[16][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][28] ), .S0(n641), .S1(n654), .Z(n1066)
         );
  MUX4D0 U714 ( .I0(\FIFO_U1/RegFile1/Storage[16][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][29] ), .S0(n640), .S1(n655), .Z(n1079)
         );
  MUX4D0 U715 ( .I0(\FIFO_U1/RegFile1/Storage[16][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][30] ), .S0(n639), .S1(n656), .Z(n1092)
         );
  MUX4D0 U716 ( .I0(\FIFO_U1/RegFile1/Storage[16][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[17][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[18][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[19][31] ), .S0(n639), .S1(n657), .Z(n1105)
         );
  MUX4D0 U717 ( .I0(\FIFO_U1/RegFile1/Storage[8][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][0] ), .S0(n646), .S1(n656), .Z(n704) );
  MUX4D0 U718 ( .I0(\FIFO_U1/RegFile1/Storage[0][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][0] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][0] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][0] ), .S0(n646), .S1(n656), .Z(n706) );
  MUX4D0 U719 ( .I0(\FIFO_U1/RegFile1/Storage[8][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][1] ), .S0(n646), .S1(n656), .Z(n717) );
  MUX4D0 U720 ( .I0(\FIFO_U1/RegFile1/Storage[0][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][1] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][1] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][1] ), .S0(n646), .S1(n656), .Z(n719) );
  MUX4D0 U721 ( .I0(\FIFO_U1/RegFile1/Storage[8][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][2] ), .S0(n645), .S1(n657), .Z(n730) );
  MUX4D0 U722 ( .I0(\FIFO_U1/RegFile1/Storage[0][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][2] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][2] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][2] ), .S0(n643), .S1(n656), .Z(n732) );
  MUX4D0 U723 ( .I0(\FIFO_U1/RegFile1/Storage[8][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][3] ), .S0(n651), .S1(n659), .Z(n743) );
  MUX4D0 U724 ( .I0(\FIFO_U1/RegFile1/Storage[0][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][3] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][3] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][3] ), .S0(n645), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n745) );
  MUX4D0 U725 ( .I0(\FIFO_U1/RegFile1/Storage[8][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][4] ), .S0(n642), .S1(n659), .Z(n756) );
  MUX4D0 U726 ( .I0(\FIFO_U1/RegFile1/Storage[0][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][4] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][4] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][4] ), .S0(n645), .S1(n657), .Z(n758) );
  MUX4D0 U727 ( .I0(\FIFO_U1/RegFile1/Storage[8][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][5] ), .S0(n647), .S1(n660), .Z(n769) );
  MUX4D0 U728 ( .I0(\FIFO_U1/RegFile1/Storage[0][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][5] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][5] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][5] ), .S0(n646), .S1(n660), .Z(n771) );
  MUX4D0 U729 ( .I0(\FIFO_U1/RegFile1/Storage[8][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][6] ), .S0(n640), .S1(n656), .Z(n782) );
  MUX4D0 U730 ( .I0(\FIFO_U1/RegFile1/Storage[0][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][6] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][6] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][6] ), .S0(n647), .S1(n660), .Z(n784) );
  MUX4D0 U731 ( .I0(\FIFO_U1/RegFile1/Storage[8][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][7] ), .S0(n647), .S1(n659), .Z(n795) );
  MUX4D0 U732 ( .I0(\FIFO_U1/RegFile1/Storage[0][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][7] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][7] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][7] ), .S0(n648), .S1(n655), .Z(n797) );
  MUX4D0 U733 ( .I0(\FIFO_U1/RegFile1/Storage[8][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][8] ), .S0(\FIFO_U1/RegFile1/N75 ), .S1(
        n658), .Z(n808) );
  MUX4D0 U734 ( .I0(\FIFO_U1/RegFile1/Storage[0][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][8] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][8] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][8] ), .S0(n647), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n810) );
  MUX4D0 U735 ( .I0(\FIFO_U1/RegFile1/Storage[8][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][9] ), .S0(n647), .S1(n654), .Z(n821) );
  MUX4D0 U736 ( .I0(\FIFO_U1/RegFile1/Storage[0][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][9] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][9] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][9] ), .S0(n639), .S1(n660), .Z(n823) );
  MUX4D0 U737 ( .I0(\FIFO_U1/RegFile1/Storage[8][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][10] ), .S0(n640), .S1(n655), .Z(n834) );
  MUX4D0 U738 ( .I0(\FIFO_U1/RegFile1/Storage[0][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][10] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][10] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][10] ), .S0(n641), .S1(
        \FIFO_U1/RegFile1/N76 ), .Z(n836) );
  MUX4D0 U739 ( .I0(\FIFO_U1/RegFile1/Storage[8][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][11] ), .S0(n640), .S1(n652), .Z(n847) );
  MUX4D0 U740 ( .I0(\FIFO_U1/RegFile1/Storage[0][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][11] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][11] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][11] ), .S0(n639), .S1(n656), .Z(n849) );
  MUX4D0 U741 ( .I0(\FIFO_U1/RegFile1/Storage[8][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][12] ), .S0(n647), .S1(n659), .Z(n860) );
  MUX4D0 U742 ( .I0(\FIFO_U1/RegFile1/Storage[0][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][12] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][12] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][12] ), .S0(n647), .S1(n654), .Z(n862) );
  MUX4D0 U743 ( .I0(\FIFO_U1/RegFile1/Storage[8][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][13] ), .S0(n639), .S1(n657), .Z(n873) );
  MUX4D0 U744 ( .I0(\FIFO_U1/RegFile1/Storage[0][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][13] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][13] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][13] ), .S0(n642), .S1(n658), .Z(n875) );
  MUX4D0 U745 ( .I0(\FIFO_U1/RegFile1/Storage[8][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][14] ), .S0(n646), .S1(n657), .Z(n886) );
  MUX4D0 U746 ( .I0(\FIFO_U1/RegFile1/Storage[0][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][14] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][14] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][14] ), .S0(n641), .S1(n660), .Z(n888) );
  MUX4D0 U747 ( .I0(\FIFO_U1/RegFile1/Storage[8][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][15] ), .S0(n648), .S1(n657), .Z(n899) );
  MUX4D0 U748 ( .I0(\FIFO_U1/RegFile1/Storage[0][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][15] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][15] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][15] ), .S0(n647), .S1(n658), .Z(n901) );
  MUX4D0 U749 ( .I0(\FIFO_U1/RegFile1/Storage[8][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][16] ), .S0(n645), .S1(n658), .Z(n912) );
  MUX4D0 U750 ( .I0(\FIFO_U1/RegFile1/Storage[0][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][16] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][16] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][16] ), .S0(n649), .S1(n659), .Z(n914) );
  MUX4D0 U751 ( .I0(\FIFO_U1/RegFile1/Storage[8][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][17] ), .S0(n645), .S1(n652), .Z(n925) );
  MUX4D0 U752 ( .I0(\FIFO_U1/RegFile1/Storage[0][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][17] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][17] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][17] ), .S0(n645), .S1(n653), .Z(n927) );
  MUX4D0 U753 ( .I0(\FIFO_U1/RegFile1/Storage[8][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][18] ), .S0(n645), .S1(n658), .Z(n938) );
  MUX4D0 U754 ( .I0(\FIFO_U1/RegFile1/Storage[0][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][18] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][18] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][18] ), .S0(n645), .S1(n655), .Z(n940) );
  MUX4D0 U755 ( .I0(\FIFO_U1/RegFile1/Storage[8][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][19] ), .S0(n648), .S1(n658), .Z(n951) );
  MUX4D0 U756 ( .I0(\FIFO_U1/RegFile1/Storage[0][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][19] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][19] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][19] ), .S0(n651), .S1(n658), .Z(n953) );
  MUX4D0 U757 ( .I0(\FIFO_U1/RegFile1/Storage[8][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][20] ), .S0(n643), .S1(n660), .Z(n964) );
  MUX4D0 U758 ( .I0(\FIFO_U1/RegFile1/Storage[0][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][20] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][20] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][20] ), .S0(n650), .S1(n652), .Z(n966) );
  MUX4D0 U759 ( .I0(\FIFO_U1/RegFile1/Storage[8][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][21] ), .S0(n644), .S1(n658), .Z(n977) );
  MUX4D0 U760 ( .I0(\FIFO_U1/RegFile1/Storage[0][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][21] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][21] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][21] ), .S0(n644), .S1(n652), .Z(n979) );
  MUX4D0 U761 ( .I0(\FIFO_U1/RegFile1/Storage[8][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][22] ), .S0(n644), .S1(n655), .Z(n990) );
  MUX4D0 U762 ( .I0(\FIFO_U1/RegFile1/Storage[0][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][22] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][22] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][22] ), .S0(n643), .S1(n657), .Z(n992) );
  MUX4D0 U763 ( .I0(\FIFO_U1/RegFile1/Storage[8][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][23] ), .S0(n643), .S1(n652), .Z(n1003)
         );
  MUX4D0 U764 ( .I0(\FIFO_U1/RegFile1/Storage[0][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][23] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][23] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][23] ), .S0(n643), .S1(n652), .Z(n1005) );
  MUX4D0 U765 ( .I0(\FIFO_U1/RegFile1/Storage[8][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][24] ), .S0(n643), .S1(n652), .Z(n1016)
         );
  MUX4D0 U766 ( .I0(\FIFO_U1/RegFile1/Storage[0][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][24] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][24] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][24] ), .S0(n642), .S1(n653), .Z(n1018) );
  MUX4D0 U767 ( .I0(\FIFO_U1/RegFile1/Storage[8][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][25] ), .S0(n642), .S1(n653), .Z(n1029)
         );
  MUX4D0 U768 ( .I0(\FIFO_U1/RegFile1/Storage[0][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][25] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][25] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][25] ), .S0(n642), .S1(n653), .Z(n1031) );
  MUX4D0 U769 ( .I0(\FIFO_U1/RegFile1/Storage[8][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][26] ), .S0(n641), .S1(n654), .Z(n1042)
         );
  MUX4D0 U770 ( .I0(\FIFO_U1/RegFile1/Storage[0][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][26] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][26] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][26] ), .S0(n641), .S1(n654), .Z(n1044) );
  MUX4D0 U771 ( .I0(\FIFO_U1/RegFile1/Storage[8][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][27] ), .S0(n641), .S1(n654), .Z(n1055)
         );
  MUX4D0 U772 ( .I0(\FIFO_U1/RegFile1/Storage[0][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][27] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][27] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][27] ), .S0(n641), .S1(n654), .Z(n1057) );
  MUX4D0 U773 ( .I0(\FIFO_U1/RegFile1/Storage[8][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][28] ), .S0(n640), .S1(n655), .Z(n1068)
         );
  MUX4D0 U774 ( .I0(\FIFO_U1/RegFile1/Storage[0][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][28] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][28] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][28] ), .S0(n640), .S1(n655), .Z(n1070) );
  MUX4D0 U775 ( .I0(\FIFO_U1/RegFile1/Storage[8][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][29] ), .S0(n640), .S1(n655), .Z(n1081)
         );
  MUX4D0 U776 ( .I0(\FIFO_U1/RegFile1/Storage[0][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][29] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][29] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][29] ), .S0(n640), .S1(n655), .Z(n1083) );
  MUX4D0 U777 ( .I0(\FIFO_U1/RegFile1/Storage[8][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][30] ), .S0(n639), .S1(n652), .Z(n1094)
         );
  MUX4D0 U778 ( .I0(\FIFO_U1/RegFile1/Storage[0][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][30] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][30] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][30] ), .S0(n639), .S1(n655), .Z(n1096) );
  MUX4D0 U779 ( .I0(\FIFO_U1/RegFile1/Storage[8][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[9][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[10][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[11][31] ), .S0(n639), .S1(n653), .Z(n1107)
         );
  MUX4D0 U780 ( .I0(\FIFO_U1/RegFile1/Storage[0][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[1][31] ), .I2(
        \FIFO_U1/RegFile1/Storage[2][31] ), .I3(
        \FIFO_U1/RegFile1/Storage[3][31] ), .S0(n639), .S1(n653), .Z(n1109) );
  BUFFD1 U781 ( .I(n487), .Z(n636) );
  BUFFD1 U782 ( .I(n487), .Z(n637) );
  BUFFD1 U783 ( .I(n487), .Z(n638) );
  MUX3ND0 U784 ( .I0(n698), .I1(n699), .I2(n700), .S0(n653), .S1(n661), .ZN(
        n697) );
  MUX3ND0 U785 ( .I0(n707), .I1(n708), .I2(n709), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N113 ) );
  MUX3ND0 U786 ( .I0(n711), .I1(n712), .I2(n713), .S0(n652), .S1(n663), .ZN(
        n710) );
  MUX3ND0 U787 ( .I0(n720), .I1(n721), .I2(n722), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N112 ) );
  MUX3ND0 U788 ( .I0(n724), .I1(n725), .I2(n726), .S0(n653), .S1(n664), .ZN(
        n723) );
  MUX3ND0 U789 ( .I0(n733), .I1(n734), .I2(n735), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N111 ) );
  MUX3ND0 U790 ( .I0(n737), .I1(n738), .I2(n739), .S0(n659), .S1(n662), .ZN(
        n736) );
  MUX3ND0 U791 ( .I0(n746), .I1(n747), .I2(n748), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N110 ) );
  MUX3ND0 U792 ( .I0(n750), .I1(n751), .I2(n752), .S0(n658), .S1(n664), .ZN(
        n749) );
  MUX3ND0 U793 ( .I0(n759), .I1(n760), .I2(n761), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N109 ) );
  MUX3ND0 U794 ( .I0(n763), .I1(n764), .I2(n765), .S0(n659), .S1(n665), .ZN(
        n762) );
  MUX3ND0 U795 ( .I0(n772), .I1(n773), .I2(n774), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N108 ) );
  MUX3ND0 U796 ( .I0(n776), .I1(n777), .I2(n778), .S0(n657), .S1(n665), .ZN(
        n775) );
  MUX3ND0 U797 ( .I0(n785), .I1(n786), .I2(n787), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N107 ) );
  MUX3ND0 U798 ( .I0(n789), .I1(n790), .I2(n791), .S0(n655), .S1(n664), .ZN(
        n788) );
  MUX3ND0 U799 ( .I0(n798), .I1(n799), .I2(n800), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N106 ) );
  MUX3ND0 U800 ( .I0(n802), .I1(n803), .I2(n804), .S0(n656), .S1(n662), .ZN(
        n801) );
  MUX3ND0 U801 ( .I0(n811), .I1(n812), .I2(n813), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N105 ) );
  MUX3ND0 U802 ( .I0(n815), .I1(n816), .I2(n817), .S0(n655), .S1(n663), .ZN(
        n814) );
  MUX3ND0 U803 ( .I0(n824), .I1(n825), .I2(n826), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N104 ) );
  MUX3ND0 U804 ( .I0(n828), .I1(n829), .I2(n830), .S0(n654), .S1(n664), .ZN(
        n827) );
  MUX3ND0 U805 ( .I0(n837), .I1(n838), .I2(n839), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N103 ) );
  MUX3ND0 U806 ( .I0(n841), .I1(n842), .I2(n843), .S0(n654), .S1(n661), .ZN(
        n840) );
  MUX3ND0 U807 ( .I0(n850), .I1(n851), .I2(n852), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N102 ) );
  MUX3ND0 U808 ( .I0(n854), .I1(n855), .I2(n856), .S0(n657), .S1(n664), .ZN(
        n853) );
  MUX3ND0 U809 ( .I0(n863), .I1(n864), .I2(n865), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N101 ) );
  MUX3ND0 U810 ( .I0(n867), .I1(n868), .I2(n869), .S0(n659), .S1(n661), .ZN(
        n866) );
  MUX3ND0 U811 ( .I0(n876), .I1(n877), .I2(n878), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N100 ) );
  MUX3ND0 U812 ( .I0(n880), .I1(n881), .I2(n882), .S0(n655), .S1(n665), .ZN(
        n879) );
  MUX3ND0 U813 ( .I0(n889), .I1(n890), .I2(n891), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N99 ) );
  MUX3ND0 U814 ( .I0(n893), .I1(n894), .I2(n895), .S0(n654), .S1(n662), .ZN(
        n892) );
  MUX3ND0 U815 ( .I0(n902), .I1(n903), .I2(n904), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N98 ) );
  MUX3ND0 U816 ( .I0(n906), .I1(n907), .I2(n908), .S0(n653), .S1(n663), .ZN(
        n905) );
  MUX3ND0 U817 ( .I0(n915), .I1(n916), .I2(n917), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N97 ) );
  MUX3ND0 U818 ( .I0(n919), .I1(n920), .I2(n921), .S0(n655), .S1(n665), .ZN(
        n918) );
  MUX3ND0 U819 ( .I0(n928), .I1(n929), .I2(n930), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N96 ) );
  MUX3ND0 U820 ( .I0(n932), .I1(n933), .I2(n934), .S0(n655), .S1(n665), .ZN(
        n931) );
  MUX3ND0 U821 ( .I0(n941), .I1(n942), .I2(n943), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N95 ) );
  MUX3ND0 U822 ( .I0(n945), .I1(n946), .I2(n947), .S0(n660), .S1(n665), .ZN(
        n944) );
  MUX3ND0 U823 ( .I0(n954), .I1(n955), .I2(n956), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N94 ) );
  MUX3ND0 U824 ( .I0(n958), .I1(n959), .I2(n960), .S0(n652), .S1(n665), .ZN(
        n957) );
  MUX3ND0 U825 ( .I0(n967), .I1(n968), .I2(n969), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N93 ) );
  MUX3ND0 U826 ( .I0(n971), .I1(n972), .I2(n973), .S0(n657), .S1(n665), .ZN(
        n970) );
  MUX3ND0 U827 ( .I0(n980), .I1(n981), .I2(n982), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N92 ) );
  MUX3ND0 U828 ( .I0(n984), .I1(n985), .I2(n986), .S0(n652), .S1(n665), .ZN(
        n983) );
  MUX3ND0 U829 ( .I0(n993), .I1(n994), .I2(n995), .S0(\FIFO_U1/RegFile1/N78 ), 
        .S1(\FIFO_U1/RegFile1/N79 ), .ZN(\FIFO_U1/RegFile1/N91 ) );
  MUX3ND0 U830 ( .I0(n997), .I1(n998), .I2(n999), .S0(n653), .S1(n665), .ZN(
        n996) );
  MUX3ND0 U831 ( .I0(n1006), .I1(n1007), .I2(n1008), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N90 ) );
  MUX3ND0 U832 ( .I0(n1010), .I1(n1011), .I2(n1012), .S0(n654), .S1(n665), 
        .ZN(n1009) );
  MUX3ND0 U833 ( .I0(n1019), .I1(n1020), .I2(n1021), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N89 ) );
  MUX3ND0 U834 ( .I0(n1023), .I1(n1024), .I2(n1025), .S0(n657), .S1(n665), 
        .ZN(n1022) );
  MUX3ND0 U835 ( .I0(n1032), .I1(n1033), .I2(n1034), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N88 ) );
  MUX3ND0 U836 ( .I0(n1036), .I1(n1037), .I2(n1038), .S0(n656), .S1(n665), 
        .ZN(n1035) );
  MUX3ND0 U837 ( .I0(n1045), .I1(n1046), .I2(n1047), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N87 ) );
  MUX3ND0 U838 ( .I0(n1049), .I1(n1050), .I2(n1051), .S0(n658), .S1(n664), 
        .ZN(n1048) );
  MUX3ND0 U839 ( .I0(n1058), .I1(n1059), .I2(n1060), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N86 ) );
  MUX3ND0 U840 ( .I0(n1062), .I1(n1063), .I2(n1064), .S0(n656), .S1(n665), 
        .ZN(n1061) );
  MUX3ND0 U841 ( .I0(n1071), .I1(n1072), .I2(n1073), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N85 ) );
  MUX3ND0 U842 ( .I0(n1075), .I1(n1076), .I2(n1077), .S0(n657), .S1(n665), 
        .ZN(n1074) );
  MUX3ND0 U843 ( .I0(n1084), .I1(n1085), .I2(n1086), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N84 ) );
  MUX3ND0 U844 ( .I0(n1088), .I1(n1089), .I2(n1090), .S0(
        \FIFO_U1/RegFile1/N76 ), .S1(n664), .ZN(n1087) );
  MUX3ND0 U845 ( .I0(n1097), .I1(n1098), .I2(n1099), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N83 ) );
  MUX3ND0 U846 ( .I0(n1101), .I1(n1102), .I2(n1103), .S0(n652), .S1(n664), 
        .ZN(n1100) );
  MUX3ND0 U847 ( .I0(n1110), .I1(n1111), .I2(n1112), .S0(
        \FIFO_U1/RegFile1/N78 ), .S1(\FIFO_U1/RegFile1/N79 ), .ZN(
        \FIFO_U1/RegFile1/N82 ) );
  MUX2ND0 U848 ( .I0(\FIFO_U1/RegFile1/Storage[26][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][0] ), .S(n650), .ZN(n699) );
  MUX2ND0 U849 ( .I0(\FIFO_U1/RegFile1/Storage[24][0] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][0] ), .S(n648), .ZN(n698) );
  MUX3ND0 U850 ( .I0(n702), .I1(n701), .I2(n697), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n709) );
  MUX2ND0 U851 ( .I0(n704), .I1(n703), .S(n664), .ZN(n708) );
  MUX2ND0 U852 ( .I0(n706), .I1(n705), .S(n664), .ZN(n707) );
  MUX2ND0 U853 ( .I0(\FIFO_U1/RegFile1/Storage[26][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][1] ), .S(n649), .ZN(n712) );
  MUX2ND0 U854 ( .I0(\FIFO_U1/RegFile1/Storage[24][1] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][1] ), .S(n646), .ZN(n711) );
  MUX3ND0 U855 ( .I0(n715), .I1(n714), .I2(n710), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n722) );
  MUX2ND0 U856 ( .I0(n717), .I1(n716), .S(n664), .ZN(n721) );
  MUX2ND0 U857 ( .I0(n719), .I1(n718), .S(n664), .ZN(n720) );
  MUX2ND0 U858 ( .I0(\FIFO_U1/RegFile1/Storage[26][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][2] ), .S(n643), .ZN(n725) );
  MUX2ND0 U859 ( .I0(\FIFO_U1/RegFile1/Storage[24][2] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][2] ), .S(n648), .ZN(n724) );
  MUX3ND0 U860 ( .I0(n728), .I1(n727), .I2(n723), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n735) );
  MUX2ND0 U861 ( .I0(n730), .I1(n729), .S(n664), .ZN(n734) );
  MUX2ND0 U862 ( .I0(n732), .I1(n731), .S(n663), .ZN(n733) );
  MUX2ND0 U863 ( .I0(\FIFO_U1/RegFile1/Storage[26][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][3] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n738) );
  MUX2ND0 U864 ( .I0(\FIFO_U1/RegFile1/Storage[24][3] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][3] ), .S(n649), .ZN(n737) );
  MUX3ND0 U865 ( .I0(n741), .I1(n740), .I2(n736), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n748) );
  MUX2ND0 U866 ( .I0(n743), .I1(n742), .S(n664), .ZN(n747) );
  MUX2ND0 U867 ( .I0(n745), .I1(n744), .S(n664), .ZN(n746) );
  MUX2ND0 U868 ( .I0(\FIFO_U1/RegFile1/Storage[26][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][4] ), .S(n651), .ZN(n751) );
  MUX2ND0 U869 ( .I0(\FIFO_U1/RegFile1/Storage[24][4] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][4] ), .S(n650), .ZN(n750) );
  MUX3ND0 U870 ( .I0(n754), .I1(n753), .I2(n749), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n761) );
  MUX2ND0 U871 ( .I0(n756), .I1(n755), .S(n664), .ZN(n760) );
  MUX2ND0 U872 ( .I0(n758), .I1(n757), .S(n661), .ZN(n759) );
  MUX2ND0 U873 ( .I0(\FIFO_U1/RegFile1/Storage[26][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][5] ), .S(n651), .ZN(n764) );
  MUX2ND0 U874 ( .I0(\FIFO_U1/RegFile1/Storage[24][5] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][5] ), .S(n646), .ZN(n763) );
  MUX3ND0 U875 ( .I0(n767), .I1(n766), .I2(n762), .S0(n665), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n774) );
  MUX2ND0 U876 ( .I0(n769), .I1(n768), .S(n662), .ZN(n773) );
  MUX2ND0 U877 ( .I0(n771), .I1(n770), .S(n663), .ZN(n772) );
  MUX2ND0 U878 ( .I0(\FIFO_U1/RegFile1/Storage[26][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][6] ), .S(n648), .ZN(n777) );
  MUX2ND0 U879 ( .I0(\FIFO_U1/RegFile1/Storage[24][6] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][6] ), .S(n647), .ZN(n776) );
  MUX3ND0 U880 ( .I0(n780), .I1(n779), .I2(n775), .S0(n663), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n787) );
  MUX2ND0 U881 ( .I0(n782), .I1(n781), .S(n662), .ZN(n786) );
  MUX2ND0 U882 ( .I0(n784), .I1(n783), .S(n665), .ZN(n785) );
  MUX2ND0 U883 ( .I0(\FIFO_U1/RegFile1/Storage[26][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][7] ), .S(n644), .ZN(n790) );
  MUX2ND0 U884 ( .I0(\FIFO_U1/RegFile1/Storage[24][7] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][7] ), .S(n647), .ZN(n789) );
  MUX3ND0 U885 ( .I0(n793), .I1(n792), .I2(n788), .S0(n664), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n800) );
  MUX2ND0 U886 ( .I0(n795), .I1(n794), .S(n665), .ZN(n799) );
  MUX2ND0 U887 ( .I0(n797), .I1(n796), .S(n663), .ZN(n798) );
  MUX2ND0 U888 ( .I0(\FIFO_U1/RegFile1/Storage[26][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][8] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n803) );
  MUX2ND0 U889 ( .I0(\FIFO_U1/RegFile1/Storage[24][8] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][8] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n802) );
  MUX3ND0 U890 ( .I0(n806), .I1(n805), .I2(n801), .S0(n663), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n813) );
  MUX2ND0 U891 ( .I0(n808), .I1(n807), .S(n661), .ZN(n812) );
  MUX2ND0 U892 ( .I0(n810), .I1(n809), .S(n661), .ZN(n811) );
  MUX2ND0 U893 ( .I0(\FIFO_U1/RegFile1/Storage[26][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][9] ), .S(n647), .ZN(n816) );
  MUX2ND0 U894 ( .I0(\FIFO_U1/RegFile1/Storage[24][9] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][9] ), .S(n643), .ZN(n815) );
  MUX3ND0 U895 ( .I0(n819), .I1(n818), .I2(n814), .S0(n664), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n826) );
  MUX2ND0 U896 ( .I0(n821), .I1(n820), .S(n664), .ZN(n825) );
  MUX2ND0 U897 ( .I0(n823), .I1(n822), .S(n664), .ZN(n824) );
  MUX2ND0 U898 ( .I0(\FIFO_U1/RegFile1/Storage[26][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][10] ), .S(n648), .ZN(n829) );
  MUX2ND0 U899 ( .I0(\FIFO_U1/RegFile1/Storage[24][10] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][10] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n828) );
  MUX3ND0 U900 ( .I0(n832), .I1(n831), .I2(n827), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n839) );
  MUX2ND0 U901 ( .I0(n834), .I1(n833), .S(n663), .ZN(n838) );
  MUX2ND0 U902 ( .I0(n836), .I1(n835), .S(n665), .ZN(n837) );
  MUX2ND0 U903 ( .I0(\FIFO_U1/RegFile1/Storage[26][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][11] ), .S(n648), .ZN(n842) );
  MUX2ND0 U904 ( .I0(\FIFO_U1/RegFile1/Storage[24][11] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][11] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n841) );
  MUX3ND0 U905 ( .I0(n845), .I1(n844), .I2(n840), .S0(n663), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n852) );
  MUX2ND0 U906 ( .I0(n847), .I1(n846), .S(n662), .ZN(n851) );
  MUX2ND0 U907 ( .I0(n849), .I1(n848), .S(n664), .ZN(n850) );
  MUX2ND0 U908 ( .I0(\FIFO_U1/RegFile1/Storage[26][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][12] ), .S(n650), .ZN(n855) );
  MUX2ND0 U909 ( .I0(\FIFO_U1/RegFile1/Storage[24][12] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][12] ), .S(n650), .ZN(n854) );
  MUX3ND0 U910 ( .I0(n858), .I1(n857), .I2(n853), .S0(n665), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n865) );
  MUX2ND0 U911 ( .I0(n860), .I1(n859), .S(n665), .ZN(n864) );
  MUX2ND0 U912 ( .I0(n862), .I1(n861), .S(n661), .ZN(n863) );
  MUX2ND0 U913 ( .I0(\FIFO_U1/RegFile1/Storage[26][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][13] ), .S(n651), .ZN(n868) );
  MUX2ND0 U914 ( .I0(\FIFO_U1/RegFile1/Storage[24][13] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][13] ), .S(n649), .ZN(n867) );
  MUX3ND0 U915 ( .I0(n871), .I1(n870), .I2(n866), .S0(n665), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n878) );
  MUX2ND0 U916 ( .I0(n873), .I1(n872), .S(n665), .ZN(n877) );
  MUX2ND0 U917 ( .I0(n875), .I1(n874), .S(n663), .ZN(n876) );
  MUX2ND0 U918 ( .I0(\FIFO_U1/RegFile1/Storage[26][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][14] ), .S(n648), .ZN(n881) );
  MUX2ND0 U919 ( .I0(\FIFO_U1/RegFile1/Storage[24][14] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][14] ), .S(n651), .ZN(n880) );
  MUX3ND0 U920 ( .I0(n884), .I1(n883), .I2(n879), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n891) );
  MUX2ND0 U921 ( .I0(n886), .I1(n885), .S(n662), .ZN(n890) );
  MUX2ND0 U922 ( .I0(n888), .I1(n887), .S(n663), .ZN(n889) );
  MUX2ND0 U923 ( .I0(\FIFO_U1/RegFile1/Storage[26][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][15] ), .S(n640), .ZN(n894) );
  MUX2ND0 U924 ( .I0(\FIFO_U1/RegFile1/Storage[24][15] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][15] ), .S(n650), .ZN(n893) );
  MUX3ND0 U925 ( .I0(n897), .I1(n896), .I2(n892), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n904) );
  MUX2ND0 U926 ( .I0(n899), .I1(n898), .S(n661), .ZN(n903) );
  MUX2ND0 U927 ( .I0(n901), .I1(n900), .S(n663), .ZN(n902) );
  MUX2ND0 U928 ( .I0(\FIFO_U1/RegFile1/Storage[26][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][16] ), .S(n649), .ZN(n907) );
  MUX2ND0 U929 ( .I0(\FIFO_U1/RegFile1/Storage[24][16] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][16] ), .S(n650), .ZN(n906) );
  MUX3ND0 U930 ( .I0(n910), .I1(n909), .I2(n905), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n917) );
  MUX2ND0 U931 ( .I0(n912), .I1(n911), .S(n661), .ZN(n916) );
  MUX2ND0 U932 ( .I0(n914), .I1(n913), .S(n663), .ZN(n915) );
  MUX2ND0 U933 ( .I0(\FIFO_U1/RegFile1/Storage[26][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][17] ), .S(n639), .ZN(n920) );
  MUX2ND0 U934 ( .I0(\FIFO_U1/RegFile1/Storage[24][17] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][17] ), .S(n647), .ZN(n919) );
  MUX3ND0 U935 ( .I0(n923), .I1(n922), .I2(n918), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n930) );
  MUX2ND0 U936 ( .I0(n925), .I1(n924), .S(n663), .ZN(n929) );
  MUX2ND0 U937 ( .I0(n927), .I1(n926), .S(n662), .ZN(n928) );
  MUX2ND0 U938 ( .I0(\FIFO_U1/RegFile1/Storage[26][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][18] ), .S(n651), .ZN(n933) );
  MUX2ND0 U939 ( .I0(\FIFO_U1/RegFile1/Storage[24][18] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][18] ), .S(n643), .ZN(n932) );
  MUX3ND0 U940 ( .I0(n936), .I1(n935), .I2(n931), .S0(n664), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n943) );
  MUX2ND0 U941 ( .I0(n938), .I1(n937), .S(n663), .ZN(n942) );
  MUX2ND0 U942 ( .I0(n940), .I1(n939), .S(n663), .ZN(n941) );
  MUX2ND0 U943 ( .I0(\FIFO_U1/RegFile1/Storage[26][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][19] ), .S(n644), .ZN(n946) );
  MUX2ND0 U944 ( .I0(\FIFO_U1/RegFile1/Storage[24][19] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][19] ), .S(n640), .ZN(n945) );
  MUX3ND0 U945 ( .I0(n949), .I1(n948), .I2(n944), .S0(n663), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n956) );
  MUX2ND0 U946 ( .I0(n951), .I1(n950), .S(n661), .ZN(n955) );
  MUX2ND0 U947 ( .I0(n953), .I1(n952), .S(n663), .ZN(n954) );
  MUX2ND0 U948 ( .I0(\FIFO_U1/RegFile1/Storage[26][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][20] ), .S(n650), .ZN(n959) );
  MUX2ND0 U949 ( .I0(\FIFO_U1/RegFile1/Storage[24][20] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][20] ), .S(n649), .ZN(n958) );
  MUX3ND0 U950 ( .I0(n962), .I1(n961), .I2(n957), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n969) );
  MUX2ND0 U951 ( .I0(n964), .I1(n963), .S(n665), .ZN(n968) );
  MUX2ND0 U952 ( .I0(n966), .I1(n965), .S(n662), .ZN(n967) );
  MUX2ND0 U953 ( .I0(\FIFO_U1/RegFile1/Storage[26][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][21] ), .S(n641), .ZN(n972) );
  MUX2ND0 U954 ( .I0(\FIFO_U1/RegFile1/Storage[24][21] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][21] ), .S(n641), .ZN(n971) );
  MUX3ND0 U955 ( .I0(n975), .I1(n974), .I2(n970), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n982) );
  MUX2ND0 U956 ( .I0(n977), .I1(n976), .S(n664), .ZN(n981) );
  MUX2ND0 U957 ( .I0(n979), .I1(n978), .S(n662), .ZN(n980) );
  MUX2ND0 U958 ( .I0(\FIFO_U1/RegFile1/Storage[26][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][22] ), .S(n642), .ZN(n985) );
  MUX2ND0 U959 ( .I0(\FIFO_U1/RegFile1/Storage[24][22] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][22] ), .S(n647), .ZN(n984) );
  MUX3ND0 U960 ( .I0(n988), .I1(n987), .I2(n983), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n995) );
  MUX2ND0 U961 ( .I0(n990), .I1(n989), .S(n662), .ZN(n994) );
  MUX2ND0 U962 ( .I0(n992), .I1(n991), .S(n663), .ZN(n993) );
  MUX2ND0 U963 ( .I0(\FIFO_U1/RegFile1/Storage[26][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][23] ), .S(n642), .ZN(n998) );
  MUX2ND0 U964 ( .I0(\FIFO_U1/RegFile1/Storage[24][23] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][23] ), .S(n650), .ZN(n997) );
  MUX3ND0 U965 ( .I0(n1001), .I1(n1000), .I2(n996), .S0(n665), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1008) );
  MUX2ND0 U966 ( .I0(n1003), .I1(n1002), .S(n661), .ZN(n1007) );
  MUX2ND0 U967 ( .I0(n1005), .I1(n1004), .S(n662), .ZN(n1006) );
  MUX2ND0 U968 ( .I0(\FIFO_U1/RegFile1/Storage[26][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][24] ), .S(n648), .ZN(n1011) );
  MUX2ND0 U969 ( .I0(\FIFO_U1/RegFile1/Storage[24][24] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][24] ), .S(n651), .ZN(n1010) );
  MUX3ND0 U970 ( .I0(n1014), .I1(n1013), .I2(n1009), .S0(n662), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1021) );
  MUX2ND0 U971 ( .I0(n1016), .I1(n1015), .S(n662), .ZN(n1020) );
  MUX2ND0 U972 ( .I0(n1018), .I1(n1017), .S(n663), .ZN(n1019) );
  MUX2ND0 U973 ( .I0(\FIFO_U1/RegFile1/Storage[26][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][25] ), .S(n651), .ZN(n1024) );
  MUX2ND0 U974 ( .I0(\FIFO_U1/RegFile1/Storage[24][25] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][25] ), .S(n649), .ZN(n1023) );
  MUX3ND0 U975 ( .I0(n1027), .I1(n1026), .I2(n1022), .S0(n663), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1034) );
  MUX2ND0 U976 ( .I0(n1029), .I1(n1028), .S(n665), .ZN(n1033) );
  MUX2ND0 U977 ( .I0(n1031), .I1(n1030), .S(n662), .ZN(n1032) );
  MUX2ND0 U978 ( .I0(\FIFO_U1/RegFile1/Storage[26][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][26] ), .S(n649), .ZN(n1037) );
  MUX2ND0 U979 ( .I0(\FIFO_U1/RegFile1/Storage[24][26] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][26] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n1036) );
  MUX3ND0 U980 ( .I0(n1040), .I1(n1039), .I2(n1035), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1047) );
  MUX2ND0 U981 ( .I0(n1042), .I1(n1041), .S(n662), .ZN(n1046) );
  MUX2ND0 U982 ( .I0(n1044), .I1(n1043), .S(n663), .ZN(n1045) );
  MUX2ND0 U983 ( .I0(\FIFO_U1/RegFile1/Storage[26][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][27] ), .S(n651), .ZN(n1050) );
  MUX2ND0 U984 ( .I0(\FIFO_U1/RegFile1/Storage[24][27] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][27] ), .S(n648), .ZN(n1049) );
  MUX3ND0 U985 ( .I0(n1053), .I1(n1052), .I2(n1048), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1060) );
  MUX2ND0 U986 ( .I0(n1055), .I1(n1054), .S(n663), .ZN(n1059) );
  MUX2ND0 U987 ( .I0(n1057), .I1(n1056), .S(n662), .ZN(n1058) );
  MUX2ND0 U988 ( .I0(\FIFO_U1/RegFile1/Storage[26][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][28] ), .S(n649), .ZN(n1063) );
  MUX2ND0 U989 ( .I0(\FIFO_U1/RegFile1/Storage[24][28] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][28] ), .S(n647), .ZN(n1062) );
  MUX3ND0 U990 ( .I0(n1066), .I1(n1065), .I2(n1061), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1073) );
  MUX2ND0 U991 ( .I0(n1068), .I1(n1067), .S(n662), .ZN(n1072) );
  MUX2ND0 U992 ( .I0(n1070), .I1(n1069), .S(n664), .ZN(n1071) );
  MUX2ND0 U993 ( .I0(\FIFO_U1/RegFile1/Storage[26][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][29] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n1076) );
  MUX2ND0 U994 ( .I0(\FIFO_U1/RegFile1/Storage[24][29] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][29] ), .S(\FIFO_U1/RegFile1/N75 ), .ZN(
        n1075) );
  MUX3ND0 U995 ( .I0(n1079), .I1(n1078), .I2(n1074), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1086) );
  MUX2ND0 U996 ( .I0(n1081), .I1(n1080), .S(n664), .ZN(n1085) );
  MUX2ND0 U997 ( .I0(n1083), .I1(n1082), .S(n662), .ZN(n1084) );
  MUX2ND0 U998 ( .I0(\FIFO_U1/RegFile1/Storage[26][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][30] ), .S(n650), .ZN(n1089) );
  MUX2ND0 U999 ( .I0(\FIFO_U1/RegFile1/Storage[24][30] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][30] ), .S(n639), .ZN(n1088) );
  MUX3ND0 U1000 ( .I0(n1092), .I1(n1091), .I2(n1087), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1099) );
  MUX2ND0 U1001 ( .I0(n1094), .I1(n1093), .S(n662), .ZN(n1098) );
  MUX2ND0 U1002 ( .I0(n1096), .I1(n1095), .S(n665), .ZN(n1097) );
  MUX2ND0 U1003 ( .I0(\FIFO_U1/RegFile1/Storage[26][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[27][31] ), .S(n651), .ZN(n1102) );
  MUX2ND0 U1004 ( .I0(\FIFO_U1/RegFile1/Storage[24][31] ), .I1(
        \FIFO_U1/RegFile1/Storage[25][31] ), .S(n649), .ZN(n1101) );
  MUX3ND0 U1005 ( .I0(n1105), .I1(n1104), .I2(n1100), .S0(n661), .S1(
        \FIFO_U1/RegFile1/N78 ), .ZN(n1112) );
  MUX2ND0 U1006 ( .I0(n1107), .I1(n1106), .S(n663), .ZN(n1111) );
  MUX2ND0 U1007 ( .I0(n1109), .I1(n1108), .S(n664), .ZN(n1110) );
  MUX2D0 U1008 ( .I0(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[4] ), .I1(
        \SerialRx_U1/PLL_RxU1/VFO1/N53 ), .S(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .Z(n489) );
  XNR2D0 U1009 ( .A1(SerialClk), .A2(n1113), .ZN(n488) );
  MUX2ND0 U1010 ( .I0(n561), .I1(n375), .S(\DesDecoder_U1/N44 ), .ZN(n486) );
  MUX2ND0 U1011 ( .I0(n560), .I1(n341), .S(\DesDecoder_U1/N44 ), .ZN(n485) );
  MUX2ND0 U1012 ( .I0(n559), .I1(n339), .S(\DesDecoder_U1/N44 ), .ZN(n484) );
  MUX2ND0 U1013 ( .I0(n558), .I1(n337), .S(\DesDecoder_U1/N44 ), .ZN(n483) );
  MUX2ND0 U1014 ( .I0(n557), .I1(n335), .S(\DesDecoder_U1/N44 ), .ZN(n482) );
  MUX2ND0 U1015 ( .I0(n556), .I1(n333), .S(\DesDecoder_U1/N44 ), .ZN(n481) );
  MUX2ND0 U1016 ( .I0(n555), .I1(n331), .S(\DesDecoder_U1/N44 ), .ZN(n480) );
  MUX2ND0 U1017 ( .I0(n554), .I1(n329), .S(\DesDecoder_U1/N44 ), .ZN(n479) );
  MUX2ND0 U1018 ( .I0(n553), .I1(n327), .S(\DesDecoder_U1/N44 ), .ZN(n478) );
  MUX2ND0 U1019 ( .I0(n552), .I1(n325), .S(\DesDecoder_U1/N44 ), .ZN(n477) );
  MUX2ND0 U1020 ( .I0(n551), .I1(n323), .S(\DesDecoder_U1/N44 ), .ZN(n476) );
  MUX2ND0 U1021 ( .I0(n550), .I1(n321), .S(\DesDecoder_U1/N44 ), .ZN(n475) );
  MUX2ND0 U1022 ( .I0(n549), .I1(n319), .S(\DesDecoder_U1/N44 ), .ZN(n474) );
  MUX2ND0 U1023 ( .I0(n548), .I1(n317), .S(\DesDecoder_U1/N44 ), .ZN(n473) );
  MUX2ND0 U1024 ( .I0(n547), .I1(n315), .S(\DesDecoder_U1/N44 ), .ZN(n472) );
  MUX2ND0 U1025 ( .I0(n546), .I1(n313), .S(\DesDecoder_U1/N44 ), .ZN(n471) );
  MUX2ND0 U1026 ( .I0(n545), .I1(n311), .S(\DesDecoder_U1/N44 ), .ZN(n470) );
  MUX2ND0 U1027 ( .I0(n544), .I1(n309), .S(\DesDecoder_U1/N44 ), .ZN(n469) );
  MUX2ND0 U1028 ( .I0(n543), .I1(n307), .S(\DesDecoder_U1/N44 ), .ZN(n468) );
  MUX2ND0 U1029 ( .I0(n542), .I1(n305), .S(\DesDecoder_U1/N44 ), .ZN(n467) );
  MUX2ND0 U1030 ( .I0(n541), .I1(n303), .S(\DesDecoder_U1/N44 ), .ZN(n466) );
  MUX2ND0 U1031 ( .I0(n540), .I1(n301), .S(\DesDecoder_U1/N44 ), .ZN(n465) );
  MUX2ND0 U1032 ( .I0(n539), .I1(n299), .S(\DesDecoder_U1/N44 ), .ZN(n464) );
  MUX2ND0 U1033 ( .I0(n538), .I1(n297), .S(\DesDecoder_U1/N44 ), .ZN(n463) );
  MUX2ND0 U1034 ( .I0(n537), .I1(n295), .S(\DesDecoder_U1/N44 ), .ZN(n462) );
  MUX2ND0 U1035 ( .I0(n536), .I1(n293), .S(\DesDecoder_U1/N44 ), .ZN(n461) );
  MUX2ND0 U1036 ( .I0(n535), .I1(n291), .S(\DesDecoder_U1/N44 ), .ZN(n460) );
  MUX2ND0 U1037 ( .I0(n534), .I1(n289), .S(\DesDecoder_U1/N44 ), .ZN(n459) );
  MUX2ND0 U1038 ( .I0(n533), .I1(n287), .S(\DesDecoder_U1/N44 ), .ZN(n458) );
  MUX2ND0 U1039 ( .I0(n532), .I1(n285), .S(\DesDecoder_U1/N44 ), .ZN(n457) );
  MUX2ND0 U1040 ( .I0(n531), .I1(n283), .S(\DesDecoder_U1/N44 ), .ZN(n456) );
  MUX2ND0 U1041 ( .I0(n530), .I1(n281), .S(\DesDecoder_U1/N44 ), .ZN(n455) );
  MUX2D0 U1042 ( .I0(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[0] ), .I1(
        \SerialRx_U1/PLL_RxU1/VFO1/N45 ), .S(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .Z(n454) );
  MUX2D0 U1043 ( .I0(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] ), .I1(
        \SerialRx_U1/PLL_RxU1/VFO1/N47 ), .S(\SerialRx_U1/PLL_RxU1/VFO1/N54 ), 
        .Z(n453) );
  MUX2ND0 U1044 ( .I0(n279), .I1(n530), .S(n1242), .ZN(n452) );
  MUX2ND0 U1045 ( .I0(n278), .I1(n531), .S(n1242), .ZN(n451) );
  MUX2ND0 U1046 ( .I0(n277), .I1(n532), .S(n1242), .ZN(n450) );
  MUX2ND0 U1047 ( .I0(n276), .I1(n533), .S(n1242), .ZN(n449) );
  MUX2ND0 U1048 ( .I0(n275), .I1(n534), .S(n1242), .ZN(n448) );
  MUX2ND0 U1049 ( .I0(n274), .I1(n535), .S(n1242), .ZN(n447) );
  MUX2ND0 U1050 ( .I0(n273), .I1(n536), .S(n1242), .ZN(n446) );
  MUX2ND0 U1051 ( .I0(n272), .I1(n537), .S(n1242), .ZN(n445) );
  MUX2ND0 U1052 ( .I0(n271), .I1(n538), .S(n1242), .ZN(n444) );
  MUX2ND0 U1053 ( .I0(n270), .I1(n539), .S(n1242), .ZN(n443) );
  MUX2ND0 U1054 ( .I0(n269), .I1(n540), .S(n1242), .ZN(n442) );
  MUX2ND0 U1055 ( .I0(n268), .I1(n541), .S(n1242), .ZN(n441) );
  MUX2ND0 U1056 ( .I0(n267), .I1(n542), .S(n1242), .ZN(n440) );
  MUX2ND0 U1057 ( .I0(n266), .I1(n543), .S(n1242), .ZN(n439) );
  MUX2ND0 U1058 ( .I0(n265), .I1(n544), .S(n1242), .ZN(n438) );
  MUX2ND0 U1059 ( .I0(n264), .I1(n545), .S(n1242), .ZN(n437) );
  MUX2ND0 U1060 ( .I0(n263), .I1(n546), .S(n1242), .ZN(n436) );
  MUX2ND0 U1061 ( .I0(n262), .I1(n547), .S(n1242), .ZN(n435) );
  MUX2ND0 U1062 ( .I0(n261), .I1(n548), .S(n1242), .ZN(n434) );
  MUX2ND0 U1063 ( .I0(n260), .I1(n549), .S(n1242), .ZN(n433) );
  MUX2ND0 U1064 ( .I0(n259), .I1(n550), .S(n1242), .ZN(n432) );
  MUX2ND0 U1065 ( .I0(n258), .I1(n551), .S(n1242), .ZN(n431) );
  MUX2ND0 U1066 ( .I0(n257), .I1(n552), .S(n1242), .ZN(n430) );
  MUX2ND0 U1067 ( .I0(n256), .I1(n553), .S(n1242), .ZN(n429) );
  MUX2ND0 U1068 ( .I0(n255), .I1(n554), .S(n1242), .ZN(n428) );
  MUX2ND0 U1069 ( .I0(n254), .I1(n555), .S(n1242), .ZN(n427) );
  MUX2ND0 U1070 ( .I0(n253), .I1(n556), .S(n1242), .ZN(n426) );
  MUX2ND0 U1071 ( .I0(n252), .I1(n557), .S(n1242), .ZN(n425) );
  MUX2ND0 U1072 ( .I0(n251), .I1(n558), .S(n1242), .ZN(n424) );
  MUX2ND0 U1073 ( .I0(n250), .I1(n559), .S(n1242), .ZN(n423) );
  MUX2ND0 U1074 ( .I0(n249), .I1(n560), .S(n1242), .ZN(n422) );
  MUX2ND0 U1075 ( .I0(n248), .I1(n561), .S(n1242), .ZN(n421) );
  AO21D0 U1076 ( .A1(DecoderParClk), .A2(n1247), .B(n1242), .Z(n420) );
  CKND0 U1077 ( .CLK(\FIFO_U1/RegFile1/N32 ), .CN(n418) );
  CKND0 U1078 ( .CLK(\FIFO_U1/RegFile1/N33 ), .CN(n417) );
  CKND0 U1079 ( .CLK(\FIFO_U1/RegFile1/N34 ), .CN(n416) );
  CKND0 U1080 ( .CLK(\FIFO_U1/RegFile1/N35 ), .CN(n415) );
  CKND0 U1081 ( .CLK(\FIFO_U1/RegFile1/N36 ), .CN(n414) );
  CKND0 U1082 ( .CLK(\FIFO_U1/RegFile1/N37 ), .CN(n413) );
  CKND0 U1083 ( .CLK(\FIFO_U1/RegFile1/N38 ), .CN(n412) );
  CKND0 U1084 ( .CLK(\FIFO_U1/RegFile1/N39 ), .CN(n411) );
  CKND0 U1085 ( .CLK(\FIFO_U1/RegFile1/N40 ), .CN(n410) );
  CKND0 U1086 ( .CLK(\FIFO_U1/RegFile1/N41 ), .CN(n409) );
  CKND0 U1087 ( .CLK(\FIFO_U1/RegFile1/N42 ), .CN(n408) );
  CKND0 U1088 ( .CLK(\FIFO_U1/RegFile1/N43 ), .CN(n407) );
  CKND0 U1089 ( .CLK(\FIFO_U1/RegFile1/N44 ), .CN(n406) );
  CKND0 U1090 ( .CLK(\FIFO_U1/RegFile1/N45 ), .CN(n405) );
  CKND0 U1091 ( .CLK(\FIFO_U1/RegFile1/N46 ), .CN(n404) );
  CKND0 U1092 ( .CLK(\FIFO_U1/RegFile1/N47 ), .CN(n403) );
  CKND0 U1093 ( .CLK(\FIFO_U1/RegFile1/N48 ), .CN(n402) );
  CKND0 U1094 ( .CLK(\FIFO_U1/RegFile1/N49 ), .CN(n401) );
  CKND0 U1095 ( .CLK(\FIFO_U1/RegFile1/N50 ), .CN(n400) );
  CKND0 U1096 ( .CLK(\FIFO_U1/RegFile1/N51 ), .CN(n399) );
  CKND0 U1097 ( .CLK(\FIFO_U1/RegFile1/N52 ), .CN(n398) );
  CKND0 U1098 ( .CLK(\FIFO_U1/RegFile1/N53 ), .CN(n397) );
  CKND0 U1099 ( .CLK(\FIFO_U1/RegFile1/N54 ), .CN(n396) );
  CKND0 U1100 ( .CLK(\FIFO_U1/RegFile1/N55 ), .CN(n395) );
  CKND0 U1101 ( .CLK(\FIFO_U1/RegFile1/N56 ), .CN(n394) );
  CKND0 U1102 ( .CLK(\FIFO_U1/RegFile1/N57 ), .CN(n393) );
  CKND0 U1103 ( .CLK(\FIFO_U1/RegFile1/N58 ), .CN(n392) );
  CKND0 U1104 ( .CLK(\FIFO_U1/RegFile1/N59 ), .CN(n391) );
  CKND0 U1105 ( .CLK(\FIFO_U1/RegFile1/N60 ), .CN(n390) );
  CKND0 U1106 ( .CLK(\FIFO_U1/RegFile1/N61 ), .CN(n389) );
  CKND0 U1107 ( .CLK(\FIFO_U1/RegFile1/N62 ), .CN(n388) );
  CKND0 U1108 ( .CLK(\FIFO_U1/RegFile1/N63 ), .CN(n387) );
  CKND0 U1109 ( .CLK(\FIFO_U1/FIFO_SM1/N0 ), .CN(n386) );
  CKND0 U1110 ( .CLK(\FIFO_U1/FIFO_SM1/N1 ), .CN(n385) );
  CKND0 U1111 ( .CLK(\FIFO_U1/FIFO_SM1/N2 ), .CN(n384) );
  CKND0 U1112 ( .CLK(\FIFO_U1/FIFO_SM1/N3 ), .CN(n383) );
  CKND0 U1113 ( .CLK(\FIFO_U1/FIFO_SM1/N4 ), .CN(n382) );
  CKND0 U1114 ( .CLK(\FIFO_U1/FIFO_SM1/N5 ), .CN(n381) );
  CKND0 U1115 ( .CLK(\FIFO_U1/FIFO_SM1/N6 ), .CN(n380) );
  CKND0 U1116 ( .CLK(\FIFO_U1/FIFO_SM1/N7 ), .CN(n379) );
  CKND0 U1117 ( .CLK(\FIFO_U1/FIFO_SM1/N8 ), .CN(n378) );
  CKND0 U1118 ( .CLK(\FIFO_U1/FIFO_SM1/N9 ), .CN(n377) );
  AN3D0 U1119 ( .A1(\SerialRx_U1/PLL_RxU1/AdjFreq [0]), .A2(n1114), .A3(
        \SerialRx_U1/PLL_RxU1/AdjFreq [1]), .Z(\U3/U2/Z_0 ) );
  OAI22D0 U1120 ( .A1(n1115), .A2(n1116), .B1(n1117), .B2(n1118), .ZN(
        \U3/U1/Z_4 ) );
  IOA22D0 U1121 ( .B1(n1117), .B2(n1119), .A1(n1120), .A2(
        \FIFO_U1/SM_ReadAddr [3]), .ZN(\U3/U1/Z_3 ) );
  OAI22D0 U1122 ( .A1(n1115), .A2(n1121), .B1(n1117), .B2(n1122), .ZN(
        \U3/U1/Z_2 ) );
  IOA22D0 U1123 ( .B1(n1117), .B2(n1123), .A1(n1120), .A2(
        \FIFO_U1/SM_ReadAddr [1]), .ZN(\U3/U1/Z_1 ) );
  IOA22D0 U1124 ( .B1(n1117), .B2(n1124), .A1(n1120), .A2(
        \FIFO_U1/SM_ReadAddr [0]), .ZN(\U3/U1/Z_0 ) );
  CKND2D0 U1125 ( .A1(n1125), .A2(n621), .ZN(n1117) );
  MUX2ND0 U1126 ( .I0(n1126), .I1(n1127), .S(\SerialRx_U1/PLL_RxU1/AdjFreq [0]), .ZN(\SerialRx_U1/PLL_RxU1/VFO1/N54 ) );
  CKND2D0 U1127 ( .A1(\SerialRx_U1/PLL_RxU1/AdjFreq [1]), .A2(n1114), .ZN(
        n1127) );
  ND3D0 U1128 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1114) );
  OAI31D0 U1129 ( .A1(n1129), .A2(n1130), .A3(n1128), .B(n1131), .ZN(n1126) );
  CKND0 U1130 ( .CLK(\SerialRx_U1/PLL_RxU1/AdjFreq [1]), .CN(n1131) );
  ND3D0 U1131 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[2] ), .A2(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] ), .A3(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n1130) );
  AN2D0 U1132 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N14 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N21 ) );
  AN2D0 U1133 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N13 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N20 ) );
  AN2D0 U1134 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N12 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N19 ) );
  AN2D0 U1135 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N11 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N18 ) );
  AN2D0 U1136 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N10 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N17 ) );
  AN2D0 U1137 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/N9 ), .A2(n1113), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/N16 ) );
  OAI21D0 U1138 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[5] ), .A2(n1129), 
        .B(n1132), .ZN(n1113) );
  AO221D0 U1139 ( .A1(n1128), .A2(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[4] ), 
        .B1(n1129), .B2(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[5] ), .C(n1133), 
        .Z(n1132) );
  OA21D0 U1140 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[4] ), .A2(n1128), 
        .B(n1134), .Z(n1133) );
  OAI22D0 U1141 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] ), .A2(n1135), 
        .B1(n1136), .B2(n1137), .ZN(n1134) );
  IOA22D0 U1142 ( .B1(n1138), .B2(n1139), .A1(n1135), .A2(
        \SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[3] ), .ZN(n1137) );
  AOI21D0 U1143 ( .A1(n1138), .A2(n1139), .B(
        \SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[2] ), .ZN(n1136) );
  CKND0 U1144 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[2] ), .CN(n1139)
         );
  OA32D0 U1145 ( .A1(n1140), .A2(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[0] ), 
        .A3(n1141), .B1(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[1] ), .B2(n1142), 
        .Z(n1138) );
  AN2D0 U1146 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[1] ), .A2(n1142), .Z(
        n1141) );
  CKND0 U1147 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[1] ), .CN(n1142)
         );
  CKND0 U1148 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[0] ), .CN(n1140)
         );
  CKND0 U1149 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/FastDivvy[3] ), .CN(n1135) );
  CKND0 U1150 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[4] ), .CN(n1128)
         );
  CKND0 U1151 ( .CLK(\SerialRx_U1/PLL_RxU1/VFO1/DivideFactor[5] ), .CN(n1129)
         );
  AN2D0 U1152 ( .A1(\SerialRx_U1/PLL_RxU1/VFO1/WireD [5]), .A2(n621), .Z(
        \SerialRx_U1/PLL_RxU1/VFO1/FastClock ) );
  CKXOR2D0 U1153 ( .A1(n1243), .A2(n1244), .Z(\SerialRx_U1/PLL_RxU1/Comp1/N8 )
         );
  XNR2D0 U1154 ( .A1(n1143), .A2(\SerialRx_U1/PLL_RxU1/Comp1/ClockInN[0] ), 
        .ZN(\SerialRx_U1/PLL_RxU1/Comp1/N6 ) );
  OAI221D0 U1155 ( .A1(n1243), .A2(n1144), .B1(n1244), .B2(n1143), .C(n1145), 
        .ZN(\SerialRx_U1/PLL_RxU1/Comp1/N20 ) );
  IAO21D0 U1156 ( .A1(\SerialRx_U1/PLL_RxU1/Comp1/N5 ), .A2(n1244), .B(
        \SerialRx_U1/PLL_RxU1/Comp1/ClockInN[1] ), .ZN(n1144) );
  OAI22D0 U1157 ( .A1(n1243), .A2(n1145), .B1(n1244), .B2(n1146), .ZN(
        \SerialRx_U1/PLL_RxU1/Comp1/N19 ) );
  INR3D0 U1158 ( .A1(n1243), .B1(\SerialRx_U1/PLL_RxU1/Comp1/ClockInN[1] ), 
        .B2(\SerialRx_U1/PLL_RxU1/Comp1/ClockInN[0] ), .ZN(n1146) );
  CKND0 U1159 ( .CLK(\SerialRx_U1/PLL_RxU1/Comp1/N9 ), .CN(n1145) );
  NR2D0 U1160 ( .A1(n1143), .A2(\SerialRx_U1/PLL_RxU1/Comp1/N5 ), .ZN(
        \SerialRx_U1/PLL_RxU1/Comp1/N9 ) );
  CKND0 U1161 ( .CLK(\SerialRx_U1/PLL_RxU1/Comp1/ClockInN[0] ), .CN(
        \SerialRx_U1/PLL_RxU1/Comp1/N5 ) );
  CKND0 U1162 ( .CLK(\SerialRx_U1/PLL_RxU1/Comp1/ClockInN[1] ), .CN(n1143) );
  INR2D0 U1163 ( .A1(FIFO_Out[6]), .B1(n1147), .ZN(N9) );
  INR2D0 U1164 ( .A1(FIFO_Out[5]), .B1(n1147), .ZN(N8) );
  INR2D0 U1165 ( .A1(FIFO_Out[4]), .B1(n1147), .ZN(N7) );
  INR2D0 U1166 ( .A1(FIFO_Out[3]), .B1(n1147), .ZN(N6) );
  INR2D0 U1167 ( .A1(FIFO_Out[2]), .B1(n1147), .ZN(N5) );
  INR2D0 U1168 ( .A1(FIFO_Out[1]), .B1(n1147), .ZN(N4) );
  NR2D0 U1169 ( .A1(FIFOEmpty), .A2(n1147), .ZN(N35) );
  INR2D0 U1170 ( .A1(FIFO_Out[31]), .B1(n1147), .ZN(N34) );
  INR2D0 U1171 ( .A1(FIFO_Out[30]), .B1(n1147), .ZN(N33) );
  INR2D0 U1172 ( .A1(FIFO_Out[29]), .B1(n1147), .ZN(N32) );
  INR2D0 U1173 ( .A1(FIFO_Out[28]), .B1(n1147), .ZN(N31) );
  INR2D0 U1174 ( .A1(FIFO_Out[27]), .B1(n1147), .ZN(N30) );
  INR2D0 U1175 ( .A1(FIFO_Out[0]), .B1(n1147), .ZN(N3) );
  INR2D0 U1176 ( .A1(FIFO_Out[26]), .B1(n1147), .ZN(N29) );
  INR2D0 U1177 ( .A1(FIFO_Out[25]), .B1(n1147), .ZN(N28) );
  INR2D0 U1178 ( .A1(FIFO_Out[24]), .B1(n1147), .ZN(N27) );
  INR2D0 U1179 ( .A1(FIFO_Out[23]), .B1(n1147), .ZN(N26) );
  INR2D0 U1180 ( .A1(FIFO_Out[22]), .B1(n1147), .ZN(N25) );
  INR2D0 U1181 ( .A1(FIFO_Out[21]), .B1(n1147), .ZN(N24) );
  INR2D0 U1182 ( .A1(FIFO_Out[20]), .B1(n1147), .ZN(N23) );
  INR2D0 U1183 ( .A1(FIFO_Out[19]), .B1(n1147), .ZN(N22) );
  INR2D0 U1184 ( .A1(FIFO_Out[18]), .B1(n1147), .ZN(N21) );
  INR2D0 U1185 ( .A1(FIFO_Out[17]), .B1(n1147), .ZN(N20) );
  INR2D0 U1186 ( .A1(FIFO_Out[16]), .B1(n1147), .ZN(N19) );
  INR2D0 U1187 ( .A1(FIFO_Out[15]), .B1(n1147), .ZN(N18) );
  INR2D0 U1188 ( .A1(FIFO_Out[14]), .B1(n1147), .ZN(N17) );
  INR2D0 U1189 ( .A1(FIFO_Out[13]), .B1(n1147), .ZN(N16) );
  INR2D0 U1190 ( .A1(FIFO_Out[12]), .B1(n1147), .ZN(N15) );
  INR2D0 U1191 ( .A1(FIFO_Out[11]), .B1(n1147), .ZN(N14) );
  INR2D0 U1192 ( .A1(FIFO_Out[10]), .B1(n1147), .ZN(N13) );
  INR2D0 U1193 ( .A1(FIFO_Out[9]), .B1(n1147), .ZN(N12) );
  INR2D0 U1194 ( .A1(FIFO_Out[8]), .B1(n1147), .ZN(N11) );
  INR2D0 U1195 ( .A1(FIFO_Out[7]), .B1(n1147), .ZN(N10) );
  ND3D0 U1196 ( .A1(n658), .A2(n663), .A3(n647), .ZN(n1152) );
  ND3D0 U1197 ( .A1(n1165), .A2(n662), .A3(n658), .ZN(n1153) );
  ND3D0 U1198 ( .A1(n1166), .A2(n663), .A3(n651), .ZN(n1154) );
  ND3D0 U1199 ( .A1(n1165), .A2(n1166), .A3(n661), .ZN(n1155) );
  ND3D0 U1200 ( .A1(n564), .A2(n655), .A3(n649), .ZN(n1156) );
  ND3D0 U1201 ( .A1(n1165), .A2(n564), .A3(n657), .ZN(n1157) );
  CKND0 U1202 ( .CLK(n1166), .CN(\FIFO_U1/RegFile1/N76 ) );
  CKND0 U1203 ( .CLK(n1165), .CN(\FIFO_U1/RegFile1/N75 ) );
  CKND2D0 U1204 ( .A1(n419), .A2(\FIFO_U1/SM_MemWriteCmd ), .ZN(n1150) );
  CKND0 U1205 ( .CLK(\FIFO_U1/RegFile1/N79 ), .CN(n1163) );
  CKND0 U1206 ( .CLK(\FIFO_U1/SM_ReadAddr [4]), .CN(n1116) );
  MUX2ND0 U1207 ( .I0(\FIFO_U1/SM_WriteAddr [3]), .I1(\FIFO_U1/SM_ReadAddr [3]), .S(n1167), .ZN(n1161) );
  ND3D0 U1208 ( .A1(n1166), .A2(n564), .A3(n1165), .ZN(n1159) );
  MUX2ND0 U1209 ( .I0(\FIFO_U1/SM_WriteAddr [0]), .I1(\FIFO_U1/SM_ReadAddr [0]), .S(n1167), .ZN(n1165) );
  CKND0 U1210 ( .CLK(\FIFO_U1/SM_ReadAddr [2]), .CN(n1121) );
  MUX2ND0 U1211 ( .I0(\FIFO_U1/SM_WriteAddr [1]), .I1(\FIFO_U1/SM_ReadAddr [1]), .S(n1167), .ZN(n1166) );
  NR2D0 U1212 ( .A1(n1148), .A2(\FIFO_U1/SM_MemWriteCmd ), .ZN(n1167) );
  CKND0 U1213 ( .CLK(\FIFO_U1/SM_MemReadCmd ), .CN(n1148) );
  NR2D0 U1214 ( .A1(n1168), .A2(n1149), .ZN(\FIFO_U1/RegFile1/ChipClock ) );
  AOI21D0 U1215 ( .A1(n1169), .A2(n1170), .B(DecoderParClk), .ZN(
        \FIFO_U1/FIFO_SM1/N211 ) );
  AN2D0 U1216 ( .A1(\FIFO_U1/FIFO_SM1/N182 ), .A2(n1168), .Z(
        \FIFO_U1/FIFO_SM1/N210 ) );
  NR2D0 U1217 ( .A1(DecoderParClk), .A2(n1171), .ZN(\FIFO_U1/FIFO_SM1/N200 )
         );
  AOI211D0 U1218 ( .A1(n1172), .A2(n1173), .B(n1174), .C(
        \FIFO_U1/FIFO_SM1/N184 ), .ZN(n1171) );
  AN2D0 U1219 ( .A1(\FIFO_U1/FIFO_SM1/N148 ), .A2(n1168), .Z(
        \FIFO_U1/FIFO_SM1/N199 ) );
  AOI21D0 U1220 ( .A1(n1176), .A2(n1177), .B(DecoderParClk), .ZN(
        \FIFO_U1/FIFO_SM1/N189 ) );
  AOI31D0 U1221 ( .A1(n1178), .A2(n1179), .A3(n1180), .B(DecoderParClk), .ZN(
        \FIFO_U1/FIFO_SM1/N188 ) );
  NR2D0 U1222 ( .A1(n1120), .A2(n1174), .ZN(n1180) );
  CKND2D0 U1223 ( .A1(n1183), .A2(Reset), .ZN(n1177) );
  CKND0 U1224 ( .CLK(n1115), .CN(n1120) );
  CKND0 U1225 ( .CLK(n1184), .CN(n1179) );
  MUX2ND0 U1226 ( .I0(n528), .I1(n1185), .S(n529), .ZN(n1178) );
  NR2D0 U1227 ( .A1(\FIFO_U1/FIFO_SM1/CurState[1] ), .A2(n528), .ZN(n1185) );
  IND2D0 U1228 ( .A1(\FIFO_U1/FIFO_SM1/N209 ), .B1(n1186), .ZN(
        \FIFO_U1/FIFO_SM1/N185 ) );
  OAI21D0 U1229 ( .A1(n1181), .A2(n1184), .B(n1168), .ZN(n1186) );
  CKND0 U1230 ( .CLK(DecoderParClk), .CN(n1168) );
  OAI22D0 U1231 ( .A1(n1187), .A2(n1169), .B1(n1188), .B2(n1189), .ZN(n1184)
         );
  NR2D0 U1232 ( .A1(n1188), .A2(n1190), .ZN(n1181) );
  AOI211D0 U1233 ( .A1(n1191), .A2(n1175), .B(n1192), .C(n1193), .ZN(n1115) );
  OAI211D0 U1234 ( .A1(n1187), .A2(n1169), .B(n1194), .C(n1195), .ZN(
        \FIFO_U1/FIFO_SM1/N184 ) );
  NR2D0 U1235 ( .A1(n1193), .A2(n1192), .ZN(n1195) );
  NR2D0 U1236 ( .A1(n1189), .A2(n1187), .ZN(n1192) );
  NR2D0 U1237 ( .A1(n1170), .A2(n1173), .ZN(\FIFO_U1/FIFO_SM1/N182 ) );
  CKND0 U1238 ( .CLK(n1188), .CN(n1173) );
  OAI22D0 U1239 ( .A1(n1196), .A2(n1197), .B1(n1118), .B2(n1198), .ZN(
        \FIFO_U1/FIFO_SM1/N179 ) );
  CKND0 U1240 ( .CLK(\FIFO_U1/FIFO_SM1/N126 ), .CN(n1197) );
  OAI22D0 U1241 ( .A1(n1196), .A2(n1199), .B1(n1119), .B2(n1198), .ZN(
        \FIFO_U1/FIFO_SM1/N176 ) );
  CKND0 U1242 ( .CLK(\FIFO_U1/FIFO_SM1/N125 ), .CN(n1199) );
  OAI22D0 U1243 ( .A1(n1196), .A2(n1200), .B1(n1122), .B2(n1198), .ZN(
        \FIFO_U1/FIFO_SM1/N173 ) );
  CKND0 U1244 ( .CLK(\FIFO_U1/SM_WriteAddr [2]), .CN(n1122) );
  CKND0 U1245 ( .CLK(\FIFO_U1/FIFO_SM1/N124 ), .CN(n1200) );
  OAI22D0 U1246 ( .A1(n1196), .A2(n1201), .B1(n1123), .B2(n1198), .ZN(
        \FIFO_U1/FIFO_SM1/N170 ) );
  CKND0 U1247 ( .CLK(\FIFO_U1/SM_WriteAddr [1]), .CN(n1123) );
  CKND0 U1248 ( .CLK(\FIFO_U1/FIFO_SM1/N123 ), .CN(n1201) );
  OAI22D0 U1249 ( .A1(n1196), .A2(n1202), .B1(n1124), .B2(n1198), .ZN(
        \FIFO_U1/FIFO_SM1/N167 ) );
  CKND2D0 U1250 ( .A1(n1183), .A2(n621), .ZN(n1198) );
  CKND0 U1251 ( .CLK(\FIFO_U1/SM_WriteAddr [0]), .CN(n1124) );
  CKND0 U1252 ( .CLK(\FIFO_U1/FIFO_SM1/N122 ), .CN(n1202) );
  AN2D0 U1253 ( .A1(n1176), .A2(n1203), .Z(n1196) );
  CKND2D0 U1254 ( .A1(n1182), .A2(n1204), .ZN(\FIFO_U1/FIFO_SM1/N165 ) );
  OAI21D0 U1255 ( .A1(n1172), .A2(n1205), .B(n1187), .ZN(n1204) );
  AO222D0 U1256 ( .A1(\FIFO_U1/SM_ReadAddr [4]), .A2(n1175), .B1(
        \FIFO_U1/FIFO_SM1/N126 ), .B2(n1125), .C1(\FIFO_U1/FIFO_SM1/N76 ), 
        .C2(n1205), .Z(\FIFO_U1/FIFO_SM1/N162 ) );
  AO222D0 U1257 ( .A1(\FIFO_U1/SM_ReadAddr [3]), .A2(n1175), .B1(
        \FIFO_U1/FIFO_SM1/N125 ), .B2(n1125), .C1(\FIFO_U1/FIFO_SM1/N75 ), 
        .C2(n1205), .Z(\FIFO_U1/FIFO_SM1/N159 ) );
  AO222D0 U1258 ( .A1(\FIFO_U1/SM_ReadAddr [2]), .A2(n1175), .B1(
        \FIFO_U1/FIFO_SM1/N124 ), .B2(n1125), .C1(\FIFO_U1/FIFO_SM1/N74 ), 
        .C2(n1205), .Z(\FIFO_U1/FIFO_SM1/N156 ) );
  AO222D0 U1259 ( .A1(\FIFO_U1/SM_ReadAddr [1]), .A2(n1175), .B1(
        \FIFO_U1/FIFO_SM1/N123 ), .B2(n1125), .C1(\FIFO_U1/FIFO_SM1/N73 ), 
        .C2(n1205), .Z(\FIFO_U1/FIFO_SM1/N153 ) );
  AO222D0 U1260 ( .A1(\FIFO_U1/SM_ReadAddr [0]), .A2(n1175), .B1(
        \FIFO_U1/FIFO_SM1/N122 ), .B2(n1125), .C1(\FIFO_U1/FIFO_SM1/N72 ), 
        .C2(n1205), .Z(\FIFO_U1/FIFO_SM1/N150 ) );
  NR2D0 U1261 ( .A1(n1194), .A2(n1191), .ZN(\FIFO_U1/FIFO_SM1/N148 ) );
  OAI21D0 U1262 ( .A1(n1191), .A2(n1206), .B(n1194), .ZN(
        \FIFO_U1/FIFO_SM1/N146 ) );
  CKND0 U1263 ( .CLK(n1175), .CN(n1194) );
  IAO21D0 U1264 ( .A1(n1207), .A2(n1203), .B(n1172), .ZN(n1206) );
  IND4D0 U1265 ( .A1(n1193), .B1(n1189), .B2(n1182), .B3(n1208), .ZN(
        \FIFO_U1/FIFO_SM1/N144 ) );
  MAOI22D0 U1266 ( .A1(n1209), .A2(n1207), .B1(n1169), .B2(n1191), .ZN(n1208)
         );
  ND3D0 U1267 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1207) );
  NR3D0 U1268 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
  CKXOR2D0 U1269 ( .A1(\FIFO_U1/SM_ReadAddr [3]), .A2(\FIFO_U1/FIFO_SM1/N91 ), 
        .Z(n1215) );
  CKXOR2D0 U1270 ( .A1(\FIFO_U1/SM_ReadAddr [1]), .A2(\FIFO_U1/FIFO_SM1/N89 ), 
        .Z(n1214) );
  CKXOR2D0 U1271 ( .A1(\FIFO_U1/SM_ReadAddr [0]), .A2(\FIFO_U1/FIFO_SM1/N88 ), 
        .Z(n1213) );
  XNR2D0 U1272 ( .A1(\FIFO_U1/FIFO_SM1/N90 ), .A2(\FIFO_U1/SM_ReadAddr [2]), 
        .ZN(n1211) );
  XNR2D0 U1273 ( .A1(\FIFO_U1/FIFO_SM1/N92 ), .A2(\FIFO_U1/SM_ReadAddr [4]), 
        .ZN(n1210) );
  CKND0 U1274 ( .CLK(n1125), .CN(n1182) );
  NR2D0 U1275 ( .A1(n1170), .A2(n1188), .ZN(n1125) );
  CKND2D0 U1276 ( .A1(n1247), .A2(n1147), .ZN(n1188) );
  CKND0 U1277 ( .CLK(n1183), .CN(n1170) );
  NR3D0 U1278 ( .A1(n1246), .A2(n1245), .A3(\FIFO_U1/FIFO_SM1/CurState[1] ), 
        .ZN(n1183) );
  CKND0 U1279 ( .CLK(n1172), .CN(n1189) );
  NR2D0 U1280 ( .A1(n1187), .A2(n1203), .ZN(n1193) );
  CKND0 U1281 ( .CLK(n1191), .CN(n1187) );
  OAI211D0 U1282 ( .A1(n1191), .A2(n1190), .B(n1216), .C(n1176), .ZN(
        \FIFO_U1/FIFO_SM1/N142 ) );
  NR2D0 U1283 ( .A1(n1172), .A2(n1175), .ZN(n1176) );
  NR3D0 U1284 ( .A1(n528), .A2(n1217), .A3(n529), .ZN(n1175) );
  NR3D0 U1285 ( .A1(n528), .A2(\FIFO_U1/FIFO_SM1/CurState[1] ), .A3(n529), 
        .ZN(n1172) );
  OAI31D0 U1286 ( .A1(n1218), .A2(n1219), .A3(n1220), .B(n1209), .ZN(n1216) );
  XNR2D0 U1287 ( .A1(n1118), .A2(\FIFO_U1/FIFO_SM1/N109 ), .ZN(n1220) );
  CKND0 U1288 ( .CLK(\FIFO_U1/SM_WriteAddr [4]), .CN(n1118) );
  XNR2D0 U1289 ( .A1(n1119), .A2(\FIFO_U1/FIFO_SM1/N108 ), .ZN(n1219) );
  CKND0 U1290 ( .CLK(\FIFO_U1/SM_WriteAddr [3]), .CN(n1119) );
  ND3D0 U1291 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1218) );
  XNR2D0 U1292 ( .A1(\FIFO_U1/FIFO_SM1/N106 ), .A2(\FIFO_U1/SM_WriteAddr [1]), 
        .ZN(n1223) );
  XNR2D0 U1293 ( .A1(\FIFO_U1/FIFO_SM1/N107 ), .A2(\FIFO_U1/SM_WriteAddr [2]), 
        .ZN(n1222) );
  XNR2D0 U1294 ( .A1(\FIFO_U1/FIFO_SM1/N105 ), .A2(\FIFO_U1/SM_WriteAddr [0]), 
        .ZN(n1221) );
  CKND0 U1295 ( .CLK(n1205), .CN(n1190) );
  CKND2D0 U1296 ( .A1(n1203), .A2(n1169), .ZN(n1205) );
  ND3D0 U1297 ( .A1(n529), .A2(n528), .A3(\FIFO_U1/FIFO_SM1/CurState[1] ), 
        .ZN(n1169) );
  CKND0 U1298 ( .CLK(n1209), .CN(n1203) );
  NR3D0 U1299 ( .A1(n1217), .A2(n1246), .A3(n528), .ZN(n1209) );
  CKND0 U1300 ( .CLK(\FIFO_U1/FIFO_SM1/CurState[1] ), .CN(n1217) );
  NR2D0 U1301 ( .A1(n1147), .A2(n1247), .ZN(n1191) );
  INR2D0 U1302 ( .A1(\DesDecoder_U1/N53 ), .B1(n1224), .ZN(\DesDecoder_U1/N70 ) );
  CKND2D0 U1303 ( .A1(n1225), .A2(n621), .ZN(\DesDecoder_U1/N69 ) );
  INR2D0 U1304 ( .A1(\DesDecoder_U1/N52 ), .B1(n1224), .ZN(\DesDecoder_U1/N68 ) );
  INR2D0 U1305 ( .A1(\DesDecoder_U1/N51 ), .B1(n1224), .ZN(\DesDecoder_U1/N67 ) );
  NR2D0 U1306 ( .A1(n1224), .A2(n1226), .ZN(\DesDecoder_U1/N66 ) );
  NR2D0 U1307 ( .A1(n1224), .A2(n1227), .ZN(\DesDecoder_U1/N65 ) );
  NR2D0 U1308 ( .A1(DecoderParClk), .A2(n1224), .ZN(\DesDecoder_U1/N63 ) );
  IND3D0 U1309 ( .A1(n1248), .B1(n621), .B2(SerValid), .ZN(n1224) );
  OAI21D0 U1310 ( .A1(n1228), .A2(n1225), .B(n621), .ZN(\DesDecoder_U1/N62 )
         );
  CKND0 U1311 ( .CLK(Reset), .CN(n491) );
  CKND0 U1312 ( .CLK(SerValid), .CN(n1225) );
  AOI31D0 U1313 ( .A1(n1227), .A2(n1226), .A3(n1229), .B(n1248), .ZN(n1228) );
  NR3D0 U1314 ( .A1(\DesDecoder_U1/N51 ), .A2(\DesDecoder_U1/N53 ), .A3(
        \DesDecoder_U1/N52 ), .ZN(n1229) );
  CKND0 U1315 ( .CLK(\DesDecoder_U1/N50 ), .CN(n1226) );
  CKND0 U1316 ( .CLK(\DesDecoder_U1/N49 ), .CN(n1227) );
  NR2D0 U1317 ( .A1(n1230), .A2(n1231), .ZN(\DesDecoder_U1/N12 ) );
  CKND2D0 U1318 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
  NR4D0 U1319 ( .A1(\DesDecoder_U1/FrameSR[7] ), .A2(
        \DesDecoder_U1/FrameSR[6] ), .A3(\DesDecoder_U1/FrameSR[5] ), .A4(
        \DesDecoder_U1/FrameSR[4] ), .ZN(n1233) );
  NR4D0 U1320 ( .A1(\DesDecoder_U1/FrameSR[3] ), .A2(
        \DesDecoder_U1/FrameSR[2] ), .A3(\DesDecoder_U1/FrameSR[1] ), .A4(
        \DesDecoder_U1/FrameSR[0] ), .ZN(n1232) );
  NR4D0 U1321 ( .A1(n1238), .A2(\DesDecoder_U1/FrameSR[50] ), .A3(n374), .A4(
        \DesDecoder_U1/FrameSR[49] ), .ZN(n1237) );
  ND3D0 U1322 ( .A1(\DesDecoder_U1/FrameSR[52] ), .A2(
        \DesDecoder_U1/FrameSR[51] ), .A3(\DesDecoder_U1/FrameSR[36] ), .ZN(
        n1238) );
  NR4D0 U1323 ( .A1(n1239), .A2(\DesDecoder_U1/FrameSR[21] ), .A3(
        \DesDecoder_U1/FrameSR[33] ), .A4(\DesDecoder_U1/FrameSR[20] ), .ZN(
        n1236) );
  ND3D0 U1324 ( .A1(n360), .A2(n356), .A3(n361), .ZN(n1239) );
  NR4D0 U1325 ( .A1(n1240), .A2(\DesDecoder_U1/FrameSR[39] ), .A3(
        \DesDecoder_U1/FrameSR[54] ), .A4(\DesDecoder_U1/FrameSR[37] ), .ZN(
        n1235) );
  ND3D0 U1326 ( .A1(n1253), .A2(n368), .A3(n1252), .ZN(n1240) );
  NR4D0 U1327 ( .A1(n1241), .A2(\DesDecoder_U1/FrameSR[17] ), .A3(
        \DesDecoder_U1/FrameSR[23] ), .A4(\DesDecoder_U1/FrameSR[16] ), .ZN(
        n1234) );
  ND3D0 U1328 ( .A1(n1250), .A2(n1251), .A3(n1249), .ZN(n1241) );
endmodule


module Deserializer_DW01_incdec_0 ( A, INC_DEC, SUM );
  input [5:0] A;
  output [5:0] SUM;
  input INC_DEC;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[1] ,
         \carry[0] ;

  XOR3D1 U1_5 ( .A1(A[5]), .A2(INC_DEC), .A3(\carry[5] ), .Z(SUM[5]) );
  FA1D0 U1_2 ( .A(A[2]), .B(INC_DEC), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  FA1D0 U1_3 ( .A(A[3]), .B(INC_DEC), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  FA1D0 U1_4 ( .A(A[4]), .B(INC_DEC), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  FA1D0 U1_1 ( .A(A[1]), .B(INC_DEC), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  FA1D0 U1_0 ( .A(A[0]), .B(INC_DEC), .CI(\carry[0] ), .CO(\carry[1] ), .S(
        SUM[0]) );
  CKND0 U1 ( .CLK(INC_DEC), .CN(\carry[0] ) );
endmodule


module Deserializer_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_3 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_4 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_5 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module Deserializer_DW01_inc_6 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

