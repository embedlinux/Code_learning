
module DesDecoder ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, Reset
 );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   n3149, SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41,
         N42, N43, N47, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n60, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n298,
         n299, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3009, n3011, n3013, n3015, n3017, n3019,
         n3021, n3023, n3025, n3027, n3029, n3031, n3033, n3035, n3037, n3039,
         n3041, n3043, n3045, n3047, n3049, n3051, n3053, n3055, n3057, n3059,
         n3061, n3063, n3065, n3067, n3069, n3071, n3073, n3074, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148;
  wire   [3:0] ParValidTimer;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  OA21D1 U131 ( .A1(n58), .A2(n298), .B(n2432), .Z(N43) );
  OR2D1 U133 ( .A1(n2364), .A2(n2418), .Z(n60) );
  DesDecoder_DW01_inc_0 \ClkGen/add_204  ( .A({Count32[4:2], n2364, n2418}), 
        .SUM({N34, N33, N32, N31, N30}) );
  EDFCNQD1 ParClkr_reg ( .D(n301), .E(n306), .CP(SerClock), .CDN(n3134), .Q(
        n3149) );
  DFNCND1 \FrameSR_reg[51]  ( .D(n321), .CPN(n3145), .CDN(n261), .Q(
        FrameSR[51]), .QN(n140) );
  DFNCND1 \FrameSR_reg[52]  ( .D(n339), .CPN(n3145), .CDN(n3138), .Q(
        FrameSR[52]), .QN(n139) );
  DFNCND1 \FrameSR_reg[36]  ( .D(n357), .CPN(n3146), .CDN(n3140), .Q(
        FrameSR[36]), .QN(n155) );
  DFNCND1 \FrameSR_reg[16]  ( .D(n375), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[16]), .QN(n175) );
  DFNCND1 \FrameSR_reg[23]  ( .D(n393), .CPN(n3147), .CDN(n3135), .Q(
        FrameSR[23]), .QN(n168) );
  DFNCND1 \FrameSR_reg[38]  ( .D(n411), .CPN(n3146), .CDN(n261), .Q(
        FrameSR[38]), .QN(n153) );
  DFNCND1 \FrameSR_reg[54]  ( .D(n429), .CPN(n3144), .CDN(n261), .Q(
        FrameSR[54]), .QN(n137) );
  DFNCND1 \FrameSR_reg[17]  ( .D(n447), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[17]), .QN(n174) );
  DFNCND1 \FrameSR_reg[32]  ( .D(n465), .CPN(n3146), .CDN(n3136), .Q(
        FrameSR[32]), .QN(n159) );
  DFNCND1 \FrameSR_reg[39]  ( .D(n483), .CPN(n3146), .CDN(n3139), .Q(
        FrameSR[39]), .QN(n152) );
  DFNCND1 \FrameSR_reg[55]  ( .D(n501), .CPN(n3144), .CDN(n3139), .Q(
        FrameSR[55]), .QN(n136) );
  DFNCND1 \FrameSR_reg[8]  ( .D(n519), .CPN(n3146), .CDN(n3134), .Q(FrameSR[8]), .QN(n183) );
  DFNCND1 \FrameSR_reg[9]  ( .D(n536), .CPN(n3148), .CDN(n3134), .Q(FrameSR[9]), .QN(n182) );
  DFNCND1 \FrameSR_reg[10]  ( .D(n555), .CPN(n3148), .CDN(n3134), .Q(
        FrameSR[10]), .QN(n181) );
  DFNCND1 \FrameSR_reg[11]  ( .D(n573), .CPN(n3148), .CDN(n3134), .Q(
        FrameSR[11]), .QN(n180) );
  DFNCND1 \FrameSR_reg[12]  ( .D(n591), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[12]), .QN(n179) );
  DFNCND1 \FrameSR_reg[13]  ( .D(n609), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[13]), .QN(n178) );
  DFNCND1 \FrameSR_reg[14]  ( .D(n627), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[14]), .QN(n177) );
  DFNCND1 \FrameSR_reg[15]  ( .D(n645), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[15]), .QN(n176) );
  DFNCND1 \FrameSR_reg[24]  ( .D(n663), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[24]), .QN(n167) );
  DFNCND1 \FrameSR_reg[25]  ( .D(n681), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[25]), .QN(n166) );
  DFNCND1 \FrameSR_reg[26]  ( .D(n699), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[26]), .QN(n165) );
  DFNCND1 \FrameSR_reg[27]  ( .D(n717), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[27]), .QN(n164) );
  DFNCND1 \FrameSR_reg[28]  ( .D(n735), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[28]), .QN(n163) );
  DFNCND1 \FrameSR_reg[29]  ( .D(n753), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[29]), .QN(n162) );
  DFNCND1 \FrameSR_reg[30]  ( .D(n771), .CPN(n3147), .CDN(n3136), .Q(
        FrameSR[30]), .QN(n161) );
  DFNCND1 \FrameSR_reg[31]  ( .D(n789), .CPN(n3146), .CDN(n3136), .Q(
        FrameSR[31]), .QN(n160) );
  DFNCND1 \FrameSR_reg[40]  ( .D(n807), .CPN(n3146), .CDN(n261), .Q(
        FrameSR[40]), .QN(n151) );
  DFNCND1 \FrameSR_reg[41]  ( .D(n825), .CPN(n3146), .CDN(n3140), .Q(
        FrameSR[41]), .QN(n150) );
  DFNCND1 \FrameSR_reg[42]  ( .D(n843), .CPN(n3145), .CDN(n261), .Q(
        FrameSR[42]), .QN(n149) );
  DFNCND1 \FrameSR_reg[43]  ( .D(n861), .CPN(n3145), .CDN(n3139), .Q(
        FrameSR[43]), .QN(n148) );
  DFNCND1 \FrameSR_reg[44]  ( .D(n879), .CPN(n3145), .CDN(n3139), .Q(
        FrameSR[44]), .QN(n147) );
  DFNCND1 \FrameSR_reg[45]  ( .D(n897), .CPN(n3145), .CDN(n3140), .Q(
        FrameSR[45]), .QN(n146) );
  DFNCND1 \FrameSR_reg[46]  ( .D(n915), .CPN(n3145), .CDN(n261), .Q(
        FrameSR[46]), .QN(n145) );
  DFNCND1 \FrameSR_reg[47]  ( .D(n933), .CPN(n3145), .CDN(n3139), .Q(
        FrameSR[47]), .QN(n144) );
  DFNCND1 \FrameSR_reg[56]  ( .D(n951), .CPN(n3144), .CDN(n3136), .Q(
        FrameSR[56]), .QN(n135) );
  DFNCND1 \FrameSR_reg[57]  ( .D(n969), .CPN(n3144), .CDN(n3136), .Q(
        FrameSR[57]), .QN(n134) );
  DFNCND1 \FrameSR_reg[58]  ( .D(n987), .CPN(n3144), .CDN(n3140), .Q(
        FrameSR[58]), .QN(n133) );
  DFNCND1 \FrameSR_reg[59]  ( .D(n1005), .CPN(n3144), .CDN(n261), .Q(
        FrameSR[59]), .QN(n132) );
  DFNCND1 \FrameSR_reg[60]  ( .D(n1023), .CPN(n3144), .CDN(n3135), .Q(
        FrameSR[60]), .QN(n131) );
  DFNCND1 \FrameSR_reg[61]  ( .D(n1041), .CPN(n3144), .CDN(n3137), .Q(
        FrameSR[61]), .QN(n130) );
  DFNCND1 \FrameSR_reg[62]  ( .D(n1059), .CPN(n3144), .CDN(n3139), .Q(
        FrameSR[62]), .QN(n129) );
  DFNCND1 \FrameSR_reg[63]  ( .D(n1077), .CPN(n3144), .CDN(n3134), .QN(n128)
         );
  DFNCND1 \FrameSR_reg[22]  ( .D(n1095), .CPN(n3147), .CDN(n3135), .Q(
        FrameSR[22]), .QN(n169) );
  DFNCND1 \FrameSR_reg[37]  ( .D(n1113), .CPN(n3146), .CDN(n3139), .Q(
        FrameSR[37]), .QN(n154) );
  DFNCND1 \FrameSR_reg[53]  ( .D(n1131), .CPN(n3144), .CDN(n3139), .Q(
        FrameSR[53]), .QN(n138) );
  DFNCND1 \Decoder_reg[31]  ( .D(n1149), .CPN(n3148), .CDN(n3139), .QN(n13) );
  DFNCND1 \Decoder_reg[30]  ( .D(n1166), .CPN(n3143), .CDN(n3137), .QN(n14) );
  DFNCND1 \Decoder_reg[29]  ( .D(n1183), .CPN(n3143), .CDN(n3140), .QN(n15) );
  DFNCND1 \Decoder_reg[28]  ( .D(n1200), .CPN(n3142), .CDN(n261), .QN(n16) );
  DFNCND1 \Decoder_reg[27]  ( .D(n1217), .CPN(n3143), .CDN(n3139), .QN(n17) );
  DFNCND1 \Decoder_reg[26]  ( .D(n1234), .CPN(n3142), .CDN(n261), .QN(n18) );
  DFNCND1 \Decoder_reg[25]  ( .D(n1251), .CPN(n3142), .CDN(n3140), .QN(n19) );
  DFNCND1 \Decoder_reg[24]  ( .D(n1268), .CPN(SerClock), .CDN(n3140), .QN(n20)
         );
  DFNCND1 \Decoder_reg[23]  ( .D(n1285), .CPN(n3142), .CDN(n261), .QN(n21) );
  DFNCND1 \Decoder_reg[22]  ( .D(n1302), .CPN(n3143), .CDN(n3137), .QN(n22) );
  DFNCND1 \Decoder_reg[21]  ( .D(n1319), .CPN(n3142), .CDN(n3134), .QN(n23) );
  DFNCND1 \Decoder_reg[20]  ( .D(n1336), .CPN(n3142), .CDN(n3135), .QN(n24) );
  DFNCND1 \Decoder_reg[19]  ( .D(n1353), .CPN(n3148), .CDN(n3138), .QN(n25) );
  DFNCND1 \Decoder_reg[18]  ( .D(n1370), .CPN(n3143), .CDN(n3136), .QN(n26) );
  DFNCND1 \Decoder_reg[17]  ( .D(n1387), .CPN(n3147), .CDN(n3140), .QN(n27) );
  DFNCND1 \Decoder_reg[16]  ( .D(n1404), .CPN(SerClock), .CDN(n3139), .QN(n28)
         );
  DFNCND1 \Decoder_reg[15]  ( .D(n1420), .CPN(n3143), .CDN(n261), .QN(n29) );
  DFNCND1 \Decoder_reg[14]  ( .D(n1436), .CPN(n3142), .CDN(n3137), .QN(n30) );
  DFNCND1 \Decoder_reg[13]  ( .D(n1453), .CPN(n3144), .CDN(n3135), .QN(n31) );
  DFNCND1 \Decoder_reg[12]  ( .D(n1469), .CPN(n3146), .CDN(n3138), .QN(n32) );
  DFNCND1 \Decoder_reg[11]  ( .D(n1486), .CPN(SerClock), .CDN(n3137), .QN(n33)
         );
  DFNCND1 \Decoder_reg[10]  ( .D(n1502), .CPN(n3143), .CDN(n3137), .QN(n34) );
  DFNCND1 \Decoder_reg[9]  ( .D(n1518), .CPN(n3143), .CDN(n3137), .QN(n35) );
  DFNCND1 \Decoder_reg[8]  ( .D(n1534), .CPN(n3142), .CDN(n3137), .QN(n36) );
  DFNCND1 \Decoder_reg[7]  ( .D(n1551), .CPN(n3145), .CDN(n3137), .QN(n37) );
  DFNCND1 \Decoder_reg[6]  ( .D(n1567), .CPN(SerClock), .CDN(n3137), .QN(n38)
         );
  DFNCND1 \Decoder_reg[5]  ( .D(n1583), .CPN(n3146), .CDN(n3137), .QN(n39) );
  DFNCND1 \Decoder_reg[4]  ( .D(n1600), .CPN(SerClock), .CDN(n3137), .QN(n40)
         );
  DFNCND1 \Decoder_reg[3]  ( .D(n1616), .CPN(n3143), .CDN(n3137), .QN(n41) );
  DFNCND1 \Decoder_reg[2]  ( .D(n1632), .CPN(n3142), .CDN(n3137), .QN(n42) );
  DFNCND1 \Decoder_reg[1]  ( .D(n1649), .CPN(n3147), .CDN(n3137), .QN(n43) );
  DFNCND1 \Decoder_reg[0]  ( .D(n1666), .CPN(n3144), .CDN(n3137), .QN(n44) );
  EDFCNQD1 \Count32_reg[4]  ( .D(n1683), .E(n2432), .CP(n3143), .CDN(n3138), 
        .Q(Count32[4]) );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n1697), .CPN(n3146), .CDN(n261), .QN(
        n262) );
  DFNCND1 \FrameSR_reg[0]  ( .D(n1710), .CPN(n3146), .CDN(n3134), .Q(
        FrameSR[0]) );
  DFNCND1 \FrameSR_reg[4]  ( .D(n2040), .CPN(n3147), .CDN(n3134), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(n2057), .CPN(n3147), .CDN(n3135), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(n2075), .CPN(n3146), .CDN(n3136), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(n2093), .CPN(n3145), .CDN(n3134), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(n2111), .CPN(n3144), .CDN(n3134), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(n2129), .CPN(n3147), .CDN(n3134), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(n2147), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(n2165), .CPN(n3146), .CDN(n3136), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(n2183), .CPN(n3145), .CDN(n3137), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(n2201), .CPN(n3143), .CDN(n3134), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(n2219), .CPN(n3142), .CDN(n3134), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(n2237), .CPN(n3148), .CDN(n3134), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(n2255), .CPN(SerClock), .CDN(n3134), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(n2273), .CPN(n3147), .CDN(n3135), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(n2291), .CPN(n3146), .CDN(n3136), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(n2309), .CPN(n3145), .CDN(n3140), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(n2327), .CPN(n3148), .CDN(n3135), .Q(
        FrameSR[19]) );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n2345), .CPN(n3148), .CDN(n3140), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(n2359), .E(n2432), .CP(n3143), .CDN(n3135), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n2373), .CPN(n3142), .CDN(n3139), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(n2386), .E(n2432), .CP(n3145), .CDN(n3140), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(n2401), .E(n2432), .CP(SerClock), .CDN(n3139), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(n2416), .E(n2432), .CP(n3144), .CDN(n3136), 
        .Q(Count32[0]) );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n2446), .CPN(n3147), .CDN(n3136), .QN(
        n264) );
  DFNCND1 UnLoad_reg ( .D(n2464), .CPN(SerClock), .CDN(n261), .Q(n299), .QN(
        n263) );
  DFNCND1 doParSync_reg ( .D(n2465), .CPN(SerClock), .CDN(n3139), .Q(n298), 
        .QN(n2) );
  DFNCND1 ParValidr_reg ( .D(n2480), .CPN(n3143), .CDN(n3138), .QN(n3098) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n2495), .CPN(n3145), .CDN(n3140), .QN(n3099)
         );
  DFNCND1 \ParOutr_reg[1]  ( .D(n2511), .CPN(n3144), .CDN(n3137), .QN(n3100)
         );
  DFNCND1 \ParOutr_reg[2]  ( .D(n2527), .CPN(n3142), .CDN(n3136), .QN(n3101)
         );
  DFNCND1 \ParOutr_reg[3]  ( .D(n2543), .CPN(n3146), .CDN(n3138), .QN(n3102)
         );
  DFNCND1 \ParOutr_reg[4]  ( .D(n2559), .CPN(SerClock), .CDN(n3135), .QN(n3103) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n2575), .CPN(n3143), .CDN(n3134), .QN(n3104)
         );
  DFNCND1 \ParOutr_reg[6]  ( .D(n2591), .CPN(SerClock), .CDN(n3140), .QN(n3105) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n2607), .CPN(n3142), .CDN(n261), .QN(n3106) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n2623), .CPN(n3145), .CDN(n3139), .QN(n3107)
         );
  DFNCND1 \ParOutr_reg[9]  ( .D(n2639), .CPN(n3146), .CDN(n3139), .QN(n3108)
         );
  DFNCND1 \ParOutr_reg[10]  ( .D(n2655), .CPN(n3147), .CDN(n3138), .QN(n3109)
         );
  DFNCND1 \ParOutr_reg[11]  ( .D(n2671), .CPN(n3142), .CDN(n3138), .QN(n3110)
         );
  DFNCND1 \ParOutr_reg[12]  ( .D(n2687), .CPN(SerClock), .CDN(n3138), .QN(
        n3111) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n2703), .CPN(SerClock), .CDN(n3138), .QN(
        n3112) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n2719), .CPN(n3142), .CDN(n3138), .QN(n3113)
         );
  DFNCND1 \ParOutr_reg[15]  ( .D(n2735), .CPN(n3148), .CDN(n3138), .QN(n3114)
         );
  DFNCND1 \ParOutr_reg[16]  ( .D(n2751), .CPN(n3147), .CDN(n3138), .QN(n3115)
         );
  DFNCND1 \ParOutr_reg[17]  ( .D(n2767), .CPN(n3146), .CDN(n3138), .QN(n3116)
         );
  DFNCND1 \ParOutr_reg[18]  ( .D(n2783), .CPN(n3145), .CDN(n3138), .QN(n3117)
         );
  DFNCND1 \ParOutr_reg[19]  ( .D(n2799), .CPN(n3148), .CDN(n3138), .QN(n3118)
         );
  DFNCND1 \ParOutr_reg[20]  ( .D(n2815), .CPN(n3144), .CDN(n3138), .QN(n3119)
         );
  DFNCND1 \ParOutr_reg[21]  ( .D(n2831), .CPN(n3148), .CDN(n3138), .QN(n3120)
         );
  DFNCND1 \ParOutr_reg[22]  ( .D(n2847), .CPN(n3143), .CDN(n3140), .QN(n3121)
         );
  DFNCND1 \ParOutr_reg[23]  ( .D(n2863), .CPN(SerClock), .CDN(n3135), .QN(
        n3122) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n2879), .CPN(n3145), .CDN(n3139), .QN(n3123)
         );
  DFNCND1 \ParOutr_reg[25]  ( .D(n2895), .CPN(n3143), .CDN(n261), .QN(n3124)
         );
  DFNCND1 \ParOutr_reg[26]  ( .D(n2911), .CPN(n3144), .CDN(n261), .QN(n3125)
         );
  DFNCND1 \ParOutr_reg[27]  ( .D(n2927), .CPN(n3143), .CDN(n3140), .QN(n3126)
         );
  DFNCND1 \ParOutr_reg[28]  ( .D(n2943), .CPN(n3145), .CDN(n3134), .QN(n3127)
         );
  DFNCND1 \ParOutr_reg[29]  ( .D(n2959), .CPN(n3142), .CDN(n3139), .QN(n3128)
         );
  DFNCND1 \ParOutr_reg[30]  ( .D(n2975), .CPN(n3148), .CDN(n3140), .QN(n3129)
         );
  DFNCND1 \ParOutr_reg[31]  ( .D(n2991), .CPN(n3147), .CDN(n261), .QN(n3130)
         );
  CKBD0 U141 ( .CLK(n1405), .C(n1419) );
  CKBD0 U142 ( .CLK(n1629), .C(n1628) );
  CKBD0 U143 ( .CLK(n1421), .C(n1435) );
  CKBD0 U144 ( .CLK(n1609), .C(n1608) );
  CKBD0 U145 ( .CLK(n1454), .C(n1468) );
  CKBD0 U146 ( .CLK(n1579), .C(n1578) );
  CKBD0 U147 ( .CLK(n1566), .C(n1565) );
  CKBD0 U148 ( .CLK(n1529), .C(n1528) );
  CKBD0 U149 ( .CLK(n1516), .C(n1515) );
  CKBD0 U150 ( .CLK(n240), .C(n1487) );
  IND2D1 U151 ( .A1(n46), .B1(n47), .ZN(n45) );
  XOR2D0 U152 ( .A1(n2444), .A2(n9), .Z(n8) );
  CKBD0 U153 ( .CLK(n2347), .C(n2345) );
  CKBD0 U154 ( .CLK(n2481), .C(n2480) );
  CKBD0 U155 ( .CLK(n2992), .C(n3006) );
  CKBD0 U156 ( .CLK(n2680), .C(n2679) );
  NR2D1 U157 ( .A1(n47), .A2(n46), .ZN(N47) );
  CKNXD12 U158 ( .I(n3071), .ZN(n3073) );
  CKNXD16 U159 ( .I(n2492), .ZN(ParValid) );
  BUFFD0 U160 ( .I(N37), .Z(n301) );
  BUFFD0 U161 ( .I(n303), .Z(n302) );
  BUFFD0 U162 ( .I(n304), .Z(n303) );
  BUFFD0 U163 ( .I(n305), .Z(n304) );
  BUFFD0 U164 ( .I(n3073), .Z(n305) );
  NR2XD0 U165 ( .A1(n302), .A2(n298), .ZN(N37) );
  BUFFD0 U166 ( .I(n307), .Z(n306) );
  BUFFD0 U167 ( .I(n308), .Z(n307) );
  BUFFD0 U168 ( .I(n309), .Z(n308) );
  BUFFD0 U169 ( .I(n310), .Z(n309) );
  BUFFD0 U170 ( .I(n311), .Z(n310) );
  BUFFD0 U171 ( .I(n312), .Z(n311) );
  BUFFD0 U172 ( .I(n313), .Z(n312) );
  BUFFD0 U173 ( .I(n314), .Z(n313) );
  BUFFD0 U174 ( .I(n315), .Z(n314) );
  BUFFD0 U175 ( .I(n316), .Z(n315) );
  BUFFD0 U176 ( .I(n317), .Z(n316) );
  BUFFD0 U177 ( .I(n318), .Z(n317) );
  BUFFD0 U178 ( .I(n319), .Z(n318) );
  BUFFD0 U179 ( .I(n320), .Z(n319) );
  BUFFD0 U180 ( .I(N43), .Z(n320) );
  BUFFD0 U181 ( .I(n322), .Z(n321) );
  BUFFD0 U182 ( .I(n323), .Z(n322) );
  BUFFD0 U183 ( .I(n324), .Z(n323) );
  BUFFD0 U184 ( .I(n325), .Z(n324) );
  BUFFD0 U185 ( .I(n326), .Z(n325) );
  BUFFD0 U186 ( .I(n327), .Z(n326) );
  BUFFD0 U187 ( .I(n328), .Z(n327) );
  BUFFD0 U188 ( .I(n329), .Z(n328) );
  BUFFD0 U189 ( .I(n330), .Z(n329) );
  BUFFD0 U190 ( .I(n331), .Z(n330) );
  BUFFD0 U191 ( .I(n332), .Z(n331) );
  BUFFD0 U192 ( .I(n333), .Z(n332) );
  BUFFD0 U193 ( .I(n334), .Z(n333) );
  BUFFD0 U194 ( .I(n335), .Z(n334) );
  BUFFD0 U195 ( .I(n336), .Z(n335) );
  BUFFD0 U196 ( .I(n337), .Z(n336) );
  BUFFD0 U197 ( .I(n338), .Z(n337) );
  BUFFD0 U198 ( .I(FrameSR[50]), .Z(n338) );
  CKBD0 U199 ( .CLK(FrameSR[51]), .C(n356) );
  BUFFD0 U200 ( .I(n340), .Z(n339) );
  BUFFD0 U201 ( .I(n341), .Z(n340) );
  BUFFD0 U202 ( .I(n342), .Z(n341) );
  BUFFD0 U203 ( .I(n343), .Z(n342) );
  BUFFD0 U204 ( .I(n344), .Z(n343) );
  BUFFD0 U205 ( .I(n345), .Z(n344) );
  BUFFD0 U206 ( .I(n346), .Z(n345) );
  BUFFD0 U207 ( .I(n347), .Z(n346) );
  BUFFD0 U208 ( .I(n348), .Z(n347) );
  BUFFD0 U209 ( .I(n349), .Z(n348) );
  BUFFD0 U210 ( .I(n350), .Z(n349) );
  BUFFD0 U211 ( .I(n351), .Z(n350) );
  BUFFD0 U212 ( .I(n352), .Z(n351) );
  BUFFD0 U213 ( .I(n353), .Z(n352) );
  BUFFD0 U214 ( .I(n354), .Z(n353) );
  BUFFD0 U215 ( .I(n355), .Z(n354) );
  BUFFD0 U216 ( .I(n356), .Z(n355) );
  BUFFD0 U217 ( .I(n358), .Z(n357) );
  BUFFD0 U218 ( .I(n359), .Z(n358) );
  BUFFD0 U219 ( .I(n360), .Z(n359) );
  BUFFD0 U220 ( .I(n361), .Z(n360) );
  BUFFD0 U221 ( .I(n362), .Z(n361) );
  BUFFD0 U222 ( .I(n363), .Z(n362) );
  BUFFD0 U223 ( .I(n364), .Z(n363) );
  BUFFD0 U224 ( .I(n365), .Z(n364) );
  BUFFD0 U225 ( .I(n366), .Z(n365) );
  BUFFD0 U226 ( .I(n367), .Z(n366) );
  BUFFD0 U227 ( .I(n368), .Z(n367) );
  BUFFD0 U228 ( .I(n369), .Z(n368) );
  BUFFD0 U229 ( .I(n370), .Z(n369) );
  BUFFD0 U230 ( .I(n371), .Z(n370) );
  BUFFD0 U231 ( .I(n372), .Z(n371) );
  BUFFD0 U232 ( .I(n373), .Z(n372) );
  BUFFD0 U233 ( .I(n374), .Z(n373) );
  BUFFD0 U234 ( .I(FrameSR[35]), .Z(n374) );
  CKBD0 U235 ( .CLK(FrameSR[15]), .C(n392) );
  BUFFD0 U236 ( .I(n376), .Z(n375) );
  BUFFD0 U237 ( .I(n377), .Z(n376) );
  BUFFD0 U238 ( .I(n378), .Z(n377) );
  BUFFD0 U239 ( .I(n379), .Z(n378) );
  BUFFD0 U240 ( .I(n380), .Z(n379) );
  BUFFD0 U241 ( .I(n381), .Z(n380) );
  BUFFD0 U242 ( .I(n382), .Z(n381) );
  BUFFD0 U243 ( .I(n383), .Z(n382) );
  BUFFD0 U244 ( .I(n384), .Z(n383) );
  BUFFD0 U245 ( .I(n385), .Z(n384) );
  BUFFD0 U246 ( .I(n386), .Z(n385) );
  BUFFD0 U247 ( .I(n387), .Z(n386) );
  BUFFD0 U248 ( .I(n388), .Z(n387) );
  BUFFD0 U249 ( .I(n389), .Z(n388) );
  BUFFD0 U250 ( .I(n390), .Z(n389) );
  BUFFD0 U251 ( .I(n391), .Z(n390) );
  BUFFD0 U252 ( .I(n392), .Z(n391) );
  CKBD0 U253 ( .CLK(FrameSR[22]), .C(n410) );
  BUFFD0 U254 ( .I(n394), .Z(n393) );
  BUFFD0 U255 ( .I(n395), .Z(n394) );
  BUFFD0 U256 ( .I(n396), .Z(n395) );
  BUFFD0 U257 ( .I(n397), .Z(n396) );
  BUFFD0 U258 ( .I(n398), .Z(n397) );
  BUFFD0 U259 ( .I(n399), .Z(n398) );
  BUFFD0 U260 ( .I(n400), .Z(n399) );
  BUFFD0 U261 ( .I(n401), .Z(n400) );
  BUFFD0 U262 ( .I(n402), .Z(n401) );
  BUFFD0 U263 ( .I(n403), .Z(n402) );
  BUFFD0 U264 ( .I(n404), .Z(n403) );
  BUFFD0 U265 ( .I(n405), .Z(n404) );
  BUFFD0 U266 ( .I(n406), .Z(n405) );
  BUFFD0 U267 ( .I(n407), .Z(n406) );
  BUFFD0 U268 ( .I(n408), .Z(n407) );
  BUFFD0 U269 ( .I(n409), .Z(n408) );
  BUFFD0 U270 ( .I(n410), .Z(n409) );
  CKBD0 U271 ( .CLK(FrameSR[37]), .C(n428) );
  BUFFD0 U272 ( .I(n412), .Z(n411) );
  BUFFD0 U273 ( .I(n413), .Z(n412) );
  BUFFD0 U274 ( .I(n414), .Z(n413) );
  BUFFD0 U275 ( .I(n415), .Z(n414) );
  BUFFD0 U276 ( .I(n416), .Z(n415) );
  BUFFD0 U277 ( .I(n417), .Z(n416) );
  BUFFD0 U278 ( .I(n418), .Z(n417) );
  BUFFD0 U279 ( .I(n419), .Z(n418) );
  BUFFD0 U280 ( .I(n420), .Z(n419) );
  BUFFD0 U281 ( .I(n421), .Z(n420) );
  BUFFD0 U282 ( .I(n422), .Z(n421) );
  BUFFD0 U283 ( .I(n423), .Z(n422) );
  BUFFD0 U284 ( .I(n424), .Z(n423) );
  BUFFD0 U285 ( .I(n425), .Z(n424) );
  BUFFD0 U286 ( .I(n426), .Z(n425) );
  BUFFD0 U287 ( .I(n427), .Z(n426) );
  BUFFD0 U288 ( .I(n428), .Z(n427) );
  CKBD0 U289 ( .CLK(FrameSR[53]), .C(n446) );
  BUFFD0 U290 ( .I(n430), .Z(n429) );
  BUFFD0 U291 ( .I(n431), .Z(n430) );
  BUFFD0 U292 ( .I(n432), .Z(n431) );
  BUFFD0 U293 ( .I(n433), .Z(n432) );
  BUFFD0 U294 ( .I(n434), .Z(n433) );
  BUFFD0 U295 ( .I(n435), .Z(n434) );
  BUFFD0 U296 ( .I(n436), .Z(n435) );
  BUFFD0 U297 ( .I(n437), .Z(n436) );
  BUFFD0 U298 ( .I(n438), .Z(n437) );
  BUFFD0 U299 ( .I(n439), .Z(n438) );
  BUFFD0 U300 ( .I(n440), .Z(n439) );
  BUFFD0 U301 ( .I(n441), .Z(n440) );
  BUFFD0 U302 ( .I(n442), .Z(n441) );
  BUFFD0 U303 ( .I(n443), .Z(n442) );
  BUFFD0 U304 ( .I(n444), .Z(n443) );
  BUFFD0 U305 ( .I(n445), .Z(n444) );
  BUFFD0 U306 ( .I(n446), .Z(n445) );
  CKBD0 U307 ( .CLK(FrameSR[16]), .C(n464) );
  BUFFD0 U308 ( .I(n448), .Z(n447) );
  BUFFD0 U309 ( .I(n449), .Z(n448) );
  BUFFD0 U310 ( .I(n450), .Z(n449) );
  BUFFD0 U311 ( .I(n451), .Z(n450) );
  BUFFD0 U312 ( .I(n452), .Z(n451) );
  BUFFD0 U313 ( .I(n453), .Z(n452) );
  BUFFD0 U314 ( .I(n454), .Z(n453) );
  BUFFD0 U315 ( .I(n455), .Z(n454) );
  BUFFD0 U316 ( .I(n456), .Z(n455) );
  BUFFD0 U317 ( .I(n457), .Z(n456) );
  BUFFD0 U318 ( .I(n458), .Z(n457) );
  BUFFD0 U319 ( .I(n459), .Z(n458) );
  BUFFD0 U320 ( .I(n460), .Z(n459) );
  BUFFD0 U321 ( .I(n461), .Z(n460) );
  BUFFD0 U322 ( .I(n462), .Z(n461) );
  BUFFD0 U323 ( .I(n463), .Z(n462) );
  BUFFD0 U324 ( .I(n464), .Z(n463) );
  CKBD0 U325 ( .CLK(FrameSR[31]), .C(n482) );
  BUFFD0 U326 ( .I(n466), .Z(n465) );
  BUFFD0 U327 ( .I(n467), .Z(n466) );
  BUFFD0 U328 ( .I(n468), .Z(n467) );
  BUFFD0 U329 ( .I(n469), .Z(n468) );
  BUFFD0 U330 ( .I(n470), .Z(n469) );
  BUFFD0 U331 ( .I(n471), .Z(n470) );
  BUFFD0 U332 ( .I(n472), .Z(n471) );
  BUFFD0 U333 ( .I(n473), .Z(n472) );
  BUFFD0 U334 ( .I(n474), .Z(n473) );
  BUFFD0 U335 ( .I(n475), .Z(n474) );
  BUFFD0 U336 ( .I(n476), .Z(n475) );
  BUFFD0 U337 ( .I(n477), .Z(n476) );
  BUFFD0 U338 ( .I(n478), .Z(n477) );
  BUFFD0 U339 ( .I(n479), .Z(n478) );
  BUFFD0 U340 ( .I(n480), .Z(n479) );
  BUFFD0 U341 ( .I(n481), .Z(n480) );
  BUFFD0 U342 ( .I(n482), .Z(n481) );
  CKBD0 U343 ( .CLK(FrameSR[38]), .C(n500) );
  BUFFD0 U344 ( .I(n484), .Z(n483) );
  BUFFD0 U345 ( .I(n485), .Z(n484) );
  BUFFD0 U346 ( .I(n486), .Z(n485) );
  BUFFD0 U347 ( .I(n487), .Z(n486) );
  BUFFD0 U348 ( .I(n488), .Z(n487) );
  BUFFD0 U349 ( .I(n489), .Z(n488) );
  BUFFD0 U350 ( .I(n490), .Z(n489) );
  BUFFD0 U351 ( .I(n491), .Z(n490) );
  BUFFD0 U352 ( .I(n492), .Z(n491) );
  BUFFD0 U353 ( .I(n493), .Z(n492) );
  BUFFD0 U354 ( .I(n494), .Z(n493) );
  BUFFD0 U355 ( .I(n495), .Z(n494) );
  BUFFD0 U356 ( .I(n496), .Z(n495) );
  BUFFD0 U357 ( .I(n497), .Z(n496) );
  BUFFD0 U358 ( .I(n498), .Z(n497) );
  BUFFD0 U359 ( .I(n499), .Z(n498) );
  BUFFD0 U360 ( .I(n500), .Z(n499) );
  CKBD0 U361 ( .CLK(FrameSR[54]), .C(n518) );
  BUFFD0 U362 ( .I(n502), .Z(n501) );
  BUFFD0 U363 ( .I(n503), .Z(n502) );
  BUFFD0 U364 ( .I(n504), .Z(n503) );
  BUFFD0 U365 ( .I(n505), .Z(n504) );
  BUFFD0 U366 ( .I(n506), .Z(n505) );
  BUFFD0 U367 ( .I(n507), .Z(n506) );
  BUFFD0 U368 ( .I(n508), .Z(n507) );
  BUFFD0 U369 ( .I(n509), .Z(n508) );
  BUFFD0 U370 ( .I(n510), .Z(n509) );
  BUFFD0 U371 ( .I(n511), .Z(n510) );
  BUFFD0 U372 ( .I(n512), .Z(n511) );
  BUFFD0 U373 ( .I(n513), .Z(n512) );
  BUFFD0 U374 ( .I(n514), .Z(n513) );
  BUFFD0 U375 ( .I(n515), .Z(n514) );
  BUFFD0 U376 ( .I(n516), .Z(n515) );
  BUFFD0 U377 ( .I(n517), .Z(n516) );
  BUFFD0 U378 ( .I(n518), .Z(n517) );
  BUFFD0 U379 ( .I(n520), .Z(n519) );
  BUFFD0 U380 ( .I(n521), .Z(n520) );
  BUFFD0 U381 ( .I(n522), .Z(n521) );
  BUFFD0 U382 ( .I(n523), .Z(n522) );
  BUFFD0 U383 ( .I(n524), .Z(n523) );
  BUFFD0 U384 ( .I(n525), .Z(n524) );
  BUFFD0 U385 ( .I(n526), .Z(n525) );
  BUFFD0 U386 ( .I(n527), .Z(n526) );
  BUFFD0 U387 ( .I(n528), .Z(n527) );
  BUFFD0 U388 ( .I(n529), .Z(n528) );
  BUFFD0 U389 ( .I(n530), .Z(n529) );
  BUFFD0 U390 ( .I(n531), .Z(n530) );
  BUFFD0 U391 ( .I(n532), .Z(n531) );
  BUFFD0 U392 ( .I(n533), .Z(n532) );
  BUFFD0 U393 ( .I(n534), .Z(n533) );
  BUFFD0 U394 ( .I(n535), .Z(n534) );
  BUFFD0 U395 ( .I(n2462), .Z(n535) );
  BUFFD0 U396 ( .I(n537), .Z(n536) );
  BUFFD0 U397 ( .I(n538), .Z(n537) );
  BUFFD0 U398 ( .I(n539), .Z(n538) );
  BUFFD0 U399 ( .I(n540), .Z(n539) );
  BUFFD0 U400 ( .I(n541), .Z(n540) );
  BUFFD0 U401 ( .I(n542), .Z(n541) );
  BUFFD0 U402 ( .I(n543), .Z(n542) );
  BUFFD0 U403 ( .I(n544), .Z(n543) );
  BUFFD0 U404 ( .I(n545), .Z(n544) );
  BUFFD0 U405 ( .I(n546), .Z(n545) );
  BUFFD0 U406 ( .I(n547), .Z(n546) );
  BUFFD0 U407 ( .I(n548), .Z(n547) );
  BUFFD0 U408 ( .I(n549), .Z(n548) );
  BUFFD0 U409 ( .I(n550), .Z(n549) );
  BUFFD0 U410 ( .I(n551), .Z(n550) );
  BUFFD0 U411 ( .I(n552), .Z(n551) );
  BUFFD0 U412 ( .I(n553), .Z(n552) );
  BUFFD0 U413 ( .I(n554), .Z(n553) );
  BUFFD0 U414 ( .I(FrameSR[8]), .Z(n554) );
  CKBD0 U415 ( .CLK(FrameSR[9]), .C(n572) );
  BUFFD0 U416 ( .I(n556), .Z(n555) );
  BUFFD0 U417 ( .I(n557), .Z(n556) );
  BUFFD0 U418 ( .I(n558), .Z(n557) );
  BUFFD0 U419 ( .I(n559), .Z(n558) );
  BUFFD0 U420 ( .I(n560), .Z(n559) );
  BUFFD0 U421 ( .I(n561), .Z(n560) );
  BUFFD0 U422 ( .I(n562), .Z(n561) );
  BUFFD0 U423 ( .I(n563), .Z(n562) );
  BUFFD0 U424 ( .I(n564), .Z(n563) );
  BUFFD0 U425 ( .I(n565), .Z(n564) );
  BUFFD0 U426 ( .I(n566), .Z(n565) );
  BUFFD0 U427 ( .I(n567), .Z(n566) );
  BUFFD0 U428 ( .I(n568), .Z(n567) );
  BUFFD0 U429 ( .I(n569), .Z(n568) );
  BUFFD0 U430 ( .I(n570), .Z(n569) );
  BUFFD0 U431 ( .I(n571), .Z(n570) );
  BUFFD0 U432 ( .I(n572), .Z(n571) );
  CKBD0 U433 ( .CLK(FrameSR[10]), .C(n590) );
  BUFFD0 U434 ( .I(n574), .Z(n573) );
  BUFFD0 U435 ( .I(n575), .Z(n574) );
  BUFFD0 U436 ( .I(n576), .Z(n575) );
  BUFFD0 U437 ( .I(n577), .Z(n576) );
  BUFFD0 U438 ( .I(n578), .Z(n577) );
  BUFFD0 U439 ( .I(n579), .Z(n578) );
  BUFFD0 U440 ( .I(n580), .Z(n579) );
  BUFFD0 U441 ( .I(n581), .Z(n580) );
  BUFFD0 U442 ( .I(n582), .Z(n581) );
  BUFFD0 U443 ( .I(n583), .Z(n582) );
  BUFFD0 U444 ( .I(n584), .Z(n583) );
  BUFFD0 U445 ( .I(n585), .Z(n584) );
  BUFFD0 U446 ( .I(n586), .Z(n585) );
  BUFFD0 U447 ( .I(n587), .Z(n586) );
  BUFFD0 U448 ( .I(n588), .Z(n587) );
  BUFFD0 U449 ( .I(n589), .Z(n588) );
  BUFFD0 U450 ( .I(n590), .Z(n589) );
  CKBD0 U451 ( .CLK(FrameSR[11]), .C(n608) );
  BUFFD0 U452 ( .I(n592), .Z(n591) );
  BUFFD0 U453 ( .I(n593), .Z(n592) );
  BUFFD0 U454 ( .I(n594), .Z(n593) );
  BUFFD0 U455 ( .I(n595), .Z(n594) );
  BUFFD0 U456 ( .I(n596), .Z(n595) );
  BUFFD0 U457 ( .I(n597), .Z(n596) );
  BUFFD0 U458 ( .I(n598), .Z(n597) );
  BUFFD0 U459 ( .I(n599), .Z(n598) );
  BUFFD0 U460 ( .I(n600), .Z(n599) );
  BUFFD0 U461 ( .I(n601), .Z(n600) );
  BUFFD0 U462 ( .I(n602), .Z(n601) );
  BUFFD0 U463 ( .I(n603), .Z(n602) );
  BUFFD0 U464 ( .I(n604), .Z(n603) );
  BUFFD0 U465 ( .I(n605), .Z(n604) );
  BUFFD0 U466 ( .I(n606), .Z(n605) );
  BUFFD0 U467 ( .I(n607), .Z(n606) );
  BUFFD0 U468 ( .I(n608), .Z(n607) );
  CKBD0 U469 ( .CLK(FrameSR[12]), .C(n626) );
  BUFFD0 U470 ( .I(n610), .Z(n609) );
  BUFFD0 U471 ( .I(n611), .Z(n610) );
  BUFFD0 U472 ( .I(n612), .Z(n611) );
  BUFFD0 U473 ( .I(n613), .Z(n612) );
  BUFFD0 U474 ( .I(n614), .Z(n613) );
  BUFFD0 U475 ( .I(n615), .Z(n614) );
  BUFFD0 U476 ( .I(n616), .Z(n615) );
  BUFFD0 U477 ( .I(n617), .Z(n616) );
  BUFFD0 U478 ( .I(n618), .Z(n617) );
  BUFFD0 U479 ( .I(n619), .Z(n618) );
  BUFFD0 U480 ( .I(n620), .Z(n619) );
  BUFFD0 U481 ( .I(n621), .Z(n620) );
  BUFFD0 U482 ( .I(n622), .Z(n621) );
  BUFFD0 U483 ( .I(n623), .Z(n622) );
  BUFFD0 U484 ( .I(n624), .Z(n623) );
  BUFFD0 U485 ( .I(n625), .Z(n624) );
  BUFFD0 U486 ( .I(n626), .Z(n625) );
  CKBD0 U487 ( .CLK(FrameSR[13]), .C(n644) );
  BUFFD0 U488 ( .I(n628), .Z(n627) );
  BUFFD0 U489 ( .I(n629), .Z(n628) );
  BUFFD0 U490 ( .I(n630), .Z(n629) );
  BUFFD0 U491 ( .I(n631), .Z(n630) );
  BUFFD0 U492 ( .I(n632), .Z(n631) );
  BUFFD0 U493 ( .I(n633), .Z(n632) );
  BUFFD0 U494 ( .I(n634), .Z(n633) );
  BUFFD0 U495 ( .I(n635), .Z(n634) );
  BUFFD0 U496 ( .I(n636), .Z(n635) );
  BUFFD0 U497 ( .I(n637), .Z(n636) );
  BUFFD0 U498 ( .I(n638), .Z(n637) );
  BUFFD0 U499 ( .I(n639), .Z(n638) );
  BUFFD0 U500 ( .I(n640), .Z(n639) );
  BUFFD0 U501 ( .I(n641), .Z(n640) );
  BUFFD0 U502 ( .I(n642), .Z(n641) );
  BUFFD0 U503 ( .I(n643), .Z(n642) );
  BUFFD0 U504 ( .I(n644), .Z(n643) );
  CKBD0 U505 ( .CLK(FrameSR[14]), .C(n662) );
  BUFFD0 U506 ( .I(n646), .Z(n645) );
  BUFFD0 U507 ( .I(n647), .Z(n646) );
  BUFFD0 U508 ( .I(n648), .Z(n647) );
  BUFFD0 U509 ( .I(n649), .Z(n648) );
  BUFFD0 U510 ( .I(n650), .Z(n649) );
  BUFFD0 U511 ( .I(n651), .Z(n650) );
  BUFFD0 U512 ( .I(n652), .Z(n651) );
  BUFFD0 U513 ( .I(n653), .Z(n652) );
  BUFFD0 U514 ( .I(n654), .Z(n653) );
  BUFFD0 U515 ( .I(n655), .Z(n654) );
  BUFFD0 U516 ( .I(n656), .Z(n655) );
  BUFFD0 U517 ( .I(n657), .Z(n656) );
  BUFFD0 U518 ( .I(n658), .Z(n657) );
  BUFFD0 U519 ( .I(n659), .Z(n658) );
  BUFFD0 U520 ( .I(n660), .Z(n659) );
  BUFFD0 U521 ( .I(n661), .Z(n660) );
  BUFFD0 U522 ( .I(n662), .Z(n661) );
  CKBD0 U523 ( .CLK(FrameSR[23]), .C(n680) );
  BUFFD0 U524 ( .I(n664), .Z(n663) );
  BUFFD0 U525 ( .I(n665), .Z(n664) );
  BUFFD0 U526 ( .I(n666), .Z(n665) );
  BUFFD0 U527 ( .I(n667), .Z(n666) );
  BUFFD0 U528 ( .I(n668), .Z(n667) );
  BUFFD0 U529 ( .I(n669), .Z(n668) );
  BUFFD0 U530 ( .I(n670), .Z(n669) );
  BUFFD0 U531 ( .I(n671), .Z(n670) );
  BUFFD0 U532 ( .I(n672), .Z(n671) );
  BUFFD0 U533 ( .I(n673), .Z(n672) );
  BUFFD0 U534 ( .I(n674), .Z(n673) );
  BUFFD0 U535 ( .I(n675), .Z(n674) );
  BUFFD0 U536 ( .I(n676), .Z(n675) );
  BUFFD0 U537 ( .I(n677), .Z(n676) );
  BUFFD0 U538 ( .I(n678), .Z(n677) );
  BUFFD0 U539 ( .I(n679), .Z(n678) );
  BUFFD0 U540 ( .I(n680), .Z(n679) );
  CKBD0 U541 ( .CLK(FrameSR[24]), .C(n698) );
  BUFFD0 U542 ( .I(n682), .Z(n681) );
  BUFFD0 U543 ( .I(n683), .Z(n682) );
  BUFFD0 U544 ( .I(n684), .Z(n683) );
  BUFFD0 U545 ( .I(n685), .Z(n684) );
  BUFFD0 U546 ( .I(n686), .Z(n685) );
  BUFFD0 U547 ( .I(n687), .Z(n686) );
  BUFFD0 U548 ( .I(n688), .Z(n687) );
  BUFFD0 U549 ( .I(n689), .Z(n688) );
  BUFFD0 U550 ( .I(n690), .Z(n689) );
  BUFFD0 U551 ( .I(n691), .Z(n690) );
  BUFFD0 U552 ( .I(n692), .Z(n691) );
  BUFFD0 U553 ( .I(n693), .Z(n692) );
  BUFFD0 U554 ( .I(n694), .Z(n693) );
  BUFFD0 U555 ( .I(n695), .Z(n694) );
  BUFFD0 U556 ( .I(n696), .Z(n695) );
  BUFFD0 U557 ( .I(n697), .Z(n696) );
  BUFFD0 U558 ( .I(n698), .Z(n697) );
  CKBD0 U559 ( .CLK(FrameSR[25]), .C(n716) );
  BUFFD0 U560 ( .I(n700), .Z(n699) );
  BUFFD0 U561 ( .I(n701), .Z(n700) );
  BUFFD0 U562 ( .I(n702), .Z(n701) );
  BUFFD0 U563 ( .I(n703), .Z(n702) );
  BUFFD0 U564 ( .I(n704), .Z(n703) );
  BUFFD0 U565 ( .I(n705), .Z(n704) );
  BUFFD0 U566 ( .I(n706), .Z(n705) );
  BUFFD0 U567 ( .I(n707), .Z(n706) );
  BUFFD0 U568 ( .I(n708), .Z(n707) );
  BUFFD0 U569 ( .I(n709), .Z(n708) );
  BUFFD0 U570 ( .I(n710), .Z(n709) );
  BUFFD0 U571 ( .I(n711), .Z(n710) );
  BUFFD0 U572 ( .I(n712), .Z(n711) );
  BUFFD0 U573 ( .I(n713), .Z(n712) );
  BUFFD0 U574 ( .I(n714), .Z(n713) );
  BUFFD0 U575 ( .I(n715), .Z(n714) );
  BUFFD0 U576 ( .I(n716), .Z(n715) );
  CKBD0 U577 ( .CLK(FrameSR[26]), .C(n734) );
  BUFFD0 U578 ( .I(n718), .Z(n717) );
  BUFFD0 U579 ( .I(n719), .Z(n718) );
  BUFFD0 U580 ( .I(n720), .Z(n719) );
  BUFFD0 U581 ( .I(n721), .Z(n720) );
  BUFFD0 U582 ( .I(n722), .Z(n721) );
  BUFFD0 U583 ( .I(n723), .Z(n722) );
  BUFFD0 U584 ( .I(n724), .Z(n723) );
  BUFFD0 U585 ( .I(n725), .Z(n724) );
  BUFFD0 U586 ( .I(n726), .Z(n725) );
  BUFFD0 U587 ( .I(n727), .Z(n726) );
  BUFFD0 U588 ( .I(n728), .Z(n727) );
  BUFFD0 U589 ( .I(n729), .Z(n728) );
  BUFFD0 U590 ( .I(n730), .Z(n729) );
  BUFFD0 U591 ( .I(n731), .Z(n730) );
  BUFFD0 U592 ( .I(n732), .Z(n731) );
  BUFFD0 U593 ( .I(n733), .Z(n732) );
  BUFFD0 U594 ( .I(n734), .Z(n733) );
  CKBD0 U595 ( .CLK(FrameSR[27]), .C(n752) );
  BUFFD0 U596 ( .I(n736), .Z(n735) );
  BUFFD0 U597 ( .I(n737), .Z(n736) );
  BUFFD0 U598 ( .I(n738), .Z(n737) );
  BUFFD0 U599 ( .I(n739), .Z(n738) );
  BUFFD0 U600 ( .I(n740), .Z(n739) );
  BUFFD0 U601 ( .I(n741), .Z(n740) );
  BUFFD0 U602 ( .I(n742), .Z(n741) );
  BUFFD0 U603 ( .I(n743), .Z(n742) );
  BUFFD0 U604 ( .I(n744), .Z(n743) );
  BUFFD0 U605 ( .I(n745), .Z(n744) );
  BUFFD0 U606 ( .I(n746), .Z(n745) );
  BUFFD0 U607 ( .I(n747), .Z(n746) );
  BUFFD0 U608 ( .I(n748), .Z(n747) );
  BUFFD0 U609 ( .I(n749), .Z(n748) );
  BUFFD0 U610 ( .I(n750), .Z(n749) );
  BUFFD0 U611 ( .I(n751), .Z(n750) );
  BUFFD0 U612 ( .I(n752), .Z(n751) );
  CKBD0 U613 ( .CLK(FrameSR[28]), .C(n770) );
  BUFFD0 U614 ( .I(n754), .Z(n753) );
  BUFFD0 U615 ( .I(n755), .Z(n754) );
  BUFFD0 U616 ( .I(n756), .Z(n755) );
  BUFFD0 U617 ( .I(n757), .Z(n756) );
  BUFFD0 U618 ( .I(n758), .Z(n757) );
  BUFFD0 U619 ( .I(n759), .Z(n758) );
  BUFFD0 U620 ( .I(n760), .Z(n759) );
  BUFFD0 U621 ( .I(n761), .Z(n760) );
  BUFFD0 U622 ( .I(n762), .Z(n761) );
  BUFFD0 U623 ( .I(n763), .Z(n762) );
  BUFFD0 U624 ( .I(n764), .Z(n763) );
  BUFFD0 U625 ( .I(n765), .Z(n764) );
  BUFFD0 U626 ( .I(n766), .Z(n765) );
  BUFFD0 U627 ( .I(n767), .Z(n766) );
  BUFFD0 U628 ( .I(n768), .Z(n767) );
  BUFFD0 U629 ( .I(n769), .Z(n768) );
  BUFFD0 U630 ( .I(n770), .Z(n769) );
  CKBD0 U631 ( .CLK(FrameSR[29]), .C(n788) );
  BUFFD0 U632 ( .I(n772), .Z(n771) );
  BUFFD0 U633 ( .I(n773), .Z(n772) );
  BUFFD0 U634 ( .I(n774), .Z(n773) );
  BUFFD0 U635 ( .I(n775), .Z(n774) );
  BUFFD0 U636 ( .I(n776), .Z(n775) );
  BUFFD0 U637 ( .I(n777), .Z(n776) );
  BUFFD0 U638 ( .I(n778), .Z(n777) );
  BUFFD0 U639 ( .I(n779), .Z(n778) );
  BUFFD0 U640 ( .I(n780), .Z(n779) );
  BUFFD0 U641 ( .I(n781), .Z(n780) );
  BUFFD0 U642 ( .I(n782), .Z(n781) );
  BUFFD0 U643 ( .I(n783), .Z(n782) );
  BUFFD0 U644 ( .I(n784), .Z(n783) );
  BUFFD0 U645 ( .I(n785), .Z(n784) );
  BUFFD0 U646 ( .I(n786), .Z(n785) );
  BUFFD0 U647 ( .I(n787), .Z(n786) );
  BUFFD0 U648 ( .I(n788), .Z(n787) );
  CKBD0 U649 ( .CLK(FrameSR[30]), .C(n806) );
  BUFFD0 U650 ( .I(n790), .Z(n789) );
  BUFFD0 U651 ( .I(n791), .Z(n790) );
  BUFFD0 U652 ( .I(n792), .Z(n791) );
  BUFFD0 U653 ( .I(n793), .Z(n792) );
  BUFFD0 U654 ( .I(n794), .Z(n793) );
  BUFFD0 U655 ( .I(n795), .Z(n794) );
  BUFFD0 U656 ( .I(n796), .Z(n795) );
  BUFFD0 U657 ( .I(n797), .Z(n796) );
  BUFFD0 U658 ( .I(n798), .Z(n797) );
  BUFFD0 U659 ( .I(n799), .Z(n798) );
  BUFFD0 U660 ( .I(n800), .Z(n799) );
  BUFFD0 U661 ( .I(n801), .Z(n800) );
  BUFFD0 U662 ( .I(n802), .Z(n801) );
  BUFFD0 U663 ( .I(n803), .Z(n802) );
  BUFFD0 U664 ( .I(n804), .Z(n803) );
  BUFFD0 U665 ( .I(n805), .Z(n804) );
  BUFFD0 U666 ( .I(n806), .Z(n805) );
  CKBD0 U667 ( .CLK(FrameSR[39]), .C(n824) );
  BUFFD0 U668 ( .I(n808), .Z(n807) );
  BUFFD0 U669 ( .I(n809), .Z(n808) );
  BUFFD0 U670 ( .I(n810), .Z(n809) );
  BUFFD0 U671 ( .I(n811), .Z(n810) );
  BUFFD0 U672 ( .I(n812), .Z(n811) );
  BUFFD0 U673 ( .I(n813), .Z(n812) );
  BUFFD0 U674 ( .I(n814), .Z(n813) );
  BUFFD0 U675 ( .I(n815), .Z(n814) );
  BUFFD0 U676 ( .I(n816), .Z(n815) );
  BUFFD0 U677 ( .I(n817), .Z(n816) );
  BUFFD0 U678 ( .I(n818), .Z(n817) );
  BUFFD0 U679 ( .I(n819), .Z(n818) );
  BUFFD0 U680 ( .I(n820), .Z(n819) );
  BUFFD0 U681 ( .I(n821), .Z(n820) );
  BUFFD0 U682 ( .I(n822), .Z(n821) );
  BUFFD0 U683 ( .I(n823), .Z(n822) );
  BUFFD0 U684 ( .I(n824), .Z(n823) );
  CKBD0 U685 ( .CLK(FrameSR[40]), .C(n842) );
  BUFFD0 U686 ( .I(n826), .Z(n825) );
  BUFFD0 U687 ( .I(n827), .Z(n826) );
  BUFFD0 U688 ( .I(n828), .Z(n827) );
  BUFFD0 U689 ( .I(n829), .Z(n828) );
  BUFFD0 U690 ( .I(n830), .Z(n829) );
  BUFFD0 U691 ( .I(n831), .Z(n830) );
  BUFFD0 U692 ( .I(n832), .Z(n831) );
  BUFFD0 U693 ( .I(n833), .Z(n832) );
  BUFFD0 U694 ( .I(n834), .Z(n833) );
  BUFFD0 U695 ( .I(n835), .Z(n834) );
  BUFFD0 U696 ( .I(n836), .Z(n835) );
  BUFFD0 U697 ( .I(n837), .Z(n836) );
  BUFFD0 U698 ( .I(n838), .Z(n837) );
  BUFFD0 U699 ( .I(n839), .Z(n838) );
  BUFFD0 U700 ( .I(n840), .Z(n839) );
  BUFFD0 U701 ( .I(n841), .Z(n840) );
  BUFFD0 U702 ( .I(n842), .Z(n841) );
  CKBD0 U703 ( .CLK(FrameSR[41]), .C(n860) );
  BUFFD0 U704 ( .I(n844), .Z(n843) );
  BUFFD0 U705 ( .I(n845), .Z(n844) );
  BUFFD0 U706 ( .I(n846), .Z(n845) );
  BUFFD0 U707 ( .I(n847), .Z(n846) );
  BUFFD0 U708 ( .I(n848), .Z(n847) );
  BUFFD0 U709 ( .I(n849), .Z(n848) );
  BUFFD0 U710 ( .I(n850), .Z(n849) );
  BUFFD0 U711 ( .I(n851), .Z(n850) );
  BUFFD0 U712 ( .I(n852), .Z(n851) );
  BUFFD0 U713 ( .I(n853), .Z(n852) );
  BUFFD0 U714 ( .I(n854), .Z(n853) );
  BUFFD0 U715 ( .I(n855), .Z(n854) );
  BUFFD0 U716 ( .I(n856), .Z(n855) );
  BUFFD0 U717 ( .I(n857), .Z(n856) );
  BUFFD0 U718 ( .I(n858), .Z(n857) );
  BUFFD0 U719 ( .I(n859), .Z(n858) );
  BUFFD0 U720 ( .I(n860), .Z(n859) );
  CKBD0 U721 ( .CLK(FrameSR[42]), .C(n878) );
  BUFFD0 U722 ( .I(n862), .Z(n861) );
  BUFFD0 U723 ( .I(n863), .Z(n862) );
  BUFFD0 U724 ( .I(n864), .Z(n863) );
  BUFFD0 U725 ( .I(n865), .Z(n864) );
  BUFFD0 U726 ( .I(n866), .Z(n865) );
  BUFFD0 U727 ( .I(n867), .Z(n866) );
  BUFFD0 U728 ( .I(n868), .Z(n867) );
  BUFFD0 U729 ( .I(n869), .Z(n868) );
  BUFFD0 U730 ( .I(n870), .Z(n869) );
  BUFFD0 U731 ( .I(n871), .Z(n870) );
  BUFFD0 U732 ( .I(n872), .Z(n871) );
  BUFFD0 U733 ( .I(n873), .Z(n872) );
  BUFFD0 U734 ( .I(n874), .Z(n873) );
  BUFFD0 U735 ( .I(n875), .Z(n874) );
  BUFFD0 U736 ( .I(n876), .Z(n875) );
  BUFFD0 U737 ( .I(n877), .Z(n876) );
  BUFFD0 U738 ( .I(n878), .Z(n877) );
  CKBD0 U739 ( .CLK(FrameSR[43]), .C(n896) );
  BUFFD0 U740 ( .I(n880), .Z(n879) );
  BUFFD0 U741 ( .I(n881), .Z(n880) );
  BUFFD0 U742 ( .I(n882), .Z(n881) );
  BUFFD0 U743 ( .I(n883), .Z(n882) );
  BUFFD0 U744 ( .I(n884), .Z(n883) );
  BUFFD0 U745 ( .I(n885), .Z(n884) );
  BUFFD0 U746 ( .I(n886), .Z(n885) );
  BUFFD0 U747 ( .I(n887), .Z(n886) );
  BUFFD0 U748 ( .I(n888), .Z(n887) );
  BUFFD0 U749 ( .I(n889), .Z(n888) );
  BUFFD0 U750 ( .I(n890), .Z(n889) );
  BUFFD0 U751 ( .I(n891), .Z(n890) );
  BUFFD0 U752 ( .I(n892), .Z(n891) );
  BUFFD0 U753 ( .I(n893), .Z(n892) );
  BUFFD0 U754 ( .I(n894), .Z(n893) );
  BUFFD0 U755 ( .I(n895), .Z(n894) );
  BUFFD0 U756 ( .I(n896), .Z(n895) );
  CKBD0 U757 ( .CLK(FrameSR[44]), .C(n914) );
  BUFFD0 U758 ( .I(n898), .Z(n897) );
  BUFFD0 U759 ( .I(n899), .Z(n898) );
  BUFFD0 U760 ( .I(n900), .Z(n899) );
  BUFFD0 U761 ( .I(n901), .Z(n900) );
  BUFFD0 U762 ( .I(n902), .Z(n901) );
  BUFFD0 U763 ( .I(n903), .Z(n902) );
  BUFFD0 U764 ( .I(n904), .Z(n903) );
  BUFFD0 U765 ( .I(n905), .Z(n904) );
  BUFFD0 U766 ( .I(n906), .Z(n905) );
  BUFFD0 U767 ( .I(n907), .Z(n906) );
  BUFFD0 U768 ( .I(n908), .Z(n907) );
  BUFFD0 U769 ( .I(n909), .Z(n908) );
  BUFFD0 U770 ( .I(n910), .Z(n909) );
  BUFFD0 U771 ( .I(n911), .Z(n910) );
  BUFFD0 U772 ( .I(n912), .Z(n911) );
  BUFFD0 U773 ( .I(n913), .Z(n912) );
  BUFFD0 U774 ( .I(n914), .Z(n913) );
  CKBD0 U775 ( .CLK(FrameSR[45]), .C(n932) );
  BUFFD0 U776 ( .I(n916), .Z(n915) );
  BUFFD0 U777 ( .I(n917), .Z(n916) );
  BUFFD0 U778 ( .I(n918), .Z(n917) );
  BUFFD0 U779 ( .I(n919), .Z(n918) );
  BUFFD0 U780 ( .I(n920), .Z(n919) );
  BUFFD0 U781 ( .I(n921), .Z(n920) );
  BUFFD0 U782 ( .I(n922), .Z(n921) );
  BUFFD0 U783 ( .I(n923), .Z(n922) );
  BUFFD0 U784 ( .I(n924), .Z(n923) );
  BUFFD0 U785 ( .I(n925), .Z(n924) );
  BUFFD0 U786 ( .I(n926), .Z(n925) );
  BUFFD0 U787 ( .I(n927), .Z(n926) );
  BUFFD0 U788 ( .I(n928), .Z(n927) );
  BUFFD0 U789 ( .I(n929), .Z(n928) );
  BUFFD0 U790 ( .I(n930), .Z(n929) );
  BUFFD0 U791 ( .I(n931), .Z(n930) );
  BUFFD0 U792 ( .I(n932), .Z(n931) );
  CKBD0 U793 ( .CLK(FrameSR[46]), .C(n950) );
  BUFFD0 U794 ( .I(n934), .Z(n933) );
  BUFFD0 U795 ( .I(n935), .Z(n934) );
  BUFFD0 U796 ( .I(n936), .Z(n935) );
  BUFFD0 U797 ( .I(n937), .Z(n936) );
  BUFFD0 U798 ( .I(n938), .Z(n937) );
  BUFFD0 U799 ( .I(n939), .Z(n938) );
  BUFFD0 U800 ( .I(n940), .Z(n939) );
  BUFFD0 U801 ( .I(n941), .Z(n940) );
  BUFFD0 U802 ( .I(n942), .Z(n941) );
  BUFFD0 U803 ( .I(n943), .Z(n942) );
  BUFFD0 U804 ( .I(n944), .Z(n943) );
  BUFFD0 U805 ( .I(n945), .Z(n944) );
  BUFFD0 U806 ( .I(n946), .Z(n945) );
  BUFFD0 U807 ( .I(n947), .Z(n946) );
  BUFFD0 U808 ( .I(n948), .Z(n947) );
  BUFFD0 U809 ( .I(n949), .Z(n948) );
  BUFFD0 U810 ( .I(n950), .Z(n949) );
  CKBD0 U811 ( .CLK(FrameSR[55]), .C(n968) );
  BUFFD0 U812 ( .I(n952), .Z(n951) );
  BUFFD0 U813 ( .I(n953), .Z(n952) );
  BUFFD0 U814 ( .I(n954), .Z(n953) );
  BUFFD0 U815 ( .I(n955), .Z(n954) );
  BUFFD0 U816 ( .I(n956), .Z(n955) );
  BUFFD0 U817 ( .I(n957), .Z(n956) );
  BUFFD0 U818 ( .I(n958), .Z(n957) );
  BUFFD0 U819 ( .I(n959), .Z(n958) );
  BUFFD0 U820 ( .I(n960), .Z(n959) );
  BUFFD0 U821 ( .I(n961), .Z(n960) );
  BUFFD0 U822 ( .I(n962), .Z(n961) );
  BUFFD0 U823 ( .I(n963), .Z(n962) );
  BUFFD0 U824 ( .I(n964), .Z(n963) );
  BUFFD0 U825 ( .I(n965), .Z(n964) );
  BUFFD0 U826 ( .I(n966), .Z(n965) );
  BUFFD0 U827 ( .I(n967), .Z(n966) );
  BUFFD0 U828 ( .I(n968), .Z(n967) );
  CKBD0 U829 ( .CLK(FrameSR[56]), .C(n986) );
  BUFFD0 U830 ( .I(n970), .Z(n969) );
  BUFFD0 U831 ( .I(n971), .Z(n970) );
  BUFFD0 U832 ( .I(n972), .Z(n971) );
  BUFFD0 U833 ( .I(n973), .Z(n972) );
  BUFFD0 U834 ( .I(n974), .Z(n973) );
  BUFFD0 U835 ( .I(n975), .Z(n974) );
  BUFFD0 U836 ( .I(n976), .Z(n975) );
  BUFFD0 U837 ( .I(n977), .Z(n976) );
  BUFFD0 U838 ( .I(n978), .Z(n977) );
  BUFFD0 U839 ( .I(n979), .Z(n978) );
  BUFFD0 U840 ( .I(n980), .Z(n979) );
  BUFFD0 U841 ( .I(n981), .Z(n980) );
  BUFFD0 U842 ( .I(n982), .Z(n981) );
  BUFFD0 U843 ( .I(n983), .Z(n982) );
  BUFFD0 U844 ( .I(n984), .Z(n983) );
  BUFFD0 U845 ( .I(n985), .Z(n984) );
  BUFFD0 U846 ( .I(n986), .Z(n985) );
  CKBD0 U847 ( .CLK(FrameSR[57]), .C(n1004) );
  BUFFD0 U848 ( .I(n988), .Z(n987) );
  BUFFD0 U849 ( .I(n989), .Z(n988) );
  BUFFD0 U850 ( .I(n990), .Z(n989) );
  BUFFD0 U851 ( .I(n991), .Z(n990) );
  BUFFD0 U852 ( .I(n992), .Z(n991) );
  BUFFD0 U853 ( .I(n993), .Z(n992) );
  BUFFD0 U854 ( .I(n994), .Z(n993) );
  BUFFD0 U855 ( .I(n995), .Z(n994) );
  BUFFD0 U856 ( .I(n996), .Z(n995) );
  BUFFD0 U857 ( .I(n997), .Z(n996) );
  BUFFD0 U858 ( .I(n998), .Z(n997) );
  BUFFD0 U859 ( .I(n999), .Z(n998) );
  BUFFD0 U860 ( .I(n1000), .Z(n999) );
  BUFFD0 U861 ( .I(n1001), .Z(n1000) );
  BUFFD0 U862 ( .I(n1002), .Z(n1001) );
  BUFFD0 U863 ( .I(n1003), .Z(n1002) );
  BUFFD0 U864 ( .I(n1004), .Z(n1003) );
  CKBD0 U865 ( .CLK(FrameSR[58]), .C(n1022) );
  BUFFD0 U866 ( .I(n1006), .Z(n1005) );
  BUFFD0 U867 ( .I(n1007), .Z(n1006) );
  BUFFD0 U868 ( .I(n1008), .Z(n1007) );
  BUFFD0 U869 ( .I(n1009), .Z(n1008) );
  BUFFD0 U870 ( .I(n1010), .Z(n1009) );
  BUFFD0 U871 ( .I(n1011), .Z(n1010) );
  BUFFD0 U872 ( .I(n1012), .Z(n1011) );
  BUFFD0 U873 ( .I(n1013), .Z(n1012) );
  BUFFD0 U874 ( .I(n1014), .Z(n1013) );
  BUFFD0 U875 ( .I(n1015), .Z(n1014) );
  BUFFD0 U876 ( .I(n1016), .Z(n1015) );
  BUFFD0 U877 ( .I(n1017), .Z(n1016) );
  BUFFD0 U878 ( .I(n1018), .Z(n1017) );
  BUFFD0 U879 ( .I(n1019), .Z(n1018) );
  BUFFD0 U880 ( .I(n1020), .Z(n1019) );
  BUFFD0 U881 ( .I(n1021), .Z(n1020) );
  BUFFD0 U882 ( .I(n1022), .Z(n1021) );
  CKBD0 U883 ( .CLK(FrameSR[59]), .C(n1040) );
  BUFFD0 U884 ( .I(n1024), .Z(n1023) );
  BUFFD0 U885 ( .I(n1025), .Z(n1024) );
  BUFFD0 U886 ( .I(n1026), .Z(n1025) );
  BUFFD0 U887 ( .I(n1027), .Z(n1026) );
  BUFFD0 U888 ( .I(n1028), .Z(n1027) );
  BUFFD0 U889 ( .I(n1029), .Z(n1028) );
  BUFFD0 U890 ( .I(n1030), .Z(n1029) );
  BUFFD0 U891 ( .I(n1031), .Z(n1030) );
  BUFFD0 U892 ( .I(n1032), .Z(n1031) );
  BUFFD0 U893 ( .I(n1033), .Z(n1032) );
  BUFFD0 U894 ( .I(n1034), .Z(n1033) );
  BUFFD0 U895 ( .I(n1035), .Z(n1034) );
  BUFFD0 U896 ( .I(n1036), .Z(n1035) );
  BUFFD0 U897 ( .I(n1037), .Z(n1036) );
  BUFFD0 U898 ( .I(n1038), .Z(n1037) );
  BUFFD0 U899 ( .I(n1039), .Z(n1038) );
  BUFFD0 U900 ( .I(n1040), .Z(n1039) );
  CKBD0 U901 ( .CLK(FrameSR[60]), .C(n1058) );
  BUFFD0 U902 ( .I(n1042), .Z(n1041) );
  BUFFD0 U903 ( .I(n1043), .Z(n1042) );
  BUFFD0 U904 ( .I(n1044), .Z(n1043) );
  BUFFD0 U905 ( .I(n1045), .Z(n1044) );
  BUFFD0 U906 ( .I(n1046), .Z(n1045) );
  BUFFD0 U907 ( .I(n1047), .Z(n1046) );
  BUFFD0 U908 ( .I(n1048), .Z(n1047) );
  BUFFD0 U909 ( .I(n1049), .Z(n1048) );
  BUFFD0 U910 ( .I(n1050), .Z(n1049) );
  BUFFD0 U911 ( .I(n1051), .Z(n1050) );
  BUFFD0 U912 ( .I(n1052), .Z(n1051) );
  BUFFD0 U913 ( .I(n1053), .Z(n1052) );
  BUFFD0 U914 ( .I(n1054), .Z(n1053) );
  BUFFD0 U915 ( .I(n1055), .Z(n1054) );
  BUFFD0 U916 ( .I(n1056), .Z(n1055) );
  BUFFD0 U917 ( .I(n1057), .Z(n1056) );
  BUFFD0 U918 ( .I(n1058), .Z(n1057) );
  CKBD0 U919 ( .CLK(FrameSR[61]), .C(n1076) );
  BUFFD0 U920 ( .I(n1060), .Z(n1059) );
  BUFFD0 U921 ( .I(n1061), .Z(n1060) );
  BUFFD0 U922 ( .I(n1062), .Z(n1061) );
  BUFFD0 U923 ( .I(n1063), .Z(n1062) );
  BUFFD0 U924 ( .I(n1064), .Z(n1063) );
  BUFFD0 U925 ( .I(n1065), .Z(n1064) );
  BUFFD0 U926 ( .I(n1066), .Z(n1065) );
  BUFFD0 U927 ( .I(n1067), .Z(n1066) );
  BUFFD0 U928 ( .I(n1068), .Z(n1067) );
  BUFFD0 U929 ( .I(n1069), .Z(n1068) );
  BUFFD0 U930 ( .I(n1070), .Z(n1069) );
  BUFFD0 U931 ( .I(n1071), .Z(n1070) );
  BUFFD0 U932 ( .I(n1072), .Z(n1071) );
  BUFFD0 U933 ( .I(n1073), .Z(n1072) );
  BUFFD0 U934 ( .I(n1074), .Z(n1073) );
  BUFFD0 U935 ( .I(n1075), .Z(n1074) );
  BUFFD0 U936 ( .I(n1076), .Z(n1075) );
  CKBD0 U937 ( .CLK(FrameSR[62]), .C(n1094) );
  BUFFD0 U938 ( .I(n1078), .Z(n1077) );
  BUFFD0 U939 ( .I(n1079), .Z(n1078) );
  BUFFD0 U940 ( .I(n1080), .Z(n1079) );
  BUFFD0 U941 ( .I(n1081), .Z(n1080) );
  BUFFD0 U942 ( .I(n1082), .Z(n1081) );
  BUFFD0 U943 ( .I(n1083), .Z(n1082) );
  BUFFD0 U944 ( .I(n1084), .Z(n1083) );
  BUFFD0 U945 ( .I(n1085), .Z(n1084) );
  BUFFD0 U946 ( .I(n1086), .Z(n1085) );
  BUFFD0 U947 ( .I(n1087), .Z(n1086) );
  BUFFD0 U948 ( .I(n1088), .Z(n1087) );
  BUFFD0 U949 ( .I(n1089), .Z(n1088) );
  BUFFD0 U950 ( .I(n1090), .Z(n1089) );
  BUFFD0 U951 ( .I(n1091), .Z(n1090) );
  BUFFD0 U952 ( .I(n1092), .Z(n1091) );
  BUFFD0 U953 ( .I(n1093), .Z(n1092) );
  BUFFD0 U954 ( .I(n1094), .Z(n1093) );
  BUFFD0 U955 ( .I(n1096), .Z(n1095) );
  BUFFD0 U956 ( .I(n1097), .Z(n1096) );
  BUFFD0 U957 ( .I(n1098), .Z(n1097) );
  BUFFD0 U958 ( .I(n1099), .Z(n1098) );
  BUFFD0 U959 ( .I(n1100), .Z(n1099) );
  BUFFD0 U960 ( .I(n1101), .Z(n1100) );
  BUFFD0 U961 ( .I(n1102), .Z(n1101) );
  BUFFD0 U962 ( .I(n1103), .Z(n1102) );
  BUFFD0 U963 ( .I(n1104), .Z(n1103) );
  BUFFD0 U964 ( .I(n1105), .Z(n1104) );
  BUFFD0 U965 ( .I(n1106), .Z(n1105) );
  BUFFD0 U966 ( .I(n1107), .Z(n1106) );
  BUFFD0 U967 ( .I(n1108), .Z(n1107) );
  BUFFD0 U968 ( .I(n1109), .Z(n1108) );
  BUFFD0 U969 ( .I(n1110), .Z(n1109) );
  BUFFD0 U970 ( .I(n1111), .Z(n1110) );
  BUFFD0 U971 ( .I(n1112), .Z(n1111) );
  BUFFD0 U972 ( .I(FrameSR[21]), .Z(n1112) );
  CKBD0 U973 ( .CLK(FrameSR[36]), .C(n1130) );
  BUFFD0 U974 ( .I(n1114), .Z(n1113) );
  BUFFD0 U975 ( .I(n1115), .Z(n1114) );
  BUFFD0 U976 ( .I(n1116), .Z(n1115) );
  BUFFD0 U977 ( .I(n1117), .Z(n1116) );
  BUFFD0 U978 ( .I(n1118), .Z(n1117) );
  BUFFD0 U979 ( .I(n1119), .Z(n1118) );
  BUFFD0 U980 ( .I(n1120), .Z(n1119) );
  BUFFD0 U981 ( .I(n1121), .Z(n1120) );
  BUFFD0 U982 ( .I(n1122), .Z(n1121) );
  BUFFD0 U983 ( .I(n1123), .Z(n1122) );
  BUFFD0 U984 ( .I(n1124), .Z(n1123) );
  BUFFD0 U985 ( .I(n1125), .Z(n1124) );
  BUFFD0 U986 ( .I(n1126), .Z(n1125) );
  BUFFD0 U987 ( .I(n1127), .Z(n1126) );
  BUFFD0 U988 ( .I(n1128), .Z(n1127) );
  BUFFD0 U989 ( .I(n1129), .Z(n1128) );
  BUFFD0 U990 ( .I(n1130), .Z(n1129) );
  CKBD0 U991 ( .CLK(FrameSR[52]), .C(n1148) );
  BUFFD0 U992 ( .I(n1132), .Z(n1131) );
  BUFFD0 U993 ( .I(n1133), .Z(n1132) );
  BUFFD0 U994 ( .I(n1134), .Z(n1133) );
  BUFFD0 U995 ( .I(n1135), .Z(n1134) );
  BUFFD0 U996 ( .I(n1136), .Z(n1135) );
  BUFFD0 U997 ( .I(n1137), .Z(n1136) );
  BUFFD0 U998 ( .I(n1138), .Z(n1137) );
  BUFFD0 U999 ( .I(n1139), .Z(n1138) );
  BUFFD0 U1000 ( .I(n1140), .Z(n1139) );
  BUFFD0 U1001 ( .I(n1141), .Z(n1140) );
  BUFFD0 U1002 ( .I(n1142), .Z(n1141) );
  BUFFD0 U1003 ( .I(n1143), .Z(n1142) );
  BUFFD0 U1004 ( .I(n1144), .Z(n1143) );
  BUFFD0 U1005 ( .I(n1145), .Z(n1144) );
  BUFFD0 U1006 ( .I(n1146), .Z(n1145) );
  BUFFD0 U1007 ( .I(n1147), .Z(n1146) );
  BUFFD0 U1008 ( .I(n1148), .Z(n1147) );
  BUFFD0 U1009 ( .I(n1151), .Z(n1149) );
  BUFFD0 U1010 ( .I(n260), .Z(n1150) );
  BUFFD0 U1011 ( .I(n1152), .Z(n1151) );
  BUFFD0 U1012 ( .I(n1153), .Z(n1152) );
  BUFFD0 U1013 ( .I(n1154), .Z(n1153) );
  BUFFD0 U1014 ( .I(n1155), .Z(n1154) );
  BUFFD0 U1015 ( .I(n1156), .Z(n1155) );
  BUFFD0 U1016 ( .I(n1157), .Z(n1156) );
  BUFFD0 U1017 ( .I(n1158), .Z(n1157) );
  BUFFD0 U1018 ( .I(n1159), .Z(n1158) );
  BUFFD0 U1019 ( .I(n1160), .Z(n1159) );
  BUFFD0 U1020 ( .I(n1161), .Z(n1160) );
  BUFFD0 U1021 ( .I(n1162), .Z(n1161) );
  BUFFD0 U1022 ( .I(n1163), .Z(n1162) );
  BUFFD0 U1023 ( .I(n1164), .Z(n1163) );
  BUFFD0 U1024 ( .I(n1165), .Z(n1164) );
  BUFFD0 U1025 ( .I(n1150), .Z(n1165) );
  BUFFD0 U1026 ( .I(n1168), .Z(n1166) );
  BUFFD0 U1027 ( .I(n259), .Z(n1167) );
  BUFFD0 U1028 ( .I(n1169), .Z(n1168) );
  BUFFD0 U1029 ( .I(n1170), .Z(n1169) );
  BUFFD0 U1030 ( .I(n1171), .Z(n1170) );
  BUFFD0 U1031 ( .I(n1172), .Z(n1171) );
  BUFFD0 U1032 ( .I(n1173), .Z(n1172) );
  BUFFD0 U1033 ( .I(n1174), .Z(n1173) );
  BUFFD0 U1034 ( .I(n1175), .Z(n1174) );
  BUFFD0 U1035 ( .I(n1176), .Z(n1175) );
  BUFFD0 U1036 ( .I(n1177), .Z(n1176) );
  BUFFD0 U1037 ( .I(n1178), .Z(n1177) );
  BUFFD0 U1038 ( .I(n1179), .Z(n1178) );
  BUFFD0 U1039 ( .I(n1180), .Z(n1179) );
  BUFFD0 U1040 ( .I(n1181), .Z(n1180) );
  BUFFD0 U1041 ( .I(n1182), .Z(n1181) );
  BUFFD0 U1042 ( .I(n1167), .Z(n1182) );
  BUFFD0 U1043 ( .I(n1185), .Z(n1183) );
  BUFFD0 U1044 ( .I(n258), .Z(n1184) );
  BUFFD0 U1045 ( .I(n1186), .Z(n1185) );
  BUFFD0 U1046 ( .I(n1187), .Z(n1186) );
  BUFFD0 U1047 ( .I(n1188), .Z(n1187) );
  BUFFD0 U1048 ( .I(n1189), .Z(n1188) );
  BUFFD0 U1049 ( .I(n1190), .Z(n1189) );
  BUFFD0 U1050 ( .I(n1191), .Z(n1190) );
  BUFFD0 U1051 ( .I(n1192), .Z(n1191) );
  BUFFD0 U1052 ( .I(n1193), .Z(n1192) );
  BUFFD0 U1053 ( .I(n1194), .Z(n1193) );
  BUFFD0 U1054 ( .I(n1195), .Z(n1194) );
  BUFFD0 U1055 ( .I(n1196), .Z(n1195) );
  BUFFD0 U1056 ( .I(n1197), .Z(n1196) );
  BUFFD0 U1057 ( .I(n1198), .Z(n1197) );
  BUFFD0 U1058 ( .I(n1199), .Z(n1198) );
  BUFFD0 U1059 ( .I(n1184), .Z(n1199) );
  BUFFD0 U1060 ( .I(n1202), .Z(n1200) );
  BUFFD0 U1061 ( .I(n257), .Z(n1201) );
  BUFFD0 U1062 ( .I(n1203), .Z(n1202) );
  BUFFD0 U1063 ( .I(n1204), .Z(n1203) );
  BUFFD0 U1064 ( .I(n1205), .Z(n1204) );
  BUFFD0 U1065 ( .I(n1206), .Z(n1205) );
  BUFFD0 U1066 ( .I(n1207), .Z(n1206) );
  BUFFD0 U1067 ( .I(n1208), .Z(n1207) );
  BUFFD0 U1068 ( .I(n1209), .Z(n1208) );
  BUFFD0 U1069 ( .I(n1210), .Z(n1209) );
  BUFFD0 U1070 ( .I(n1211), .Z(n1210) );
  BUFFD0 U1071 ( .I(n1212), .Z(n1211) );
  BUFFD0 U1072 ( .I(n1213), .Z(n1212) );
  BUFFD0 U1073 ( .I(n1214), .Z(n1213) );
  BUFFD0 U1074 ( .I(n1215), .Z(n1214) );
  BUFFD0 U1075 ( .I(n1216), .Z(n1215) );
  BUFFD0 U1076 ( .I(n1201), .Z(n1216) );
  BUFFD0 U1077 ( .I(n1219), .Z(n1217) );
  BUFFD0 U1078 ( .I(n256), .Z(n1218) );
  BUFFD0 U1079 ( .I(n1220), .Z(n1219) );
  BUFFD0 U1080 ( .I(n1221), .Z(n1220) );
  BUFFD0 U1081 ( .I(n1222), .Z(n1221) );
  BUFFD0 U1082 ( .I(n1223), .Z(n1222) );
  BUFFD0 U1083 ( .I(n1224), .Z(n1223) );
  BUFFD0 U1084 ( .I(n1225), .Z(n1224) );
  BUFFD0 U1085 ( .I(n1226), .Z(n1225) );
  BUFFD0 U1086 ( .I(n1227), .Z(n1226) );
  BUFFD0 U1087 ( .I(n1228), .Z(n1227) );
  BUFFD0 U1088 ( .I(n1229), .Z(n1228) );
  BUFFD0 U1089 ( .I(n1230), .Z(n1229) );
  BUFFD0 U1090 ( .I(n1231), .Z(n1230) );
  BUFFD0 U1091 ( .I(n1232), .Z(n1231) );
  BUFFD0 U1092 ( .I(n1233), .Z(n1232) );
  BUFFD0 U1093 ( .I(n1218), .Z(n1233) );
  BUFFD0 U1094 ( .I(n1236), .Z(n1234) );
  BUFFD0 U1095 ( .I(n255), .Z(n1235) );
  BUFFD0 U1096 ( .I(n1237), .Z(n1236) );
  BUFFD0 U1097 ( .I(n1238), .Z(n1237) );
  BUFFD0 U1098 ( .I(n1239), .Z(n1238) );
  BUFFD0 U1099 ( .I(n1240), .Z(n1239) );
  BUFFD0 U1100 ( .I(n1241), .Z(n1240) );
  BUFFD0 U1101 ( .I(n1242), .Z(n1241) );
  BUFFD0 U1102 ( .I(n1243), .Z(n1242) );
  BUFFD0 U1103 ( .I(n1244), .Z(n1243) );
  BUFFD0 U1104 ( .I(n1245), .Z(n1244) );
  BUFFD0 U1105 ( .I(n1246), .Z(n1245) );
  BUFFD0 U1106 ( .I(n1247), .Z(n1246) );
  BUFFD0 U1107 ( .I(n1248), .Z(n1247) );
  BUFFD0 U1108 ( .I(n1249), .Z(n1248) );
  BUFFD0 U1109 ( .I(n1250), .Z(n1249) );
  BUFFD0 U1110 ( .I(n1235), .Z(n1250) );
  BUFFD0 U1111 ( .I(n1253), .Z(n1251) );
  BUFFD0 U1112 ( .I(n254), .Z(n1252) );
  BUFFD0 U1113 ( .I(n1254), .Z(n1253) );
  BUFFD0 U1114 ( .I(n1255), .Z(n1254) );
  BUFFD0 U1115 ( .I(n1256), .Z(n1255) );
  BUFFD0 U1116 ( .I(n1257), .Z(n1256) );
  BUFFD0 U1117 ( .I(n1258), .Z(n1257) );
  BUFFD0 U1118 ( .I(n1259), .Z(n1258) );
  BUFFD0 U1119 ( .I(n1260), .Z(n1259) );
  BUFFD0 U1120 ( .I(n1261), .Z(n1260) );
  BUFFD0 U1121 ( .I(n1262), .Z(n1261) );
  BUFFD0 U1122 ( .I(n1263), .Z(n1262) );
  BUFFD0 U1123 ( .I(n1264), .Z(n1263) );
  BUFFD0 U1124 ( .I(n1265), .Z(n1264) );
  BUFFD0 U1125 ( .I(n1266), .Z(n1265) );
  BUFFD0 U1126 ( .I(n1267), .Z(n1266) );
  BUFFD0 U1127 ( .I(n1252), .Z(n1267) );
  BUFFD0 U1128 ( .I(n1270), .Z(n1268) );
  BUFFD0 U1129 ( .I(n253), .Z(n1269) );
  BUFFD0 U1130 ( .I(n1271), .Z(n1270) );
  BUFFD0 U1131 ( .I(n1272), .Z(n1271) );
  BUFFD0 U1132 ( .I(n1273), .Z(n1272) );
  BUFFD0 U1133 ( .I(n1274), .Z(n1273) );
  BUFFD0 U1134 ( .I(n1275), .Z(n1274) );
  BUFFD0 U1135 ( .I(n1276), .Z(n1275) );
  BUFFD0 U1136 ( .I(n1277), .Z(n1276) );
  BUFFD0 U1137 ( .I(n1278), .Z(n1277) );
  BUFFD0 U1138 ( .I(n1279), .Z(n1278) );
  BUFFD0 U1139 ( .I(n1280), .Z(n1279) );
  BUFFD0 U1140 ( .I(n1281), .Z(n1280) );
  BUFFD0 U1141 ( .I(n1282), .Z(n1281) );
  BUFFD0 U1142 ( .I(n1283), .Z(n1282) );
  BUFFD0 U1143 ( .I(n1284), .Z(n1283) );
  BUFFD0 U1144 ( .I(n1269), .Z(n1284) );
  BUFFD0 U1145 ( .I(n1287), .Z(n1285) );
  BUFFD0 U1146 ( .I(n252), .Z(n1286) );
  BUFFD0 U1147 ( .I(n1288), .Z(n1287) );
  BUFFD0 U1148 ( .I(n1289), .Z(n1288) );
  BUFFD0 U1149 ( .I(n1290), .Z(n1289) );
  BUFFD0 U1150 ( .I(n1291), .Z(n1290) );
  BUFFD0 U1151 ( .I(n1292), .Z(n1291) );
  BUFFD0 U1152 ( .I(n1293), .Z(n1292) );
  BUFFD0 U1153 ( .I(n1294), .Z(n1293) );
  BUFFD0 U1154 ( .I(n1295), .Z(n1294) );
  BUFFD0 U1155 ( .I(n1296), .Z(n1295) );
  BUFFD0 U1156 ( .I(n1297), .Z(n1296) );
  BUFFD0 U1157 ( .I(n1298), .Z(n1297) );
  BUFFD0 U1158 ( .I(n1299), .Z(n1298) );
  BUFFD0 U1159 ( .I(n1300), .Z(n1299) );
  BUFFD0 U1160 ( .I(n1301), .Z(n1300) );
  BUFFD0 U1161 ( .I(n1286), .Z(n1301) );
  BUFFD0 U1162 ( .I(n1304), .Z(n1302) );
  BUFFD0 U1163 ( .I(n251), .Z(n1303) );
  BUFFD0 U1164 ( .I(n1305), .Z(n1304) );
  BUFFD0 U1165 ( .I(n1306), .Z(n1305) );
  BUFFD0 U1166 ( .I(n1307), .Z(n1306) );
  BUFFD0 U1167 ( .I(n1308), .Z(n1307) );
  BUFFD0 U1168 ( .I(n1309), .Z(n1308) );
  BUFFD0 U1169 ( .I(n1310), .Z(n1309) );
  BUFFD0 U1170 ( .I(n1311), .Z(n1310) );
  BUFFD0 U1171 ( .I(n1312), .Z(n1311) );
  BUFFD0 U1172 ( .I(n1313), .Z(n1312) );
  BUFFD0 U1173 ( .I(n1314), .Z(n1313) );
  BUFFD0 U1174 ( .I(n1315), .Z(n1314) );
  BUFFD0 U1175 ( .I(n1316), .Z(n1315) );
  BUFFD0 U1176 ( .I(n1317), .Z(n1316) );
  BUFFD0 U1177 ( .I(n1318), .Z(n1317) );
  BUFFD0 U1178 ( .I(n1303), .Z(n1318) );
  BUFFD0 U1179 ( .I(n1321), .Z(n1319) );
  BUFFD0 U1180 ( .I(n250), .Z(n1320) );
  BUFFD0 U1181 ( .I(n1322), .Z(n1321) );
  BUFFD0 U1182 ( .I(n1323), .Z(n1322) );
  BUFFD0 U1183 ( .I(n1324), .Z(n1323) );
  BUFFD0 U1184 ( .I(n1325), .Z(n1324) );
  BUFFD0 U1185 ( .I(n1326), .Z(n1325) );
  BUFFD0 U1186 ( .I(n1327), .Z(n1326) );
  BUFFD0 U1187 ( .I(n1328), .Z(n1327) );
  BUFFD0 U1188 ( .I(n1329), .Z(n1328) );
  BUFFD0 U1189 ( .I(n1330), .Z(n1329) );
  BUFFD0 U1190 ( .I(n1331), .Z(n1330) );
  BUFFD0 U1191 ( .I(n1332), .Z(n1331) );
  BUFFD0 U1192 ( .I(n1333), .Z(n1332) );
  BUFFD0 U1193 ( .I(n1334), .Z(n1333) );
  BUFFD0 U1194 ( .I(n1335), .Z(n1334) );
  BUFFD0 U1195 ( .I(n1320), .Z(n1335) );
  BUFFD0 U1196 ( .I(n1338), .Z(n1336) );
  BUFFD0 U1197 ( .I(n249), .Z(n1337) );
  BUFFD0 U1198 ( .I(n1339), .Z(n1338) );
  BUFFD0 U1199 ( .I(n1340), .Z(n1339) );
  BUFFD0 U1200 ( .I(n1341), .Z(n1340) );
  BUFFD0 U1201 ( .I(n1342), .Z(n1341) );
  BUFFD0 U1202 ( .I(n1343), .Z(n1342) );
  BUFFD0 U1203 ( .I(n1344), .Z(n1343) );
  BUFFD0 U1204 ( .I(n1345), .Z(n1344) );
  BUFFD0 U1205 ( .I(n1346), .Z(n1345) );
  BUFFD0 U1206 ( .I(n1347), .Z(n1346) );
  BUFFD0 U1207 ( .I(n1348), .Z(n1347) );
  BUFFD0 U1208 ( .I(n1349), .Z(n1348) );
  BUFFD0 U1209 ( .I(n1350), .Z(n1349) );
  BUFFD0 U1210 ( .I(n1351), .Z(n1350) );
  BUFFD0 U1211 ( .I(n1352), .Z(n1351) );
  BUFFD0 U1212 ( .I(n1337), .Z(n1352) );
  BUFFD0 U1213 ( .I(n1355), .Z(n1353) );
  BUFFD0 U1214 ( .I(n248), .Z(n1354) );
  BUFFD0 U1215 ( .I(n1356), .Z(n1355) );
  BUFFD0 U1216 ( .I(n1357), .Z(n1356) );
  BUFFD0 U1217 ( .I(n1358), .Z(n1357) );
  BUFFD0 U1218 ( .I(n1359), .Z(n1358) );
  BUFFD0 U1219 ( .I(n1360), .Z(n1359) );
  BUFFD0 U1220 ( .I(n1361), .Z(n1360) );
  BUFFD0 U1221 ( .I(n1362), .Z(n1361) );
  BUFFD0 U1222 ( .I(n1363), .Z(n1362) );
  BUFFD0 U1223 ( .I(n1364), .Z(n1363) );
  BUFFD0 U1224 ( .I(n1365), .Z(n1364) );
  BUFFD0 U1225 ( .I(n1366), .Z(n1365) );
  BUFFD0 U1226 ( .I(n1367), .Z(n1366) );
  BUFFD0 U1227 ( .I(n1368), .Z(n1367) );
  BUFFD0 U1228 ( .I(n1369), .Z(n1368) );
  BUFFD0 U1229 ( .I(n1354), .Z(n1369) );
  BUFFD0 U1230 ( .I(n1372), .Z(n1370) );
  BUFFD0 U1231 ( .I(n247), .Z(n1371) );
  BUFFD0 U1232 ( .I(n1373), .Z(n1372) );
  BUFFD0 U1233 ( .I(n1374), .Z(n1373) );
  BUFFD0 U1234 ( .I(n1375), .Z(n1374) );
  BUFFD0 U1235 ( .I(n1376), .Z(n1375) );
  BUFFD0 U1236 ( .I(n1377), .Z(n1376) );
  BUFFD0 U1237 ( .I(n1378), .Z(n1377) );
  BUFFD0 U1238 ( .I(n1379), .Z(n1378) );
  BUFFD0 U1239 ( .I(n1380), .Z(n1379) );
  BUFFD0 U1240 ( .I(n1381), .Z(n1380) );
  BUFFD0 U1241 ( .I(n1382), .Z(n1381) );
  BUFFD0 U1242 ( .I(n1383), .Z(n1382) );
  BUFFD0 U1243 ( .I(n1384), .Z(n1383) );
  BUFFD0 U1244 ( .I(n1385), .Z(n1384) );
  BUFFD0 U1245 ( .I(n1386), .Z(n1385) );
  BUFFD0 U1246 ( .I(n1371), .Z(n1386) );
  BUFFD0 U1247 ( .I(n1389), .Z(n1387) );
  BUFFD0 U1248 ( .I(n246), .Z(n1388) );
  BUFFD0 U1249 ( .I(n1390), .Z(n1389) );
  BUFFD0 U1250 ( .I(n1391), .Z(n1390) );
  BUFFD0 U1251 ( .I(n1392), .Z(n1391) );
  BUFFD0 U1252 ( .I(n1393), .Z(n1392) );
  BUFFD0 U1253 ( .I(n1394), .Z(n1393) );
  BUFFD0 U1254 ( .I(n1395), .Z(n1394) );
  BUFFD0 U1255 ( .I(n1396), .Z(n1395) );
  BUFFD0 U1256 ( .I(n1397), .Z(n1396) );
  BUFFD0 U1257 ( .I(n1398), .Z(n1397) );
  BUFFD0 U1258 ( .I(n1399), .Z(n1398) );
  BUFFD0 U1259 ( .I(n1400), .Z(n1399) );
  BUFFD0 U1260 ( .I(n1401), .Z(n1400) );
  BUFFD0 U1261 ( .I(n1402), .Z(n1401) );
  BUFFD0 U1262 ( .I(n1403), .Z(n1402) );
  BUFFD0 U1263 ( .I(n1388), .Z(n1403) );
  BUFFD0 U1264 ( .I(n1406), .Z(n1404) );
  BUFFD0 U1265 ( .I(n245), .Z(n1405) );
  BUFFD0 U1266 ( .I(n1407), .Z(n1406) );
  BUFFD0 U1267 ( .I(n1408), .Z(n1407) );
  BUFFD0 U1268 ( .I(n1409), .Z(n1408) );
  BUFFD0 U1269 ( .I(n1410), .Z(n1409) );
  BUFFD0 U1270 ( .I(n1411), .Z(n1410) );
  BUFFD0 U1271 ( .I(n1412), .Z(n1411) );
  BUFFD0 U1272 ( .I(n1413), .Z(n1412) );
  BUFFD0 U1273 ( .I(n1414), .Z(n1413) );
  BUFFD0 U1274 ( .I(n1415), .Z(n1414) );
  BUFFD0 U1275 ( .I(n1416), .Z(n1415) );
  BUFFD0 U1276 ( .I(n1417), .Z(n1416) );
  BUFFD0 U1277 ( .I(n1418), .Z(n1417) );
  BUFFD0 U1278 ( .I(n1419), .Z(n1418) );
  BUFFD0 U1279 ( .I(n1422), .Z(n1420) );
  BUFFD0 U1280 ( .I(n244), .Z(n1421) );
  BUFFD0 U1281 ( .I(n1423), .Z(n1422) );
  BUFFD0 U1282 ( .I(n1424), .Z(n1423) );
  BUFFD0 U1283 ( .I(n1425), .Z(n1424) );
  BUFFD0 U1284 ( .I(n1426), .Z(n1425) );
  BUFFD0 U1285 ( .I(n1427), .Z(n1426) );
  BUFFD0 U1286 ( .I(n1428), .Z(n1427) );
  BUFFD0 U1287 ( .I(n1429), .Z(n1428) );
  BUFFD0 U1288 ( .I(n1430), .Z(n1429) );
  BUFFD0 U1289 ( .I(n1431), .Z(n1430) );
  BUFFD0 U1290 ( .I(n1432), .Z(n1431) );
  BUFFD0 U1291 ( .I(n1433), .Z(n1432) );
  BUFFD0 U1292 ( .I(n1434), .Z(n1433) );
  BUFFD0 U1293 ( .I(n1435), .Z(n1434) );
  BUFFD0 U1294 ( .I(n1438), .Z(n1436) );
  BUFFD0 U1295 ( .I(n243), .Z(n1437) );
  BUFFD0 U1296 ( .I(n1439), .Z(n1438) );
  BUFFD0 U1297 ( .I(n1440), .Z(n1439) );
  BUFFD0 U1298 ( .I(n1441), .Z(n1440) );
  BUFFD0 U1299 ( .I(n1442), .Z(n1441) );
  BUFFD0 U1300 ( .I(n1443), .Z(n1442) );
  BUFFD0 U1301 ( .I(n1444), .Z(n1443) );
  BUFFD0 U1302 ( .I(n1445), .Z(n1444) );
  BUFFD0 U1303 ( .I(n1446), .Z(n1445) );
  BUFFD0 U1304 ( .I(n1447), .Z(n1446) );
  BUFFD0 U1305 ( .I(n1448), .Z(n1447) );
  BUFFD0 U1306 ( .I(n1449), .Z(n1448) );
  BUFFD0 U1307 ( .I(n1450), .Z(n1449) );
  BUFFD0 U1308 ( .I(n1451), .Z(n1450) );
  BUFFD0 U1309 ( .I(n1452), .Z(n1451) );
  BUFFD0 U1310 ( .I(n1437), .Z(n1452) );
  BUFFD0 U1311 ( .I(n1455), .Z(n1453) );
  BUFFD0 U1312 ( .I(n242), .Z(n1454) );
  BUFFD0 U1313 ( .I(n1456), .Z(n1455) );
  BUFFD0 U1314 ( .I(n1457), .Z(n1456) );
  BUFFD0 U1315 ( .I(n1458), .Z(n1457) );
  BUFFD0 U1316 ( .I(n1459), .Z(n1458) );
  BUFFD0 U1317 ( .I(n1460), .Z(n1459) );
  BUFFD0 U1318 ( .I(n1461), .Z(n1460) );
  BUFFD0 U1319 ( .I(n1462), .Z(n1461) );
  BUFFD0 U1320 ( .I(n1463), .Z(n1462) );
  BUFFD0 U1321 ( .I(n1464), .Z(n1463) );
  BUFFD0 U1322 ( .I(n1465), .Z(n1464) );
  BUFFD0 U1323 ( .I(n1466), .Z(n1465) );
  BUFFD0 U1324 ( .I(n1467), .Z(n1466) );
  BUFFD0 U1325 ( .I(n1468), .Z(n1467) );
  BUFFD0 U1326 ( .I(n1471), .Z(n1469) );
  BUFFD0 U1327 ( .I(n241), .Z(n1470) );
  BUFFD0 U1328 ( .I(n1472), .Z(n1471) );
  BUFFD0 U1329 ( .I(n1473), .Z(n1472) );
  BUFFD0 U1330 ( .I(n1474), .Z(n1473) );
  BUFFD0 U1331 ( .I(n1475), .Z(n1474) );
  BUFFD0 U1332 ( .I(n1476), .Z(n1475) );
  BUFFD0 U1333 ( .I(n1477), .Z(n1476) );
  BUFFD0 U1334 ( .I(n1478), .Z(n1477) );
  BUFFD0 U1335 ( .I(n1479), .Z(n1478) );
  BUFFD0 U1336 ( .I(n1480), .Z(n1479) );
  BUFFD0 U1337 ( .I(n1481), .Z(n1480) );
  BUFFD0 U1338 ( .I(n1482), .Z(n1481) );
  BUFFD0 U1339 ( .I(n1483), .Z(n1482) );
  BUFFD0 U1340 ( .I(n1484), .Z(n1483) );
  BUFFD0 U1341 ( .I(n1485), .Z(n1484) );
  BUFFD0 U1342 ( .I(n1470), .Z(n1485) );
  BUFFD0 U1343 ( .I(n1488), .Z(n1486) );
  BUFFD0 U1344 ( .I(n1489), .Z(n1488) );
  BUFFD0 U1345 ( .I(n1490), .Z(n1489) );
  BUFFD0 U1346 ( .I(n1491), .Z(n1490) );
  BUFFD0 U1347 ( .I(n1492), .Z(n1491) );
  BUFFD0 U1348 ( .I(n1493), .Z(n1492) );
  BUFFD0 U1349 ( .I(n1494), .Z(n1493) );
  BUFFD0 U1350 ( .I(n1495), .Z(n1494) );
  BUFFD0 U1351 ( .I(n1496), .Z(n1495) );
  BUFFD0 U1352 ( .I(n1497), .Z(n1496) );
  BUFFD0 U1353 ( .I(n1498), .Z(n1497) );
  BUFFD0 U1354 ( .I(n1499), .Z(n1498) );
  BUFFD0 U1355 ( .I(n1500), .Z(n1499) );
  BUFFD0 U1356 ( .I(n1501), .Z(n1500) );
  BUFFD0 U1357 ( .I(n1487), .Z(n1501) );
  BUFFD0 U1358 ( .I(n1504), .Z(n1502) );
  BUFFD0 U1359 ( .I(n239), .Z(n1503) );
  BUFFD0 U1360 ( .I(n1505), .Z(n1504) );
  BUFFD0 U1361 ( .I(n1506), .Z(n1505) );
  BUFFD0 U1362 ( .I(n1507), .Z(n1506) );
  BUFFD0 U1363 ( .I(n1508), .Z(n1507) );
  BUFFD0 U1364 ( .I(n1509), .Z(n1508) );
  BUFFD0 U1365 ( .I(n1510), .Z(n1509) );
  BUFFD0 U1366 ( .I(n1511), .Z(n1510) );
  BUFFD0 U1367 ( .I(n1512), .Z(n1511) );
  BUFFD0 U1368 ( .I(n1513), .Z(n1512) );
  BUFFD0 U1369 ( .I(n1514), .Z(n1513) );
  BUFFD0 U1370 ( .I(n1515), .Z(n1514) );
  BUFFD0 U1371 ( .I(n1517), .Z(n1516) );
  BUFFD0 U1372 ( .I(n1503), .Z(n1517) );
  BUFFD0 U1373 ( .I(n1520), .Z(n1518) );
  BUFFD0 U1374 ( .I(n238), .Z(n1519) );
  BUFFD0 U1375 ( .I(n1521), .Z(n1520) );
  BUFFD0 U1376 ( .I(n1522), .Z(n1521) );
  BUFFD0 U1377 ( .I(n1523), .Z(n1522) );
  BUFFD0 U1378 ( .I(n1524), .Z(n1523) );
  BUFFD0 U1379 ( .I(n1525), .Z(n1524) );
  BUFFD0 U1380 ( .I(n1526), .Z(n1525) );
  BUFFD0 U1381 ( .I(n1527), .Z(n1526) );
  BUFFD0 U1382 ( .I(n1528), .Z(n1527) );
  BUFFD0 U1383 ( .I(n1530), .Z(n1529) );
  BUFFD0 U1384 ( .I(n1531), .Z(n1530) );
  BUFFD0 U1385 ( .I(n1532), .Z(n1531) );
  BUFFD0 U1386 ( .I(n1533), .Z(n1532) );
  BUFFD0 U1387 ( .I(n1519), .Z(n1533) );
  BUFFD0 U1388 ( .I(n1536), .Z(n1534) );
  BUFFD0 U1389 ( .I(n237), .Z(n1535) );
  BUFFD0 U1390 ( .I(n1537), .Z(n1536) );
  BUFFD0 U1391 ( .I(n1538), .Z(n1537) );
  BUFFD0 U1392 ( .I(n1539), .Z(n1538) );
  BUFFD0 U1393 ( .I(n1540), .Z(n1539) );
  BUFFD0 U1394 ( .I(n1541), .Z(n1540) );
  BUFFD0 U1395 ( .I(n1542), .Z(n1541) );
  BUFFD0 U1396 ( .I(n1543), .Z(n1542) );
  BUFFD0 U1397 ( .I(n1544), .Z(n1543) );
  BUFFD0 U1398 ( .I(n1545), .Z(n1544) );
  BUFFD0 U1399 ( .I(n1546), .Z(n1545) );
  BUFFD0 U1400 ( .I(n1547), .Z(n1546) );
  BUFFD0 U1401 ( .I(n1548), .Z(n1547) );
  BUFFD0 U1402 ( .I(n1549), .Z(n1548) );
  BUFFD0 U1403 ( .I(n1550), .Z(n1549) );
  BUFFD0 U1404 ( .I(n1535), .Z(n1550) );
  BUFFD0 U1405 ( .I(n1553), .Z(n1551) );
  BUFFD0 U1406 ( .I(n236), .Z(n1552) );
  BUFFD0 U1407 ( .I(n1554), .Z(n1553) );
  BUFFD0 U1408 ( .I(n1555), .Z(n1554) );
  BUFFD0 U1409 ( .I(n1556), .Z(n1555) );
  BUFFD0 U1410 ( .I(n1557), .Z(n1556) );
  BUFFD0 U1411 ( .I(n1558), .Z(n1557) );
  BUFFD0 U1412 ( .I(n1559), .Z(n1558) );
  BUFFD0 U1413 ( .I(n1560), .Z(n1559) );
  BUFFD0 U1414 ( .I(n1561), .Z(n1560) );
  BUFFD0 U1415 ( .I(n1562), .Z(n1561) );
  BUFFD0 U1416 ( .I(n1563), .Z(n1562) );
  BUFFD0 U1417 ( .I(n1564), .Z(n1563) );
  BUFFD0 U1418 ( .I(n1565), .Z(n1564) );
  BUFFD0 U1419 ( .I(n1552), .Z(n1566) );
  BUFFD0 U1420 ( .I(n1569), .Z(n1567) );
  BUFFD0 U1421 ( .I(n235), .Z(n1568) );
  BUFFD0 U1422 ( .I(n1570), .Z(n1569) );
  BUFFD0 U1423 ( .I(n1571), .Z(n1570) );
  BUFFD0 U1424 ( .I(n1572), .Z(n1571) );
  BUFFD0 U1425 ( .I(n1573), .Z(n1572) );
  BUFFD0 U1426 ( .I(n1574), .Z(n1573) );
  BUFFD0 U1427 ( .I(n1575), .Z(n1574) );
  BUFFD0 U1428 ( .I(n1576), .Z(n1575) );
  BUFFD0 U1429 ( .I(n1577), .Z(n1576) );
  BUFFD0 U1430 ( .I(n1578), .Z(n1577) );
  BUFFD0 U1431 ( .I(n1580), .Z(n1579) );
  BUFFD0 U1432 ( .I(n1581), .Z(n1580) );
  BUFFD0 U1433 ( .I(n1582), .Z(n1581) );
  BUFFD0 U1434 ( .I(n1568), .Z(n1582) );
  BUFFD0 U1435 ( .I(n1585), .Z(n1583) );
  BUFFD0 U1436 ( .I(n234), .Z(n1584) );
  BUFFD0 U1437 ( .I(n1586), .Z(n1585) );
  BUFFD0 U1438 ( .I(n1587), .Z(n1586) );
  BUFFD0 U1439 ( .I(n1588), .Z(n1587) );
  BUFFD0 U1440 ( .I(n1589), .Z(n1588) );
  BUFFD0 U1441 ( .I(n1590), .Z(n1589) );
  BUFFD0 U1442 ( .I(n1591), .Z(n1590) );
  BUFFD0 U1443 ( .I(n1592), .Z(n1591) );
  BUFFD0 U1444 ( .I(n1593), .Z(n1592) );
  BUFFD0 U1445 ( .I(n1594), .Z(n1593) );
  BUFFD0 U1446 ( .I(n1595), .Z(n1594) );
  BUFFD0 U1447 ( .I(n1596), .Z(n1595) );
  BUFFD0 U1448 ( .I(n1597), .Z(n1596) );
  BUFFD0 U1449 ( .I(n1598), .Z(n1597) );
  BUFFD0 U1450 ( .I(n1599), .Z(n1598) );
  BUFFD0 U1451 ( .I(n1584), .Z(n1599) );
  BUFFD0 U1452 ( .I(n1602), .Z(n1600) );
  BUFFD0 U1453 ( .I(n233), .Z(n1601) );
  BUFFD0 U1454 ( .I(n1603), .Z(n1602) );
  BUFFD0 U1455 ( .I(n1604), .Z(n1603) );
  BUFFD0 U1456 ( .I(n1605), .Z(n1604) );
  BUFFD0 U1457 ( .I(n1606), .Z(n1605) );
  BUFFD0 U1458 ( .I(n1607), .Z(n1606) );
  BUFFD0 U1459 ( .I(n1608), .Z(n1607) );
  BUFFD0 U1460 ( .I(n1610), .Z(n1609) );
  BUFFD0 U1461 ( .I(n1611), .Z(n1610) );
  BUFFD0 U1462 ( .I(n1612), .Z(n1611) );
  BUFFD0 U1463 ( .I(n1613), .Z(n1612) );
  BUFFD0 U1464 ( .I(n1614), .Z(n1613) );
  BUFFD0 U1465 ( .I(n1615), .Z(n1614) );
  BUFFD0 U1466 ( .I(n1601), .Z(n1615) );
  BUFFD0 U1467 ( .I(n1618), .Z(n1616) );
  BUFFD0 U1468 ( .I(n232), .Z(n1617) );
  BUFFD0 U1469 ( .I(n1619), .Z(n1618) );
  BUFFD0 U1470 ( .I(n1620), .Z(n1619) );
  BUFFD0 U1471 ( .I(n1621), .Z(n1620) );
  BUFFD0 U1472 ( .I(n1622), .Z(n1621) );
  BUFFD0 U1473 ( .I(n1623), .Z(n1622) );
  BUFFD0 U1474 ( .I(n1624), .Z(n1623) );
  BUFFD0 U1475 ( .I(n1625), .Z(n1624) );
  BUFFD0 U1476 ( .I(n1626), .Z(n1625) );
  BUFFD0 U1477 ( .I(n1627), .Z(n1626) );
  BUFFD0 U1478 ( .I(n1628), .Z(n1627) );
  BUFFD0 U1479 ( .I(n1630), .Z(n1629) );
  BUFFD0 U1480 ( .I(n1631), .Z(n1630) );
  BUFFD0 U1481 ( .I(n1617), .Z(n1631) );
  BUFFD0 U1482 ( .I(n1634), .Z(n1632) );
  BUFFD0 U1483 ( .I(n231), .Z(n1633) );
  BUFFD0 U1484 ( .I(n1635), .Z(n1634) );
  BUFFD0 U1485 ( .I(n1636), .Z(n1635) );
  BUFFD0 U1486 ( .I(n1637), .Z(n1636) );
  BUFFD0 U1487 ( .I(n1638), .Z(n1637) );
  BUFFD0 U1488 ( .I(n1639), .Z(n1638) );
  BUFFD0 U1489 ( .I(n1640), .Z(n1639) );
  BUFFD0 U1490 ( .I(n1641), .Z(n1640) );
  BUFFD0 U1491 ( .I(n1642), .Z(n1641) );
  BUFFD0 U1492 ( .I(n1643), .Z(n1642) );
  BUFFD0 U1493 ( .I(n1644), .Z(n1643) );
  BUFFD0 U1494 ( .I(n1645), .Z(n1644) );
  BUFFD0 U1495 ( .I(n1646), .Z(n1645) );
  BUFFD0 U1496 ( .I(n1647), .Z(n1646) );
  BUFFD0 U1497 ( .I(n1648), .Z(n1647) );
  BUFFD0 U1498 ( .I(n1633), .Z(n1648) );
  BUFFD0 U1499 ( .I(n1651), .Z(n1649) );
  BUFFD0 U1500 ( .I(n230), .Z(n1650) );
  BUFFD0 U1501 ( .I(n1652), .Z(n1651) );
  BUFFD0 U1502 ( .I(n1653), .Z(n1652) );
  BUFFD0 U1503 ( .I(n1654), .Z(n1653) );
  BUFFD0 U1504 ( .I(n1655), .Z(n1654) );
  BUFFD0 U1505 ( .I(n1656), .Z(n1655) );
  BUFFD0 U1506 ( .I(n1657), .Z(n1656) );
  BUFFD0 U1507 ( .I(n1658), .Z(n1657) );
  BUFFD0 U1508 ( .I(n1659), .Z(n1658) );
  BUFFD0 U1509 ( .I(n1660), .Z(n1659) );
  BUFFD0 U1510 ( .I(n1661), .Z(n1660) );
  BUFFD0 U1511 ( .I(n1662), .Z(n1661) );
  BUFFD0 U1512 ( .I(n1663), .Z(n1662) );
  BUFFD0 U1513 ( .I(n1664), .Z(n1663) );
  BUFFD0 U1514 ( .I(n1665), .Z(n1664) );
  BUFFD0 U1515 ( .I(n1650), .Z(n1665) );
  BUFFD0 U1516 ( .I(n1667), .Z(n1666) );
  BUFFD0 U1517 ( .I(n1668), .Z(n1667) );
  BUFFD0 U1518 ( .I(n1669), .Z(n1668) );
  BUFFD0 U1519 ( .I(n1670), .Z(n1669) );
  BUFFD0 U1520 ( .I(n1671), .Z(n1670) );
  BUFFD0 U1521 ( .I(n1672), .Z(n1671) );
  BUFFD0 U1522 ( .I(n1673), .Z(n1672) );
  BUFFD0 U1523 ( .I(n1674), .Z(n1673) );
  BUFFD0 U1524 ( .I(n1675), .Z(n1674) );
  BUFFD0 U1525 ( .I(n1676), .Z(n1675) );
  BUFFD0 U1526 ( .I(n1677), .Z(n1676) );
  BUFFD0 U1527 ( .I(n1678), .Z(n1677) );
  BUFFD0 U1528 ( .I(n1679), .Z(n1678) );
  BUFFD0 U1529 ( .I(n1680), .Z(n1679) );
  BUFFD0 U1530 ( .I(n1682), .Z(n1680) );
  BUFFD0 U1531 ( .I(n183), .Z(n1681) );
  BUFFD0 U1532 ( .I(n229), .Z(n1682) );
  CKAN2D0 U1533 ( .A1(N34), .A2(n2), .Z(N42) );
  BUFFD0 U1534 ( .I(n1684), .Z(n1683) );
  BUFFD0 U1535 ( .I(n1685), .Z(n1684) );
  BUFFD0 U1536 ( .I(n1686), .Z(n1685) );
  BUFFD0 U1537 ( .I(n1687), .Z(n1686) );
  BUFFD0 U1538 ( .I(n1688), .Z(n1687) );
  BUFFD0 U1539 ( .I(n1689), .Z(n1688) );
  BUFFD0 U1540 ( .I(n1690), .Z(n1689) );
  BUFFD0 U1541 ( .I(n1691), .Z(n1690) );
  BUFFD0 U1542 ( .I(n1692), .Z(n1691) );
  BUFFD0 U1543 ( .I(n1693), .Z(n1692) );
  BUFFD0 U1544 ( .I(n1694), .Z(n1693) );
  BUFFD0 U1545 ( .I(n1695), .Z(n1694) );
  BUFFD0 U1546 ( .I(n1696), .Z(n1695) );
  BUFFD0 U1547 ( .I(N42), .Z(n1696) );
  BUFFD0 U1548 ( .I(n1699), .Z(n1697) );
  BUFFD0 U1549 ( .I(n1701), .Z(n1698) );
  BUFFD0 U1550 ( .I(n1700), .Z(n1699) );
  BUFFD0 U1551 ( .I(n1702), .Z(n1700) );
  BUFFD0 U1552 ( .I(n1703), .Z(n1701) );
  BUFFD0 U1553 ( .I(n1704), .Z(n1702) );
  BUFFD0 U1554 ( .I(n1705), .Z(n1703) );
  BUFFD0 U1555 ( .I(n1706), .Z(n1704) );
  BUFFD0 U1556 ( .I(n1707), .Z(n1705) );
  BUFFD0 U1557 ( .I(n1708), .Z(n1706) );
  BUFFD0 U1558 ( .I(n1709), .Z(n1707) );
  BUFFD0 U1559 ( .I(n194), .Z(n1708) );
  BUFFD0 U1560 ( .I(n8), .Z(n1709) );
  BUFFD0 U1561 ( .I(n1711), .Z(n1710) );
  BUFFD0 U1562 ( .I(n1712), .Z(n1711) );
  BUFFD0 U1563 ( .I(n1713), .Z(n1712) );
  BUFFD0 U1564 ( .I(n1714), .Z(n1713) );
  BUFFD0 U1565 ( .I(n1715), .Z(n1714) );
  BUFFD0 U1566 ( .I(n1716), .Z(n1715) );
  BUFFD0 U1567 ( .I(n1717), .Z(n1716) );
  BUFFD0 U1568 ( .I(n1718), .Z(n1717) );
  BUFFD0 U1569 ( .I(n1719), .Z(n1718) );
  BUFFD0 U1570 ( .I(n1720), .Z(n1719) );
  BUFFD0 U1571 ( .I(n1721), .Z(n1720) );
  BUFFD0 U1572 ( .I(n1722), .Z(n1721) );
  BUFFD0 U1573 ( .I(n1723), .Z(n1722) );
  BUFFD0 U1574 ( .I(n1724), .Z(n1723) );
  BUFFD0 U1575 ( .I(n1725), .Z(n1724) );
  BUFFD0 U1576 ( .I(n1726), .Z(n1725) );
  BUFFD0 U1577 ( .I(n1727), .Z(n1726) );
  BUFFD0 U1578 ( .I(n1728), .Z(n1727) );
  BUFFD0 U1579 ( .I(n1729), .Z(n1728) );
  BUFFD0 U1580 ( .I(n1730), .Z(n1729) );
  BUFFD0 U1581 ( .I(n1731), .Z(n1730) );
  BUFFD0 U1582 ( .I(n1732), .Z(n1731) );
  BUFFD0 U1583 ( .I(n1733), .Z(n1732) );
  BUFFD0 U1584 ( .I(n1734), .Z(n1733) );
  BUFFD0 U1585 ( .I(n1735), .Z(n1734) );
  BUFFD0 U1586 ( .I(n1736), .Z(n1735) );
  BUFFD0 U1587 ( .I(n1737), .Z(n1736) );
  BUFFD0 U1588 ( .I(n1738), .Z(n1737) );
  BUFFD0 U1589 ( .I(n1739), .Z(n1738) );
  BUFFD0 U1590 ( .I(n1740), .Z(n1739) );
  BUFFD0 U1591 ( .I(n1741), .Z(n1740) );
  BUFFD0 U1592 ( .I(n1742), .Z(n1741) );
  BUFFD0 U1593 ( .I(n1743), .Z(n1742) );
  BUFFD0 U1594 ( .I(n1744), .Z(n1743) );
  BUFFD0 U1595 ( .I(n1745), .Z(n1744) );
  BUFFD0 U1596 ( .I(n1746), .Z(n1745) );
  BUFFD0 U1597 ( .I(n1747), .Z(n1746) );
  BUFFD0 U1598 ( .I(n1748), .Z(n1747) );
  BUFFD0 U1599 ( .I(n1749), .Z(n1748) );
  BUFFD0 U1600 ( .I(n1750), .Z(n1749) );
  BUFFD0 U1601 ( .I(n1751), .Z(n1750) );
  BUFFD0 U1602 ( .I(n1752), .Z(n1751) );
  BUFFD0 U1603 ( .I(n1753), .Z(n1752) );
  BUFFD0 U1604 ( .I(n1754), .Z(n1753) );
  BUFFD0 U1605 ( .I(n1755), .Z(n1754) );
  BUFFD0 U1606 ( .I(n1756), .Z(n1755) );
  BUFFD0 U1607 ( .I(n1757), .Z(n1756) );
  BUFFD0 U1608 ( .I(n1758), .Z(n1757) );
  BUFFD0 U1609 ( .I(n1759), .Z(n1758) );
  BUFFD0 U1610 ( .I(n1760), .Z(n1759) );
  BUFFD0 U1611 ( .I(n1761), .Z(n1760) );
  BUFFD0 U1612 ( .I(n1762), .Z(n1761) );
  BUFFD0 U1613 ( .I(n1763), .Z(n1762) );
  BUFFD0 U1614 ( .I(n1764), .Z(n1763) );
  BUFFD0 U1615 ( .I(n1765), .Z(n1764) );
  BUFFD0 U1616 ( .I(n1766), .Z(n1765) );
  BUFFD0 U1617 ( .I(n1767), .Z(n1766) );
  BUFFD0 U1618 ( .I(n1768), .Z(n1767) );
  BUFFD0 U1619 ( .I(n1769), .Z(n1768) );
  BUFFD0 U1620 ( .I(n1770), .Z(n1769) );
  BUFFD0 U1621 ( .I(n1771), .Z(n1770) );
  BUFFD0 U1622 ( .I(n1772), .Z(n1771) );
  BUFFD0 U1623 ( .I(n1773), .Z(n1772) );
  BUFFD0 U1624 ( .I(n1774), .Z(n1773) );
  BUFFD0 U1625 ( .I(n1775), .Z(n1774) );
  BUFFD0 U1626 ( .I(n1776), .Z(n1775) );
  BUFFD0 U1627 ( .I(n1777), .Z(n1776) );
  BUFFD0 U1628 ( .I(n1778), .Z(n1777) );
  BUFFD0 U1629 ( .I(n1779), .Z(n1778) );
  BUFFD0 U1630 ( .I(n1780), .Z(n1779) );
  BUFFD0 U1631 ( .I(n1781), .Z(n1780) );
  BUFFD0 U1632 ( .I(n1782), .Z(n1781) );
  BUFFD0 U1633 ( .I(n1783), .Z(n1782) );
  BUFFD0 U1634 ( .I(n1784), .Z(n1783) );
  BUFFD0 U1635 ( .I(n1785), .Z(n1784) );
  BUFFD0 U1636 ( .I(n1786), .Z(n1785) );
  BUFFD0 U1637 ( .I(n1787), .Z(n1786) );
  BUFFD0 U1638 ( .I(n1788), .Z(n1787) );
  BUFFD0 U1639 ( .I(n1789), .Z(n1788) );
  BUFFD0 U1640 ( .I(n1790), .Z(n1789) );
  BUFFD0 U1641 ( .I(n1791), .Z(n1790) );
  BUFFD0 U1642 ( .I(n1792), .Z(n1791) );
  BUFFD0 U1643 ( .I(n1793), .Z(n1792) );
  BUFFD0 U1644 ( .I(n1794), .Z(n1793) );
  BUFFD0 U1645 ( .I(n1795), .Z(n1794) );
  BUFFD0 U1646 ( .I(n1796), .Z(n1795) );
  BUFFD0 U1647 ( .I(n1797), .Z(n1796) );
  BUFFD0 U1648 ( .I(n1798), .Z(n1797) );
  BUFFD0 U1649 ( .I(n1799), .Z(n1798) );
  BUFFD0 U1650 ( .I(n1800), .Z(n1799) );
  BUFFD0 U1651 ( .I(n1801), .Z(n1800) );
  BUFFD0 U1652 ( .I(n1802), .Z(n1801) );
  BUFFD0 U1653 ( .I(n1803), .Z(n1802) );
  BUFFD0 U1654 ( .I(n1804), .Z(n1803) );
  BUFFD0 U1655 ( .I(n1805), .Z(n1804) );
  BUFFD0 U1656 ( .I(n1806), .Z(n1805) );
  BUFFD0 U1657 ( .I(n1807), .Z(n1806) );
  BUFFD0 U1658 ( .I(n1808), .Z(n1807) );
  BUFFD0 U1659 ( .I(n1809), .Z(n1808) );
  BUFFD0 U1660 ( .I(n1810), .Z(n1809) );
  BUFFD0 U1661 ( .I(n1811), .Z(n1810) );
  BUFFD0 U1662 ( .I(n1812), .Z(n1811) );
  BUFFD0 U1663 ( .I(n1813), .Z(n1812) );
  BUFFD0 U1664 ( .I(n1814), .Z(n1813) );
  BUFFD0 U1665 ( .I(n1815), .Z(n1814) );
  BUFFD0 U1666 ( .I(n1816), .Z(n1815) );
  BUFFD0 U1667 ( .I(n1817), .Z(n1816) );
  BUFFD0 U1668 ( .I(n1818), .Z(n1817) );
  BUFFD0 U1669 ( .I(n1819), .Z(n1818) );
  BUFFD0 U1670 ( .I(n1820), .Z(n1819) );
  BUFFD0 U1671 ( .I(n1821), .Z(n1820) );
  BUFFD0 U1672 ( .I(n1822), .Z(n1821) );
  BUFFD0 U1673 ( .I(n1823), .Z(n1822) );
  BUFFD0 U1674 ( .I(n1824), .Z(n1823) );
  BUFFD0 U1675 ( .I(n1825), .Z(n1824) );
  BUFFD0 U1676 ( .I(n1826), .Z(n1825) );
  BUFFD0 U1677 ( .I(n1827), .Z(n1826) );
  BUFFD0 U1678 ( .I(n1828), .Z(n1827) );
  BUFFD0 U1679 ( .I(n1829), .Z(n1828) );
  BUFFD0 U1680 ( .I(n1830), .Z(n1829) );
  BUFFD0 U1681 ( .I(n1831), .Z(n1830) );
  BUFFD0 U1682 ( .I(n1832), .Z(n1831) );
  BUFFD0 U1683 ( .I(n1833), .Z(n1832) );
  BUFFD0 U1684 ( .I(n1834), .Z(n1833) );
  BUFFD0 U1685 ( .I(n1835), .Z(n1834) );
  BUFFD0 U1686 ( .I(n1836), .Z(n1835) );
  BUFFD0 U1687 ( .I(n1837), .Z(n1836) );
  BUFFD0 U1688 ( .I(n1838), .Z(n1837) );
  BUFFD0 U1689 ( .I(n1839), .Z(n1838) );
  BUFFD0 U1690 ( .I(n1840), .Z(n1839) );
  BUFFD0 U1691 ( .I(n1841), .Z(n1840) );
  BUFFD0 U1692 ( .I(n1842), .Z(n1841) );
  BUFFD0 U1693 ( .I(n1843), .Z(n1842) );
  BUFFD0 U1694 ( .I(n1844), .Z(n1843) );
  BUFFD0 U1695 ( .I(n1845), .Z(n1844) );
  BUFFD0 U1696 ( .I(n1846), .Z(n1845) );
  BUFFD0 U1697 ( .I(n1847), .Z(n1846) );
  BUFFD0 U1698 ( .I(n1848), .Z(n1847) );
  BUFFD0 U1699 ( .I(n1849), .Z(n1848) );
  BUFFD0 U1700 ( .I(n1850), .Z(n1849) );
  BUFFD0 U1701 ( .I(n1851), .Z(n1850) );
  BUFFD0 U1702 ( .I(n1852), .Z(n1851) );
  BUFFD0 U1703 ( .I(n1853), .Z(n1852) );
  BUFFD0 U1704 ( .I(n1854), .Z(n1853) );
  BUFFD0 U1705 ( .I(n1855), .Z(n1854) );
  BUFFD0 U1706 ( .I(n1856), .Z(n1855) );
  BUFFD0 U1707 ( .I(n1857), .Z(n1856) );
  BUFFD0 U1708 ( .I(n1858), .Z(n1857) );
  BUFFD0 U1709 ( .I(n1859), .Z(n1858) );
  BUFFD0 U1710 ( .I(n1860), .Z(n1859) );
  BUFFD0 U1711 ( .I(n1861), .Z(n1860) );
  BUFFD0 U1712 ( .I(n1862), .Z(n1861) );
  BUFFD0 U1713 ( .I(n1863), .Z(n1862) );
  BUFFD0 U1714 ( .I(n1864), .Z(n1863) );
  BUFFD0 U1715 ( .I(n1865), .Z(n1864) );
  BUFFD0 U1716 ( .I(n1866), .Z(n1865) );
  BUFFD0 U1717 ( .I(n1867), .Z(n1866) );
  BUFFD0 U1718 ( .I(n1868), .Z(n1867) );
  BUFFD0 U1719 ( .I(n1869), .Z(n1868) );
  BUFFD0 U1720 ( .I(n1870), .Z(n1869) );
  BUFFD0 U1721 ( .I(n1871), .Z(n1870) );
  BUFFD0 U1722 ( .I(n1872), .Z(n1871) );
  BUFFD0 U1723 ( .I(n1873), .Z(n1872) );
  BUFFD0 U1724 ( .I(n1874), .Z(n1873) );
  BUFFD0 U1725 ( .I(n1875), .Z(n1874) );
  BUFFD0 U1726 ( .I(n1876), .Z(n1875) );
  BUFFD0 U1727 ( .I(n1877), .Z(n1876) );
  BUFFD0 U1728 ( .I(n1878), .Z(n1877) );
  BUFFD0 U1729 ( .I(n1879), .Z(n1878) );
  BUFFD0 U1730 ( .I(n1880), .Z(n1879) );
  BUFFD0 U1731 ( .I(n1881), .Z(n1880) );
  BUFFD0 U1732 ( .I(n1882), .Z(n1881) );
  BUFFD0 U1733 ( .I(n1883), .Z(n1882) );
  BUFFD0 U1734 ( .I(n1884), .Z(n1883) );
  BUFFD0 U1735 ( .I(n1885), .Z(n1884) );
  BUFFD0 U1736 ( .I(n1886), .Z(n1885) );
  BUFFD0 U1737 ( .I(n1887), .Z(n1886) );
  BUFFD0 U1738 ( .I(n1888), .Z(n1887) );
  BUFFD0 U1739 ( .I(n1889), .Z(n1888) );
  BUFFD0 U1740 ( .I(n1890), .Z(n1889) );
  BUFFD0 U1741 ( .I(n1891), .Z(n1890) );
  BUFFD0 U1742 ( .I(n1892), .Z(n1891) );
  BUFFD0 U1743 ( .I(n1893), .Z(n1892) );
  BUFFD0 U1744 ( .I(n1894), .Z(n1893) );
  BUFFD0 U1745 ( .I(n1895), .Z(n1894) );
  BUFFD0 U1746 ( .I(n1896), .Z(n1895) );
  BUFFD0 U1747 ( .I(n1897), .Z(n1896) );
  BUFFD0 U1748 ( .I(n1898), .Z(n1897) );
  BUFFD0 U1749 ( .I(n1899), .Z(n1898) );
  BUFFD0 U1750 ( .I(n1900), .Z(n1899) );
  BUFFD0 U1751 ( .I(n1901), .Z(n1900) );
  BUFFD0 U1752 ( .I(n1902), .Z(n1901) );
  BUFFD0 U1753 ( .I(n1903), .Z(n1902) );
  BUFFD0 U1754 ( .I(n1904), .Z(n1903) );
  BUFFD0 U1755 ( .I(n1905), .Z(n1904) );
  BUFFD0 U1756 ( .I(n1906), .Z(n1905) );
  BUFFD0 U1757 ( .I(n1907), .Z(n1906) );
  BUFFD0 U1758 ( .I(n1908), .Z(n1907) );
  BUFFD0 U1759 ( .I(n1909), .Z(n1908) );
  BUFFD0 U1760 ( .I(n1910), .Z(n1909) );
  BUFFD0 U1761 ( .I(n1911), .Z(n1910) );
  BUFFD0 U1762 ( .I(n1912), .Z(n1911) );
  BUFFD0 U1763 ( .I(n1913), .Z(n1912) );
  BUFFD0 U1764 ( .I(n1914), .Z(n1913) );
  BUFFD0 U1765 ( .I(n1915), .Z(n1914) );
  BUFFD0 U1766 ( .I(n1916), .Z(n1915) );
  BUFFD0 U1767 ( .I(n1917), .Z(n1916) );
  BUFFD0 U1768 ( .I(n1918), .Z(n1917) );
  BUFFD0 U1769 ( .I(n1919), .Z(n1918) );
  BUFFD0 U1770 ( .I(n1920), .Z(n1919) );
  BUFFD0 U1771 ( .I(n1921), .Z(n1920) );
  BUFFD0 U1772 ( .I(n1922), .Z(n1921) );
  BUFFD0 U1773 ( .I(n1923), .Z(n1922) );
  BUFFD0 U1774 ( .I(n1924), .Z(n1923) );
  BUFFD0 U1775 ( .I(n1925), .Z(n1924) );
  BUFFD0 U1776 ( .I(n1926), .Z(n1925) );
  BUFFD0 U1777 ( .I(n1927), .Z(n1926) );
  BUFFD0 U1778 ( .I(n1928), .Z(n1927) );
  BUFFD0 U1779 ( .I(n1929), .Z(n1928) );
  BUFFD0 U1780 ( .I(n1930), .Z(n1929) );
  BUFFD0 U1781 ( .I(n1931), .Z(n1930) );
  BUFFD0 U1782 ( .I(n1932), .Z(n1931) );
  BUFFD0 U1783 ( .I(n1933), .Z(n1932) );
  BUFFD0 U1784 ( .I(n1934), .Z(n1933) );
  BUFFD0 U1785 ( .I(n1935), .Z(n1934) );
  BUFFD0 U1786 ( .I(n1936), .Z(n1935) );
  BUFFD0 U1787 ( .I(n1937), .Z(n1936) );
  BUFFD0 U1788 ( .I(n1938), .Z(n1937) );
  BUFFD0 U1789 ( .I(n1939), .Z(n1938) );
  BUFFD0 U1790 ( .I(n1940), .Z(n1939) );
  BUFFD0 U1791 ( .I(n1941), .Z(n1940) );
  BUFFD0 U1792 ( .I(n1942), .Z(n1941) );
  BUFFD0 U1793 ( .I(n1943), .Z(n1942) );
  BUFFD0 U1794 ( .I(n1944), .Z(n1943) );
  BUFFD0 U1795 ( .I(n1945), .Z(n1944) );
  BUFFD0 U1796 ( .I(n1946), .Z(n1945) );
  BUFFD0 U1797 ( .I(n1947), .Z(n1946) );
  BUFFD0 U1798 ( .I(n1948), .Z(n1947) );
  BUFFD0 U1799 ( .I(n1949), .Z(n1948) );
  BUFFD0 U1800 ( .I(n1950), .Z(n1949) );
  BUFFD0 U1801 ( .I(n1951), .Z(n1950) );
  BUFFD0 U1802 ( .I(n1952), .Z(n1951) );
  BUFFD0 U1803 ( .I(n1953), .Z(n1952) );
  BUFFD0 U1804 ( .I(n1954), .Z(n1953) );
  BUFFD0 U1805 ( .I(n1955), .Z(n1954) );
  BUFFD0 U1806 ( .I(n1956), .Z(n1955) );
  BUFFD0 U1807 ( .I(n1957), .Z(n1956) );
  BUFFD0 U1808 ( .I(n1958), .Z(n1957) );
  BUFFD0 U1809 ( .I(n1959), .Z(n1958) );
  BUFFD0 U1810 ( .I(n1960), .Z(n1959) );
  BUFFD0 U1811 ( .I(n1961), .Z(n1960) );
  BUFFD0 U1812 ( .I(n1962), .Z(n1961) );
  BUFFD0 U1813 ( .I(n1963), .Z(n1962) );
  BUFFD0 U1814 ( .I(n1964), .Z(n1963) );
  BUFFD0 U1815 ( .I(n1965), .Z(n1964) );
  BUFFD0 U1816 ( .I(n1966), .Z(n1965) );
  BUFFD0 U1817 ( .I(n1967), .Z(n1966) );
  BUFFD0 U1818 ( .I(n1968), .Z(n1967) );
  BUFFD0 U1819 ( .I(n1969), .Z(n1968) );
  BUFFD0 U1820 ( .I(n1970), .Z(n1969) );
  BUFFD0 U1821 ( .I(n1971), .Z(n1970) );
  BUFFD0 U1822 ( .I(n1972), .Z(n1971) );
  BUFFD0 U1823 ( .I(n1973), .Z(n1972) );
  BUFFD0 U1824 ( .I(n1974), .Z(n1973) );
  BUFFD0 U1825 ( .I(n1975), .Z(n1974) );
  BUFFD0 U1826 ( .I(n1976), .Z(n1975) );
  BUFFD0 U1827 ( .I(n1977), .Z(n1976) );
  BUFFD0 U1828 ( .I(n1978), .Z(n1977) );
  BUFFD0 U1829 ( .I(n1979), .Z(n1978) );
  BUFFD0 U1830 ( .I(n1980), .Z(n1979) );
  BUFFD0 U1831 ( .I(n1981), .Z(n1980) );
  BUFFD0 U1832 ( .I(n1982), .Z(n1981) );
  BUFFD0 U1833 ( .I(n1983), .Z(n1982) );
  BUFFD0 U1834 ( .I(n1984), .Z(n1983) );
  BUFFD0 U1835 ( .I(n1985), .Z(n1984) );
  BUFFD0 U1836 ( .I(n1986), .Z(n1985) );
  BUFFD0 U1837 ( .I(n1987), .Z(n1986) );
  BUFFD0 U1838 ( .I(n1988), .Z(n1987) );
  BUFFD0 U1839 ( .I(n1989), .Z(n1988) );
  BUFFD0 U1840 ( .I(n1990), .Z(n1989) );
  BUFFD0 U1841 ( .I(n1991), .Z(n1990) );
  BUFFD0 U1842 ( .I(n1992), .Z(n1991) );
  BUFFD0 U1843 ( .I(n1993), .Z(n1992) );
  BUFFD0 U1844 ( .I(n1994), .Z(n1993) );
  BUFFD0 U1845 ( .I(n1995), .Z(n1994) );
  BUFFD0 U1846 ( .I(n1996), .Z(n1995) );
  BUFFD0 U1847 ( .I(n1997), .Z(n1996) );
  BUFFD0 U1848 ( .I(n1998), .Z(n1997) );
  BUFFD0 U1849 ( .I(n1999), .Z(n1998) );
  BUFFD0 U1850 ( .I(n2000), .Z(n1999) );
  BUFFD0 U1851 ( .I(n2001), .Z(n2000) );
  BUFFD0 U1852 ( .I(n2002), .Z(n2001) );
  BUFFD0 U1853 ( .I(n2003), .Z(n2002) );
  BUFFD0 U1854 ( .I(n2004), .Z(n2003) );
  BUFFD0 U1855 ( .I(n2005), .Z(n2004) );
  BUFFD0 U1856 ( .I(n2006), .Z(n2005) );
  BUFFD0 U1857 ( .I(n2007), .Z(n2006) );
  BUFFD0 U1858 ( .I(n2008), .Z(n2007) );
  BUFFD0 U1859 ( .I(n2009), .Z(n2008) );
  BUFFD0 U1860 ( .I(n2010), .Z(n2009) );
  BUFFD0 U1861 ( .I(n2011), .Z(n2010) );
  BUFFD0 U1862 ( .I(n2012), .Z(n2011) );
  BUFFD0 U1863 ( .I(n2013), .Z(n2012) );
  BUFFD0 U1864 ( .I(n2014), .Z(n2013) );
  BUFFD0 U1865 ( .I(n2015), .Z(n2014) );
  BUFFD0 U1866 ( .I(n2016), .Z(n2015) );
  BUFFD0 U1867 ( .I(n2017), .Z(n2016) );
  BUFFD0 U1868 ( .I(n2018), .Z(n2017) );
  BUFFD0 U1869 ( .I(n2019), .Z(n2018) );
  BUFFD0 U1870 ( .I(n2020), .Z(n2019) );
  BUFFD0 U1871 ( .I(n2021), .Z(n2020) );
  BUFFD0 U1872 ( .I(n2022), .Z(n2021) );
  BUFFD0 U1873 ( .I(n2023), .Z(n2022) );
  BUFFD0 U1874 ( .I(n2024), .Z(n2023) );
  BUFFD0 U1875 ( .I(n2025), .Z(n2024) );
  BUFFD0 U1876 ( .I(n2026), .Z(n2025) );
  BUFFD0 U1877 ( .I(n2027), .Z(n2026) );
  BUFFD0 U1878 ( .I(n2028), .Z(n2027) );
  BUFFD0 U1879 ( .I(n2029), .Z(n2028) );
  BUFFD0 U1880 ( .I(n2030), .Z(n2029) );
  BUFFD0 U1881 ( .I(n2031), .Z(n2030) );
  BUFFD0 U1882 ( .I(n2032), .Z(n2031) );
  BUFFD0 U1883 ( .I(n2033), .Z(n2032) );
  BUFFD0 U1884 ( .I(n2034), .Z(n2033) );
  BUFFD0 U1885 ( .I(n2035), .Z(n2034) );
  BUFFD0 U1886 ( .I(n2036), .Z(n2035) );
  BUFFD0 U1887 ( .I(n2037), .Z(n2036) );
  BUFFD0 U1888 ( .I(n2039), .Z(n2037) );
  INVD0 U1889 ( .I(n2038), .ZN(n2039) );
  CKNXD16 U1890 ( .I(SerIn), .ZN(n2038) );
  BUFFD0 U1891 ( .I(n2041), .Z(n2040) );
  BUFFD0 U1892 ( .I(n2042), .Z(n2041) );
  BUFFD0 U1893 ( .I(n2043), .Z(n2042) );
  BUFFD0 U1894 ( .I(n2044), .Z(n2043) );
  BUFFD0 U1895 ( .I(n2045), .Z(n2044) );
  BUFFD0 U1896 ( .I(n2046), .Z(n2045) );
  BUFFD0 U1897 ( .I(n2047), .Z(n2046) );
  BUFFD0 U1898 ( .I(n2048), .Z(n2047) );
  BUFFD0 U1899 ( .I(n2049), .Z(n2048) );
  BUFFD0 U1900 ( .I(n2050), .Z(n2049) );
  BUFFD0 U1901 ( .I(n2051), .Z(n2050) );
  BUFFD0 U1902 ( .I(n2052), .Z(n2051) );
  BUFFD0 U1903 ( .I(n2053), .Z(n2052) );
  BUFFD0 U1904 ( .I(n2054), .Z(n2053) );
  BUFFD0 U1905 ( .I(n2055), .Z(n2054) );
  BUFFD0 U1906 ( .I(n2056), .Z(n2055) );
  BUFFD0 U1907 ( .I(n2461), .Z(n2056) );
  BUFFD0 U1908 ( .I(n2058), .Z(n2057) );
  BUFFD0 U1909 ( .I(n2059), .Z(n2058) );
  BUFFD0 U1910 ( .I(n2060), .Z(n2059) );
  BUFFD0 U1911 ( .I(n2061), .Z(n2060) );
  BUFFD0 U1912 ( .I(n2062), .Z(n2061) );
  BUFFD0 U1913 ( .I(n2063), .Z(n2062) );
  BUFFD0 U1914 ( .I(n2064), .Z(n2063) );
  BUFFD0 U1915 ( .I(n2065), .Z(n2064) );
  BUFFD0 U1916 ( .I(n2066), .Z(n2065) );
  BUFFD0 U1917 ( .I(n2067), .Z(n2066) );
  BUFFD0 U1918 ( .I(n2068), .Z(n2067) );
  BUFFD0 U1919 ( .I(n2069), .Z(n2068) );
  BUFFD0 U1920 ( .I(n2070), .Z(n2069) );
  BUFFD0 U1921 ( .I(n2071), .Z(n2070) );
  BUFFD0 U1922 ( .I(n2072), .Z(n2071) );
  BUFFD0 U1923 ( .I(n2073), .Z(n2072) );
  BUFFD0 U1924 ( .I(n2074), .Z(n2073) );
  BUFFD0 U1925 ( .I(FrameSR[19]), .Z(n2074) );
  BUFFD0 U1926 ( .I(n2076), .Z(n2075) );
  BUFFD0 U1927 ( .I(n2077), .Z(n2076) );
  BUFFD0 U1928 ( .I(n2078), .Z(n2077) );
  BUFFD0 U1929 ( .I(n2079), .Z(n2078) );
  BUFFD0 U1930 ( .I(n2080), .Z(n2079) );
  BUFFD0 U1931 ( .I(n2081), .Z(n2080) );
  BUFFD0 U1932 ( .I(n2082), .Z(n2081) );
  BUFFD0 U1933 ( .I(n2083), .Z(n2082) );
  BUFFD0 U1934 ( .I(n2084), .Z(n2083) );
  BUFFD0 U1935 ( .I(n2085), .Z(n2084) );
  BUFFD0 U1936 ( .I(n2086), .Z(n2085) );
  BUFFD0 U1937 ( .I(n2087), .Z(n2086) );
  BUFFD0 U1938 ( .I(n2088), .Z(n2087) );
  BUFFD0 U1939 ( .I(n2089), .Z(n2088) );
  BUFFD0 U1940 ( .I(n2090), .Z(n2089) );
  BUFFD0 U1941 ( .I(n2091), .Z(n2090) );
  BUFFD0 U1942 ( .I(n2092), .Z(n2091) );
  BUFFD0 U1943 ( .I(FrameSR[33]), .Z(n2092) );
  BUFFD0 U1944 ( .I(n2094), .Z(n2093) );
  BUFFD0 U1945 ( .I(n2095), .Z(n2094) );
  BUFFD0 U1946 ( .I(n2096), .Z(n2095) );
  BUFFD0 U1947 ( .I(n2097), .Z(n2096) );
  BUFFD0 U1948 ( .I(n2098), .Z(n2097) );
  BUFFD0 U1949 ( .I(n2099), .Z(n2098) );
  BUFFD0 U1950 ( .I(n2100), .Z(n2099) );
  BUFFD0 U1951 ( .I(n2101), .Z(n2100) );
  BUFFD0 U1952 ( .I(n2102), .Z(n2101) );
  BUFFD0 U1953 ( .I(n2103), .Z(n2102) );
  BUFFD0 U1954 ( .I(n2104), .Z(n2103) );
  BUFFD0 U1955 ( .I(n2105), .Z(n2104) );
  BUFFD0 U1956 ( .I(n2106), .Z(n2105) );
  BUFFD0 U1957 ( .I(n2107), .Z(n2106) );
  BUFFD0 U1958 ( .I(n2108), .Z(n2107) );
  BUFFD0 U1959 ( .I(n2109), .Z(n2108) );
  BUFFD0 U1960 ( .I(n2110), .Z(n2109) );
  BUFFD0 U1961 ( .I(FrameSR[48]), .Z(n2110) );
  BUFFD0 U1962 ( .I(n2112), .Z(n2111) );
  BUFFD0 U1963 ( .I(n2113), .Z(n2112) );
  BUFFD0 U1964 ( .I(n2114), .Z(n2113) );
  BUFFD0 U1965 ( .I(n2115), .Z(n2114) );
  BUFFD0 U1966 ( .I(n2116), .Z(n2115) );
  BUFFD0 U1967 ( .I(n2118), .Z(n2116) );
  BUFFD0 U1968 ( .I(FrameSR[1]), .Z(n2117) );
  BUFFD0 U1969 ( .I(n2119), .Z(n2118) );
  BUFFD0 U1970 ( .I(n2120), .Z(n2119) );
  BUFFD0 U1971 ( .I(n2121), .Z(n2120) );
  BUFFD0 U1972 ( .I(n2122), .Z(n2121) );
  BUFFD0 U1973 ( .I(n2123), .Z(n2122) );
  BUFFD0 U1974 ( .I(n2124), .Z(n2123) );
  BUFFD0 U1975 ( .I(n2125), .Z(n2124) );
  BUFFD0 U1976 ( .I(n2126), .Z(n2125) );
  BUFFD0 U1977 ( .I(n2127), .Z(n2126) );
  BUFFD0 U1978 ( .I(n2128), .Z(n2127) );
  BUFFD0 U1979 ( .I(n2117), .Z(n2128) );
  BUFFD0 U1980 ( .I(n2130), .Z(n2129) );
  BUFFD0 U1981 ( .I(n2131), .Z(n2130) );
  BUFFD0 U1982 ( .I(n2132), .Z(n2131) );
  BUFFD0 U1983 ( .I(n2133), .Z(n2132) );
  BUFFD0 U1984 ( .I(n2134), .Z(n2133) );
  BUFFD0 U1985 ( .I(n2136), .Z(n2134) );
  BUFFD0 U1986 ( .I(FrameSR[5]), .Z(n2135) );
  BUFFD0 U1987 ( .I(n2137), .Z(n2136) );
  BUFFD0 U1988 ( .I(n2138), .Z(n2137) );
  BUFFD0 U1989 ( .I(n2139), .Z(n2138) );
  BUFFD0 U1990 ( .I(n2140), .Z(n2139) );
  BUFFD0 U1991 ( .I(n2141), .Z(n2140) );
  BUFFD0 U1992 ( .I(n2142), .Z(n2141) );
  BUFFD0 U1993 ( .I(n2143), .Z(n2142) );
  BUFFD0 U1994 ( .I(n2144), .Z(n2143) );
  BUFFD0 U1995 ( .I(n2145), .Z(n2144) );
  BUFFD0 U1996 ( .I(n2146), .Z(n2145) );
  BUFFD0 U1997 ( .I(n2135), .Z(n2146) );
  CKBD0 U1998 ( .CLK(FrameSR[17]), .C(n2164) );
  BUFFD0 U1999 ( .I(n2148), .Z(n2147) );
  BUFFD0 U2000 ( .I(n2149), .Z(n2148) );
  BUFFD0 U2001 ( .I(n2150), .Z(n2149) );
  BUFFD0 U2002 ( .I(n2151), .Z(n2150) );
  BUFFD0 U2003 ( .I(n2152), .Z(n2151) );
  BUFFD0 U2004 ( .I(n2153), .Z(n2152) );
  BUFFD0 U2005 ( .I(n2154), .Z(n2153) );
  BUFFD0 U2006 ( .I(n2155), .Z(n2154) );
  BUFFD0 U2007 ( .I(n2156), .Z(n2155) );
  BUFFD0 U2008 ( .I(n2157), .Z(n2156) );
  BUFFD0 U2009 ( .I(n2158), .Z(n2157) );
  BUFFD0 U2010 ( .I(n2159), .Z(n2158) );
  BUFFD0 U2011 ( .I(n2160), .Z(n2159) );
  BUFFD0 U2012 ( .I(n2161), .Z(n2160) );
  BUFFD0 U2013 ( .I(n2162), .Z(n2161) );
  BUFFD0 U2014 ( .I(n2163), .Z(n2162) );
  BUFFD0 U2015 ( .I(n2164), .Z(n2163) );
  CKBD0 U2016 ( .CLK(FrameSR[32]), .C(n2182) );
  BUFFD0 U2017 ( .I(n2166), .Z(n2165) );
  BUFFD0 U2018 ( .I(n2167), .Z(n2166) );
  BUFFD0 U2019 ( .I(n2168), .Z(n2167) );
  BUFFD0 U2020 ( .I(n2169), .Z(n2168) );
  BUFFD0 U2021 ( .I(n2170), .Z(n2169) );
  BUFFD0 U2022 ( .I(n2171), .Z(n2170) );
  BUFFD0 U2023 ( .I(n2172), .Z(n2171) );
  BUFFD0 U2024 ( .I(n2173), .Z(n2172) );
  BUFFD0 U2025 ( .I(n2174), .Z(n2173) );
  BUFFD0 U2026 ( .I(n2175), .Z(n2174) );
  BUFFD0 U2027 ( .I(n2176), .Z(n2175) );
  BUFFD0 U2028 ( .I(n2177), .Z(n2176) );
  BUFFD0 U2029 ( .I(n2178), .Z(n2177) );
  BUFFD0 U2030 ( .I(n2179), .Z(n2178) );
  BUFFD0 U2031 ( .I(n2180), .Z(n2179) );
  BUFFD0 U2032 ( .I(n2181), .Z(n2180) );
  BUFFD0 U2033 ( .I(n2182), .Z(n2181) );
  CKBD0 U2034 ( .CLK(FrameSR[47]), .C(n2200) );
  BUFFD0 U2035 ( .I(n2184), .Z(n2183) );
  BUFFD0 U2036 ( .I(n2185), .Z(n2184) );
  BUFFD0 U2037 ( .I(n2186), .Z(n2185) );
  BUFFD0 U2038 ( .I(n2187), .Z(n2186) );
  BUFFD0 U2039 ( .I(n2188), .Z(n2187) );
  BUFFD0 U2040 ( .I(n2189), .Z(n2188) );
  BUFFD0 U2041 ( .I(n2190), .Z(n2189) );
  BUFFD0 U2042 ( .I(n2191), .Z(n2190) );
  BUFFD0 U2043 ( .I(n2192), .Z(n2191) );
  BUFFD0 U2044 ( .I(n2193), .Z(n2192) );
  BUFFD0 U2045 ( .I(n2194), .Z(n2193) );
  BUFFD0 U2046 ( .I(n2195), .Z(n2194) );
  BUFFD0 U2047 ( .I(n2196), .Z(n2195) );
  BUFFD0 U2048 ( .I(n2197), .Z(n2196) );
  BUFFD0 U2049 ( .I(n2198), .Z(n2197) );
  BUFFD0 U2050 ( .I(n2199), .Z(n2198) );
  BUFFD0 U2051 ( .I(n2200), .Z(n2199) );
  BUFFD0 U2052 ( .I(n2202), .Z(n2201) );
  BUFFD0 U2053 ( .I(n2203), .Z(n2202) );
  BUFFD0 U2054 ( .I(n2204), .Z(n2203) );
  BUFFD0 U2055 ( .I(n2205), .Z(n2204) );
  BUFFD0 U2056 ( .I(n2206), .Z(n2205) );
  BUFFD0 U2057 ( .I(n2208), .Z(n2206) );
  BUFFD0 U2058 ( .I(FrameSR[0]), .Z(n2207) );
  BUFFD0 U2059 ( .I(n2209), .Z(n2208) );
  BUFFD0 U2060 ( .I(n2210), .Z(n2209) );
  BUFFD0 U2061 ( .I(n2211), .Z(n2210) );
  BUFFD0 U2062 ( .I(n2212), .Z(n2211) );
  BUFFD0 U2063 ( .I(n2213), .Z(n2212) );
  BUFFD0 U2064 ( .I(n2214), .Z(n2213) );
  BUFFD0 U2065 ( .I(n2215), .Z(n2214) );
  BUFFD0 U2066 ( .I(n2216), .Z(n2215) );
  BUFFD0 U2067 ( .I(n2217), .Z(n2216) );
  BUFFD0 U2068 ( .I(n2218), .Z(n2217) );
  BUFFD0 U2069 ( .I(n2207), .Z(n2218) );
  BUFFD0 U2070 ( .I(n2220), .Z(n2219) );
  BUFFD0 U2071 ( .I(n2221), .Z(n2220) );
  BUFFD0 U2072 ( .I(n2222), .Z(n2221) );
  BUFFD0 U2073 ( .I(n2223), .Z(n2222) );
  BUFFD0 U2074 ( .I(n2224), .Z(n2223) );
  BUFFD0 U2075 ( .I(n2226), .Z(n2224) );
  BUFFD0 U2076 ( .I(FrameSR[2]), .Z(n2225) );
  BUFFD0 U2077 ( .I(n2227), .Z(n2226) );
  BUFFD0 U2078 ( .I(n2228), .Z(n2227) );
  BUFFD0 U2079 ( .I(n2229), .Z(n2228) );
  BUFFD0 U2080 ( .I(n2230), .Z(n2229) );
  BUFFD0 U2081 ( .I(n2231), .Z(n2230) );
  BUFFD0 U2082 ( .I(n2232), .Z(n2231) );
  BUFFD0 U2083 ( .I(n2233), .Z(n2232) );
  BUFFD0 U2084 ( .I(n2234), .Z(n2233) );
  BUFFD0 U2085 ( .I(n2235), .Z(n2234) );
  BUFFD0 U2086 ( .I(n2236), .Z(n2235) );
  BUFFD0 U2087 ( .I(n2225), .Z(n2236) );
  BUFFD0 U2088 ( .I(n2238), .Z(n2237) );
  BUFFD0 U2089 ( .I(n2239), .Z(n2238) );
  BUFFD0 U2090 ( .I(n2240), .Z(n2239) );
  BUFFD0 U2091 ( .I(n2241), .Z(n2240) );
  BUFFD0 U2092 ( .I(n2242), .Z(n2241) );
  BUFFD0 U2093 ( .I(n2244), .Z(n2242) );
  BUFFD0 U2094 ( .I(FrameSR[4]), .Z(n2243) );
  BUFFD0 U2095 ( .I(n2245), .Z(n2244) );
  BUFFD0 U2096 ( .I(n2246), .Z(n2245) );
  BUFFD0 U2097 ( .I(n2247), .Z(n2246) );
  BUFFD0 U2098 ( .I(n2248), .Z(n2247) );
  BUFFD0 U2099 ( .I(n2249), .Z(n2248) );
  BUFFD0 U2100 ( .I(n2250), .Z(n2249) );
  BUFFD0 U2101 ( .I(n2251), .Z(n2250) );
  BUFFD0 U2102 ( .I(n2252), .Z(n2251) );
  BUFFD0 U2103 ( .I(n2253), .Z(n2252) );
  BUFFD0 U2104 ( .I(n2254), .Z(n2253) );
  BUFFD0 U2105 ( .I(n2243), .Z(n2254) );
  BUFFD0 U2106 ( .I(n2256), .Z(n2255) );
  BUFFD0 U2107 ( .I(n2257), .Z(n2256) );
  BUFFD0 U2108 ( .I(n2258), .Z(n2257) );
  BUFFD0 U2109 ( .I(n2259), .Z(n2258) );
  BUFFD0 U2110 ( .I(n2260), .Z(n2259) );
  BUFFD0 U2111 ( .I(n2262), .Z(n2260) );
  BUFFD0 U2112 ( .I(FrameSR[6]), .Z(n2261) );
  BUFFD0 U2113 ( .I(n2263), .Z(n2262) );
  BUFFD0 U2114 ( .I(n2264), .Z(n2263) );
  BUFFD0 U2115 ( .I(n2265), .Z(n2264) );
  BUFFD0 U2116 ( .I(n2266), .Z(n2265) );
  BUFFD0 U2117 ( .I(n2267), .Z(n2266) );
  BUFFD0 U2118 ( .I(n2268), .Z(n2267) );
  BUFFD0 U2119 ( .I(n2269), .Z(n2268) );
  BUFFD0 U2120 ( .I(n2270), .Z(n2269) );
  BUFFD0 U2121 ( .I(n2271), .Z(n2270) );
  BUFFD0 U2122 ( .I(n2272), .Z(n2271) );
  BUFFD0 U2123 ( .I(n2261), .Z(n2272) );
  BUFFD0 U2124 ( .I(n2274), .Z(n2273) );
  BUFFD0 U2125 ( .I(n2275), .Z(n2274) );
  BUFFD0 U2126 ( .I(n2276), .Z(n2275) );
  BUFFD0 U2127 ( .I(n2277), .Z(n2276) );
  BUFFD0 U2128 ( .I(n2278), .Z(n2277) );
  BUFFD0 U2129 ( .I(n2279), .Z(n2278) );
  BUFFD0 U2130 ( .I(n2280), .Z(n2279) );
  BUFFD0 U2131 ( .I(n2281), .Z(n2280) );
  BUFFD0 U2132 ( .I(n2282), .Z(n2281) );
  BUFFD0 U2133 ( .I(n2283), .Z(n2282) );
  BUFFD0 U2134 ( .I(n2284), .Z(n2283) );
  BUFFD0 U2135 ( .I(n2285), .Z(n2284) );
  BUFFD0 U2136 ( .I(n2286), .Z(n2285) );
  BUFFD0 U2137 ( .I(n2287), .Z(n2286) );
  BUFFD0 U2138 ( .I(n2288), .Z(n2287) );
  BUFFD0 U2139 ( .I(n2289), .Z(n2288) );
  BUFFD0 U2140 ( .I(n2290), .Z(n2289) );
  BUFFD0 U2141 ( .I(FrameSR[20]), .Z(n2290) );
  BUFFD0 U2142 ( .I(n2292), .Z(n2291) );
  BUFFD0 U2143 ( .I(n2293), .Z(n2292) );
  BUFFD0 U2144 ( .I(n2294), .Z(n2293) );
  BUFFD0 U2145 ( .I(n2295), .Z(n2294) );
  BUFFD0 U2146 ( .I(n2296), .Z(n2295) );
  BUFFD0 U2147 ( .I(n2297), .Z(n2296) );
  BUFFD0 U2148 ( .I(n2298), .Z(n2297) );
  BUFFD0 U2149 ( .I(n2299), .Z(n2298) );
  BUFFD0 U2150 ( .I(n2300), .Z(n2299) );
  BUFFD0 U2151 ( .I(n2301), .Z(n2300) );
  BUFFD0 U2152 ( .I(n2302), .Z(n2301) );
  BUFFD0 U2153 ( .I(n2303), .Z(n2302) );
  BUFFD0 U2154 ( .I(n2304), .Z(n2303) );
  BUFFD0 U2155 ( .I(n2305), .Z(n2304) );
  BUFFD0 U2156 ( .I(n2306), .Z(n2305) );
  BUFFD0 U2157 ( .I(n2307), .Z(n2306) );
  BUFFD0 U2158 ( .I(n2308), .Z(n2307) );
  BUFFD0 U2159 ( .I(FrameSR[34]), .Z(n2308) );
  BUFFD0 U2160 ( .I(n2310), .Z(n2309) );
  BUFFD0 U2161 ( .I(n2311), .Z(n2310) );
  BUFFD0 U2162 ( .I(n2312), .Z(n2311) );
  BUFFD0 U2163 ( .I(n2313), .Z(n2312) );
  BUFFD0 U2164 ( .I(n2314), .Z(n2313) );
  BUFFD0 U2165 ( .I(n2315), .Z(n2314) );
  BUFFD0 U2166 ( .I(n2316), .Z(n2315) );
  BUFFD0 U2167 ( .I(n2317), .Z(n2316) );
  BUFFD0 U2168 ( .I(n2318), .Z(n2317) );
  BUFFD0 U2169 ( .I(n2319), .Z(n2318) );
  BUFFD0 U2170 ( .I(n2320), .Z(n2319) );
  BUFFD0 U2171 ( .I(n2321), .Z(n2320) );
  BUFFD0 U2172 ( .I(n2322), .Z(n2321) );
  BUFFD0 U2173 ( .I(n2323), .Z(n2322) );
  BUFFD0 U2174 ( .I(n2324), .Z(n2323) );
  BUFFD0 U2175 ( .I(n2325), .Z(n2324) );
  BUFFD0 U2176 ( .I(n2326), .Z(n2325) );
  BUFFD0 U2177 ( .I(FrameSR[49]), .Z(n2326) );
  BUFFD0 U2178 ( .I(n2328), .Z(n2327) );
  BUFFD0 U2179 ( .I(n2329), .Z(n2328) );
  BUFFD0 U2180 ( .I(n2330), .Z(n2329) );
  BUFFD0 U2181 ( .I(n2331), .Z(n2330) );
  BUFFD0 U2182 ( .I(n2332), .Z(n2331) );
  BUFFD0 U2183 ( .I(n2333), .Z(n2332) );
  BUFFD0 U2184 ( .I(n2334), .Z(n2333) );
  BUFFD0 U2185 ( .I(n2335), .Z(n2334) );
  BUFFD0 U2186 ( .I(n2336), .Z(n2335) );
  BUFFD0 U2187 ( .I(n2337), .Z(n2336) );
  BUFFD0 U2188 ( .I(n2338), .Z(n2337) );
  BUFFD0 U2189 ( .I(n2339), .Z(n2338) );
  BUFFD0 U2190 ( .I(n2340), .Z(n2339) );
  BUFFD0 U2191 ( .I(n2341), .Z(n2340) );
  BUFFD0 U2192 ( .I(n2342), .Z(n2341) );
  BUFFD0 U2193 ( .I(n2343), .Z(n2342) );
  BUFFD0 U2194 ( .I(n2344), .Z(n2343) );
  BUFFD0 U2195 ( .I(FrameSR[18]), .Z(n2344) );
  BUFFD0 U2196 ( .I(n2349), .Z(n2346) );
  BUFFD0 U2197 ( .I(n2348), .Z(n2347) );
  BUFFD0 U2198 ( .I(n2350), .Z(n2348) );
  BUFFD0 U2199 ( .I(n11), .Z(n2349) );
  BUFFD0 U2200 ( .I(n2351), .Z(n2350) );
  BUFFD0 U2201 ( .I(n2352), .Z(n2351) );
  BUFFD0 U2202 ( .I(n2353), .Z(n2352) );
  BUFFD0 U2203 ( .I(n2354), .Z(n2353) );
  BUFFD0 U2204 ( .I(n2355), .Z(n2354) );
  BUFFD0 U2205 ( .I(n2356), .Z(n2355) );
  BUFFD0 U2206 ( .I(n2357), .Z(n2356) );
  BUFFD0 U2207 ( .I(n2358), .Z(n2357) );
  BUFFD0 U2208 ( .I(n195), .Z(n2358) );
  CKAN2D0 U2209 ( .A1(N31), .A2(n2), .Z(N39) );
  BUFFD0 U2210 ( .I(n2360), .Z(n2359) );
  BUFFD0 U2211 ( .I(n2361), .Z(n2360) );
  BUFFD0 U2212 ( .I(n2362), .Z(n2361) );
  BUFFD0 U2213 ( .I(n2363), .Z(n2362) );
  BUFFD0 U2214 ( .I(n2371), .Z(n2363) );
  BUFFD0 U2215 ( .I(n2365), .Z(n2364) );
  BUFFD0 U2216 ( .I(n2366), .Z(n2365) );
  BUFFD0 U2217 ( .I(n2367), .Z(n2366) );
  BUFFD0 U2218 ( .I(n2368), .Z(n2367) );
  BUFFD0 U2219 ( .I(n2369), .Z(n2368) );
  BUFFD0 U2220 ( .I(n2370), .Z(n2369) );
  BUFFD0 U2221 ( .I(n2372), .Z(n2370) );
  BUFFD0 U2222 ( .I(N39), .Z(n2371) );
  BUFFD0 U2223 ( .I(Count32[1]), .Z(n2372) );
  BUFFD0 U2224 ( .I(n2374), .Z(n2373) );
  BUFFD0 U2225 ( .I(n2376), .Z(n2374) );
  BUFFD0 U2226 ( .I(n2377), .Z(n2375) );
  BUFFD0 U2227 ( .I(n2378), .Z(n2376) );
  BUFFD0 U2228 ( .I(n2379), .Z(n2377) );
  BUFFD0 U2229 ( .I(n2382), .Z(n2378) );
  BUFFD0 U2230 ( .I(n2380), .Z(n2379) );
  BUFFD0 U2231 ( .I(n2381), .Z(n2380) );
  INVD0 U2232 ( .I(n3133), .ZN(n3132) );
  BUFFD0 U2233 ( .I(n263), .Z(n3133) );
  BUFFD0 U2234 ( .I(n2385), .Z(n2381) );
  BUFFD0 U2235 ( .I(n2383), .Z(n2382) );
  BUFFD0 U2236 ( .I(n2384), .Z(n2383) );
  BUFFD0 U2237 ( .I(n196), .Z(n2384) );
  BUFFD0 U2238 ( .I(n12), .Z(n2385) );
  CKBD0 U2239 ( .CLK(ParValidTimer[0]), .C(n2445) );
  CKXOR2D0 U2240 ( .A1(n2443), .A2(n6), .Z(n12) );
  BUFFD0 U2241 ( .I(n2387), .Z(n2386) );
  BUFFD0 U2242 ( .I(n2388), .Z(n2387) );
  BUFFD0 U2243 ( .I(n2389), .Z(n2388) );
  BUFFD0 U2244 ( .I(n2390), .Z(n2389) );
  BUFFD0 U2245 ( .I(n2391), .Z(n2390) );
  BUFFD0 U2246 ( .I(n2392), .Z(n2391) );
  BUFFD0 U2247 ( .I(n2393), .Z(n2392) );
  BUFFD0 U2248 ( .I(n2394), .Z(n2393) );
  BUFFD0 U2249 ( .I(n2395), .Z(n2394) );
  BUFFD0 U2250 ( .I(n2396), .Z(n2395) );
  BUFFD0 U2251 ( .I(n2397), .Z(n2396) );
  BUFFD0 U2252 ( .I(n2398), .Z(n2397) );
  BUFFD0 U2253 ( .I(n2399), .Z(n2398) );
  BUFFD0 U2254 ( .I(n2400), .Z(n2399) );
  BUFFD0 U2255 ( .I(N41), .Z(n2400) );
  BUFFD0 U2256 ( .I(n2402), .Z(n2401) );
  BUFFD0 U2257 ( .I(n2403), .Z(n2402) );
  BUFFD0 U2258 ( .I(n2404), .Z(n2403) );
  BUFFD0 U2259 ( .I(n2405), .Z(n2404) );
  BUFFD0 U2260 ( .I(n2406), .Z(n2405) );
  BUFFD0 U2261 ( .I(n2407), .Z(n2406) );
  BUFFD0 U2262 ( .I(n2408), .Z(n2407) );
  BUFFD0 U2263 ( .I(n2409), .Z(n2408) );
  BUFFD0 U2264 ( .I(n2410), .Z(n2409) );
  BUFFD0 U2265 ( .I(n2411), .Z(n2410) );
  BUFFD0 U2266 ( .I(n2412), .Z(n2411) );
  BUFFD0 U2267 ( .I(n2413), .Z(n2412) );
  BUFFD0 U2268 ( .I(n2414), .Z(n2413) );
  BUFFD0 U2269 ( .I(n2415), .Z(n2414) );
  BUFFD0 U2270 ( .I(N40), .Z(n2415) );
  BUFFD0 U2271 ( .I(n2417), .Z(n2416) );
  BUFFD0 U2272 ( .I(n2419), .Z(n2417) );
  BUFFD0 U2273 ( .I(n2420), .Z(n2418) );
  BUFFD0 U2274 ( .I(n2421), .Z(n2419) );
  BUFFD0 U2275 ( .I(n2422), .Z(n2420) );
  BUFFD0 U2276 ( .I(n2424), .Z(n2421) );
  BUFFD0 U2277 ( .I(n2423), .Z(n2422) );
  BUFFD0 U2278 ( .I(n2425), .Z(n2423) );
  BUFFD0 U2279 ( .I(N38), .Z(n2424) );
  BUFFD0 U2280 ( .I(n2426), .Z(n2425) );
  BUFFD0 U2281 ( .I(n2427), .Z(n2426) );
  BUFFD0 U2282 ( .I(n2428), .Z(n2427) );
  BUFFD0 U2283 ( .I(n2429), .Z(n2428) );
  BUFFD0 U2284 ( .I(Count32[0]), .Z(n2429) );
  CKNXD16 U2285 ( .I(SerValid), .ZN(n2430) );
  INVD1 U2286 ( .I(n2430), .ZN(n2431) );
  BUFFD0 U2287 ( .I(n2433), .Z(n2432) );
  BUFFD0 U2288 ( .I(n2434), .Z(n2433) );
  BUFFD0 U2289 ( .I(n2435), .Z(n2434) );
  BUFFD0 U2290 ( .I(n2436), .Z(n2435) );
  BUFFD0 U2291 ( .I(n2437), .Z(n2436) );
  BUFFD0 U2292 ( .I(n2438), .Z(n2437) );
  BUFFD0 U2293 ( .I(n2439), .Z(n2438) );
  BUFFD0 U2294 ( .I(n2440), .Z(n2439) );
  BUFFD0 U2295 ( .I(n2441), .Z(n2440) );
  BUFFD0 U2296 ( .I(n2442), .Z(n2441) );
  BUFFD0 U2297 ( .I(SerValid), .Z(n2442) );
  BUFFD0 U2298 ( .I(n264), .Z(n2443) );
  BUFFD0 U2299 ( .I(n262), .Z(n2444) );
  BUFFD0 U2300 ( .I(n2447), .Z(n2446) );
  BUFFD0 U2301 ( .I(n2448), .Z(n2447) );
  BUFFD0 U2302 ( .I(n2449), .Z(n2448) );
  BUFFD0 U2303 ( .I(n2450), .Z(n2449) );
  BUFFD0 U2304 ( .I(n2451), .Z(n2450) );
  BUFFD0 U2305 ( .I(n2452), .Z(n2451) );
  BUFFD0 U2306 ( .I(n2453), .Z(n2452) );
  BUFFD0 U2307 ( .I(n2454), .Z(n2453) );
  BUFFD0 U2308 ( .I(n2455), .Z(n2454) );
  BUFFD0 U2309 ( .I(n2456), .Z(n2455) );
  BUFFD0 U2310 ( .I(n2457), .Z(n2456) );
  BUFFD0 U2311 ( .I(n2458), .Z(n2457) );
  BUFFD0 U2312 ( .I(n2459), .Z(n2458) );
  BUFFD0 U2313 ( .I(n193), .Z(n2459) );
  CKBD0 U2314 ( .CLK(ParValidTimer[1]), .C(n2460) );
  BUFFD0 U2315 ( .I(FrameSR[3]), .Z(n2461) );
  BUFFD0 U2316 ( .I(FrameSR[7]), .Z(n2462) );
  BUFFD0 U2317 ( .I(n45), .Z(n2463) );
  BUFFD0 U2318 ( .I(n3141), .Z(n2464) );
  AN4D0 U2319 ( .A1(n50), .A2(n51), .A3(n52), .A4(n53), .Z(n47) );
  BUFFD0 U2320 ( .I(n2466), .Z(n2465) );
  BUFFD0 U2321 ( .I(n2467), .Z(n2466) );
  BUFFD0 U2322 ( .I(n2468), .Z(n2467) );
  BUFFD0 U2323 ( .I(n2469), .Z(n2468) );
  BUFFD0 U2324 ( .I(n2470), .Z(n2469) );
  BUFFD0 U2325 ( .I(n2471), .Z(n2470) );
  BUFFD0 U2326 ( .I(n2472), .Z(n2471) );
  BUFFD0 U2327 ( .I(n2473), .Z(n2472) );
  BUFFD0 U2328 ( .I(n2474), .Z(n2473) );
  BUFFD0 U2329 ( .I(n2475), .Z(n2474) );
  BUFFD0 U2330 ( .I(n2476), .Z(n2475) );
  BUFFD0 U2331 ( .I(n2477), .Z(n2476) );
  BUFFD0 U2332 ( .I(n2478), .Z(n2477) );
  BUFFD0 U2333 ( .I(N47), .Z(n2478) );
  BUFFD0 U2334 ( .I(n192), .Z(n2479) );
  BUFFD0 U2335 ( .I(n2482), .Z(n2481) );
  BUFFD0 U2336 ( .I(n2483), .Z(n2482) );
  BUFFD0 U2337 ( .I(n2484), .Z(n2483) );
  BUFFD0 U2338 ( .I(n2485), .Z(n2484) );
  BUFFD0 U2339 ( .I(n2486), .Z(n2485) );
  BUFFD0 U2340 ( .I(n2487), .Z(n2486) );
  BUFFD0 U2341 ( .I(n2488), .Z(n2487) );
  BUFFD0 U2342 ( .I(n2489), .Z(n2488) );
  BUFFD0 U2343 ( .I(n2490), .Z(n2489) );
  BUFFD0 U2344 ( .I(n2491), .Z(n2490) );
  BUFFD0 U2345 ( .I(n2493), .Z(n2491) );
  CKBD0 U2346 ( .CLK(n3098), .C(n2492) );
  BUFFD0 U2347 ( .I(n2494), .Z(n2493) );
  BUFFD0 U2348 ( .I(n2479), .Z(n2494) );
  OAI21D0 U2349 ( .A1(n3), .A2(n2492), .B(n3133), .ZN(n192) );
  BUFFD0 U2350 ( .I(n2497), .Z(n2495) );
  BUFFD0 U2351 ( .I(n228), .Z(n2496) );
  BUFFD0 U2352 ( .I(n2498), .Z(n2497) );
  BUFFD0 U2353 ( .I(n2499), .Z(n2498) );
  BUFFD0 U2354 ( .I(n2500), .Z(n2499) );
  BUFFD0 U2355 ( .I(n2501), .Z(n2500) );
  BUFFD0 U2356 ( .I(n2502), .Z(n2501) );
  BUFFD0 U2357 ( .I(n2503), .Z(n2502) );
  BUFFD0 U2358 ( .I(n2504), .Z(n2503) );
  BUFFD0 U2359 ( .I(n2505), .Z(n2504) );
  BUFFD0 U2360 ( .I(n2506), .Z(n2505) );
  BUFFD0 U2361 ( .I(n2507), .Z(n2506) );
  BUFFD0 U2362 ( .I(n2508), .Z(n2507) );
  BUFFD0 U2363 ( .I(n2509), .Z(n2508) );
  BUFFD0 U2364 ( .I(n2510), .Z(n2509) );
  BUFFD0 U2365 ( .I(n2496), .Z(n2510) );
  BUFFD0 U2366 ( .I(n2513), .Z(n2511) );
  BUFFD0 U2367 ( .I(n227), .Z(n2512) );
  BUFFD0 U2368 ( .I(n2514), .Z(n2513) );
  BUFFD0 U2369 ( .I(n2515), .Z(n2514) );
  BUFFD0 U2370 ( .I(n2516), .Z(n2515) );
  BUFFD0 U2371 ( .I(n2517), .Z(n2516) );
  BUFFD0 U2372 ( .I(n2518), .Z(n2517) );
  BUFFD0 U2373 ( .I(n2519), .Z(n2518) );
  BUFFD0 U2374 ( .I(n2520), .Z(n2519) );
  BUFFD0 U2375 ( .I(n2521), .Z(n2520) );
  BUFFD0 U2376 ( .I(n2522), .Z(n2521) );
  BUFFD0 U2377 ( .I(n2523), .Z(n2522) );
  BUFFD0 U2378 ( .I(n2524), .Z(n2523) );
  BUFFD0 U2379 ( .I(n2525), .Z(n2524) );
  BUFFD0 U2380 ( .I(n2526), .Z(n2525) );
  BUFFD0 U2381 ( .I(n2512), .Z(n2526) );
  BUFFD0 U2382 ( .I(n2529), .Z(n2527) );
  BUFFD0 U2383 ( .I(n226), .Z(n2528) );
  BUFFD0 U2384 ( .I(n2530), .Z(n2529) );
  BUFFD0 U2385 ( .I(n2531), .Z(n2530) );
  BUFFD0 U2386 ( .I(n2532), .Z(n2531) );
  BUFFD0 U2387 ( .I(n2533), .Z(n2532) );
  BUFFD0 U2388 ( .I(n2534), .Z(n2533) );
  BUFFD0 U2389 ( .I(n2535), .Z(n2534) );
  BUFFD0 U2390 ( .I(n2536), .Z(n2535) );
  BUFFD0 U2391 ( .I(n2537), .Z(n2536) );
  BUFFD0 U2392 ( .I(n2538), .Z(n2537) );
  BUFFD0 U2393 ( .I(n2539), .Z(n2538) );
  BUFFD0 U2394 ( .I(n2540), .Z(n2539) );
  BUFFD0 U2395 ( .I(n2541), .Z(n2540) );
  BUFFD0 U2396 ( .I(n2542), .Z(n2541) );
  BUFFD0 U2397 ( .I(n2528), .Z(n2542) );
  BUFFD0 U2398 ( .I(n2545), .Z(n2543) );
  BUFFD0 U2399 ( .I(n225), .Z(n2544) );
  BUFFD0 U2400 ( .I(n2546), .Z(n2545) );
  BUFFD0 U2401 ( .I(n2547), .Z(n2546) );
  BUFFD0 U2402 ( .I(n2548), .Z(n2547) );
  BUFFD0 U2403 ( .I(n2549), .Z(n2548) );
  BUFFD0 U2404 ( .I(n2550), .Z(n2549) );
  BUFFD0 U2405 ( .I(n2551), .Z(n2550) );
  BUFFD0 U2406 ( .I(n2552), .Z(n2551) );
  BUFFD0 U2407 ( .I(n2553), .Z(n2552) );
  BUFFD0 U2408 ( .I(n2554), .Z(n2553) );
  BUFFD0 U2409 ( .I(n2555), .Z(n2554) );
  BUFFD0 U2410 ( .I(n2556), .Z(n2555) );
  BUFFD0 U2411 ( .I(n2557), .Z(n2556) );
  BUFFD0 U2412 ( .I(n2558), .Z(n2557) );
  BUFFD0 U2413 ( .I(n2544), .Z(n2558) );
  BUFFD0 U2414 ( .I(n2561), .Z(n2559) );
  BUFFD0 U2415 ( .I(n224), .Z(n2560) );
  BUFFD0 U2416 ( .I(n2562), .Z(n2561) );
  BUFFD0 U2417 ( .I(n2563), .Z(n2562) );
  BUFFD0 U2418 ( .I(n2564), .Z(n2563) );
  BUFFD0 U2419 ( .I(n2565), .Z(n2564) );
  BUFFD0 U2420 ( .I(n2566), .Z(n2565) );
  BUFFD0 U2421 ( .I(n2567), .Z(n2566) );
  BUFFD0 U2422 ( .I(n2568), .Z(n2567) );
  BUFFD0 U2423 ( .I(n2569), .Z(n2568) );
  BUFFD0 U2424 ( .I(n2570), .Z(n2569) );
  BUFFD0 U2425 ( .I(n2571), .Z(n2570) );
  BUFFD0 U2426 ( .I(n2572), .Z(n2571) );
  BUFFD0 U2427 ( .I(n2573), .Z(n2572) );
  BUFFD0 U2428 ( .I(n2574), .Z(n2573) );
  BUFFD0 U2429 ( .I(n2560), .Z(n2574) );
  BUFFD0 U2430 ( .I(n2577), .Z(n2575) );
  BUFFD0 U2431 ( .I(n223), .Z(n2576) );
  BUFFD0 U2432 ( .I(n2578), .Z(n2577) );
  BUFFD0 U2433 ( .I(n2579), .Z(n2578) );
  BUFFD0 U2434 ( .I(n2580), .Z(n2579) );
  BUFFD0 U2435 ( .I(n2581), .Z(n2580) );
  BUFFD0 U2436 ( .I(n2582), .Z(n2581) );
  BUFFD0 U2437 ( .I(n2583), .Z(n2582) );
  BUFFD0 U2438 ( .I(n2584), .Z(n2583) );
  BUFFD0 U2439 ( .I(n2585), .Z(n2584) );
  BUFFD0 U2440 ( .I(n2586), .Z(n2585) );
  BUFFD0 U2441 ( .I(n2587), .Z(n2586) );
  BUFFD0 U2442 ( .I(n2588), .Z(n2587) );
  BUFFD0 U2443 ( .I(n2589), .Z(n2588) );
  BUFFD0 U2444 ( .I(n2590), .Z(n2589) );
  BUFFD0 U2445 ( .I(n2576), .Z(n2590) );
  BUFFD0 U2446 ( .I(n2593), .Z(n2591) );
  BUFFD0 U2447 ( .I(n222), .Z(n2592) );
  BUFFD0 U2448 ( .I(n2594), .Z(n2593) );
  BUFFD0 U2449 ( .I(n2595), .Z(n2594) );
  BUFFD0 U2450 ( .I(n2596), .Z(n2595) );
  BUFFD0 U2451 ( .I(n2597), .Z(n2596) );
  BUFFD0 U2452 ( .I(n2598), .Z(n2597) );
  BUFFD0 U2453 ( .I(n2599), .Z(n2598) );
  BUFFD0 U2454 ( .I(n2600), .Z(n2599) );
  BUFFD0 U2455 ( .I(n2601), .Z(n2600) );
  BUFFD0 U2456 ( .I(n2602), .Z(n2601) );
  BUFFD0 U2457 ( .I(n2603), .Z(n2602) );
  BUFFD0 U2458 ( .I(n2604), .Z(n2603) );
  BUFFD0 U2459 ( .I(n2605), .Z(n2604) );
  BUFFD0 U2460 ( .I(n2606), .Z(n2605) );
  BUFFD0 U2461 ( .I(n2592), .Z(n2606) );
  BUFFD0 U2462 ( .I(n2609), .Z(n2607) );
  BUFFD0 U2463 ( .I(n221), .Z(n2608) );
  BUFFD0 U2464 ( .I(n2610), .Z(n2609) );
  BUFFD0 U2465 ( .I(n2611), .Z(n2610) );
  BUFFD0 U2466 ( .I(n2612), .Z(n2611) );
  BUFFD0 U2467 ( .I(n2613), .Z(n2612) );
  BUFFD0 U2468 ( .I(n2614), .Z(n2613) );
  BUFFD0 U2469 ( .I(n2615), .Z(n2614) );
  BUFFD0 U2470 ( .I(n2616), .Z(n2615) );
  BUFFD0 U2471 ( .I(n2617), .Z(n2616) );
  BUFFD0 U2472 ( .I(n2618), .Z(n2617) );
  BUFFD0 U2473 ( .I(n2619), .Z(n2618) );
  BUFFD0 U2474 ( .I(n2620), .Z(n2619) );
  BUFFD0 U2475 ( .I(n2621), .Z(n2620) );
  BUFFD0 U2476 ( .I(n2622), .Z(n2621) );
  BUFFD0 U2477 ( .I(n2608), .Z(n2622) );
  BUFFD0 U2478 ( .I(n2625), .Z(n2623) );
  BUFFD0 U2479 ( .I(n220), .Z(n2624) );
  BUFFD0 U2480 ( .I(n2626), .Z(n2625) );
  BUFFD0 U2481 ( .I(n2627), .Z(n2626) );
  BUFFD0 U2482 ( .I(n2628), .Z(n2627) );
  BUFFD0 U2483 ( .I(n2629), .Z(n2628) );
  BUFFD0 U2484 ( .I(n2630), .Z(n2629) );
  BUFFD0 U2485 ( .I(n2631), .Z(n2630) );
  BUFFD0 U2486 ( .I(n2632), .Z(n2631) );
  BUFFD0 U2487 ( .I(n2633), .Z(n2632) );
  BUFFD0 U2488 ( .I(n2634), .Z(n2633) );
  BUFFD0 U2489 ( .I(n2635), .Z(n2634) );
  BUFFD0 U2490 ( .I(n2636), .Z(n2635) );
  BUFFD0 U2491 ( .I(n2637), .Z(n2636) );
  BUFFD0 U2492 ( .I(n2638), .Z(n2637) );
  BUFFD0 U2493 ( .I(n2624), .Z(n2638) );
  BUFFD0 U2494 ( .I(n2641), .Z(n2639) );
  BUFFD0 U2495 ( .I(n219), .Z(n2640) );
  BUFFD0 U2496 ( .I(n2642), .Z(n2641) );
  BUFFD0 U2497 ( .I(n2643), .Z(n2642) );
  BUFFD0 U2498 ( .I(n2644), .Z(n2643) );
  BUFFD0 U2499 ( .I(n2645), .Z(n2644) );
  BUFFD0 U2500 ( .I(n2646), .Z(n2645) );
  BUFFD0 U2501 ( .I(n2647), .Z(n2646) );
  BUFFD0 U2502 ( .I(n2648), .Z(n2647) );
  BUFFD0 U2503 ( .I(n2649), .Z(n2648) );
  BUFFD0 U2504 ( .I(n2650), .Z(n2649) );
  BUFFD0 U2505 ( .I(n2651), .Z(n2650) );
  BUFFD0 U2506 ( .I(n2652), .Z(n2651) );
  BUFFD0 U2507 ( .I(n2653), .Z(n2652) );
  BUFFD0 U2508 ( .I(n2654), .Z(n2653) );
  BUFFD0 U2509 ( .I(n2640), .Z(n2654) );
  BUFFD0 U2510 ( .I(n2657), .Z(n2655) );
  BUFFD0 U2511 ( .I(n218), .Z(n2656) );
  BUFFD0 U2512 ( .I(n2658), .Z(n2657) );
  BUFFD0 U2513 ( .I(n2659), .Z(n2658) );
  BUFFD0 U2514 ( .I(n2660), .Z(n2659) );
  BUFFD0 U2515 ( .I(n2661), .Z(n2660) );
  BUFFD0 U2516 ( .I(n2662), .Z(n2661) );
  BUFFD0 U2517 ( .I(n2663), .Z(n2662) );
  BUFFD0 U2518 ( .I(n2664), .Z(n2663) );
  BUFFD0 U2519 ( .I(n2665), .Z(n2664) );
  BUFFD0 U2520 ( .I(n2666), .Z(n2665) );
  BUFFD0 U2521 ( .I(n2667), .Z(n2666) );
  BUFFD0 U2522 ( .I(n2668), .Z(n2667) );
  BUFFD0 U2523 ( .I(n2669), .Z(n2668) );
  BUFFD0 U2524 ( .I(n2670), .Z(n2669) );
  BUFFD0 U2525 ( .I(n2656), .Z(n2670) );
  BUFFD0 U2526 ( .I(n2673), .Z(n2671) );
  BUFFD0 U2527 ( .I(n217), .Z(n2672) );
  BUFFD0 U2528 ( .I(n2674), .Z(n2673) );
  BUFFD0 U2529 ( .I(n2675), .Z(n2674) );
  BUFFD0 U2530 ( .I(n2676), .Z(n2675) );
  BUFFD0 U2531 ( .I(n2677), .Z(n2676) );
  BUFFD0 U2532 ( .I(n2678), .Z(n2677) );
  BUFFD0 U2533 ( .I(n2679), .Z(n2678) );
  BUFFD0 U2534 ( .I(n2681), .Z(n2680) );
  BUFFD0 U2535 ( .I(n2682), .Z(n2681) );
  BUFFD0 U2536 ( .I(n2683), .Z(n2682) );
  BUFFD0 U2537 ( .I(n2684), .Z(n2683) );
  BUFFD0 U2538 ( .I(n2685), .Z(n2684) );
  BUFFD0 U2539 ( .I(n2686), .Z(n2685) );
  BUFFD0 U2540 ( .I(n2672), .Z(n2686) );
  BUFFD0 U2541 ( .I(n2689), .Z(n2687) );
  BUFFD0 U2542 ( .I(n216), .Z(n2688) );
  BUFFD0 U2543 ( .I(n2690), .Z(n2689) );
  BUFFD0 U2544 ( .I(n2691), .Z(n2690) );
  BUFFD0 U2545 ( .I(n2692), .Z(n2691) );
  BUFFD0 U2546 ( .I(n2693), .Z(n2692) );
  BUFFD0 U2547 ( .I(n2694), .Z(n2693) );
  BUFFD0 U2548 ( .I(n2695), .Z(n2694) );
  BUFFD0 U2549 ( .I(n2696), .Z(n2695) );
  BUFFD0 U2550 ( .I(n2697), .Z(n2696) );
  BUFFD0 U2551 ( .I(n2698), .Z(n2697) );
  BUFFD0 U2552 ( .I(n2699), .Z(n2698) );
  BUFFD0 U2553 ( .I(n2700), .Z(n2699) );
  BUFFD0 U2554 ( .I(n2701), .Z(n2700) );
  BUFFD0 U2555 ( .I(n2702), .Z(n2701) );
  BUFFD0 U2556 ( .I(n2688), .Z(n2702) );
  BUFFD0 U2557 ( .I(n2705), .Z(n2703) );
  BUFFD0 U2558 ( .I(n215), .Z(n2704) );
  BUFFD0 U2559 ( .I(n2706), .Z(n2705) );
  BUFFD0 U2560 ( .I(n2707), .Z(n2706) );
  BUFFD0 U2561 ( .I(n2708), .Z(n2707) );
  BUFFD0 U2562 ( .I(n2709), .Z(n2708) );
  BUFFD0 U2563 ( .I(n2710), .Z(n2709) );
  BUFFD0 U2564 ( .I(n2711), .Z(n2710) );
  BUFFD0 U2565 ( .I(n2712), .Z(n2711) );
  BUFFD0 U2566 ( .I(n2713), .Z(n2712) );
  BUFFD0 U2567 ( .I(n2714), .Z(n2713) );
  BUFFD0 U2568 ( .I(n2715), .Z(n2714) );
  BUFFD0 U2569 ( .I(n2716), .Z(n2715) );
  BUFFD0 U2570 ( .I(n2717), .Z(n2716) );
  BUFFD0 U2571 ( .I(n2718), .Z(n2717) );
  BUFFD0 U2572 ( .I(n2704), .Z(n2718) );
  BUFFD0 U2573 ( .I(n2721), .Z(n2719) );
  BUFFD0 U2574 ( .I(n214), .Z(n2720) );
  BUFFD0 U2575 ( .I(n2722), .Z(n2721) );
  BUFFD0 U2576 ( .I(n2723), .Z(n2722) );
  BUFFD0 U2577 ( .I(n2724), .Z(n2723) );
  BUFFD0 U2578 ( .I(n2725), .Z(n2724) );
  BUFFD0 U2579 ( .I(n2726), .Z(n2725) );
  BUFFD0 U2580 ( .I(n2727), .Z(n2726) );
  BUFFD0 U2581 ( .I(n2728), .Z(n2727) );
  BUFFD0 U2582 ( .I(n2729), .Z(n2728) );
  BUFFD0 U2583 ( .I(n2730), .Z(n2729) );
  BUFFD0 U2584 ( .I(n2731), .Z(n2730) );
  BUFFD0 U2585 ( .I(n2732), .Z(n2731) );
  BUFFD0 U2586 ( .I(n2733), .Z(n2732) );
  BUFFD0 U2587 ( .I(n2734), .Z(n2733) );
  BUFFD0 U2588 ( .I(n2720), .Z(n2734) );
  BUFFD0 U2589 ( .I(n2737), .Z(n2735) );
  BUFFD0 U2590 ( .I(n213), .Z(n2736) );
  BUFFD0 U2591 ( .I(n2738), .Z(n2737) );
  BUFFD0 U2592 ( .I(n2739), .Z(n2738) );
  BUFFD0 U2593 ( .I(n2740), .Z(n2739) );
  BUFFD0 U2594 ( .I(n2741), .Z(n2740) );
  BUFFD0 U2595 ( .I(n2742), .Z(n2741) );
  BUFFD0 U2596 ( .I(n2743), .Z(n2742) );
  BUFFD0 U2597 ( .I(n2744), .Z(n2743) );
  BUFFD0 U2598 ( .I(n2745), .Z(n2744) );
  BUFFD0 U2599 ( .I(n2746), .Z(n2745) );
  BUFFD0 U2600 ( .I(n2747), .Z(n2746) );
  BUFFD0 U2601 ( .I(n2748), .Z(n2747) );
  BUFFD0 U2602 ( .I(n2749), .Z(n2748) );
  BUFFD0 U2603 ( .I(n2750), .Z(n2749) );
  BUFFD0 U2604 ( .I(n2736), .Z(n2750) );
  BUFFD0 U2605 ( .I(n2753), .Z(n2751) );
  BUFFD0 U2606 ( .I(n212), .Z(n2752) );
  BUFFD0 U2607 ( .I(n2754), .Z(n2753) );
  BUFFD0 U2608 ( .I(n2755), .Z(n2754) );
  BUFFD0 U2609 ( .I(n2756), .Z(n2755) );
  BUFFD0 U2610 ( .I(n2757), .Z(n2756) );
  BUFFD0 U2611 ( .I(n2758), .Z(n2757) );
  BUFFD0 U2612 ( .I(n2759), .Z(n2758) );
  BUFFD0 U2613 ( .I(n2760), .Z(n2759) );
  BUFFD0 U2614 ( .I(n2761), .Z(n2760) );
  BUFFD0 U2615 ( .I(n2762), .Z(n2761) );
  BUFFD0 U2616 ( .I(n2763), .Z(n2762) );
  BUFFD0 U2617 ( .I(n2764), .Z(n2763) );
  BUFFD0 U2618 ( .I(n2765), .Z(n2764) );
  BUFFD0 U2619 ( .I(n2766), .Z(n2765) );
  BUFFD0 U2620 ( .I(n2752), .Z(n2766) );
  BUFFD0 U2621 ( .I(n2769), .Z(n2767) );
  BUFFD0 U2622 ( .I(n211), .Z(n2768) );
  BUFFD0 U2623 ( .I(n2770), .Z(n2769) );
  BUFFD0 U2624 ( .I(n2771), .Z(n2770) );
  BUFFD0 U2625 ( .I(n2772), .Z(n2771) );
  BUFFD0 U2626 ( .I(n2773), .Z(n2772) );
  BUFFD0 U2627 ( .I(n2774), .Z(n2773) );
  BUFFD0 U2628 ( .I(n2775), .Z(n2774) );
  BUFFD0 U2629 ( .I(n2776), .Z(n2775) );
  BUFFD0 U2630 ( .I(n2777), .Z(n2776) );
  BUFFD0 U2631 ( .I(n2778), .Z(n2777) );
  BUFFD0 U2632 ( .I(n2779), .Z(n2778) );
  BUFFD0 U2633 ( .I(n2780), .Z(n2779) );
  BUFFD0 U2634 ( .I(n2781), .Z(n2780) );
  BUFFD0 U2635 ( .I(n2782), .Z(n2781) );
  BUFFD0 U2636 ( .I(n2768), .Z(n2782) );
  BUFFD0 U2637 ( .I(n2785), .Z(n2783) );
  BUFFD0 U2638 ( .I(n210), .Z(n2784) );
  BUFFD0 U2639 ( .I(n2786), .Z(n2785) );
  BUFFD0 U2640 ( .I(n2787), .Z(n2786) );
  BUFFD0 U2641 ( .I(n2788), .Z(n2787) );
  BUFFD0 U2642 ( .I(n2789), .Z(n2788) );
  BUFFD0 U2643 ( .I(n2790), .Z(n2789) );
  BUFFD0 U2644 ( .I(n2791), .Z(n2790) );
  BUFFD0 U2645 ( .I(n2792), .Z(n2791) );
  BUFFD0 U2646 ( .I(n2793), .Z(n2792) );
  BUFFD0 U2647 ( .I(n2794), .Z(n2793) );
  BUFFD0 U2648 ( .I(n2795), .Z(n2794) );
  BUFFD0 U2649 ( .I(n2796), .Z(n2795) );
  BUFFD0 U2650 ( .I(n2797), .Z(n2796) );
  BUFFD0 U2651 ( .I(n2798), .Z(n2797) );
  BUFFD0 U2652 ( .I(n2784), .Z(n2798) );
  BUFFD0 U2653 ( .I(n2801), .Z(n2799) );
  BUFFD0 U2654 ( .I(n209), .Z(n2800) );
  BUFFD0 U2655 ( .I(n2802), .Z(n2801) );
  BUFFD0 U2656 ( .I(n2803), .Z(n2802) );
  BUFFD0 U2657 ( .I(n2804), .Z(n2803) );
  BUFFD0 U2658 ( .I(n2805), .Z(n2804) );
  BUFFD0 U2659 ( .I(n2806), .Z(n2805) );
  BUFFD0 U2660 ( .I(n2807), .Z(n2806) );
  BUFFD0 U2661 ( .I(n2808), .Z(n2807) );
  BUFFD0 U2662 ( .I(n2809), .Z(n2808) );
  BUFFD0 U2663 ( .I(n2810), .Z(n2809) );
  BUFFD0 U2664 ( .I(n2811), .Z(n2810) );
  BUFFD0 U2665 ( .I(n2812), .Z(n2811) );
  BUFFD0 U2666 ( .I(n2813), .Z(n2812) );
  BUFFD0 U2667 ( .I(n2814), .Z(n2813) );
  BUFFD0 U2668 ( .I(n2800), .Z(n2814) );
  BUFFD0 U2669 ( .I(n2817), .Z(n2815) );
  BUFFD0 U2670 ( .I(n208), .Z(n2816) );
  BUFFD0 U2671 ( .I(n2818), .Z(n2817) );
  BUFFD0 U2672 ( .I(n2819), .Z(n2818) );
  BUFFD0 U2673 ( .I(n2820), .Z(n2819) );
  BUFFD0 U2674 ( .I(n2821), .Z(n2820) );
  BUFFD0 U2675 ( .I(n2822), .Z(n2821) );
  BUFFD0 U2676 ( .I(n2823), .Z(n2822) );
  BUFFD0 U2677 ( .I(n2824), .Z(n2823) );
  BUFFD0 U2678 ( .I(n2825), .Z(n2824) );
  BUFFD0 U2679 ( .I(n2826), .Z(n2825) );
  BUFFD0 U2680 ( .I(n2827), .Z(n2826) );
  BUFFD0 U2681 ( .I(n2828), .Z(n2827) );
  BUFFD0 U2682 ( .I(n2829), .Z(n2828) );
  BUFFD0 U2683 ( .I(n2830), .Z(n2829) );
  BUFFD0 U2684 ( .I(n2816), .Z(n2830) );
  BUFFD0 U2685 ( .I(n2833), .Z(n2831) );
  BUFFD0 U2686 ( .I(n207), .Z(n2832) );
  BUFFD0 U2687 ( .I(n2834), .Z(n2833) );
  BUFFD0 U2688 ( .I(n2835), .Z(n2834) );
  BUFFD0 U2689 ( .I(n2836), .Z(n2835) );
  BUFFD0 U2690 ( .I(n2837), .Z(n2836) );
  BUFFD0 U2691 ( .I(n2838), .Z(n2837) );
  BUFFD0 U2692 ( .I(n2839), .Z(n2838) );
  BUFFD0 U2693 ( .I(n2840), .Z(n2839) );
  BUFFD0 U2694 ( .I(n2841), .Z(n2840) );
  BUFFD0 U2695 ( .I(n2842), .Z(n2841) );
  BUFFD0 U2696 ( .I(n2843), .Z(n2842) );
  BUFFD0 U2697 ( .I(n2844), .Z(n2843) );
  BUFFD0 U2698 ( .I(n2845), .Z(n2844) );
  BUFFD0 U2699 ( .I(n2846), .Z(n2845) );
  BUFFD0 U2700 ( .I(n2832), .Z(n2846) );
  BUFFD0 U2701 ( .I(n2849), .Z(n2847) );
  BUFFD0 U2702 ( .I(n206), .Z(n2848) );
  BUFFD0 U2703 ( .I(n2850), .Z(n2849) );
  BUFFD0 U2704 ( .I(n2851), .Z(n2850) );
  BUFFD0 U2705 ( .I(n2852), .Z(n2851) );
  BUFFD0 U2706 ( .I(n2853), .Z(n2852) );
  BUFFD0 U2707 ( .I(n2854), .Z(n2853) );
  BUFFD0 U2708 ( .I(n2855), .Z(n2854) );
  BUFFD0 U2709 ( .I(n2856), .Z(n2855) );
  BUFFD0 U2710 ( .I(n2857), .Z(n2856) );
  BUFFD0 U2711 ( .I(n2858), .Z(n2857) );
  BUFFD0 U2712 ( .I(n2859), .Z(n2858) );
  BUFFD0 U2713 ( .I(n2860), .Z(n2859) );
  BUFFD0 U2714 ( .I(n2861), .Z(n2860) );
  BUFFD0 U2715 ( .I(n2862), .Z(n2861) );
  BUFFD0 U2716 ( .I(n2848), .Z(n2862) );
  BUFFD0 U2717 ( .I(n2865), .Z(n2863) );
  BUFFD0 U2718 ( .I(n205), .Z(n2864) );
  BUFFD0 U2719 ( .I(n2866), .Z(n2865) );
  BUFFD0 U2720 ( .I(n2867), .Z(n2866) );
  BUFFD0 U2721 ( .I(n2868), .Z(n2867) );
  BUFFD0 U2722 ( .I(n2869), .Z(n2868) );
  BUFFD0 U2723 ( .I(n2870), .Z(n2869) );
  BUFFD0 U2724 ( .I(n2871), .Z(n2870) );
  BUFFD0 U2725 ( .I(n2872), .Z(n2871) );
  BUFFD0 U2726 ( .I(n2873), .Z(n2872) );
  BUFFD0 U2727 ( .I(n2874), .Z(n2873) );
  BUFFD0 U2728 ( .I(n2875), .Z(n2874) );
  BUFFD0 U2729 ( .I(n2876), .Z(n2875) );
  BUFFD0 U2730 ( .I(n2877), .Z(n2876) );
  BUFFD0 U2731 ( .I(n2878), .Z(n2877) );
  BUFFD0 U2732 ( .I(n2864), .Z(n2878) );
  BUFFD0 U2733 ( .I(n2881), .Z(n2879) );
  BUFFD0 U2734 ( .I(n204), .Z(n2880) );
  BUFFD0 U2735 ( .I(n2882), .Z(n2881) );
  BUFFD0 U2736 ( .I(n2883), .Z(n2882) );
  BUFFD0 U2737 ( .I(n2884), .Z(n2883) );
  BUFFD0 U2738 ( .I(n2885), .Z(n2884) );
  BUFFD0 U2739 ( .I(n2886), .Z(n2885) );
  BUFFD0 U2740 ( .I(n2887), .Z(n2886) );
  BUFFD0 U2741 ( .I(n2888), .Z(n2887) );
  BUFFD0 U2742 ( .I(n2889), .Z(n2888) );
  BUFFD0 U2743 ( .I(n2890), .Z(n2889) );
  BUFFD0 U2744 ( .I(n2891), .Z(n2890) );
  BUFFD0 U2745 ( .I(n2892), .Z(n2891) );
  BUFFD0 U2746 ( .I(n2893), .Z(n2892) );
  BUFFD0 U2747 ( .I(n2894), .Z(n2893) );
  BUFFD0 U2748 ( .I(n2880), .Z(n2894) );
  BUFFD0 U2749 ( .I(n2897), .Z(n2895) );
  BUFFD0 U2750 ( .I(n203), .Z(n2896) );
  BUFFD0 U2751 ( .I(n2898), .Z(n2897) );
  BUFFD0 U2752 ( .I(n2899), .Z(n2898) );
  BUFFD0 U2753 ( .I(n2900), .Z(n2899) );
  BUFFD0 U2754 ( .I(n2901), .Z(n2900) );
  BUFFD0 U2755 ( .I(n2902), .Z(n2901) );
  BUFFD0 U2756 ( .I(n2903), .Z(n2902) );
  BUFFD0 U2757 ( .I(n2904), .Z(n2903) );
  BUFFD0 U2758 ( .I(n2905), .Z(n2904) );
  BUFFD0 U2759 ( .I(n2906), .Z(n2905) );
  BUFFD0 U2760 ( .I(n2907), .Z(n2906) );
  BUFFD0 U2761 ( .I(n2908), .Z(n2907) );
  BUFFD0 U2762 ( .I(n2909), .Z(n2908) );
  BUFFD0 U2763 ( .I(n2910), .Z(n2909) );
  BUFFD0 U2764 ( .I(n2896), .Z(n2910) );
  BUFFD0 U2765 ( .I(n2913), .Z(n2911) );
  BUFFD0 U2766 ( .I(n202), .Z(n2912) );
  BUFFD0 U2767 ( .I(n2914), .Z(n2913) );
  BUFFD0 U2768 ( .I(n2915), .Z(n2914) );
  BUFFD0 U2769 ( .I(n2916), .Z(n2915) );
  BUFFD0 U2770 ( .I(n2917), .Z(n2916) );
  BUFFD0 U2771 ( .I(n2918), .Z(n2917) );
  BUFFD0 U2772 ( .I(n2919), .Z(n2918) );
  BUFFD0 U2773 ( .I(n2920), .Z(n2919) );
  BUFFD0 U2774 ( .I(n2921), .Z(n2920) );
  BUFFD0 U2775 ( .I(n2922), .Z(n2921) );
  BUFFD0 U2776 ( .I(n2923), .Z(n2922) );
  BUFFD0 U2777 ( .I(n2924), .Z(n2923) );
  BUFFD0 U2778 ( .I(n2925), .Z(n2924) );
  BUFFD0 U2779 ( .I(n2926), .Z(n2925) );
  BUFFD0 U2780 ( .I(n2912), .Z(n2926) );
  BUFFD0 U2781 ( .I(n2929), .Z(n2927) );
  BUFFD0 U2782 ( .I(n201), .Z(n2928) );
  BUFFD0 U2783 ( .I(n2930), .Z(n2929) );
  BUFFD0 U2784 ( .I(n2931), .Z(n2930) );
  BUFFD0 U2785 ( .I(n2932), .Z(n2931) );
  BUFFD0 U2786 ( .I(n2933), .Z(n2932) );
  BUFFD0 U2787 ( .I(n2934), .Z(n2933) );
  BUFFD0 U2788 ( .I(n2935), .Z(n2934) );
  BUFFD0 U2789 ( .I(n2936), .Z(n2935) );
  BUFFD0 U2790 ( .I(n2937), .Z(n2936) );
  BUFFD0 U2791 ( .I(n2938), .Z(n2937) );
  BUFFD0 U2792 ( .I(n2939), .Z(n2938) );
  BUFFD0 U2793 ( .I(n2940), .Z(n2939) );
  BUFFD0 U2794 ( .I(n2941), .Z(n2940) );
  BUFFD0 U2795 ( .I(n2942), .Z(n2941) );
  BUFFD0 U2796 ( .I(n2928), .Z(n2942) );
  BUFFD0 U2797 ( .I(n2945), .Z(n2943) );
  BUFFD0 U2798 ( .I(n200), .Z(n2944) );
  BUFFD0 U2799 ( .I(n2946), .Z(n2945) );
  BUFFD0 U2800 ( .I(n2947), .Z(n2946) );
  BUFFD0 U2801 ( .I(n2948), .Z(n2947) );
  BUFFD0 U2802 ( .I(n2949), .Z(n2948) );
  BUFFD0 U2803 ( .I(n2950), .Z(n2949) );
  BUFFD0 U2804 ( .I(n2951), .Z(n2950) );
  BUFFD0 U2805 ( .I(n2952), .Z(n2951) );
  BUFFD0 U2806 ( .I(n2953), .Z(n2952) );
  BUFFD0 U2807 ( .I(n2954), .Z(n2953) );
  BUFFD0 U2808 ( .I(n2955), .Z(n2954) );
  BUFFD0 U2809 ( .I(n2956), .Z(n2955) );
  BUFFD0 U2810 ( .I(n2957), .Z(n2956) );
  BUFFD0 U2811 ( .I(n2958), .Z(n2957) );
  BUFFD0 U2812 ( .I(n2944), .Z(n2958) );
  BUFFD0 U2813 ( .I(n2961), .Z(n2959) );
  BUFFD0 U2814 ( .I(n199), .Z(n2960) );
  BUFFD0 U2815 ( .I(n2962), .Z(n2961) );
  BUFFD0 U2816 ( .I(n2963), .Z(n2962) );
  BUFFD0 U2817 ( .I(n2964), .Z(n2963) );
  BUFFD0 U2818 ( .I(n2965), .Z(n2964) );
  BUFFD0 U2819 ( .I(n2966), .Z(n2965) );
  BUFFD0 U2820 ( .I(n2967), .Z(n2966) );
  BUFFD0 U2821 ( .I(n2968), .Z(n2967) );
  BUFFD0 U2822 ( .I(n2969), .Z(n2968) );
  BUFFD0 U2823 ( .I(n2970), .Z(n2969) );
  BUFFD0 U2824 ( .I(n2971), .Z(n2970) );
  BUFFD0 U2825 ( .I(n2972), .Z(n2971) );
  BUFFD0 U2826 ( .I(n2973), .Z(n2972) );
  BUFFD0 U2827 ( .I(n2974), .Z(n2973) );
  BUFFD0 U2828 ( .I(n2960), .Z(n2974) );
  BUFFD0 U2829 ( .I(n2977), .Z(n2975) );
  BUFFD0 U2830 ( .I(n198), .Z(n2976) );
  BUFFD0 U2831 ( .I(n2978), .Z(n2977) );
  BUFFD0 U2832 ( .I(n2979), .Z(n2978) );
  BUFFD0 U2833 ( .I(n2980), .Z(n2979) );
  BUFFD0 U2834 ( .I(n2981), .Z(n2980) );
  BUFFD0 U2835 ( .I(n2982), .Z(n2981) );
  BUFFD0 U2836 ( .I(n2983), .Z(n2982) );
  BUFFD0 U2837 ( .I(n2984), .Z(n2983) );
  BUFFD0 U2838 ( .I(n2985), .Z(n2984) );
  BUFFD0 U2839 ( .I(n2986), .Z(n2985) );
  BUFFD0 U2840 ( .I(n2987), .Z(n2986) );
  BUFFD0 U2841 ( .I(n2988), .Z(n2987) );
  BUFFD0 U2842 ( .I(n2989), .Z(n2988) );
  BUFFD0 U2843 ( .I(n2990), .Z(n2989) );
  BUFFD0 U2844 ( .I(n2976), .Z(n2990) );
  BUFFD0 U2845 ( .I(n2993), .Z(n2991) );
  BUFFD0 U2846 ( .I(n197), .Z(n2992) );
  BUFFD0 U2847 ( .I(n2994), .Z(n2993) );
  BUFFD0 U2848 ( .I(n2995), .Z(n2994) );
  BUFFD0 U2849 ( .I(n2996), .Z(n2995) );
  BUFFD0 U2850 ( .I(n2997), .Z(n2996) );
  BUFFD0 U2851 ( .I(n2998), .Z(n2997) );
  BUFFD0 U2852 ( .I(n2999), .Z(n2998) );
  BUFFD0 U2853 ( .I(n3000), .Z(n2999) );
  BUFFD0 U2854 ( .I(n3001), .Z(n3000) );
  BUFFD0 U2855 ( .I(n3002), .Z(n3001) );
  BUFFD0 U2856 ( .I(n3003), .Z(n3002) );
  BUFFD0 U2857 ( .I(n3004), .Z(n3003) );
  BUFFD0 U2858 ( .I(n3005), .Z(n3004) );
  BUFFD0 U2859 ( .I(n3006), .Z(n3005) );
  CKBD0 U2860 ( .CLK(n3130), .C(n3007) );
  CKNXD16 U2861 ( .I(n3007), .ZN(ParOut[31]) );
  CKBD0 U2862 ( .CLK(n3129), .C(n3009) );
  CKNXD16 U2863 ( .I(n3009), .ZN(ParOut[30]) );
  CKBD0 U2864 ( .CLK(n3128), .C(n3011) );
  CKNXD16 U2865 ( .I(n3011), .ZN(ParOut[29]) );
  CKBD0 U2866 ( .CLK(n3127), .C(n3013) );
  CKNXD16 U2867 ( .I(n3013), .ZN(ParOut[28]) );
  CKBD0 U2868 ( .CLK(n3126), .C(n3015) );
  CKNXD16 U2869 ( .I(n3015), .ZN(ParOut[27]) );
  CKBD0 U2870 ( .CLK(n3125), .C(n3017) );
  CKNXD16 U2871 ( .I(n3017), .ZN(ParOut[26]) );
  CKBD0 U2872 ( .CLK(n3124), .C(n3019) );
  CKNXD16 U2873 ( .I(n3019), .ZN(ParOut[25]) );
  CKBD0 U2874 ( .CLK(n3123), .C(n3021) );
  CKNXD16 U2875 ( .I(n3021), .ZN(ParOut[24]) );
  CKBD0 U2876 ( .CLK(n3122), .C(n3023) );
  CKNXD16 U2877 ( .I(n3023), .ZN(ParOut[23]) );
  CKBD0 U2878 ( .CLK(n3121), .C(n3025) );
  CKNXD16 U2879 ( .I(n3025), .ZN(ParOut[22]) );
  CKBD0 U2880 ( .CLK(n3120), .C(n3027) );
  CKNXD16 U2881 ( .I(n3027), .ZN(ParOut[21]) );
  CKBD0 U2882 ( .CLK(n3119), .C(n3029) );
  CKNXD16 U2883 ( .I(n3029), .ZN(ParOut[20]) );
  CKBD0 U2884 ( .CLK(n3118), .C(n3031) );
  CKNXD16 U2885 ( .I(n3031), .ZN(ParOut[19]) );
  CKBD0 U2886 ( .CLK(n3117), .C(n3033) );
  CKNXD16 U2887 ( .I(n3033), .ZN(ParOut[18]) );
  CKBD0 U2888 ( .CLK(n3116), .C(n3035) );
  CKNXD16 U2889 ( .I(n3035), .ZN(ParOut[17]) );
  CKBD0 U2890 ( .CLK(n3115), .C(n3037) );
  CKNXD16 U2891 ( .I(n3037), .ZN(ParOut[16]) );
  CKBD0 U2892 ( .CLK(n3114), .C(n3039) );
  CKNXD16 U2893 ( .I(n3039), .ZN(ParOut[15]) );
  CKBD0 U2894 ( .CLK(n3113), .C(n3041) );
  CKNXD16 U2895 ( .I(n3041), .ZN(ParOut[14]) );
  CKBD0 U2896 ( .CLK(n3112), .C(n3043) );
  CKNXD16 U2897 ( .I(n3043), .ZN(ParOut[13]) );
  CKBD0 U2898 ( .CLK(n3111), .C(n3045) );
  CKNXD16 U2899 ( .I(n3045), .ZN(ParOut[12]) );
  CKBD0 U2900 ( .CLK(n3110), .C(n3047) );
  CKNXD16 U2901 ( .I(n3047), .ZN(ParOut[11]) );
  CKBD0 U2902 ( .CLK(n3109), .C(n3049) );
  CKNXD16 U2903 ( .I(n3049), .ZN(ParOut[10]) );
  CKBD0 U2904 ( .CLK(n3108), .C(n3051) );
  CKNXD16 U2905 ( .I(n3051), .ZN(ParOut[9]) );
  CKBD0 U2906 ( .CLK(n3107), .C(n3053) );
  CKNXD16 U2907 ( .I(n3053), .ZN(ParOut[8]) );
  CKBD0 U2908 ( .CLK(n3106), .C(n3055) );
  CKNXD16 U2909 ( .I(n3055), .ZN(ParOut[7]) );
  CKBD0 U2910 ( .CLK(n3105), .C(n3057) );
  CKNXD16 U2911 ( .I(n3057), .ZN(ParOut[6]) );
  CKBD0 U2912 ( .CLK(n3104), .C(n3059) );
  CKNXD16 U2913 ( .I(n3059), .ZN(ParOut[5]) );
  CKBD0 U2914 ( .CLK(n3103), .C(n3061) );
  CKNXD16 U2915 ( .I(n3061), .ZN(ParOut[4]) );
  CKBD0 U2916 ( .CLK(n3102), .C(n3063) );
  CKNXD16 U2917 ( .I(n3063), .ZN(ParOut[3]) );
  CKBD0 U2918 ( .CLK(n3101), .C(n3065) );
  CKNXD16 U2919 ( .I(n3065), .ZN(ParOut[2]) );
  CKBD0 U2920 ( .CLK(n3100), .C(n3067) );
  CKNXD16 U2921 ( .I(n3067), .ZN(ParOut[1]) );
  CKBD0 U2922 ( .CLK(n3099), .C(n3069) );
  CKNXD16 U2923 ( .I(n3069), .ZN(ParOut[0]) );
  CKBD0 U2924 ( .CLK(n3131), .C(n3071) );
  CKNXD16 U2925 ( .I(n3071), .ZN(ParClk) );
  INVD1 U2926 ( .I(n2463), .ZN(n3141) );
  BUFFD1 U2927 ( .I(n3139), .Z(n3137) );
  BUFFD1 U2928 ( .I(n3140), .Z(n3136) );
  BUFFD1 U2929 ( .I(n3140), .Z(n3135) );
  BUFFD1 U2930 ( .I(n3140), .Z(n3134) );
  BUFFD1 U2931 ( .I(n3140), .Z(n3138) );
  BUFFD1 U2932 ( .I(n3143), .Z(n3144) );
  BUFFD1 U2933 ( .I(SerClock), .Z(n3145) );
  BUFFD1 U2934 ( .I(n3142), .Z(n3146) );
  BUFFD1 U2935 ( .I(n3142), .Z(n3147) );
  BUFFD1 U2936 ( .I(n3142), .Z(n3148) );
  BUFFD1 U2937 ( .I(SerClock), .Z(n3142) );
  BUFFD1 U2938 ( .I(n261), .Z(n3139) );
  BUFFD1 U2939 ( .I(n261), .Z(n3140) );
  BUFFD1 U2940 ( .I(SerClock), .Z(n3143) );
  NR2D1 U2941 ( .A1(n3149), .A2(n264), .ZN(n3) );
  NR4D0 U2942 ( .A1(n60), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n58) );
  AN2D1 U2943 ( .A1(N33), .A2(n2), .Z(N41) );
  AN2D1 U2944 ( .A1(N32), .A2(n2), .Z(N40) );
  AN2D1 U2945 ( .A1(N30), .A2(n2), .Z(N38) );
  NR4D0 U2946 ( .A1(n57), .A2(n139), .A3(n155), .A4(n140), .ZN(n50) );
  ND3D1 U2947 ( .A1(n175), .A2(n174), .A3(n2068), .ZN(n57) );
  OAI22D0 U2948 ( .A1(n2463), .A2(n1681), .B1(n2464), .B2(n44), .ZN(n229) );
  OAI22D0 U2949 ( .A1(n2463), .A2(n182), .B1(n3141), .B2(n43), .ZN(n230) );
  OAI22D0 U2950 ( .A1(n2463), .A2(n181), .B1(n3141), .B2(n42), .ZN(n231) );
  OAI22D0 U2951 ( .A1(n2463), .A2(n180), .B1(n2464), .B2(n41), .ZN(n232) );
  OAI22D0 U2952 ( .A1(n2463), .A2(n179), .B1(n2464), .B2(n40), .ZN(n233) );
  OAI22D0 U2953 ( .A1(n2463), .A2(n178), .B1(n2464), .B2(n39), .ZN(n234) );
  OAI22D0 U2954 ( .A1(n45), .A2(n177), .B1(n2464), .B2(n38), .ZN(n235) );
  OAI22D0 U2955 ( .A1(n45), .A2(n176), .B1(n2464), .B2(n37), .ZN(n236) );
  OAI22D0 U2956 ( .A1(n45), .A2(n167), .B1(n2464), .B2(n36), .ZN(n237) );
  OAI22D0 U2957 ( .A1(n45), .A2(n166), .B1(n2464), .B2(n35), .ZN(n238) );
  OAI22D0 U2958 ( .A1(n45), .A2(n165), .B1(n2464), .B2(n34), .ZN(n239) );
  OAI22D0 U2959 ( .A1(n45), .A2(n164), .B1(n3141), .B2(n33), .ZN(n240) );
  OAI22D0 U2960 ( .A1(n45), .A2(n163), .B1(n3141), .B2(n32), .ZN(n241) );
  OAI22D0 U2961 ( .A1(n45), .A2(n162), .B1(n3141), .B2(n31), .ZN(n242) );
  OAI22D0 U2962 ( .A1(n45), .A2(n161), .B1(n3141), .B2(n30), .ZN(n243) );
  OAI22D0 U2963 ( .A1(n2463), .A2(n160), .B1(n3141), .B2(n29), .ZN(n244) );
  OAI22D0 U2964 ( .A1(n2463), .A2(n151), .B1(n3141), .B2(n28), .ZN(n245) );
  OAI22D0 U2965 ( .A1(n2463), .A2(n150), .B1(n3141), .B2(n27), .ZN(n246) );
  OAI22D0 U2966 ( .A1(n45), .A2(n149), .B1(n3141), .B2(n26), .ZN(n247) );
  OAI22D0 U2967 ( .A1(n45), .A2(n148), .B1(n3141), .B2(n25), .ZN(n248) );
  OAI22D0 U2968 ( .A1(n2463), .A2(n147), .B1(n3141), .B2(n24), .ZN(n249) );
  OAI22D0 U2969 ( .A1(n45), .A2(n146), .B1(n3141), .B2(n23), .ZN(n250) );
  OAI22D0 U2970 ( .A1(n2463), .A2(n145), .B1(n3141), .B2(n22), .ZN(n251) );
  OAI22D0 U2971 ( .A1(n45), .A2(n144), .B1(n3141), .B2(n21), .ZN(n252) );
  OAI22D0 U2972 ( .A1(n45), .A2(n135), .B1(n2464), .B2(n20), .ZN(n253) );
  OAI22D0 U2973 ( .A1(n45), .A2(n134), .B1(n2464), .B2(n19), .ZN(n254) );
  OAI22D0 U2974 ( .A1(n2463), .A2(n133), .B1(n2464), .B2(n18), .ZN(n255) );
  OAI22D0 U2975 ( .A1(n45), .A2(n132), .B1(n2464), .B2(n17), .ZN(n256) );
  OAI22D0 U2976 ( .A1(n2463), .A2(n131), .B1(n3141), .B2(n16), .ZN(n257) );
  OAI22D0 U2977 ( .A1(n45), .A2(n130), .B1(n3141), .B2(n15), .ZN(n258) );
  OAI22D0 U2978 ( .A1(n45), .A2(n129), .B1(n3141), .B2(n14), .ZN(n259) );
  OAI22D0 U2979 ( .A1(n45), .A2(n128), .B1(n3141), .B2(n13), .ZN(n260) );
  OAI22D0 U2980 ( .A1(n3132), .A2(n3099), .B1(n263), .B2(n44), .ZN(n228) );
  OAI22D0 U2981 ( .A1(n299), .A2(n3100), .B1(n263), .B2(n43), .ZN(n227) );
  OAI22D0 U2982 ( .A1(n299), .A2(n3101), .B1(n3133), .B2(n42), .ZN(n226) );
  OAI22D0 U2983 ( .A1(n299), .A2(n3102), .B1(n3133), .B2(n41), .ZN(n225) );
  OAI22D0 U2984 ( .A1(n299), .A2(n3103), .B1(n3133), .B2(n40), .ZN(n224) );
  OAI22D0 U2985 ( .A1(n299), .A2(n3104), .B1(n263), .B2(n39), .ZN(n223) );
  OAI22D0 U2986 ( .A1(n299), .A2(n3105), .B1(n3133), .B2(n38), .ZN(n222) );
  OAI22D0 U2987 ( .A1(n299), .A2(n3106), .B1(n263), .B2(n37), .ZN(n221) );
  OAI22D0 U2988 ( .A1(n299), .A2(n3107), .B1(n263), .B2(n36), .ZN(n220) );
  OAI22D0 U2989 ( .A1(n299), .A2(n3108), .B1(n263), .B2(n35), .ZN(n219) );
  OAI22D0 U2990 ( .A1(n3132), .A2(n3109), .B1(n263), .B2(n34), .ZN(n218) );
  OAI22D0 U2991 ( .A1(n3132), .A2(n3110), .B1(n3133), .B2(n33), .ZN(n217) );
  OAI22D0 U2992 ( .A1(n3132), .A2(n3111), .B1(n263), .B2(n32), .ZN(n216) );
  OAI22D0 U2993 ( .A1(n3132), .A2(n3112), .B1(n263), .B2(n31), .ZN(n215) );
  OAI22D0 U2994 ( .A1(n3132), .A2(n3113), .B1(n263), .B2(n30), .ZN(n214) );
  OAI22D0 U2995 ( .A1(n3132), .A2(n3114), .B1(n3133), .B2(n29), .ZN(n213) );
  OAI22D0 U2996 ( .A1(n3132), .A2(n3115), .B1(n3133), .B2(n28), .ZN(n212) );
  OAI22D0 U2997 ( .A1(n299), .A2(n3116), .B1(n3133), .B2(n27), .ZN(n211) );
  OAI22D0 U2998 ( .A1(n299), .A2(n3117), .B1(n3133), .B2(n26), .ZN(n210) );
  OAI22D0 U2999 ( .A1(n299), .A2(n3118), .B1(n3133), .B2(n25), .ZN(n209) );
  OAI22D0 U3000 ( .A1(n299), .A2(n3119), .B1(n3133), .B2(n24), .ZN(n208) );
  OAI22D0 U3001 ( .A1(n299), .A2(n3120), .B1(n263), .B2(n23), .ZN(n207) );
  OAI22D0 U3002 ( .A1(n299), .A2(n3121), .B1(n263), .B2(n22), .ZN(n206) );
  OAI22D0 U3003 ( .A1(n299), .A2(n3122), .B1(n263), .B2(n21), .ZN(n205) );
  OAI22D0 U3004 ( .A1(n299), .A2(n3123), .B1(n263), .B2(n20), .ZN(n204) );
  OAI22D0 U3005 ( .A1(n299), .A2(n3124), .B1(n263), .B2(n19), .ZN(n203) );
  OAI22D0 U3006 ( .A1(n299), .A2(n3125), .B1(n263), .B2(n18), .ZN(n202) );
  OAI22D0 U3007 ( .A1(n299), .A2(n3126), .B1(n3133), .B2(n17), .ZN(n201) );
  OAI22D0 U3008 ( .A1(n3132), .A2(n3127), .B1(n263), .B2(n16), .ZN(n200) );
  OAI22D0 U3009 ( .A1(n3132), .A2(n3128), .B1(n263), .B2(n15), .ZN(n199) );
  OAI22D0 U3010 ( .A1(n3132), .A2(n3129), .B1(n263), .B2(n14), .ZN(n198) );
  OAI22D0 U3011 ( .A1(n3132), .A2(n3130), .B1(n3133), .B2(n13), .ZN(n197) );
  ND2D1 U3012 ( .A1(n48), .A2(n49), .ZN(n46) );
  NR4D0 U3013 ( .A1(n2051), .A2(n2230), .A3(n2122), .A4(n2212), .ZN(n48) );
  NR4D0 U3014 ( .A1(n2462), .A2(n2266), .A3(n2140), .A4(n2248), .ZN(n49) );
  ND2D1 U3015 ( .A1(n2443), .A2(n2445), .ZN(n10) );
  NR4D0 U3016 ( .A1(n56), .A2(n2339), .A3(FrameSR[21]), .A4(n2285), .ZN(n51)
         );
  NR4D0 U3017 ( .A1(n55), .A2(n2087), .A3(FrameSR[35]), .A4(n2304), .ZN(n52)
         );
  NR4D0 U3018 ( .A1(n54), .A2(n2105), .A3(FrameSR[50]), .A4(n2322), .ZN(n53)
         );
  NR2D1 U3019 ( .A1(n2346), .A2(n3132), .ZN(n195) );
  XOR2D1 U3020 ( .A1(n2460), .A2(n10), .Z(n11) );
  INVD1 U3021 ( .I(n2460), .ZN(n7) );
  ND3D1 U3022 ( .A1(n137), .A2(n136), .A3(n138), .ZN(n54) );
  ND3D1 U3023 ( .A1(n153), .A2(n152), .A3(n154), .ZN(n55) );
  ND3D1 U3024 ( .A1(n168), .A2(n159), .A3(n169), .ZN(n56) );
  INVD1 U3025 ( .I(n2445), .ZN(n6) );
  INR2D1 U3026 ( .A1(n3074), .B1(n3132), .ZN(n193) );
  OAI31D0 U3027 ( .A1(n6), .A2(n2444), .A3(n7), .B(n2443), .ZN(n3074) );
  NR2D1 U3028 ( .A1(n2375), .A2(n3132), .ZN(n196) );
  NR2D1 U3029 ( .A1(n3132), .A2(n1698), .ZN(n194) );
  NR2D1 U3030 ( .A1(n7), .A2(n10), .ZN(n9) );
  AN2D1 U3031 ( .A1(SerClk), .A2(n2431), .Z(SerClock) );
  INVD1 U3032 ( .I(Reset), .ZN(n261) );
  CKND0 U3033 ( .CLK(n3149), .CN(n3131) );
endmodule


module DesDecoder_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

