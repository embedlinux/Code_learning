
module FullDup ( OutParDataA, OutParDataB, InParDataA, InParDataB, InParValidA, 
        InParValidB, ClockA, ClockB, Reset );
  output [31:0] OutParDataA;
  output [31:0] OutParDataB;
  input [31:0] InParDataA;
  input [31:0] InParDataB;
  input InParValidA, InParValidB, ClockA, ClockB, Reset;
  wire   \*Logic1* , SerLine1, SerLine2, n1, n2, n3, n4, n5;

  SerDes_DWid32_RxLogDepth4_TxLogDepth3 SerDes_U1 ( .ParOutRxClk(OutParDataB), 
        .SerLineXfer(SerLine1), .ParDataIn(InParDataA), .InParClk(n3), 
        .InParValid(InParValidA), .OutParClk(n2), .RxRequest(\*Logic1* ), 
        .TxRequest(InParValidA), .Reset(n4) );
  SerDes_DWid32_RxLogDepth3_TxLogDepth4 SerDes_U2 ( .ParOutRxClk(OutParDataA), 
        .SerLineXfer(SerLine2), .ParDataIn(InParDataB), .InParClk(n2), 
        .InParValid(InParValidB), .OutParClk(n3), .RxRequest(\*Logic1* ), 
        .TxRequest(InParValidB), .Reset(n4) );
  INVD1 U2 ( .I(n5), .ZN(n4) );
  INVD1 U3 ( .I(n1), .ZN(n5) );
  BUFFD1 U4 ( .I(Reset), .Z(n1) );
  BUFFD1 U5 ( .I(ClockB), .Z(n2) );
  BUFFD1 U6 ( .I(ClockA), .Z(n3) );
  TIEH U7 ( .Z(\*Logic1* ) );
endmodule


module SerDes_DWid32_RxLogDepth4_TxLogDepth3 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4;

  Serializer_DWid32_AWid3 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n4), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid4_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n3), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD2 U1 ( .I(OutParClk), .Z(n3) );
  INVD1 U2 ( .I(n2), .ZN(n1) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  BUFFD1 U4 ( .I(InParClk), .Z(n4) );
endmodule


module SerDes_DWid32_RxLogDepth3_TxLogDepth4 ( ParOutRxClk, SerLineXfer, 
        ParDataIn, InParClk, InParValid, OutParClk, RxRequest, TxRequest, 
        Reset );
  output [31:0] ParOutRxClk;
  input [31:0] ParDataIn;
  input InParClk, InParValid, OutParClk, RxRequest, TxRequest, Reset;
  output SerLineXfer;
  wire   SerLineValid, Tx_F_Empty, Tx_F_Full, Rx_F_Empty, Rx_F_Full, n1, n2,
         n3, n4;

  Serializer_DWid32_AWid4 Ser_U1 ( .SerOut(SerLineXfer), .SerValid(
        SerLineValid), .FIFOEmpty(Tx_F_Empty), .FIFOFull(Tx_F_Full), .ParIn(
        ParDataIn), .InParValid(InParValid), .ParInClk(n3), .SendSerial(
        TxRequest), .Reset(n1) );
  Deserializer_AWid3_DWid32 Des_U1 ( .ParOut(ParOutRxClk), .FIFOEmpty(
        Rx_F_Empty), .FIFOFull(Rx_F_Full), .ParOutClk(n4), .SerialIn(
        SerLineXfer), .ReadReq(RxRequest), .SerValid(SerLineValid), .Reset(n1)
         );
  BUFFD2 U1 ( .I(OutParClk), .Z(n4) );
  INVD1 U2 ( .I(n2), .ZN(n1) );
  INVD1 U3 ( .I(Reset), .ZN(n2) );
  BUFFD1 U4 ( .I(InParClk), .Z(n3) );
endmodule


module Serializer_DWid32_AWid3 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid3_DWid32_0 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(F_ReadReq), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n1) );
  SerEncoder_DWid32_0 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n1) );
  SerialTx_0 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n1) );
  INVD1 U1 ( .I(n3), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n3) );
  AN3D1 U3 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U4 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U5 ( .A1(n1), .A2(FIFOEmpty), .ZN(F_Valid) );
  INR2D1 U6 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
endmodule


module Deserializer_AWid4_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n4, n6,
         n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34,
         n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62,
         n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid4_DWid32_0 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n98)
         );
  DesDecoder_DWid32_0 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n98) );
  SerialRx_0 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n98) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n102), .Q(n104) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n101), .Q(n105) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n101), .Q(n106) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n101), .Q(n107) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n101), .Q(n108) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n101), .Q(n109) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n101), .Q(n110) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n101), .Q(n111) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n101), .Q(n112) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n101), .Q(n113) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n101), .Q(n114) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n101), .Q(n115) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n101), .Q(n116) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n101), .Q(n117) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n100), .Q(n118) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n100), .Q(n119) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n100), .Q(n120) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n100), .Q(n121) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n100), .Q(n122) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n100), .Q(n123) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n100), .Q(n124) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n100), .Q(n125) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n100), .Q(n126) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n100), .Q(n127) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n100), .Q(n128) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n100), .Q(n129) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n100), .Q(n130) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n99), .Q(n131) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n99), .Q(n132) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n99), .Q(n133) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n99), .Q(n134) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n99), .Q(n135) );
  DFCNQD1 ParValidr_reg ( .D(N35), .CP(ParOutClk), .CDN(n102), .Q(ParValid) );
  CKBD0 U3 ( .CLK(n97), .C(n1) );
  CKNXD16 U4 ( .I(n1), .ZN(ParOut[31]) );
  CKBD0 U5 ( .CLK(n96), .C(n4) );
  CKNXD16 U6 ( .I(n4), .ZN(ParOut[30]) );
  CKBD0 U7 ( .CLK(n95), .C(n6) );
  CKNXD16 U8 ( .I(n6), .ZN(ParOut[29]) );
  CKBD0 U9 ( .CLK(n94), .C(n8) );
  CKNXD16 U10 ( .I(n8), .ZN(ParOut[28]) );
  CKBD0 U11 ( .CLK(n93), .C(n10) );
  CKNXD16 U12 ( .I(n10), .ZN(ParOut[27]) );
  CKBD0 U13 ( .CLK(n92), .C(n12) );
  CKNXD16 U14 ( .I(n12), .ZN(ParOut[26]) );
  CKBD0 U15 ( .CLK(n91), .C(n14) );
  CKNXD16 U16 ( .I(n14), .ZN(ParOut[25]) );
  CKBD0 U17 ( .CLK(n90), .C(n16) );
  CKNXD16 U18 ( .I(n16), .ZN(ParOut[24]) );
  CKBD0 U19 ( .CLK(n89), .C(n18) );
  CKNXD16 U20 ( .I(n18), .ZN(ParOut[23]) );
  CKBD0 U21 ( .CLK(n88), .C(n20) );
  CKNXD16 U22 ( .I(n20), .ZN(ParOut[22]) );
  CKBD0 U23 ( .CLK(n87), .C(n22) );
  CKNXD16 U24 ( .I(n22), .ZN(ParOut[21]) );
  CKBD0 U25 ( .CLK(n86), .C(n24) );
  CKNXD16 U26 ( .I(n24), .ZN(ParOut[20]) );
  CKBD0 U27 ( .CLK(n85), .C(n26) );
  CKNXD16 U28 ( .I(n26), .ZN(ParOut[19]) );
  CKBD0 U29 ( .CLK(n84), .C(n28) );
  CKNXD16 U30 ( .I(n28), .ZN(ParOut[18]) );
  CKBD0 U31 ( .CLK(n83), .C(n30) );
  CKNXD16 U32 ( .I(n30), .ZN(ParOut[17]) );
  CKBD0 U33 ( .CLK(n82), .C(n32) );
  CKNXD16 U34 ( .I(n32), .ZN(ParOut[16]) );
  CKBD0 U35 ( .CLK(n81), .C(n34) );
  CKNXD16 U36 ( .I(n34), .ZN(ParOut[15]) );
  CKBD0 U37 ( .CLK(n80), .C(n36) );
  CKNXD16 U38 ( .I(n36), .ZN(ParOut[14]) );
  CKBD0 U39 ( .CLK(n79), .C(n38) );
  CKNXD16 U40 ( .I(n38), .ZN(ParOut[13]) );
  CKBD0 U41 ( .CLK(n78), .C(n40) );
  CKNXD16 U42 ( .I(n40), .ZN(ParOut[12]) );
  CKBD0 U43 ( .CLK(n77), .C(n42) );
  CKNXD16 U44 ( .I(n42), .ZN(ParOut[11]) );
  CKBD0 U45 ( .CLK(n76), .C(n44) );
  CKNXD16 U46 ( .I(n44), .ZN(ParOut[10]) );
  CKBD0 U47 ( .CLK(n75), .C(n46) );
  CKNXD16 U48 ( .I(n46), .ZN(ParOut[9]) );
  CKBD0 U49 ( .CLK(n74), .C(n48) );
  CKNXD16 U50 ( .I(n48), .ZN(ParOut[8]) );
  CKBD0 U51 ( .CLK(n73), .C(n50) );
  CKNXD16 U52 ( .I(n50), .ZN(ParOut[7]) );
  CKBD0 U53 ( .CLK(n72), .C(n52) );
  CKNXD16 U54 ( .I(n52), .ZN(ParOut[6]) );
  CKBD0 U55 ( .CLK(n71), .C(n54) );
  CKNXD16 U56 ( .I(n54), .ZN(ParOut[5]) );
  CKBD0 U57 ( .CLK(n70), .C(n56) );
  CKNXD16 U58 ( .I(n56), .ZN(ParOut[4]) );
  CKBD0 U59 ( .CLK(n69), .C(n58) );
  CKNXD16 U60 ( .I(n58), .ZN(ParOut[3]) );
  CKBD0 U61 ( .CLK(n68), .C(n60) );
  CKNXD16 U62 ( .I(n60), .ZN(ParOut[2]) );
  CKBD0 U63 ( .CLK(n67), .C(n62) );
  CKNXD16 U64 ( .I(n62), .ZN(ParOut[1]) );
  CKBD0 U65 ( .CLK(n66), .C(n64) );
  CKNXD16 U66 ( .I(n64), .ZN(ParOut[0]) );
  INVD1 U67 ( .I(n99), .ZN(n98) );
  BUFFD1 U68 ( .I(n103), .Z(n99) );
  BUFFD1 U69 ( .I(n103), .Z(n100) );
  BUFFD1 U70 ( .I(n103), .Z(n101) );
  BUFFD1 U71 ( .I(n103), .Z(n102) );
  INVD1 U72 ( .I(Reset), .ZN(n103) );
  NR2D1 U73 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  INVD0 U74 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U75 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U76 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U77 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U78 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U79 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U80 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U81 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U82 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U83 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U84 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U85 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U86 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U87 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U88 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U89 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U90 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U91 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U92 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U93 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U94 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U95 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U96 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U97 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U98 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U99 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U100 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U101 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U102 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U103 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U104 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U105 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U106 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U107 ( .CLK(n135), .CN(n66) );
  CKND0 U108 ( .CLK(n134), .CN(n67) );
  CKND0 U109 ( .CLK(n133), .CN(n68) );
  CKND0 U110 ( .CLK(n132), .CN(n69) );
  CKND0 U111 ( .CLK(n131), .CN(n70) );
  CKND0 U112 ( .CLK(n130), .CN(n71) );
  CKND0 U113 ( .CLK(n129), .CN(n72) );
  CKND0 U114 ( .CLK(n128), .CN(n73) );
  CKND0 U115 ( .CLK(n127), .CN(n74) );
  CKND0 U116 ( .CLK(n126), .CN(n75) );
  CKND0 U117 ( .CLK(n125), .CN(n76) );
  CKND0 U118 ( .CLK(n124), .CN(n77) );
  CKND0 U119 ( .CLK(n123), .CN(n78) );
  CKND0 U120 ( .CLK(n122), .CN(n79) );
  CKND0 U121 ( .CLK(n121), .CN(n80) );
  CKND0 U122 ( .CLK(n120), .CN(n81) );
  CKND0 U123 ( .CLK(n119), .CN(n82) );
  CKND0 U124 ( .CLK(n118), .CN(n83) );
  CKND0 U125 ( .CLK(n117), .CN(n84) );
  CKND0 U126 ( .CLK(n116), .CN(n85) );
  CKND0 U127 ( .CLK(n115), .CN(n86) );
  CKND0 U128 ( .CLK(n114), .CN(n87) );
  CKND0 U129 ( .CLK(n113), .CN(n88) );
  CKND0 U130 ( .CLK(n112), .CN(n89) );
  CKND0 U131 ( .CLK(n111), .CN(n90) );
  CKND0 U132 ( .CLK(n110), .CN(n91) );
  CKND0 U133 ( .CLK(n109), .CN(n92) );
  CKND0 U134 ( .CLK(n108), .CN(n93) );
  CKND0 U135 ( .CLK(n107), .CN(n94) );
  CKND0 U136 ( .CLK(n106), .CN(n95) );
  CKND0 U137 ( .CLK(n105), .CN(n96) );
  CKND0 U138 ( .CLK(n104), .CN(n97) );
endmodule


module Serializer_DWid32_AWid4 ( SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk, 
        ParIn, InParValid, ParInClk, SendSerial, Reset );
  input [31:0] ParIn;
  input InParValid, ParInClk, SendSerial, Reset;
  output SerOut, SerValid, FIFOEmpty, FIFOFull, SerClk;
  wire   F_Valid, SerEncReadReq, F_ReadReq, F_WriteReq, EncD_ToTx, n2, n1, n3;
  wire   [31:0] FIFO_Out;

  FIFOTop_AWid4_DWid32_1 FIFO_Tx1 ( .Dout(FIFO_Out), .Din(ParIn), .Full(
        FIFOFull), .Empty(FIFOEmpty), .ReadIn(F_ReadReq), .WriteIn(F_WriteReq), 
        .ClkR(ParInClk), .ClkW(ParInClk), .Reseter(n1) );
  SerEncoder_DWid32_1 SerEnc_Tx1 ( .SerOut(EncD_ToTx), .SerValid(SerValid), 
        .FIFO_ReadReq(SerEncReadReq), .ParIn(FIFO_Out), .F_Empty(FIFOEmpty), 
        .ParClk(ParInClk), .SerClk(SerClk), .ParValid(F_Valid), .Reset(n1) );
  SerialTx_1 SerTx_Tx1 ( .SerOut(SerOut), .SerClk(SerClk), .SerIn(EncD_ToTx), 
        .ParClk(ParInClk), .Reset(n1) );
  INVD1 U1 ( .I(n3), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n3) );
  AN3D1 U3 ( .A1(n2), .A2(SendSerial), .A3(SerEncReadReq), .Z(F_ReadReq) );
  INVD1 U4 ( .I(FIFOEmpty), .ZN(n2) );
  NR2D1 U5 ( .A1(n1), .A2(FIFOEmpty), .ZN(F_Valid) );
  INR2D1 U6 ( .A1(InParValid), .B1(FIFOFull), .ZN(F_WriteReq) );
endmodule


module Deserializer_AWid3_DWid32 ( ParOut, ParValid, DecoderParClk, FIFOEmpty, 
        FIFOFull, ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, ParValidDecode, SerialClk, SerRxToDecode, n3, n1, n4, n6,
         n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34,
         n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62,
         n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid3_DWid32_1 FIFO_Rx1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), 
        .Full(FIFOFull), .Empty(FIFOEmpty), .ReadIn(ReadReq), .WriteIn(
        ParValidDecode), .ClkR(ParOutClk), .ClkW(DecoderParClk), .Reseter(n98)
         );
  DesDecoder_DWid32_1 DesDec_Rx1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(DecoderParClk), .SerIn(SerRxToDecode), 
        .SerClk(SerialClk), .SerValid(SerValid), .Reset(n98) );
  SerialRx_1 SerRx_Rx1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(DecoderParClk), .Reset(n98) );
  DFCNQD1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n102), .Q(n104) );
  DFCNQD1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n101), .Q(n105) );
  DFCNQD1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n101), .Q(n106) );
  DFCNQD1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n101), .Q(n107) );
  DFCNQD1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n101), .Q(n108) );
  DFCNQD1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n101), .Q(n109) );
  DFCNQD1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n101), .Q(n110) );
  DFCNQD1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n101), .Q(n111) );
  DFCNQD1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n101), .Q(n112) );
  DFCNQD1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n101), .Q(n113) );
  DFCNQD1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n101), .Q(n114) );
  DFCNQD1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n101), .Q(n115) );
  DFCNQD1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n101), .Q(n116) );
  DFCNQD1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n101), .Q(n117) );
  DFCNQD1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n100), .Q(n118) );
  DFCNQD1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n100), .Q(n119) );
  DFCNQD1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n100), .Q(n120) );
  DFCNQD1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n100), .Q(n121) );
  DFCNQD1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n100), .Q(n122) );
  DFCNQD1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n100), .Q(n123) );
  DFCNQD1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n100), .Q(n124) );
  DFCNQD1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n100), .Q(n125) );
  DFCNQD1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n100), .Q(n126) );
  DFCNQD1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n100), .Q(n127) );
  DFCNQD1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n100), .Q(n128) );
  DFCNQD1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n100), .Q(n129) );
  DFCNQD1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n100), .Q(n130) );
  DFCNQD1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n99), .Q(n131) );
  DFCNQD1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n99), .Q(n132) );
  DFCNQD1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n99), .Q(n133) );
  DFCNQD1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n99), .Q(n134) );
  DFCNQD1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n99), .Q(n135) );
  DFCNQD1 ParValidr_reg ( .D(N35), .CP(ParOutClk), .CDN(n102), .Q(ParValid) );
  CKBD0 U3 ( .CLK(n97), .C(n1) );
  CKNXD16 U4 ( .I(n1), .ZN(ParOut[31]) );
  CKBD0 U5 ( .CLK(n96), .C(n4) );
  CKNXD16 U6 ( .I(n4), .ZN(ParOut[30]) );
  CKBD0 U7 ( .CLK(n95), .C(n6) );
  CKNXD16 U8 ( .I(n6), .ZN(ParOut[29]) );
  CKBD0 U9 ( .CLK(n94), .C(n8) );
  CKNXD16 U10 ( .I(n8), .ZN(ParOut[28]) );
  CKBD0 U11 ( .CLK(n93), .C(n10) );
  CKNXD16 U12 ( .I(n10), .ZN(ParOut[27]) );
  CKBD0 U13 ( .CLK(n92), .C(n12) );
  CKNXD16 U14 ( .I(n12), .ZN(ParOut[26]) );
  CKBD0 U15 ( .CLK(n91), .C(n14) );
  CKNXD16 U16 ( .I(n14), .ZN(ParOut[25]) );
  CKBD0 U17 ( .CLK(n90), .C(n16) );
  CKNXD16 U18 ( .I(n16), .ZN(ParOut[24]) );
  CKBD0 U19 ( .CLK(n89), .C(n18) );
  CKNXD16 U20 ( .I(n18), .ZN(ParOut[23]) );
  CKBD0 U21 ( .CLK(n88), .C(n20) );
  CKNXD16 U22 ( .I(n20), .ZN(ParOut[22]) );
  CKBD0 U23 ( .CLK(n87), .C(n22) );
  CKNXD16 U24 ( .I(n22), .ZN(ParOut[21]) );
  CKBD0 U25 ( .CLK(n86), .C(n24) );
  CKNXD16 U26 ( .I(n24), .ZN(ParOut[20]) );
  CKBD0 U27 ( .CLK(n85), .C(n26) );
  CKNXD16 U28 ( .I(n26), .ZN(ParOut[19]) );
  CKBD0 U29 ( .CLK(n84), .C(n28) );
  CKNXD16 U30 ( .I(n28), .ZN(ParOut[18]) );
  CKBD0 U31 ( .CLK(n83), .C(n30) );
  CKNXD16 U32 ( .I(n30), .ZN(ParOut[17]) );
  CKBD0 U33 ( .CLK(n82), .C(n32) );
  CKNXD16 U34 ( .I(n32), .ZN(ParOut[16]) );
  CKBD0 U35 ( .CLK(n81), .C(n34) );
  CKNXD16 U36 ( .I(n34), .ZN(ParOut[15]) );
  CKBD0 U37 ( .CLK(n80), .C(n36) );
  CKNXD16 U38 ( .I(n36), .ZN(ParOut[14]) );
  CKBD0 U39 ( .CLK(n79), .C(n38) );
  CKNXD16 U40 ( .I(n38), .ZN(ParOut[13]) );
  CKBD0 U41 ( .CLK(n78), .C(n40) );
  CKNXD16 U42 ( .I(n40), .ZN(ParOut[12]) );
  CKBD0 U43 ( .CLK(n77), .C(n42) );
  CKNXD16 U44 ( .I(n42), .ZN(ParOut[11]) );
  CKBD0 U45 ( .CLK(n76), .C(n44) );
  CKNXD16 U46 ( .I(n44), .ZN(ParOut[10]) );
  CKBD0 U47 ( .CLK(n75), .C(n46) );
  CKNXD16 U48 ( .I(n46), .ZN(ParOut[9]) );
  CKBD0 U49 ( .CLK(n74), .C(n48) );
  CKNXD16 U50 ( .I(n48), .ZN(ParOut[8]) );
  CKBD0 U51 ( .CLK(n73), .C(n50) );
  CKNXD16 U52 ( .I(n50), .ZN(ParOut[7]) );
  CKBD0 U53 ( .CLK(n72), .C(n52) );
  CKNXD16 U54 ( .I(n52), .ZN(ParOut[6]) );
  CKBD0 U55 ( .CLK(n71), .C(n54) );
  CKNXD16 U56 ( .I(n54), .ZN(ParOut[5]) );
  CKBD0 U57 ( .CLK(n70), .C(n56) );
  CKNXD16 U58 ( .I(n56), .ZN(ParOut[4]) );
  CKBD0 U59 ( .CLK(n69), .C(n58) );
  CKNXD16 U60 ( .I(n58), .ZN(ParOut[3]) );
  CKBD0 U61 ( .CLK(n68), .C(n60) );
  CKNXD16 U62 ( .I(n60), .ZN(ParOut[2]) );
  CKBD0 U63 ( .CLK(n67), .C(n62) );
  CKNXD16 U64 ( .I(n62), .ZN(ParOut[1]) );
  CKBD0 U65 ( .CLK(n66), .C(n64) );
  CKNXD16 U66 ( .I(n64), .ZN(ParOut[0]) );
  INVD1 U67 ( .I(n99), .ZN(n98) );
  BUFFD1 U68 ( .I(n103), .Z(n99) );
  BUFFD1 U69 ( .I(n103), .Z(n100) );
  BUFFD1 U70 ( .I(n103), .Z(n101) );
  BUFFD1 U71 ( .I(n103), .Z(n102) );
  INVD1 U72 ( .I(Reset), .ZN(n103) );
  NR2D1 U73 ( .A1(FIFOEmpty), .A2(n3), .ZN(N35) );
  INVD0 U74 ( .I(ReadReq), .ZN(n3) );
  CKAN2D0 U75 ( .A1(FIFO_Out[0]), .A2(ReadReq), .Z(N3) );
  CKAN2D0 U76 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  CKAN2D0 U77 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  CKAN2D0 U78 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  CKAN2D0 U79 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  CKAN2D0 U80 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  CKAN2D0 U81 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  CKAN2D0 U82 ( .A1(FIFO_Out[7]), .A2(ReadReq), .Z(N10) );
  CKAN2D0 U83 ( .A1(FIFO_Out[8]), .A2(ReadReq), .Z(N11) );
  CKAN2D0 U84 ( .A1(FIFO_Out[9]), .A2(ReadReq), .Z(N12) );
  CKAN2D0 U85 ( .A1(FIFO_Out[10]), .A2(ReadReq), .Z(N13) );
  CKAN2D0 U86 ( .A1(FIFO_Out[11]), .A2(ReadReq), .Z(N14) );
  CKAN2D0 U87 ( .A1(FIFO_Out[12]), .A2(ReadReq), .Z(N15) );
  CKAN2D0 U88 ( .A1(FIFO_Out[13]), .A2(ReadReq), .Z(N16) );
  CKAN2D0 U89 ( .A1(FIFO_Out[14]), .A2(ReadReq), .Z(N17) );
  CKAN2D0 U90 ( .A1(FIFO_Out[15]), .A2(ReadReq), .Z(N18) );
  CKAN2D0 U91 ( .A1(FIFO_Out[16]), .A2(ReadReq), .Z(N19) );
  CKAN2D0 U92 ( .A1(FIFO_Out[17]), .A2(ReadReq), .Z(N20) );
  CKAN2D0 U93 ( .A1(FIFO_Out[18]), .A2(ReadReq), .Z(N21) );
  CKAN2D0 U94 ( .A1(FIFO_Out[19]), .A2(ReadReq), .Z(N22) );
  CKAN2D0 U95 ( .A1(FIFO_Out[20]), .A2(ReadReq), .Z(N23) );
  CKAN2D0 U96 ( .A1(FIFO_Out[21]), .A2(ReadReq), .Z(N24) );
  CKAN2D0 U97 ( .A1(FIFO_Out[22]), .A2(ReadReq), .Z(N25) );
  CKAN2D0 U98 ( .A1(FIFO_Out[23]), .A2(ReadReq), .Z(N26) );
  CKAN2D0 U99 ( .A1(FIFO_Out[24]), .A2(ReadReq), .Z(N27) );
  CKAN2D0 U100 ( .A1(FIFO_Out[25]), .A2(ReadReq), .Z(N28) );
  CKAN2D0 U101 ( .A1(FIFO_Out[26]), .A2(ReadReq), .Z(N29) );
  CKAN2D0 U102 ( .A1(FIFO_Out[27]), .A2(ReadReq), .Z(N30) );
  CKAN2D0 U103 ( .A1(FIFO_Out[28]), .A2(ReadReq), .Z(N31) );
  CKAN2D0 U104 ( .A1(FIFO_Out[29]), .A2(ReadReq), .Z(N32) );
  CKAN2D0 U105 ( .A1(FIFO_Out[30]), .A2(ReadReq), .Z(N33) );
  CKAN2D0 U106 ( .A1(FIFO_Out[31]), .A2(ReadReq), .Z(N34) );
  CKND0 U107 ( .CLK(n135), .CN(n66) );
  CKND0 U108 ( .CLK(n134), .CN(n67) );
  CKND0 U109 ( .CLK(n133), .CN(n68) );
  CKND0 U110 ( .CLK(n132), .CN(n69) );
  CKND0 U111 ( .CLK(n131), .CN(n70) );
  CKND0 U112 ( .CLK(n130), .CN(n71) );
  CKND0 U113 ( .CLK(n129), .CN(n72) );
  CKND0 U114 ( .CLK(n128), .CN(n73) );
  CKND0 U115 ( .CLK(n127), .CN(n74) );
  CKND0 U116 ( .CLK(n126), .CN(n75) );
  CKND0 U117 ( .CLK(n125), .CN(n76) );
  CKND0 U118 ( .CLK(n124), .CN(n77) );
  CKND0 U119 ( .CLK(n123), .CN(n78) );
  CKND0 U120 ( .CLK(n122), .CN(n79) );
  CKND0 U121 ( .CLK(n121), .CN(n80) );
  CKND0 U122 ( .CLK(n120), .CN(n81) );
  CKND0 U123 ( .CLK(n119), .CN(n82) );
  CKND0 U124 ( .CLK(n118), .CN(n83) );
  CKND0 U125 ( .CLK(n117), .CN(n84) );
  CKND0 U126 ( .CLK(n116), .CN(n85) );
  CKND0 U127 ( .CLK(n115), .CN(n86) );
  CKND0 U128 ( .CLK(n114), .CN(n87) );
  CKND0 U129 ( .CLK(n113), .CN(n88) );
  CKND0 U130 ( .CLK(n112), .CN(n89) );
  CKND0 U131 ( .CLK(n111), .CN(n90) );
  CKND0 U132 ( .CLK(n110), .CN(n91) );
  CKND0 U133 ( .CLK(n109), .CN(n92) );
  CKND0 U134 ( .CLK(n108), .CN(n93) );
  CKND0 U135 ( .CLK(n107), .CN(n94) );
  CKND0 U136 ( .CLK(n106), .CN(n95) );
  CKND0 U137 ( .CLK(n105), .CN(n96) );
  CKND0 U138 ( .CLK(n104), .CN(n97) );
endmodule


module FIFOTop_AWid3_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid3_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD1 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_0 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_0_DW01_dec_0 \ShifterBlock/sub_132  ( .A({\Sh_N[5] , N6, 
        N5, N4, N3, N2}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n26), .CP(n36), .CDN(n48), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n40), .CP(ParClk), .CDN(n45), .Q(HalfParClkr)
         );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(n39), .CDN(n45), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n39), .CDN(n45), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n39), .CDN(n46), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n38), .CDN(n46), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n38), .CDN(n46), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(n38), .CDN(n46), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(n38), .CDN(n47), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(n38), .CDN(n47), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(n37), .CDN(n47), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n37), .CDN(n47), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n37), .CDN(n47), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(n37), .CDN(n47), .Q(InBuf[9]) );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n36), .CDN(n48), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(n36), .CDN(n48), .Q(InBuf[5]) );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n36), .CDN(n48), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(n36), .CDN(n48), .Q(InBuf[1]) );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(n39), .CDN(n45), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n39), .CDN(n46), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(n39), .CDN(n46), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(n38), .CDN(n46), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(n38), .CDN(n46), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n38), .CDN(n46), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n38), .CDN(n46), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(n37), .CDN(n47), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(n37), .CDN(n47), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(n37), .CDN(n47), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(n37), .CDN(n47), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(n37), .CDN(n48), .Q(InBuf[8]) );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n36), .CDN(n48), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(n36), .CDN(n48), .Q(InBuf[4]) );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n36), .CDN(n48), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(n36), .CDN(n48), .Q(InBuf[0]) );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n45), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n45), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n45), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n45), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n45), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n45), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(N31), .CP(SerClk), .CDN(n47), .Q(SerOut) );
  BUFFD1 U3 ( .I(n42), .Z(n49) );
  INVD1 U4 ( .I(n50), .ZN(n48) );
  BUFFD1 U5 ( .I(n42), .Z(n50) );
  INVD1 U6 ( .I(n51), .ZN(n47) );
  BUFFD1 U7 ( .I(n43), .Z(n51) );
  INVD1 U8 ( .I(n52), .ZN(n46) );
  BUFFD1 U9 ( .I(n43), .Z(n52) );
  BUFFD1 U10 ( .I(Reset), .Z(n42) );
  BUFFD1 U11 ( .I(Reset), .Z(n43) );
  INVD1 U12 ( .I(n53), .ZN(n45) );
  BUFFD1 U13 ( .I(n44), .Z(n53) );
  BUFFD1 U14 ( .I(Reset), .Z(n44) );
  INVD1 U15 ( .I(n31), .ZN(n26) );
  INVD1 U16 ( .I(n31), .ZN(n27) );
  INVD1 U17 ( .I(n30), .ZN(n28) );
  INVD1 U18 ( .I(n40), .ZN(n36) );
  INVD1 U19 ( .I(n40), .ZN(n37) );
  INVD1 U20 ( .I(n41), .ZN(n38) );
  INVD1 U21 ( .I(n41), .ZN(n39) );
  INVD1 U22 ( .I(n30), .ZN(n29) );
  INVD1 U23 ( .I(n55), .ZN(n54) );
  INVD1 U24 ( .I(n33), .ZN(n31) );
  INVD1 U25 ( .I(n34), .ZN(n40) );
  INVD1 U26 ( .I(n33), .ZN(n30) );
  INVD1 U27 ( .I(n34), .ZN(n41) );
  ND2D1 U28 ( .A1(N3), .A2(N2), .ZN(n56) );
  AN2D1 U29 ( .A1(N4), .A2(n54), .Z(N26) );
  MUX2D0 U30 ( .I0(n6), .I1(n7), .S(N4), .Z(n22) );
  MUX4ND0 U31 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n6) );
  MUX4ND0 U32 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n7) );
  MUX2D0 U33 ( .I0(n8), .I1(n9), .S(N4), .Z(n20) );
  MUX4ND0 U34 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n8) );
  MUX4ND0 U35 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n9) );
  MUX2D0 U36 ( .I0(n10), .I1(n11), .S(N4), .Z(n18) );
  MUX4ND0 U37 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n10) );
  MUX4ND0 U38 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n11) );
  MUX2D0 U39 ( .I0(n12), .I1(n13), .S(N4), .Z(n24) );
  MUX4ND0 U40 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n12) );
  MUX4ND0 U41 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n13) );
  NR2D1 U42 ( .A1(n56), .A2(N4), .ZN(N24) );
  INVD1 U43 ( .I(n32), .ZN(n33) );
  INVD1 U44 ( .I(N85), .ZN(n32) );
  INVD1 U45 ( .I(n35), .ZN(n34) );
  INVD1 U46 ( .I(HalfParClkr), .ZN(n35) );
  MUX2ND0 U47 ( .I0(n14), .I1(n15), .S(N6), .ZN(N29) );
  MUX2ND0 U48 ( .I0(n16), .I1(n17), .S(N6), .ZN(N27) );
  MUX2ND0 U49 ( .I0(n15), .I1(n14), .S(N6), .ZN(N25) );
  MUX2ND0 U50 ( .I0(n17), .I1(n16), .S(N6), .ZN(N23) );
  CKND1 U51 ( .CLK(n18), .CN(n19) );
  CKND1 U52 ( .CLK(n20), .CN(n21) );
  MUX2ND0 U53 ( .I0(n21), .I1(n19), .S(N5), .ZN(n15) );
  CKND1 U54 ( .CLK(n22), .CN(n23) );
  CKND1 U55 ( .CLK(n24), .CN(n25) );
  MUX2ND0 U56 ( .I0(n25), .I1(n23), .S(N5), .ZN(n14) );
  MUX2ND0 U57 ( .I0(n19), .I1(n25), .S(N5), .ZN(n17) );
  MUX2ND0 U58 ( .I0(n23), .I1(n21), .S(N5), .ZN(n16) );
  OR2D1 U59 ( .A1(N2), .A2(N3), .Z(n55) );
  MUX2ND0 U60 ( .I0(n56), .I1(n55), .S(N4), .ZN(N28) );
  AN2D0 U61 ( .A1(ParIn[31]), .A2(n29), .Z(N84) );
  AN2D0 U62 ( .A1(ParIn[30]), .A2(n29), .Z(N83) );
  AN2D0 U63 ( .A1(ParIn[29]), .A2(n29), .Z(N82) );
  AN2D0 U64 ( .A1(ParIn[28]), .A2(n29), .Z(N81) );
  AN2D0 U65 ( .A1(ParIn[27]), .A2(n28), .Z(N80) );
  AN2D0 U66 ( .A1(ParIn[26]), .A2(n28), .Z(N79) );
  AN2D0 U67 ( .A1(ParIn[25]), .A2(n28), .Z(N78) );
  AN2D0 U68 ( .A1(ParIn[24]), .A2(n28), .Z(N77) );
  AN2D0 U69 ( .A1(ParIn[23]), .A2(n28), .Z(N76) );
  AN2D0 U70 ( .A1(ParIn[22]), .A2(n28), .Z(N75) );
  AN2D0 U71 ( .A1(ParIn[21]), .A2(n28), .Z(N74) );
  AN2D0 U72 ( .A1(ParIn[20]), .A2(n28), .Z(N73) );
  AN2D0 U73 ( .A1(ParIn[19]), .A2(n28), .Z(N72) );
  AN2D0 U74 ( .A1(ParIn[18]), .A2(n28), .Z(N71) );
  AN2D0 U75 ( .A1(ParIn[17]), .A2(n27), .Z(N70) );
  AN2D0 U76 ( .A1(ParIn[16]), .A2(n27), .Z(N69) );
  AN2D0 U77 ( .A1(ParIn[15]), .A2(n27), .Z(N68) );
  AN2D0 U78 ( .A1(ParIn[14]), .A2(n27), .Z(N67) );
  AN2D0 U79 ( .A1(ParIn[13]), .A2(n27), .Z(N66) );
  AN2D0 U80 ( .A1(ParIn[12]), .A2(n27), .Z(N65) );
  AN2D0 U81 ( .A1(ParIn[11]), .A2(n27), .Z(N64) );
  AN2D0 U82 ( .A1(ParIn[10]), .A2(n27), .Z(N63) );
  AN2D0 U83 ( .A1(ParIn[9]), .A2(n27), .Z(N62) );
  AN2D0 U84 ( .A1(ParIn[8]), .A2(n27), .Z(N61) );
  AN2D0 U85 ( .A1(ParIn[7]), .A2(n26), .Z(N60) );
  AN2D0 U86 ( .A1(ParIn[6]), .A2(n26), .Z(N59) );
  AN2D0 U87 ( .A1(ParIn[5]), .A2(n26), .Z(N58) );
  AN2D0 U88 ( .A1(ParIn[4]), .A2(n26), .Z(N57) );
  AN2D0 U89 ( .A1(ParIn[3]), .A2(n26), .Z(N56) );
  AN2D0 U90 ( .A1(ParIn[2]), .A2(n26), .Z(N55) );
  AN2D0 U91 ( .A1(ParIn[1]), .A2(n26), .Z(N54) );
  AN2D0 U92 ( .A1(ParIn[0]), .A2(n26), .Z(N53) );
  IND2D0 U93 ( .A1(n57), .B1(n58), .ZN(N31) );
  OAI21D0 U94 ( .A1(N23), .A2(n59), .B(n60), .ZN(n58) );
  MUX2ND0 U95 ( .I0(n61), .I1(n62), .S(n59), .ZN(n60) );
  MUX3ND0 U96 ( .I0(N25), .I1(n63), .I2(N24), .S0(\Sh_N[5] ), .S1(n64), .ZN(
        n62) );
  NR2D0 U97 ( .A1(\Sh_N[5] ), .A2(N5), .ZN(n64) );
  MUX2D0 U98 ( .I0(n65), .I1(N26), .S(n66), .Z(n63) );
  NR2D0 U99 ( .A1(N6), .A2(N5), .ZN(n66) );
  INR2D0 U100 ( .A1(N27), .B1(N6), .ZN(n65) );
  CKND0 U101 ( .CLK(N5), .CN(n61) );
  CKND2D0 U102 ( .A1(n67), .A2(n68), .ZN(n59) );
  MUX2ND0 U103 ( .I0(n69), .I1(n70), .S(N5), .ZN(n57) );
  CKND2D0 U104 ( .A1(N29), .A2(n71), .ZN(n70) );
  CKND2D0 U105 ( .A1(N28), .A2(n71), .ZN(n69) );
  NR2D0 U106 ( .A1(n68), .A2(n67), .ZN(n71) );
  CKND0 U107 ( .CLK(N6), .CN(n67) );
  CKND0 U108 ( .CLK(\Sh_N[5] ), .CN(n68) );
  INR3D0 U109 ( .A1(n26), .B1(n49), .B2(n40), .ZN(FIFO_ReadReq) );
  INR2D0 U110 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
endmodule


module SerialTx_0 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_0 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_0 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_0 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid4_DWid32_0 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD1 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_0 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n230, n231, n232, n84, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U17 ( .A1(n266), .A2(n32), .B1(n268), .B2(Decoder[31]), .ZN(n101)
         );
  MOAI22D1 U18 ( .A1(n266), .A2(n33), .B1(n268), .B2(Decoder[30]), .ZN(n102)
         );
  MOAI22D1 U19 ( .A1(n266), .A2(n34), .B1(n268), .B2(Decoder[29]), .ZN(n103)
         );
  MOAI22D1 U20 ( .A1(n266), .A2(n35), .B1(n268), .B2(Decoder[28]), .ZN(n104)
         );
  MOAI22D1 U21 ( .A1(n266), .A2(n36), .B1(n267), .B2(Decoder[27]), .ZN(n105)
         );
  MOAI22D1 U22 ( .A1(n266), .A2(n37), .B1(n267), .B2(Decoder[26]), .ZN(n106)
         );
  MOAI22D1 U23 ( .A1(n266), .A2(n38), .B1(n267), .B2(Decoder[25]), .ZN(n107)
         );
  MOAI22D1 U24 ( .A1(n266), .A2(n39), .B1(n267), .B2(Decoder[24]), .ZN(n108)
         );
  MOAI22D1 U25 ( .A1(n266), .A2(n40), .B1(n267), .B2(Decoder[23]), .ZN(n109)
         );
  MOAI22D1 U26 ( .A1(n266), .A2(n41), .B1(n267), .B2(Decoder[22]), .ZN(n110)
         );
  MOAI22D1 U27 ( .A1(n266), .A2(n42), .B1(n267), .B2(Decoder[21]), .ZN(n111)
         );
  MOAI22D1 U28 ( .A1(n266), .A2(n43), .B1(n266), .B2(Decoder[20]), .ZN(n112)
         );
  MOAI22D1 U29 ( .A1(n266), .A2(n44), .B1(n267), .B2(Decoder[19]), .ZN(n113)
         );
  MOAI22D1 U30 ( .A1(n266), .A2(n45), .B1(n267), .B2(Decoder[18]), .ZN(n114)
         );
  MOAI22D1 U31 ( .A1(n266), .A2(n46), .B1(n267), .B2(Decoder[17]), .ZN(n115)
         );
  MOAI22D1 U32 ( .A1(n266), .A2(n47), .B1(n267), .B2(Decoder[16]), .ZN(n116)
         );
  MOAI22D1 U33 ( .A1(n266), .A2(n48), .B1(n267), .B2(Decoder[15]), .ZN(n117)
         );
  MOAI22D1 U34 ( .A1(n266), .A2(n49), .B1(n267), .B2(Decoder[14]), .ZN(n118)
         );
  MOAI22D1 U35 ( .A1(n265), .A2(n50), .B1(n267), .B2(Decoder[13]), .ZN(n119)
         );
  MOAI22D1 U36 ( .A1(n265), .A2(n51), .B1(n267), .B2(Decoder[12]), .ZN(n120)
         );
  MOAI22D1 U37 ( .A1(n265), .A2(n52), .B1(n267), .B2(Decoder[11]), .ZN(n121)
         );
  MOAI22D1 U38 ( .A1(n265), .A2(n53), .B1(n267), .B2(Decoder[10]), .ZN(n122)
         );
  MOAI22D1 U39 ( .A1(n265), .A2(n54), .B1(n267), .B2(Decoder[9]), .ZN(n123) );
  MOAI22D1 U40 ( .A1(n265), .A2(n55), .B1(n267), .B2(Decoder[8]), .ZN(n124) );
  MOAI22D1 U41 ( .A1(n265), .A2(n56), .B1(n268), .B2(Decoder[7]), .ZN(n125) );
  MOAI22D1 U42 ( .A1(n265), .A2(n57), .B1(n267), .B2(Decoder[6]), .ZN(n126) );
  MOAI22D1 U43 ( .A1(n265), .A2(n58), .B1(n268), .B2(Decoder[5]), .ZN(n127) );
  MOAI22D1 U44 ( .A1(n265), .A2(n59), .B1(n268), .B2(Decoder[4]), .ZN(n128) );
  MOAI22D1 U45 ( .A1(n265), .A2(n60), .B1(n268), .B2(Decoder[3]), .ZN(n129) );
  MOAI22D1 U46 ( .A1(n265), .A2(n61), .B1(n268), .B2(Decoder[2]), .ZN(n130) );
  MOAI22D1 U47 ( .A1(n265), .A2(n62), .B1(n268), .B2(Decoder[1]), .ZN(n131) );
  MOAI22D1 U48 ( .A1(n266), .A2(n63), .B1(n268), .B2(Decoder[0]), .ZN(n132) );
  OR3D1 U92 ( .A1(FrameSR[55]), .A2(FrameSR[54]), .A3(FrameSR[53]), .Z(n22) );
  OR3D1 U94 ( .A1(FrameSR[39]), .A2(FrameSR[38]), .A3(FrameSR[37]), .Z(n23) );
  OR3D1 U96 ( .A1(FrameSR[32]), .A2(FrameSR[23]), .A3(FrameSR[22]), .Z(n24) );
  OA21D1 U99 ( .A1(n26), .A2(n27), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n28) );
  DesDecoder_DWid32_0_DW01_inc_0 \ClkGen/add_206  ( .A(Count32), .SUM({N34, 
        N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(FrameSR[62]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(FrameSR[21]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(FrameSR[22]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(FrameSR[36]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(FrameSR[37]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(FrameSR[52]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(FrameSR[53]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(FrameSR[31]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(FrameSR[38]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(FrameSR[54]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(FrameSR[7]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(FrameSR[8]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(FrameSR[9]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(FrameSR[10]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(FrameSR[11]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(FrameSR[12]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(FrameSR[13]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(FrameSR[14]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(FrameSR[18]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(FrameSR[23]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(FrameSR[24]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(FrameSR[25]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(FrameSR[26]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(FrameSR[27]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(FrameSR[28]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(FrameSR[29]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(FrameSR[30]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(FrameSR[39]), .CPN(n293), .CDN(n302), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(FrameSR[40]), .CPN(n293), .CDN(n302), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(FrameSR[41]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(FrameSR[42]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(FrameSR[43]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(FrameSR[44]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(FrameSR[45]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(FrameSR[46]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(FrameSR[55]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(FrameSR[56]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(FrameSR[57]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(FrameSR[58]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(FrameSR[59]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(FrameSR[60]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(FrameSR[61]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n297), .CDN(n298), .Q(FrameSR[0])
         );
  DFNCND1 \FrameSR_reg[4]  ( .D(FrameSR[3]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(FrameSR[19]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(FrameSR[33]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(FrameSR[48]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(FrameSR[1]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(FrameSR[5]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(FrameSR[17]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(FrameSR[32]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(FrameSR[47]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(FrameSR[0]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(FrameSR[2]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(FrameSR[4]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(FrameSR[6]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(FrameSR[20]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(FrameSR[34]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(FrameSR[49]), .CPN(n292), .CDN(n303), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(FrameSR[50]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(FrameSR[35]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(FrameSR[51]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(FrameSR[16]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(FrameSR[15]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(N42), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n164), .CPN(n290), .CDN(n304), .Q(Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n163), .CPN(n290), .CDN(n304), .Q(Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n162), .CPN(n290), .CDN(n304), .Q(Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n161), .CPN(n290), .CDN(n304), .Q(Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n160), .CPN(n290), .CDN(n304), .Q(Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n159), .CPN(n289), .CDN(n304), .Q(Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n158), .CPN(n289), .CDN(n305), .Q(Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n157), .CPN(n289), .CDN(n305), .Q(Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n156), .CPN(n289), .CDN(n305), .Q(Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n155), .CPN(n289), .CDN(n305), .Q(Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n154), .CPN(n289), .CDN(n305), .Q(Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n153), .CPN(n289), .CDN(n305), .Q(Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n152), .CPN(n289), .CDN(n305), .Q(Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n151), .CPN(n289), .CDN(n305), .Q(Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n150), .CPN(n288), .CDN(n305), .Q(Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n149), .CPN(n288), .CDN(n305), .Q(Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n148), .CPN(n288), .CDN(n306), .Q(Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n147), .CPN(n288), .CDN(n306), .Q(Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n146), .CPN(n288), .CDN(n306), .Q(Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n145), .CPN(n288), .CDN(n306), .Q(Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n144), .CPN(n288), .CDN(n306), .Q(Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n143), .CPN(n288), .CDN(n306), .Q(Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n142), .CPN(n288), .CDN(n306), .Q(Decoder[9])
         );
  DFNCND1 \Decoder_reg[8]  ( .D(n141), .CPN(n287), .CDN(n306), .Q(Decoder[8])
         );
  DFNCND1 \Decoder_reg[7]  ( .D(n140), .CPN(n287), .CDN(n306), .Q(Decoder[7])
         );
  DFNCND1 \Decoder_reg[6]  ( .D(n139), .CPN(n287), .CDN(n306), .Q(Decoder[6])
         );
  DFNCND1 \Decoder_reg[5]  ( .D(n138), .CPN(n287), .CDN(n307), .Q(Decoder[5])
         );
  DFNCND1 \Decoder_reg[4]  ( .D(n137), .CPN(n287), .CDN(n307), .Q(Decoder[4])
         );
  DFNCND1 \Decoder_reg[3]  ( .D(n136), .CPN(n287), .CDN(n307), .Q(Decoder[3])
         );
  DFNCND1 \Decoder_reg[2]  ( .D(n135), .CPN(n287), .CDN(n307), .Q(Decoder[2])
         );
  DFNCND1 \Decoder_reg[1]  ( .D(n134), .CPN(n287), .CDN(n307), .Q(Decoder[1])
         );
  DFNCND1 \Decoder_reg[0]  ( .D(n133), .CPN(n287), .CDN(n307), .Q(Decoder[0])
         );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n99), .CPN(n283), .CDN(n311), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(N39), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n100), .CPN(n283), .CDN(n311), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(N41), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(N40), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(N38), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[0]  ( .D(n132), .CPN(n286), .CDN(n307), .Q(ParOut[0]), 
        .QN(n63) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n131), .CPN(n286), .CDN(n307), .Q(ParOut[1]), 
        .QN(n62) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n130), .CPN(n286), .CDN(n308), .Q(ParOut[2]), 
        .QN(n61) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n129), .CPN(n286), .CDN(n308), .Q(ParOut[3]), 
        .QN(n60) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n128), .CPN(n286), .CDN(n308), .Q(ParOut[4]), 
        .QN(n59) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n127), .CPN(n286), .CDN(n308), .Q(ParOut[5]), 
        .QN(n58) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n126), .CPN(n286), .CDN(n308), .Q(ParOut[6]), 
        .QN(n57) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n125), .CPN(n285), .CDN(n308), .Q(ParOut[7]), 
        .QN(n56) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n124), .CPN(n285), .CDN(n308), .Q(ParOut[8]), 
        .QN(n55) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n123), .CPN(n285), .CDN(n308), .Q(ParOut[9]), 
        .QN(n54) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n122), .CPN(n285), .CDN(n308), .Q(ParOut[10]), 
        .QN(n53) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n121), .CPN(n285), .CDN(n308), .Q(ParOut[11]), 
        .QN(n52) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n120), .CPN(n285), .CDN(n309), .Q(ParOut[12]), 
        .QN(n51) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n119), .CPN(n285), .CDN(n309), .Q(ParOut[13]), 
        .QN(n50) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n118), .CPN(n285), .CDN(n309), .Q(ParOut[14]), 
        .QN(n49) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n117), .CPN(n285), .CDN(n309), .Q(ParOut[15]), 
        .QN(n48) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n116), .CPN(n284), .CDN(n309), .Q(ParOut[16]), 
        .QN(n47) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n115), .CPN(n284), .CDN(n309), .Q(ParOut[17]), 
        .QN(n46) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n114), .CPN(n284), .CDN(n309), .Q(ParOut[18]), 
        .QN(n45) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n113), .CPN(n284), .CDN(n309), .Q(ParOut[19]), 
        .QN(n44) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n112), .CPN(n284), .CDN(n309), .Q(ParOut[20]), 
        .QN(n43) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n111), .CPN(n284), .CDN(n309), .Q(ParOut[21]), 
        .QN(n42) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n110), .CPN(n284), .CDN(n310), .Q(ParOut[22]), 
        .QN(n41) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n109), .CPN(n284), .CDN(n310), .Q(ParOut[23]), 
        .QN(n40) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n108), .CPN(n284), .CDN(n310), .Q(ParOut[24]), 
        .QN(n39) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n107), .CPN(n283), .CDN(n310), .Q(ParOut[25]), 
        .QN(n38) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n106), .CPN(n283), .CDN(n310), .Q(ParOut[26]), 
        .QN(n37) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n105), .CPN(n283), .CDN(n310), .Q(ParOut[27]), 
        .QN(n36) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n104), .CPN(n283), .CDN(n310), .Q(ParOut[28]), 
        .QN(n35) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n103), .CPN(n283), .CDN(n310), .Q(ParOut[29]), 
        .QN(n34) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n102), .CPN(n283), .CDN(n310), .Q(ParOut[30]), 
        .QN(n33) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n101), .CPN(n283), .CDN(n310), .Q(ParOut[31]), 
        .QN(n32) );
  EDFCNQD1 ParClkr_reg ( .D(N37), .E(N43), .CP(n282), .CDN(n311), .Q(ParClk)
         );
  DFNCND1 ParValidr_reg ( .D(n96), .CPN(n282), .CDN(n311), .Q(ParValid), .QN(
        n29) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n286), .CDN(n322), .Q(n27), .QN(n2) );
  DFNCND1 UnLoad_reg ( .D(n258), .CPN(n286), .CDN(n322), .Q(n5), .QN(n231) );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n97), .CPN(n282), .CDN(n322), .QN(n232)
         );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n98), .CPN(n282), .CDN(n322), .QN(n230)
         );
  BUFFD1 U3 ( .I(n313), .Z(n309) );
  BUFFD1 U4 ( .I(n313), .Z(n308) );
  BUFFD1 U5 ( .I(n314), .Z(n307) );
  BUFFD1 U6 ( .I(n314), .Z(n306) );
  BUFFD1 U7 ( .I(n315), .Z(n305) );
  BUFFD1 U8 ( .I(n315), .Z(n304) );
  BUFFD1 U9 ( .I(n316), .Z(n303) );
  BUFFD1 U10 ( .I(n316), .Z(n302) );
  BUFFD1 U11 ( .I(n317), .Z(n301) );
  BUFFD1 U12 ( .I(n317), .Z(n300) );
  BUFFD1 U13 ( .I(n318), .Z(n299) );
  BUFFD1 U14 ( .I(n318), .Z(n298) );
  BUFFD1 U15 ( .I(n312), .Z(n311) );
  BUFFD1 U16 ( .I(n312), .Z(n310) );
  BUFFD1 U49 ( .I(n320), .Z(n313) );
  BUFFD1 U50 ( .I(n320), .Z(n314) );
  BUFFD1 U51 ( .I(n320), .Z(n315) );
  BUFFD1 U52 ( .I(n319), .Z(n316) );
  BUFFD1 U53 ( .I(n319), .Z(n317) );
  BUFFD1 U54 ( .I(n319), .Z(n318) );
  BUFFD1 U55 ( .I(n321), .Z(n312) );
  BUFFD1 U56 ( .I(n322), .Z(n321) );
  BUFFD1 U57 ( .I(n322), .Z(n320) );
  BUFFD1 U58 ( .I(n322), .Z(n319) );
  INVD1 U59 ( .I(Reset), .ZN(n322) );
  INVD1 U60 ( .I(n260), .ZN(n257) );
  INVD1 U61 ( .I(n261), .ZN(n256) );
  INVD1 U62 ( .I(n262), .ZN(n255) );
  INVD1 U63 ( .I(n259), .ZN(n258) );
  BUFFD1 U64 ( .I(n271), .Z(n282) );
  BUFFD1 U65 ( .I(n271), .Z(n283) );
  BUFFD1 U66 ( .I(n272), .Z(n284) );
  BUFFD1 U67 ( .I(n272), .Z(n285) );
  BUFFD1 U68 ( .I(n273), .Z(n286) );
  BUFFD1 U69 ( .I(n273), .Z(n287) );
  BUFFD1 U70 ( .I(n274), .Z(n288) );
  BUFFD1 U71 ( .I(n274), .Z(n289) );
  BUFFD1 U72 ( .I(n275), .Z(n290) );
  BUFFD1 U73 ( .I(n275), .Z(n291) );
  BUFFD1 U74 ( .I(n276), .Z(n292) );
  BUFFD1 U75 ( .I(n276), .Z(n293) );
  BUFFD1 U76 ( .I(n277), .Z(n294) );
  BUFFD1 U77 ( .I(n277), .Z(n295) );
  BUFFD1 U78 ( .I(n278), .Z(n296) );
  BUFFD1 U79 ( .I(n278), .Z(n297) );
  INVD1 U80 ( .I(n270), .ZN(n265) );
  INVD1 U81 ( .I(n270), .ZN(n266) );
  INVD1 U82 ( .I(n269), .ZN(n267) );
  INVD1 U83 ( .I(n269), .ZN(n268) );
  BUFFD1 U84 ( .I(n13), .Z(n259) );
  BUFFD1 U85 ( .I(n13), .Z(n260) );
  BUFFD1 U86 ( .I(n13), .Z(n261) );
  BUFFD1 U87 ( .I(n13), .Z(n262) );
  BUFFD1 U88 ( .I(n280), .Z(n273) );
  BUFFD1 U89 ( .I(n280), .Z(n274) );
  BUFFD1 U90 ( .I(n280), .Z(n275) );
  BUFFD1 U91 ( .I(n279), .Z(n276) );
  BUFFD1 U93 ( .I(n279), .Z(n277) );
  BUFFD1 U95 ( .I(n279), .Z(n278) );
  BUFFD1 U97 ( .I(n281), .Z(n271) );
  BUFFD1 U98 ( .I(n281), .Z(n272) );
  INVD1 U100 ( .I(n263), .ZN(n270) );
  INVD1 U102 ( .I(n263), .ZN(n269) );
  IND2D1 U103 ( .A1(n14), .B1(n15), .ZN(n13) );
  NR2D1 U104 ( .A1(n15), .A2(n14), .ZN(N47) );
  BUFFD1 U105 ( .I(SerClock), .Z(n280) );
  BUFFD1 U106 ( .I(SerClock), .Z(n279) );
  BUFFD1 U107 ( .I(SerClock), .Z(n281) );
  OAI21D1 U108 ( .A1(n3), .A2(n29), .B(n231), .ZN(n96) );
  NR2D1 U109 ( .A1(ParClk), .A2(n232), .ZN(n3) );
  NR2D1 U110 ( .A1(ParClk), .A2(n27), .ZN(N37) );
  NR4D0 U111 ( .A1(n28), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n26) );
  AN2D1 U112 ( .A1(N34), .A2(n2), .Z(N42) );
  AN2D1 U113 ( .A1(N33), .A2(n2), .Z(N41) );
  AN2D1 U114 ( .A1(N32), .A2(n2), .Z(N40) );
  AN2D1 U115 ( .A1(N31), .A2(n2), .Z(N39) );
  AN2D1 U116 ( .A1(N30), .A2(n2), .Z(N38) );
  ND2D1 U117 ( .A1(n232), .A2(ParValidTimer[0]), .ZN(n10) );
  INVD1 U118 ( .I(ParValidTimer[1]), .ZN(n7) );
  AO22D0 U119 ( .A1(FrameSR[8]), .A2(n257), .B1(Decoder[0]), .B2(n259), .Z(
        n133) );
  AO22D0 U120 ( .A1(FrameSR[9]), .A2(n257), .B1(Decoder[1]), .B2(n259), .Z(
        n134) );
  AO22D0 U121 ( .A1(FrameSR[10]), .A2(n257), .B1(Decoder[2]), .B2(n259), .Z(
        n135) );
  AO22D0 U122 ( .A1(FrameSR[11]), .A2(n258), .B1(Decoder[3]), .B2(n259), .Z(
        n136) );
  AO22D0 U123 ( .A1(FrameSR[12]), .A2(n258), .B1(Decoder[4]), .B2(n259), .Z(
        n137) );
  AO22D0 U124 ( .A1(FrameSR[13]), .A2(n258), .B1(Decoder[5]), .B2(n259), .Z(
        n138) );
  AO22D0 U125 ( .A1(FrameSR[14]), .A2(n258), .B1(Decoder[6]), .B2(n259), .Z(
        n139) );
  AO22D0 U126 ( .A1(FrameSR[15]), .A2(n258), .B1(Decoder[7]), .B2(n259), .Z(
        n140) );
  AO22D0 U127 ( .A1(FrameSR[24]), .A2(n255), .B1(Decoder[8]), .B2(n260), .Z(
        n141) );
  AO22D0 U128 ( .A1(FrameSR[25]), .A2(n256), .B1(Decoder[9]), .B2(n260), .Z(
        n142) );
  AO22D0 U129 ( .A1(FrameSR[26]), .A2(n256), .B1(Decoder[10]), .B2(n260), .Z(
        n143) );
  AO22D0 U130 ( .A1(FrameSR[27]), .A2(n256), .B1(Decoder[11]), .B2(n260), .Z(
        n144) );
  AO22D0 U131 ( .A1(FrameSR[28]), .A2(n257), .B1(Decoder[12]), .B2(n260), .Z(
        n145) );
  AO22D0 U132 ( .A1(FrameSR[29]), .A2(n257), .B1(Decoder[13]), .B2(n260), .Z(
        n146) );
  AO22D0 U133 ( .A1(FrameSR[30]), .A2(n257), .B1(Decoder[14]), .B2(n260), .Z(
        n147) );
  AO22D0 U134 ( .A1(FrameSR[31]), .A2(n257), .B1(Decoder[15]), .B2(n260), .Z(
        n148) );
  AO22D0 U135 ( .A1(FrameSR[40]), .A2(n257), .B1(Decoder[16]), .B2(n261), .Z(
        n149) );
  AO22D0 U136 ( .A1(FrameSR[41]), .A2(n257), .B1(Decoder[17]), .B2(n261), .Z(
        n150) );
  AO22D0 U137 ( .A1(FrameSR[42]), .A2(n255), .B1(Decoder[18]), .B2(n261), .Z(
        n151) );
  AO22D0 U138 ( .A1(FrameSR[43]), .A2(n255), .B1(Decoder[19]), .B2(n261), .Z(
        n152) );
  AO22D0 U139 ( .A1(FrameSR[44]), .A2(n255), .B1(Decoder[20]), .B2(n261), .Z(
        n153) );
  AO22D0 U140 ( .A1(FrameSR[45]), .A2(n255), .B1(Decoder[21]), .B2(n261), .Z(
        n154) );
  AO22D0 U141 ( .A1(FrameSR[46]), .A2(n256), .B1(Decoder[22]), .B2(n261), .Z(
        n155) );
  AO22D0 U142 ( .A1(FrameSR[47]), .A2(n256), .B1(Decoder[23]), .B2(n261), .Z(
        n156) );
  AO22D0 U143 ( .A1(FrameSR[56]), .A2(n256), .B1(Decoder[24]), .B2(n262), .Z(
        n157) );
  AO22D0 U144 ( .A1(FrameSR[57]), .A2(n256), .B1(Decoder[25]), .B2(n262), .Z(
        n158) );
  AO22D0 U145 ( .A1(FrameSR[58]), .A2(n256), .B1(Decoder[26]), .B2(n262), .Z(
        n159) );
  AO22D0 U146 ( .A1(FrameSR[59]), .A2(n256), .B1(Decoder[27]), .B2(n262), .Z(
        n160) );
  AO22D0 U147 ( .A1(FrameSR[60]), .A2(n255), .B1(Decoder[28]), .B2(n262), .Z(
        n161) );
  AO22D0 U148 ( .A1(FrameSR[61]), .A2(n255), .B1(Decoder[29]), .B2(n262), .Z(
        n162) );
  AO22D0 U149 ( .A1(FrameSR[62]), .A2(n255), .B1(Decoder[30]), .B2(n262), .Z(
        n163) );
  AO22D0 U150 ( .A1(FrameSR[63]), .A2(n255), .B1(Decoder[31]), .B2(n262), .Z(
        n164) );
  INVD1 U151 ( .I(ParValidTimer[0]), .ZN(n6) );
  INR2D1 U152 ( .A1(n84), .B1(n265), .ZN(n97) );
  OAI31D0 U153 ( .A1(n6), .A2(n230), .A3(n7), .B(n232), .ZN(n84) );
  NR2D1 U154 ( .A1(n11), .A2(n265), .ZN(n99) );
  XOR2D1 U155 ( .A1(ParValidTimer[1]), .A2(n10), .Z(n11) );
  NR2D1 U156 ( .A1(n12), .A2(n265), .ZN(n100) );
  XOR2D1 U157 ( .A1(n232), .A2(n6), .Z(n12) );
  INVD1 U158 ( .I(n264), .ZN(n263) );
  INVD1 U159 ( .I(n5), .ZN(n264) );
  NR2D1 U160 ( .A1(n265), .A2(n8), .ZN(n98) );
  XOR2D1 U161 ( .A1(n230), .A2(n9), .Z(n8) );
  NR2D1 U162 ( .A1(n7), .A2(n10), .ZN(n9) );
  NR4D0 U163 ( .A1(n22), .A2(FrameSR[48]), .A3(FrameSR[50]), .A4(FrameSR[49]), 
        .ZN(n21) );
  ND2D1 U164 ( .A1(n16), .A2(n17), .ZN(n14) );
  NR4D0 U165 ( .A1(FrameSR[3]), .A2(FrameSR[2]), .A3(FrameSR[1]), .A4(
        FrameSR[0]), .ZN(n16) );
  NR4D0 U166 ( .A1(FrameSR[7]), .A2(FrameSR[6]), .A3(FrameSR[5]), .A4(
        FrameSR[4]), .ZN(n17) );
  AN4D1 U167 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .Z(n15) );
  INR4D0 U168 ( .A1(FrameSR[19]), .B1(n25), .B2(FrameSR[17]), .B3(FrameSR[16]), 
        .ZN(n18) );
  NR4D0 U169 ( .A1(n24), .A2(FrameSR[18]), .A3(FrameSR[21]), .A4(FrameSR[20]), 
        .ZN(n19) );
  NR4D0 U170 ( .A1(n23), .A2(FrameSR[33]), .A3(FrameSR[35]), .A4(FrameSR[34]), 
        .ZN(n20) );
  ND3D1 U171 ( .A1(FrameSR[51]), .A2(FrameSR[36]), .A3(FrameSR[52]), .ZN(n25)
         );
  AN2D1 U172 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_0 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_3 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n178, StateClockRaw, StateClock, N46, N47, N48, N49, N63, N64, N65,
         N66, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n115, n121, n122,
         n124, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n140, n141, n142, n143, n144, n174, n175, n176, n177;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n128), .CPN(StateClock), .Q(FullFIFO), .QN(n115) );
  DFND1 EmptyFIFOr_reg ( .D(n127), .CPN(StateClock), .Q(EmptyFIFO) );
  IAO21D1 U6 ( .A1(n39), .A2(n40), .B(n176), .ZN(n38) );
  MOAI22D1 U7 ( .A1(n142), .A2(n41), .B1(n41), .B2(OldReadAr[1]), .ZN(n129) );
  MOAI22D1 U8 ( .A1(n141), .A2(n41), .B1(n41), .B2(OldReadAr[2]), .ZN(n130) );
  MOAI22D1 U9 ( .A1(n42), .A2(n43), .B1(n42), .B2(OldWriteAr[1]), .ZN(n131) );
  MOAI22D1 U10 ( .A1(n42), .A2(n44), .B1(n42), .B2(OldWriteAr[2]), .ZN(n132)
         );
  MOAI22D1 U11 ( .A1(n144), .A2(n42), .B1(n42), .B2(OldWriteAr[0]), .ZN(n133)
         );
  MOAI22D1 U70 ( .A1(n143), .A2(n41), .B1(n41), .B2(OldReadAr[0]), .ZN(n140)
         );
  DFNCND1 \NextState_reg[0]  ( .D(n137), .CPN(StateClock), .CDN(n174), .Q(
        NextState[0]), .QN(n124) );
  DFNCND1 \NextState_reg[1]  ( .D(n135), .CPN(StateClock), .CDN(n175), .Q(
        NextState[1]), .QN(n122) );
  DFNCND1 \NextState_reg[2]  ( .D(n134), .CPN(StateClock), .CDN(n174), .Q(
        NextState[2]), .QN(n121) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n175), 
        .Q(CurState[2]) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n175), 
        .Q(CurState[1]) );
  EDFCNQD1 \WriteAr_reg[2]  ( .D(N65), .E(N66), .CP(StateClock), .CDN(n175), 
        .Q(WriteAddr[2]) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n175), 
        .Q(CurState[0]) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(N64), .E(N66), .CP(StateClock), .CDN(n175), 
        .Q(WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N48), .CP(StateClock), .CDN(n177), .Q(
        ReadAddr[2]), .QN(n141) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N47), .E(N48), .CP(StateClock), .CDN(n177), .Q(
        ReadAddr[1]), .QN(n142) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N46), .E(N48), .CP(StateClock), .CDN(n177), .Q(
        ReadAddr[0]), .QN(n143) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N63), .E(N66), .CP(StateClock), .CDN(n177), 
        .Q(n178), .QN(n144) );
  DFNCND1 WriteCmdr_reg ( .D(n136), .CPN(StateClock), .CDN(n177), .Q(WriteCmd), 
        .QN(n85) );
  DFNCND1 ReadCmdr_reg ( .D(n138), .CPN(StateClock), .CDN(n177), .Q(ReadCmd)
         );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n131), .CPN(StateClock), .CDN(n177), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n132), .CPN(StateClock), .CDN(n177), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n133), .CPN(StateClock), .CDN(n177), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n130), .CPN(StateClock), .CDN(n177), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n129), .CPN(StateClock), .CDN(n177), .Q(
        OldReadAr[1]) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n140), .CPN(StateClock), .CDN(n177), .Q(
        OldReadAr[0]) );
  INVD1 U3 ( .I(n176), .ZN(n174) );
  INVD1 U4 ( .I(n176), .ZN(n175) );
  INVD1 U5 ( .I(n177), .ZN(n176) );
  INVD1 U12 ( .I(Reset), .ZN(n177) );
  INVD1 U13 ( .I(n77), .ZN(n84) );
  MAOI22D0 U14 ( .A1(ReadAddr[0]), .A2(n75), .B1(n43), .B2(n98), .ZN(n101) );
  INVD1 U15 ( .I(n40), .ZN(n35) );
  ND2D1 U16 ( .A1(n83), .A2(n37), .ZN(n86) );
  ND2D1 U17 ( .A1(WriteReq), .A2(n45), .ZN(n42) );
  ND2D1 U18 ( .A1(ReadReq), .A2(n86), .ZN(n41) );
  INVD1 U19 ( .I(n46), .ZN(n52) );
  NR2D1 U20 ( .A1(n68), .A2(n79), .ZN(n39) );
  ND2D1 U21 ( .A1(n83), .A2(n35), .ZN(n45) );
  XNR2D1 U22 ( .A1(n44), .A2(n75), .ZN(n77) );
  INVD1 U23 ( .I(n75), .ZN(n81) );
  XNR2D1 U24 ( .A1(n84), .A2(ReadAddr[2]), .ZN(n56) );
  ND3D1 U25 ( .A1(n37), .A2(n35), .A3(n112), .ZN(N66) );
  NR2D1 U26 ( .A1(ReadAddr[0]), .A2(n109), .ZN(N46) );
  NR2D1 U27 ( .A1(n99), .A2(n109), .ZN(N49) );
  NR2D1 U28 ( .A1(n113), .A2(n109), .ZN(N47) );
  XNR2D1 U29 ( .A1(ReadAddr[0]), .A2(ReadAddr[1]), .ZN(n113) );
  INVD1 U30 ( .I(ReadReq), .ZN(n106) );
  MAOI22D0 U31 ( .A1(n178), .A2(n103), .B1(n142), .B2(n98), .ZN(n102) );
  OAI222D0 U32 ( .A1(n44), .A2(ReadAddr[2]), .B1(n43), .B2(ReadAddr[1]), .C1(
        n144), .C2(ReadAddr[0]), .ZN(n73) );
  OAI33D1 U33 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n101), .B1(n44), .B2(
        WriteAddr[1]), .B3(n102), .ZN(n54) );
  OAI33D1 U34 ( .A1(ReadAddr[1]), .A2(n101), .A3(n44), .B1(n102), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n55) );
  AOI22D0 U35 ( .A1(n68), .A2(CurState[1]), .B1(n51), .B2(n39), .ZN(n83) );
  NR3D0 U36 ( .A1(CurState[1]), .A2(CurState[2]), .A3(CurState[0]), .ZN(n40)
         );
  OAI211D1 U37 ( .A1(CurState[1]), .A2(n79), .B(n83), .C(n104), .ZN(n46) );
  AOI21D1 U38 ( .A1(WriteReq), .A2(n40), .B(n105), .ZN(n104) );
  AOI21D1 U39 ( .A1(CurState[0]), .A2(n106), .B(n68), .ZN(n105) );
  ND2D1 U40 ( .A1(CurState[1]), .A2(n39), .ZN(n37) );
  INVD1 U41 ( .I(WriteAddr[2]), .ZN(n44) );
  OAI33D1 U42 ( .A1(n85), .A2(n40), .A3(n86), .B1(n87), .B2(n88), .B3(n89), 
        .ZN(n136) );
  XNR2D1 U43 ( .A1(n44), .A2(OldWriteAr[2]), .ZN(n89) );
  XNR2D1 U44 ( .A1(n43), .A2(OldWriteAr[1]), .ZN(n88) );
  INVD1 U45 ( .I(WriteAddr[1]), .ZN(n43) );
  NR2D1 U46 ( .A1(n43), .A2(n144), .ZN(n75) );
  OAI211D1 U47 ( .A1(n144), .A2(ReadAddr[1]), .B(n80), .C(n81), .ZN(n78) );
  OAI21D1 U48 ( .A1(WriteAddr[1]), .A2(n142), .B(n143), .ZN(n80) );
  OAI21D1 U49 ( .A1(WriteAddr[1]), .A2(n178), .B(n81), .ZN(n100) );
  INVD1 U50 ( .I(CurState[0]), .ZN(n79) );
  OAI32D1 U51 ( .A1(n107), .A2(n108), .A3(n106), .B1(n86), .B2(n109), .ZN(n138) );
  XNR2D1 U52 ( .A1(n142), .A2(OldReadAr[1]), .ZN(n108) );
  ND3D1 U53 ( .A1(n110), .A2(n86), .A3(n111), .ZN(n107) );
  XNR2D1 U54 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .ZN(n110) );
  XOR2D1 U55 ( .A1(n100), .A2(n142), .Z(n57) );
  INVD1 U56 ( .I(CurState[2]), .ZN(n68) );
  ND2D1 U57 ( .A1(n144), .A2(n143), .ZN(n98) );
  AOI31D0 U58 ( .A1(n65), .A2(n66), .A3(n67), .B(n68), .ZN(n64) );
  AOI22D0 U59 ( .A1(n69), .A2(ReadAddr[1]), .B1(n144), .B2(ReadAddr[0]), .ZN(
        n67) );
  OAI21D1 U60 ( .A1(n69), .A2(n73), .B(n43), .ZN(n65) );
  OAI21D1 U61 ( .A1(ReadAddr[1]), .A2(n72), .B(n73), .ZN(n66) );
  OAI22D0 U62 ( .A1(n46), .A2(n122), .B1(n52), .B2(n59), .ZN(n135) );
  AOI31D0 U63 ( .A1(n60), .A2(n61), .A3(n62), .B(n40), .ZN(n59) );
  IIND4D1 U64 ( .A1(n69), .A2(n73), .B1(n78), .B2(n79), .ZN(n61) );
  AOI31D0 U65 ( .A1(n143), .A2(CurState[0]), .A3(n63), .B(n64), .ZN(n62) );
  OAI22D0 U66 ( .A1(n46), .A2(n124), .B1(n52), .B2(n92), .ZN(n137) );
  AOI21D1 U67 ( .A1(CurState[1]), .A2(n93), .B(n39), .ZN(n92) );
  OAI21D1 U68 ( .A1(CurState[2]), .A2(n94), .B(n95), .ZN(n93) );
  AOI22D0 U69 ( .A1(n55), .A2(ReadAddr[2]), .B1(n141), .B2(n54), .ZN(n94) );
  OAI31D0 U71 ( .A1(n96), .A2(n97), .A3(n58), .B(CurState[0]), .ZN(n95) );
  XNR2D1 U72 ( .A1(WriteAddr[2]), .A2(n99), .ZN(n97) );
  INVD1 U73 ( .I(n57), .ZN(n96) );
  OAI21D1 U74 ( .A1(n46), .A2(n121), .B(n47), .ZN(n134) );
  OAI211D1 U75 ( .A1(CurState[2]), .A2(n48), .B(CurState[0]), .C(n49), .ZN(n47) );
  AOI21D1 U76 ( .A1(n50), .A2(n51), .B(n52), .ZN(n49) );
  NR4D0 U77 ( .A1(n56), .A2(n57), .A3(n51), .A4(n58), .ZN(n48) );
  INVD1 U78 ( .I(CurState[1]), .ZN(n51) );
  NR3D0 U79 ( .A1(n57), .A2(n144), .A3(n74), .ZN(n63) );
  AOI21D1 U80 ( .A1(n69), .A2(n75), .B(n76), .ZN(n74) );
  OAI32D1 U81 ( .A1(n44), .A2(n141), .A3(n75), .B1(ReadAddr[2]), .B2(n77), 
        .ZN(n76) );
  AOI31D0 U82 ( .A1(n144), .A2(CurState[0]), .A3(n82), .B(n83), .ZN(n60) );
  NR3D0 U83 ( .A1(n57), .A2(n143), .A3(n56), .ZN(n82) );
  NR2D1 U84 ( .A1(n143), .A2(n142), .ZN(n103) );
  XOR2D1 U85 ( .A1(n103), .A2(n141), .Z(n99) );
  AO22D0 U86 ( .A1(ReadAddr[2]), .A2(n54), .B1(n55), .B2(n141), .Z(n50) );
  XNR2D1 U87 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n72) );
  ND2D1 U88 ( .A1(ReadCmd), .A2(n35), .ZN(n109) );
  OAI21D1 U89 ( .A1(n144), .A2(n143), .B(n98), .ZN(n58) );
  OAI32D1 U90 ( .A1(n37), .A2(n176), .A3(ReadReq), .B1(n38), .B2(n115), .ZN(
        n128) );
  ND2D1 U91 ( .A1(WriteCmd), .A2(n37), .ZN(n112) );
  NR2D1 U92 ( .A1(WriteAddr[2]), .A2(n141), .ZN(n69) );
  OAI22D0 U93 ( .A1(n143), .A2(n37), .B1(n178), .B2(n112), .ZN(N63) );
  OAI22D0 U94 ( .A1(n141), .A2(n37), .B1(n84), .B2(n112), .ZN(N65) );
  OAI22D0 U95 ( .A1(n142), .A2(n37), .B1(n100), .B2(n112), .ZN(N64) );
  OAI31D0 U96 ( .A1(n35), .A2(WriteReq), .A3(n176), .B(n36), .ZN(n127) );
  OAI31D0 U97 ( .A1(CurState[0]), .A2(n176), .A3(CurState[2]), .B(EmptyFIFO), 
        .ZN(n36) );
  ND3D1 U98 ( .A1(n90), .A2(n45), .A3(WriteReq), .ZN(n87) );
  XNR2D1 U99 ( .A1(n178), .A2(OldWriteAr[0]), .ZN(n90) );
  IND2D1 U100 ( .A1(ReadCmd), .B1(n35), .ZN(N48) );
  XNR2D1 U101 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n111) );
  BUFFD1 U102 ( .I(n178), .Z(WriteAddr[0]) );
  ND2D1 U103 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid3_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockR, ClockW, Dreadyr, \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N87, N99, N161, N194, N227, N260, N293, N326, N359, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(n176), .A2(n175), .A3(n178), .A4(n177), .ZN(n78) );
  XOR4D1 U14 ( .A1(n180), .A2(n179), .A3(n182), .A4(n181), .Z(n77) );
  XOR4D1 U15 ( .A1(n172), .A2(n171), .A3(n174), .A4(n173), .Z(n74) );
  XOR4D1 U16 ( .A1(n165), .A2(n164), .A3(n167), .A4(n166), .Z(n71) );
  XNR4D1 U17 ( .A1(n158), .A2(n157), .A3(n160), .A4(n159), .ZN(n68) );
  XOR4D1 U21 ( .A1(n83), .A2(N74), .A3(n84), .A4(N77), .Z(n82) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n84) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n90) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n89) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n86) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n80) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n174), .E(n225), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n173), .E(n226), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n168), .E(n226), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n167), .E(n226), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n166), .E(n226), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n165), .E(n226), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n164), .E(n226), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n163), .E(n227), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n162), .E(n227), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n161), .E(n227), .CP(n275), .CDN(n321), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n160), .E(n227), .CP(n275), .CDN(n320), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n159), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n158), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n157), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n156), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n155), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n154), .E(n227), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n153), .E(n228), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n152), .E(n228), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n151), .E(n228), .CP(n276), .CDN(n320), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n174), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n173), .E(n242), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n168), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n167), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n166), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n165), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n164), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n163), .E(n243), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n162), .E(n243), .CP(n283), .CDN(n315), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n161), .E(n243), .CP(n283), .CDN(n315), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n160), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n159), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n158), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n157), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n156), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n155), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n154), .E(n243), .CP(n283), .CDN(n314), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n153), .E(n244), .CP(n284), .CDN(n314), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n152), .E(n244), .CP(n284), .CDN(n314), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n151), .E(n244), .CP(n284), .CDN(n314), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n174), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n173), .E(n194), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n168), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n167), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n166), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n165), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n164), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n163), .E(n195), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n162), .E(n195), .CP(n261), .CDN(n333), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n161), .E(n195), .CP(n261), .CDN(n333), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n160), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n159), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n158), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n157), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n156), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n155), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n154), .E(n195), .CP(n261), .CDN(n332), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n153), .E(n196), .CP(n262), .CDN(n332), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n152), .E(n196), .CP(n262), .CDN(n332), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n151), .E(n196), .CP(n262), .CDN(n332), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n174), .E(n201), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n173), .E(n202), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n168), .E(n202), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n167), .E(n202), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n166), .E(n202), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n165), .E(n202), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n164), .E(n202), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n163), .E(n203), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n162), .E(n203), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n161), .E(n203), .CP(n264), .CDN(n330), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n160), .E(n203), .CP(n264), .CDN(n329), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n159), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n158), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n157), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n156), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n155), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n154), .E(n203), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n153), .E(n204), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n152), .E(n204), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n151), .E(n204), .CP(n265), .CDN(n329), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n174), .E(n209), .CP(n267), .CDN(n328), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n173), .E(n210), .CP(n267), .CDN(n328), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n168), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n167), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n166), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n165), .E(n210), .CP(n268), .CDN(n327), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n164), .E(n210), .CP(n268), .CDN(n327), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n163), .E(n211), .CP(n268), .CDN(n327), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n162), .E(n211), .CP(n268), .CDN(n327), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n161), .E(n211), .CP(n268), .CDN(n327), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n160), .E(n211), .CP(n268), .CDN(n326), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n159), .E(n211), .CP(n268), .CDN(n326), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n158), .E(n211), .CP(n268), .CDN(n326), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n157), .E(n211), .CP(n268), .CDN(n326), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n156), .E(n211), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n155), .E(n211), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n154), .E(n211), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n153), .E(n212), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n152), .E(n212), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n151), .E(n212), .CP(n269), .CDN(n326), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n174), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n173), .E(n218), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n168), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n167), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n166), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n165), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n164), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n163), .E(n219), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n162), .E(n219), .CP(n272), .CDN(n324), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n161), .E(n219), .CP(n272), .CDN(n324), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n160), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n159), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n158), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n157), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n156), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n155), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n154), .E(n219), .CP(n272), .CDN(n323), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n153), .E(n220), .CP(n273), .CDN(n323), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n152), .E(n220), .CP(n273), .CDN(n323), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n151), .E(n220), .CP(n273), .CDN(n323), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n174), .E(n233), .CP(n278), .CDN(n319), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n173), .E(n234), .CP(n278), .CDN(n319), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n168), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n167), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n166), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n165), .E(n234), .CP(n279), .CDN(n318), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n164), .E(n234), .CP(n279), .CDN(n318), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n163), .E(n235), .CP(n279), .CDN(n318), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n162), .E(n235), .CP(n279), .CDN(n318), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n161), .E(n235), .CP(n279), .CDN(n318), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n160), .E(n235), .CP(n279), .CDN(n317), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n159), .E(n235), .CP(n279), .CDN(n317), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n158), .E(n235), .CP(n279), .CDN(n317), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n157), .E(n235), .CP(n279), .CDN(n317), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n156), .E(n235), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n155), .E(n235), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n154), .E(n235), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n153), .E(n236), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n152), .E(n236), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n151), .E(n236), .CP(n280), .CDN(n317), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n174), .E(n185), .CP(n256), .CDN(n337), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n173), .E(n186), .CP(n256), .CDN(n337), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n168), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n167), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n166), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n165), .E(n186), .CP(n257), .CDN(n336), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n164), .E(n186), .CP(n257), .CDN(n336), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n163), .E(n187), .CP(n257), .CDN(n336), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n162), .E(n187), .CP(n257), .CDN(n336), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n161), .E(n187), .CP(n257), .CDN(n336), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n160), .E(n187), .CP(n257), .CDN(n335), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n159), .E(n187), .CP(n257), .CDN(n335), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n158), .E(n187), .CP(n257), .CDN(n335), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n157), .E(n187), .CP(n257), .CDN(n335), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n156), .E(n187), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n155), .E(n187), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n154), .E(n187), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n153), .E(n188), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n152), .E(n188), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n151), .E(n188), .CP(n258), .CDN(n335), 
        .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n1), .CP(n305), .CDN(n314), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N87), .E(n225), .CP(n273), .CDN(n323), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n182), .E(n225), .CP(n273), .CDN(n322), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n181), .E(n225), .CP(n273), .CDN(n322), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n180), .E(n225), .CP(n273), .CDN(n322), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n179), .E(n225), .CP(n273), .CDN(n322), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n178), .E(n225), .CP(n273), .CDN(n322), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n177), .E(n225), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n176), .E(n225), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n175), .E(n225), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n172), .E(n226), .CP(n274), .CDN(n322), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n171), .E(n226), .CP(n274), .CDN(n321), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n170), .E(n226), .CP(n274), .CDN(n321), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n169), .E(n226), .CP(n274), .CDN(n321), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N87), .E(n241), .CP(n280), .CDN(n317), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n182), .E(n241), .CP(n280), .CDN(n316), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n181), .E(n241), .CP(n280), .CDN(n316), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n180), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n179), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n178), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n177), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n176), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n175), .E(n241), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n172), .E(n242), .CP(n281), .CDN(n316), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n171), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n170), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n169), .E(n242), .CP(n282), .CDN(n315), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N87), .E(n193), .CP(n258), .CDN(n335), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n182), .E(n193), .CP(n258), .CDN(n334), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n181), .E(n193), .CP(n258), .CDN(n334), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n180), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n179), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n178), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n177), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n176), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n175), .E(n193), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n172), .E(n194), .CP(n259), .CDN(n334), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n171), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n170), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n169), .E(n194), .CP(n260), .CDN(n333), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N87), .E(n201), .CP(n262), .CDN(n332), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n182), .E(n201), .CP(n262), .CDN(n331), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n181), .E(n201), .CP(n262), .CDN(n331), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n180), .E(n201), .CP(n262), .CDN(n331), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n179), .E(n201), .CP(n262), .CDN(n331), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n178), .E(n201), .CP(n262), .CDN(n331), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n177), .E(n201), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n176), .E(n201), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n175), .E(n201), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n172), .E(n202), .CP(n263), .CDN(n331), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n171), .E(n202), .CP(n263), .CDN(n330), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n170), .E(n202), .CP(n263), .CDN(n330), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n169), .E(n202), .CP(n263), .CDN(n330), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N87), .E(n209), .CP(n266), .CDN(n329), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n182), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n181), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n180), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n179), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n178), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n177), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n176), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n175), .E(n209), .CP(n266), .CDN(n328), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n172), .E(n210), .CP(n267), .CDN(n328), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n171), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n170), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n169), .E(n210), .CP(n267), .CDN(n327), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N87), .E(n217), .CP(n269), .CDN(n326), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n182), .E(n217), .CP(n269), .CDN(n325), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n181), .E(n217), .CP(n269), .CDN(n325), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n180), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n179), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n178), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n177), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n176), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n175), .E(n217), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n172), .E(n218), .CP(n270), .CDN(n325), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n171), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n170), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n169), .E(n218), .CP(n271), .CDN(n324), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N87), .E(n233), .CP(n277), .CDN(n320), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n182), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n181), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n180), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n179), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n178), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n177), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n176), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n175), .E(n233), .CP(n277), .CDN(n319), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n172), .E(n234), .CP(n278), .CDN(n319), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n171), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n170), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n169), .E(n234), .CP(n278), .CDN(n318), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N87), .E(n185), .CP(n255), .CDN(n338), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n182), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n181), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n180), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n179), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n178), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n177), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n176), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n175), .E(n185), .CP(n255), .CDN(n337), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n172), .E(n186), .CP(n256), .CDN(n337), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n171), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n170), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n169), .E(n186), .CP(n256), .CDN(n336), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N53), .E(n309), .CP(n302), .CDN(n341), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N54), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N55), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N56), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N57), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N58), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N59), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N60), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N61), .E(n309), .CP(n302), .CDN(n340), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N62), .E(n309), .CP(n303), .CDN(n340), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N63), .E(n309), .CP(n303), .CDN(n340), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N64), .E(n309), .CP(n303), .CDN(n340), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N65), .E(n309), .CP(n303), .CDN(n339), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N66), .E(n309), .CP(n303), .CDN(n339), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N67), .E(n309), .CP(n303), .CDN(n339), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N68), .E(n309), .CP(n303), .CDN(n339), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N69), .E(n309), .CP(n303), .CDN(n339), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N70), .E(n308), .CP(n303), .CDN(n339), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N71), .E(n308), .CP(n304), .CDN(n339), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N72), .E(n308), .CP(n304), .CDN(n339), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N73), .E(n308), .CP(n304), .CDN(n339), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N74), .E(n308), .CP(n304), .CDN(n339), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N75), .E(n308), .CP(n304), .CDN(n339), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N76), .E(n308), .CP(n304), .CDN(n338), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N77), .E(n308), .CP(n304), .CDN(n338), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N78), .E(n308), .CP(n304), .CDN(n338), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N79), .E(n308), .CP(n304), .CDN(n338), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N80), .E(n308), .CP(n305), .CDN(n338), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N81), .E(n308), .CP(n305), .CDN(n338), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N82), .E(n308), .CP(n305), .CDN(n338), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N83), .E(n308), .CP(n305), .CDN(n338), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N84), .E(n308), .CP(n305), .CDN(n338), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N85), .E(n308), .CP(n305), .CDN(n338), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKAN2D0 U3 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U4 ( .I(n313), .ZN(n129) );
  BUFFD1 U5 ( .I(n352), .Z(n320) );
  BUFFD1 U6 ( .I(n352), .Z(n321) );
  BUFFD1 U7 ( .I(n351), .Z(n322) );
  BUFFD1 U8 ( .I(n351), .Z(n323) );
  BUFFD1 U9 ( .I(n350), .Z(n324) );
  BUFFD1 U10 ( .I(n350), .Z(n325) );
  BUFFD1 U11 ( .I(n349), .Z(n326) );
  BUFFD1 U12 ( .I(n349), .Z(n327) );
  BUFFD1 U18 ( .I(n348), .Z(n328) );
  BUFFD1 U19 ( .I(n348), .Z(n329) );
  BUFFD1 U20 ( .I(n347), .Z(n330) );
  BUFFD1 U23 ( .I(n347), .Z(n331) );
  BUFFD1 U24 ( .I(n346), .Z(n332) );
  BUFFD1 U25 ( .I(n346), .Z(n333) );
  BUFFD1 U26 ( .I(n345), .Z(n334) );
  BUFFD1 U31 ( .I(n345), .Z(n335) );
  BUFFD1 U32 ( .I(n344), .Z(n336) );
  BUFFD1 U33 ( .I(n344), .Z(n337) );
  BUFFD1 U34 ( .I(n343), .Z(n338) );
  BUFFD1 U35 ( .I(n343), .Z(n339) );
  BUFFD1 U36 ( .I(n342), .Z(n340) );
  BUFFD1 U37 ( .I(n342), .Z(n341) );
  BUFFD1 U38 ( .I(n355), .Z(n314) );
  BUFFD1 U39 ( .I(n355), .Z(n315) );
  BUFFD1 U40 ( .I(n354), .Z(n316) );
  BUFFD1 U41 ( .I(n354), .Z(n317) );
  BUFFD1 U42 ( .I(n353), .Z(n318) );
  BUFFD1 U43 ( .I(n353), .Z(n319) );
  BUFFD1 U44 ( .I(n357), .Z(n352) );
  BUFFD1 U45 ( .I(n357), .Z(n351) );
  BUFFD1 U46 ( .I(n357), .Z(n350) );
  BUFFD1 U47 ( .I(n358), .Z(n349) );
  BUFFD1 U48 ( .I(n358), .Z(n348) );
  BUFFD1 U49 ( .I(n358), .Z(n347) );
  BUFFD1 U50 ( .I(n359), .Z(n346) );
  BUFFD1 U51 ( .I(n359), .Z(n345) );
  BUFFD1 U52 ( .I(n359), .Z(n344) );
  BUFFD1 U53 ( .I(n360), .Z(n343) );
  BUFFD1 U54 ( .I(n360), .Z(n342) );
  BUFFD1 U55 ( .I(n356), .Z(n354) );
  BUFFD1 U56 ( .I(n356), .Z(n353) );
  BUFFD1 U57 ( .I(n356), .Z(n355) );
  BUFFD1 U58 ( .I(n362), .Z(n357) );
  BUFFD1 U59 ( .I(n362), .Z(n358) );
  BUFFD1 U60 ( .I(n361), .Z(n359) );
  BUFFD1 U61 ( .I(n361), .Z(n360) );
  BUFFD1 U62 ( .I(n363), .Z(n356) );
  INVD1 U63 ( .I(n364), .ZN(n363) );
  INVD1 U64 ( .I(n364), .ZN(n362) );
  INVD1 U65 ( .I(n364), .ZN(n361) );
  INVD1 U66 ( .I(n365), .ZN(n364) );
  INVD1 U67 ( .I(Reset), .ZN(n365) );
  BUFFD1 U68 ( .I(n288), .Z(n278) );
  BUFFD1 U69 ( .I(n288), .Z(n277) );
  BUFFD1 U70 ( .I(n289), .Z(n276) );
  BUFFD1 U71 ( .I(n289), .Z(n275) );
  BUFFD1 U72 ( .I(n290), .Z(n274) );
  BUFFD1 U73 ( .I(n290), .Z(n273) );
  BUFFD1 U74 ( .I(n291), .Z(n272) );
  BUFFD1 U75 ( .I(n291), .Z(n271) );
  BUFFD1 U76 ( .I(n292), .Z(n270) );
  BUFFD1 U77 ( .I(n292), .Z(n269) );
  BUFFD1 U78 ( .I(n293), .Z(n268) );
  BUFFD1 U79 ( .I(n293), .Z(n267) );
  BUFFD1 U80 ( .I(n294), .Z(n266) );
  BUFFD1 U81 ( .I(n294), .Z(n265) );
  BUFFD1 U82 ( .I(n295), .Z(n264) );
  BUFFD1 U83 ( .I(n295), .Z(n263) );
  BUFFD1 U84 ( .I(n296), .Z(n262) );
  BUFFD1 U85 ( .I(n296), .Z(n261) );
  BUFFD1 U86 ( .I(n297), .Z(n260) );
  BUFFD1 U87 ( .I(n297), .Z(n259) );
  BUFFD1 U88 ( .I(n298), .Z(n258) );
  BUFFD1 U89 ( .I(n298), .Z(n257) );
  BUFFD1 U90 ( .I(n299), .Z(n256) );
  BUFFD1 U91 ( .I(n299), .Z(n255) );
  INVD1 U92 ( .I(n229), .ZN(n227) );
  INVD1 U93 ( .I(n230), .ZN(n226) );
  INVD1 U94 ( .I(n230), .ZN(n225) );
  INVD1 U95 ( .I(n221), .ZN(n219) );
  INVD1 U96 ( .I(n222), .ZN(n218) );
  INVD1 U97 ( .I(n222), .ZN(n217) );
  INVD1 U98 ( .I(n197), .ZN(n195) );
  INVD1 U99 ( .I(n198), .ZN(n194) );
  INVD1 U100 ( .I(n198), .ZN(n193) );
  INVD1 U101 ( .I(n189), .ZN(n187) );
  INVD1 U102 ( .I(n190), .ZN(n186) );
  INVD1 U103 ( .I(n190), .ZN(n185) );
  INVD1 U104 ( .I(n229), .ZN(n228) );
  INVD1 U105 ( .I(n221), .ZN(n220) );
  INVD1 U106 ( .I(n197), .ZN(n196) );
  INVD1 U107 ( .I(n189), .ZN(n188) );
  BUFFD1 U108 ( .I(n285), .Z(n283) );
  BUFFD1 U109 ( .I(n286), .Z(n282) );
  BUFFD1 U110 ( .I(n286), .Z(n281) );
  BUFFD1 U111 ( .I(n287), .Z(n280) );
  BUFFD1 U112 ( .I(n287), .Z(n279) );
  BUFFD1 U113 ( .I(n248), .Z(n288) );
  BUFFD1 U114 ( .I(n248), .Z(n289) );
  BUFFD1 U115 ( .I(n248), .Z(n290) );
  BUFFD1 U116 ( .I(n249), .Z(n291) );
  BUFFD1 U117 ( .I(n249), .Z(n292) );
  BUFFD1 U118 ( .I(n249), .Z(n293) );
  BUFFD1 U119 ( .I(n250), .Z(n294) );
  BUFFD1 U120 ( .I(n250), .Z(n295) );
  BUFFD1 U121 ( .I(n250), .Z(n296) );
  BUFFD1 U122 ( .I(n251), .Z(n297) );
  BUFFD1 U123 ( .I(n251), .Z(n298) );
  BUFFD1 U124 ( .I(n251), .Z(n299) );
  BUFFD1 U125 ( .I(n285), .Z(n284) );
  BUFFD1 U126 ( .I(n142), .Z(n147) );
  BUFFD1 U127 ( .I(n143), .Z(n146) );
  BUFFD1 U128 ( .I(n143), .Z(n145) );
  BUFFD1 U129 ( .I(n142), .Z(n148) );
  BUFFD1 U130 ( .I(n142), .Z(n149) );
  BUFFD1 U131 ( .I(n140), .Z(n138) );
  BUFFD1 U132 ( .I(n140), .Z(n137) );
  BUFFD1 U133 ( .I(n140), .Z(n136) );
  BUFFD1 U134 ( .I(n139), .Z(n135) );
  BUFFD1 U135 ( .I(n139), .Z(n134) );
  BUFFD1 U136 ( .I(n143), .Z(n144) );
  BUFFD1 U137 ( .I(n139), .Z(n133) );
  INVD1 U138 ( .I(n215), .ZN(n221) );
  INVD1 U139 ( .I(n215), .ZN(n222) );
  INVD1 U140 ( .I(n191), .ZN(n197) );
  INVD1 U141 ( .I(n191), .ZN(n198) );
  INVD1 U142 ( .I(n183), .ZN(n189) );
  INVD1 U143 ( .I(n183), .ZN(n190) );
  INVD1 U144 ( .I(n223), .ZN(n229) );
  INVD1 U145 ( .I(n223), .ZN(n230) );
  INVD1 U146 ( .I(n245), .ZN(n243) );
  INVD1 U147 ( .I(n246), .ZN(n242) );
  INVD1 U148 ( .I(n246), .ZN(n241) );
  INVD1 U149 ( .I(n237), .ZN(n235) );
  INVD1 U150 ( .I(n238), .ZN(n234) );
  INVD1 U151 ( .I(n238), .ZN(n233) );
  INVD1 U152 ( .I(n213), .ZN(n211) );
  INVD1 U153 ( .I(n214), .ZN(n210) );
  INVD1 U154 ( .I(n214), .ZN(n209) );
  INVD1 U155 ( .I(n205), .ZN(n203) );
  INVD1 U156 ( .I(n206), .ZN(n202) );
  INVD1 U157 ( .I(n206), .ZN(n201) );
  INVD1 U158 ( .I(n245), .ZN(n244) );
  INVD1 U159 ( .I(n237), .ZN(n236) );
  INVD1 U160 ( .I(n213), .ZN(n212) );
  INVD1 U161 ( .I(n205), .ZN(n204) );
  BUFFD1 U162 ( .I(n247), .Z(n285) );
  BUFFD1 U163 ( .I(n247), .Z(n286) );
  BUFFD1 U164 ( .I(n247), .Z(n287) );
  BUFFD1 U165 ( .I(n253), .Z(n248) );
  BUFFD1 U166 ( .I(n253), .Z(n249) );
  BUFFD1 U167 ( .I(n252), .Z(n250) );
  BUFFD1 U168 ( .I(n252), .Z(n251) );
  INVD1 U169 ( .I(n306), .ZN(n304) );
  INVD1 U170 ( .I(n307), .ZN(n303) );
  INVD1 U171 ( .I(n307), .ZN(n302) );
  INVD1 U172 ( .I(n306), .ZN(n305) );
  XOR3D1 U173 ( .A1(n170), .A2(n169), .A3(n76), .Z(n75) );
  XOR3D1 U174 ( .A1(n77), .A2(n168), .A3(n78), .Z(n76) );
  XOR3D1 U175 ( .A1(n71), .A2(n154), .A3(n72), .Z(n70) );
  XOR3D1 U176 ( .A1(n163), .A2(n162), .A3(n73), .Z(n72) );
  XOR3D1 U177 ( .A1(n74), .A2(n161), .A3(n75), .Z(n73) );
  XOR3D1 U178 ( .A1(n153), .A2(n152), .A3(n67), .Z(N87) );
  XOR3D1 U179 ( .A1(n151), .A2(n68), .A3(n69), .Z(n67) );
  XOR3D1 U180 ( .A1(n156), .A2(n155), .A3(n70), .Z(n69) );
  XOR3D1 U181 ( .A1(N69), .A2(N68), .A3(n85), .Z(n83) );
  XOR3D1 U182 ( .A1(N67), .A2(n86), .A3(n87), .Z(n85) );
  BUFFD1 U183 ( .I(n141), .Z(n150) );
  BUFFD1 U184 ( .I(n311), .Z(n141) );
  XOR3D1 U185 ( .A1(N62), .A2(N61), .A3(n88), .Z(n87) );
  XOR3D1 U186 ( .A1(n89), .A2(N60), .A3(n90), .Z(n88) );
  XOR3D1 U187 ( .A1(N81), .A2(N76), .A3(n79), .Z(N85) );
  XOR3D1 U188 ( .A1(N75), .A2(n80), .A3(n81), .Z(n79) );
  XOR3D1 U189 ( .A1(N79), .A2(N78), .A3(n82), .Z(n81) );
  BUFFD1 U190 ( .I(n311), .Z(n142) );
  BUFFD1 U191 ( .I(n312), .Z(n140) );
  BUFFD1 U192 ( .I(n311), .Z(n143) );
  BUFFD1 U193 ( .I(n312), .Z(n139) );
  INVD1 U194 ( .I(n129), .ZN(n131) );
  INVD1 U195 ( .I(n129), .ZN(n132) );
  INVD1 U196 ( .I(n129), .ZN(n130) );
  INVD1 U197 ( .I(AddrW[0]), .ZN(n93) );
  INVD1 U198 ( .I(n239), .ZN(n245) );
  INVD1 U199 ( .I(n239), .ZN(n246) );
  INVD1 U200 ( .I(n231), .ZN(n237) );
  INVD1 U201 ( .I(n231), .ZN(n238) );
  INVD1 U202 ( .I(n207), .ZN(n213) );
  INVD1 U203 ( .I(n207), .ZN(n214) );
  INVD1 U204 ( .I(n199), .ZN(n205) );
  INVD1 U205 ( .I(n199), .ZN(n206) );
  INVD1 U206 ( .I(n224), .ZN(n223) );
  INVD1 U207 ( .I(N194), .ZN(n224) );
  NR3D0 U208 ( .A1(n91), .A2(AddrW[0]), .A3(n66), .ZN(N194) );
  INVD1 U209 ( .I(n216), .ZN(n215) );
  INVD1 U210 ( .I(N227), .ZN(n216) );
  NR3D0 U211 ( .A1(n91), .A2(n66), .A3(n93), .ZN(N227) );
  INVD1 U212 ( .I(n192), .ZN(n191) );
  INVD1 U213 ( .I(N326), .ZN(n192) );
  NR3D0 U214 ( .A1(n91), .A2(AddrW[0]), .A3(n92), .ZN(N326) );
  INVD1 U215 ( .I(n184), .ZN(n183) );
  INVD1 U216 ( .I(N359), .ZN(n184) );
  NR3D0 U217 ( .A1(n91), .A2(n92), .A3(n93), .ZN(N359) );
  INVD1 U218 ( .I(n310), .ZN(n308) );
  INVD1 U219 ( .I(n310), .ZN(n309) );
  INVD1 U220 ( .I(n300), .ZN(n307) );
  INVD1 U221 ( .I(n300), .ZN(n306) );
  BUFFD1 U222 ( .I(ClockW), .Z(n253) );
  BUFFD1 U223 ( .I(ClockW), .Z(n252) );
  BUFFD1 U224 ( .I(n254), .Z(n247) );
  BUFFD1 U225 ( .I(ClockW), .Z(n254) );
  BUFFD1 U226 ( .I(DataI[7]), .Z(n158) );
  BUFFD1 U227 ( .I(DataI[8]), .Z(n159) );
  BUFFD1 U228 ( .I(DataI[14]), .Z(n165) );
  BUFFD1 U229 ( .I(DataI[15]), .Z(n166) );
  BUFFD1 U230 ( .I(DataI[21]), .Z(n172) );
  BUFFD1 U231 ( .I(DataI[22]), .Z(n173) );
  BUFFD1 U232 ( .I(DataI[25]), .Z(n176) );
  BUFFD1 U233 ( .I(DataI[26]), .Z(n177) );
  BUFFD1 U234 ( .I(DataI[29]), .Z(n180) );
  BUFFD1 U235 ( .I(DataI[30]), .Z(n181) );
  BUFFD1 U236 ( .I(DataI[3]), .Z(n154) );
  BUFFD1 U237 ( .I(DataI[4]), .Z(n155) );
  BUFFD1 U238 ( .I(DataI[10]), .Z(n161) );
  BUFFD1 U239 ( .I(DataI[11]), .Z(n162) );
  BUFFD1 U240 ( .I(DataI[17]), .Z(n168) );
  BUFFD1 U241 ( .I(DataI[18]), .Z(n169) );
  BUFFD1 U242 ( .I(DataI[6]), .Z(n157) );
  BUFFD1 U243 ( .I(DataI[9]), .Z(n160) );
  BUFFD1 U244 ( .I(DataI[13]), .Z(n164) );
  BUFFD1 U245 ( .I(DataI[16]), .Z(n167) );
  BUFFD1 U246 ( .I(DataI[20]), .Z(n171) );
  BUFFD1 U247 ( .I(DataI[23]), .Z(n174) );
  BUFFD1 U248 ( .I(DataI[24]), .Z(n175) );
  BUFFD1 U249 ( .I(DataI[27]), .Z(n178) );
  BUFFD1 U250 ( .I(DataI[28]), .Z(n179) );
  BUFFD1 U251 ( .I(DataI[31]), .Z(n182) );
  BUFFD1 U252 ( .I(DataI[0]), .Z(n151) );
  BUFFD1 U253 ( .I(DataI[5]), .Z(n156) );
  BUFFD1 U254 ( .I(DataI[12]), .Z(n163) );
  BUFFD1 U255 ( .I(DataI[19]), .Z(n170) );
  BUFFD1 U256 ( .I(DataI[1]), .Z(n152) );
  BUFFD1 U257 ( .I(DataI[2]), .Z(n153) );
  MUX4ND0 U258 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n150), .S1(n136), .ZN(n7)
         );
  MUX4ND0 U259 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n150), .S1(n136), .ZN(n10)
         );
  MUX4ND0 U260 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n150), .S1(n135), .ZN(n25)
         );
  MUX4ND0 U261 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n148), .S1(n135), .ZN(
        n40) );
  MUX4ND0 U262 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n149), .S1(n135), .ZN(
        n43) );
  MUX4ND0 U263 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n149), .S1(n134), .ZN(
        n61) );
  MUX4ND0 U264 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n148), .S1(n134), .ZN(
        n64) );
  MUX4ND0 U265 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n149), .S1(n134), .ZN(
        n110) );
  MUX4ND0 U266 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n150), .S1(n134), .ZN(
        n113) );
  MUX4ND0 U267 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n150), .S1(n134), .ZN(
        n122) );
  MUX4ND0 U268 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n150), .S1(n134), .ZN(
        n125) );
  MUX4ND0 U269 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n148), .S1(n135), .ZN(n22)
         );
  MUX4ND0 U270 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n149), .S1(n135), .ZN(n28)
         );
  MUX4ND0 U271 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n148), .S1(n135), .ZN(
        n52) );
  MUX4ND0 U272 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n149), .S1(n134), .ZN(
        n101) );
  MUX4ND0 U273 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n150), .S1(n134), .ZN(
        n104) );
  MUX4ND0 U274 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n150), .S1(n136), .ZN(n4)
         );
  MUX4ND0 U275 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n149), .S1(n136), .ZN(n16)
         );
  MUX4ND0 U276 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n148), .S1(n135), .ZN(
        n34) );
  MUX4ND0 U277 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n149), .S1(n135), .ZN(
        n37) );
  MUX4ND0 U278 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n148), .S1(n135), .ZN(
        n46) );
  MUX4ND0 U279 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n149), .S1(n135), .ZN(
        n58) );
  MUX4ND0 U280 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n149), .S1(n134), .ZN(
        n95) );
  MUX4ND0 U281 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n149), .S1(n134), .ZN(
        n107) );
  MUX4ND0 U282 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n150), .S1(n134), .ZN(
        n116) );
  MUX4ND0 U283 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n150), .S1(n134), .ZN(
        n119) );
  MUX4ND0 U284 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n150), .S1(n136), .ZN(n13)
         );
  MUX4ND0 U285 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n149), .S1(n136), .ZN(n19)
         );
  MUX4ND0 U286 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n148), .S1(n135), .ZN(n31)
         );
  MUX4ND0 U287 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n148), .S1(n135), .ZN(
        n49) );
  MUX4ND0 U288 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n149), .S1(n135), .ZN(
        n55) );
  MUX4ND0 U289 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n148), .S1(n134), .ZN(
        n98) );
  MUX4ND0 U290 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n150), .S1(n133), .ZN(
        n128) );
  BUFFD1 U291 ( .I(N50), .Z(n313) );
  BUFFD1 U292 ( .I(N48), .Z(n311) );
  BUFFD1 U293 ( .I(N49), .Z(n312) );
  INVD1 U294 ( .I(n240), .ZN(n239) );
  INVD1 U295 ( .I(N99), .ZN(n240) );
  NR3D0 U296 ( .A1(n66), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N99) );
  INVD1 U297 ( .I(AddrW[1]), .ZN(n91) );
  ND2D1 U298 ( .A1(AddrW[2]), .A2(Write), .ZN(n92) );
  IND2D1 U299 ( .A1(AddrW[2]), .B1(Write), .ZN(n66) );
  INVD1 U300 ( .I(n208), .ZN(n207) );
  INVD1 U301 ( .I(N260), .ZN(n208) );
  NR3D0 U302 ( .A1(n92), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N260) );
  INVD1 U303 ( .I(n232), .ZN(n231) );
  INVD1 U304 ( .I(N161), .ZN(n232) );
  NR3D0 U305 ( .A1(n93), .A2(AddrW[1]), .A3(n66), .ZN(N161) );
  INVD1 U306 ( .I(n200), .ZN(n199) );
  INVD1 U307 ( .I(N293), .ZN(n200) );
  NR3D0 U308 ( .A1(n93), .A2(AddrW[1]), .A3(n92), .ZN(N293) );
  INVD1 U309 ( .I(Read), .ZN(n310) );
  OR2D1 U310 ( .A1(n308), .A2(Dreadyr), .Z(n1) );
  CKAN2D0 U311 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  INVD1 U312 ( .I(n301), .ZN(n300) );
  INVD1 U313 ( .I(ClockR), .ZN(n301) );
  CKAN2D0 U314 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U315 ( .I0(n2), .I1(n3), .I2(n4), .S0(n138), .S1(n130), .ZN(N84) );
  MUX3ND0 U316 ( .I0(n5), .I1(n6), .I2(n7), .S0(n138), .S1(n130), .ZN(N83) );
  MUX3ND0 U317 ( .I0(n8), .I1(n9), .I2(n10), .S0(n138), .S1(n130), .ZN(N82) );
  MUX3ND0 U318 ( .I0(n11), .I1(n12), .I2(n13), .S0(n138), .S1(n130), .ZN(N81)
         );
  MUX3ND0 U319 ( .I0(n14), .I1(n15), .I2(n16), .S0(n138), .S1(n130), .ZN(N80)
         );
  MUX3ND0 U320 ( .I0(n17), .I1(n18), .I2(n19), .S0(n138), .S1(n130), .ZN(N79)
         );
  MUX3ND0 U321 ( .I0(n20), .I1(n21), .I2(n22), .S0(n138), .S1(n130), .ZN(N78)
         );
  MUX3ND0 U322 ( .I0(n23), .I1(n24), .I2(n25), .S0(n138), .S1(n131), .ZN(N77)
         );
  MUX3ND0 U323 ( .I0(n26), .I1(n27), .I2(n28), .S0(n138), .S1(n131), .ZN(N76)
         );
  MUX3ND0 U324 ( .I0(n29), .I1(n30), .I2(n31), .S0(n138), .S1(n131), .ZN(N75)
         );
  MUX3ND0 U325 ( .I0(n32), .I1(n33), .I2(n34), .S0(n138), .S1(n131), .ZN(N74)
         );
  MUX3ND0 U326 ( .I0(n35), .I1(n36), .I2(n37), .S0(n138), .S1(n131), .ZN(N73)
         );
  MUX3ND0 U327 ( .I0(n38), .I1(n39), .I2(n40), .S0(n138), .S1(n131), .ZN(N72)
         );
  MUX3ND0 U328 ( .I0(n41), .I1(n42), .I2(n43), .S0(n137), .S1(n131), .ZN(N71)
         );
  MUX3ND0 U329 ( .I0(n44), .I1(n45), .I2(n46), .S0(n137), .S1(n131), .ZN(N70)
         );
  MUX3ND0 U330 ( .I0(n47), .I1(n48), .I2(n49), .S0(n137), .S1(n131), .ZN(N69)
         );
  MUX3ND0 U331 ( .I0(n50), .I1(n51), .I2(n52), .S0(n137), .S1(n131), .ZN(N68)
         );
  MUX3ND0 U332 ( .I0(n53), .I1(n54), .I2(n55), .S0(n137), .S1(n131), .ZN(N67)
         );
  MUX3ND0 U333 ( .I0(n56), .I1(n57), .I2(n58), .S0(n137), .S1(n131), .ZN(N66)
         );
  MUX3ND0 U334 ( .I0(n59), .I1(n60), .I2(n61), .S0(n137), .S1(n131), .ZN(N65)
         );
  MUX3ND0 U335 ( .I0(n62), .I1(n63), .I2(n64), .S0(n137), .S1(n132), .ZN(N64)
         );
  MUX3ND0 U336 ( .I0(n65), .I1(n94), .I2(n95), .S0(n137), .S1(n132), .ZN(N63)
         );
  MUX3ND0 U337 ( .I0(n96), .I1(n97), .I2(n98), .S0(n137), .S1(n132), .ZN(N62)
         );
  MUX3ND0 U338 ( .I0(n99), .I1(n100), .I2(n101), .S0(n137), .S1(n132), .ZN(N61) );
  MUX3ND0 U339 ( .I0(n102), .I1(n103), .I2(n104), .S0(n137), .S1(n132), .ZN(
        N60) );
  MUX3ND0 U340 ( .I0(n105), .I1(n106), .I2(n107), .S0(n137), .S1(n132), .ZN(
        N59) );
  MUX3ND0 U341 ( .I0(n108), .I1(n109), .I2(n110), .S0(n136), .S1(n132), .ZN(
        N58) );
  MUX3ND0 U342 ( .I0(n111), .I1(n112), .I2(n113), .S0(n136), .S1(n132), .ZN(
        N57) );
  MUX3ND0 U343 ( .I0(n114), .I1(n115), .I2(n116), .S0(n136), .S1(n132), .ZN(
        N56) );
  MUX3ND0 U344 ( .I0(n117), .I1(n118), .I2(n119), .S0(n136), .S1(n132), .ZN(
        N55) );
  MUX3ND0 U345 ( .I0(n120), .I1(n121), .I2(n122), .S0(n136), .S1(n132), .ZN(
        N54) );
  MUX3ND0 U346 ( .I0(n123), .I1(n124), .I2(n125), .S0(n136), .S1(n132), .ZN(
        N53) );
  MUX3ND0 U347 ( .I0(n126), .I1(n127), .I2(n128), .S0(n136), .S1(n132), .ZN(
        N52) );
  MUX2ND0 U348 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n147), .ZN(n3)
         );
  MUX2ND0 U349 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n147), .ZN(n2)
         );
  MUX2ND0 U350 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(n146), .ZN(n6)
         );
  MUX2ND0 U351 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n147), .ZN(n5)
         );
  MUX2ND0 U352 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n148), .ZN(n9)
         );
  MUX2ND0 U353 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n147), .ZN(n8)
         );
  MUX2ND0 U354 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n148), .ZN(n12) );
  MUX2ND0 U355 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n148), .ZN(n11) );
  MUX2ND0 U356 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n147), .ZN(n15) );
  MUX2ND0 U357 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n148), .ZN(n14) );
  MUX2ND0 U358 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n147), .ZN(n18) );
  MUX2ND0 U359 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n147), .ZN(n17) );
  MUX2ND0 U360 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n148), .ZN(n21) );
  MUX2ND0 U361 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n147), .ZN(n20) );
  MUX2ND0 U362 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n147), .ZN(n24) );
  MUX2ND0 U363 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n147), .ZN(n23) );
  MUX2ND0 U364 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n147), .ZN(n27) );
  MUX2ND0 U365 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n147), .ZN(n26) );
  MUX2ND0 U366 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n147), .ZN(n30) );
  MUX2ND0 U367 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n147), .ZN(n29) );
  MUX2ND0 U368 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n147), .ZN(
        n33) );
  MUX2ND0 U369 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n147), .ZN(
        n32) );
  MUX2ND0 U370 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n147), .ZN(
        n36) );
  MUX2ND0 U371 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n147), .ZN(
        n35) );
  MUX2ND0 U372 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n147), .ZN(
        n39) );
  MUX2ND0 U373 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n146), .ZN(
        n38) );
  MUX2ND0 U374 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(n146), .ZN(
        n42) );
  MUX2ND0 U375 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n146), .ZN(
        n41) );
  MUX2ND0 U376 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(n146), .ZN(
        n45) );
  MUX2ND0 U377 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n146), .ZN(
        n44) );
  MUX2ND0 U378 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(n146), .ZN(
        n48) );
  MUX2ND0 U379 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(n146), .ZN(
        n47) );
  MUX2ND0 U380 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(n146), .ZN(
        n51) );
  MUX2ND0 U381 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(n146), .ZN(
        n50) );
  MUX2ND0 U382 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n146), .ZN(
        n54) );
  MUX2ND0 U383 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n146), .ZN(
        n53) );
  MUX2ND0 U384 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n146), .ZN(
        n57) );
  MUX2ND0 U385 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n146), .ZN(
        n56) );
  MUX2ND0 U386 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(n146), .ZN(
        n60) );
  MUX2ND0 U387 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n146), .ZN(
        n59) );
  MUX2ND0 U388 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n146), .ZN(
        n63) );
  MUX2ND0 U389 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(n146), .ZN(
        n62) );
  MUX2ND0 U390 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(n146), .ZN(
        n94) );
  MUX2ND0 U391 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(n145), .ZN(
        n65) );
  MUX2ND0 U392 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(n145), .ZN(
        n97) );
  MUX2ND0 U393 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(n145), .ZN(
        n96) );
  MUX2ND0 U394 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(n145), .ZN(
        n100) );
  MUX2ND0 U395 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(n145), .ZN(
        n99) );
  MUX2ND0 U396 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n145), .ZN(
        n103) );
  MUX2ND0 U397 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n145), .ZN(
        n102) );
  MUX2ND0 U398 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n145), .ZN(
        n106) );
  MUX2ND0 U399 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n145), .ZN(
        n105) );
  MUX2ND0 U400 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n145), .ZN(
        n109) );
  MUX2ND0 U401 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n145), .ZN(
        n108) );
  MUX2ND0 U402 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n145), .ZN(
        n112) );
  MUX2ND0 U403 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n145), .ZN(
        n111) );
  MUX2ND0 U404 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n145), .ZN(
        n115) );
  MUX2ND0 U405 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n145), .ZN(
        n114) );
  MUX2ND0 U406 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n145), .ZN(
        n118) );
  MUX2ND0 U407 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n145), .ZN(
        n117) );
  MUX2ND0 U408 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(n145), .ZN(
        n121) );
  MUX2ND0 U409 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n145), .ZN(
        n120) );
  MUX2ND0 U410 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(n145), .ZN(
        n124) );
  MUX2ND0 U411 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n144), .ZN(
        n123) );
  MUX2ND0 U412 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n147), .ZN(
        n127) );
  MUX2ND0 U413 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n146), .ZN(
        n126) );
endmodule


module PLLTop_0 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_0 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_0 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_0 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_0 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N47, N48, N49, N50, N51, N67, N68, N69,
         N70, N71, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n90, n92, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n141, n143, n144, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n190, n191,
         n192, n193, n194, n195, n196;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n151), .CPN(StateClock), .Q(FullFIFO) );
  DFND1 EmptyFIFOr_reg ( .D(n147), .CPN(StateClock), .Q(EmptyFIFO), .QN(n132)
         );
  MOAI22D1 U6 ( .A1(n165), .A2(n40), .B1(n40), .B2(OldReadAr[1]), .ZN(n149) );
  OA21D1 U11 ( .A1(n172), .A2(n190), .B(n35), .Z(n44) );
  MOAI22D1 U12 ( .A1(n168), .A2(n45), .B1(n45), .B2(OldWriteAr[2]), .ZN(n152)
         );
  MOAI22D1 U13 ( .A1(n169), .A2(n45), .B1(n45), .B2(OldWriteAr[0]), .ZN(n153)
         );
  MOAI22D1 U14 ( .A1(n45), .A2(n46), .B1(n45), .B2(OldWriteAr[1]), .ZN(n154)
         );
  MOAI22D1 U15 ( .A1(n167), .A2(n45), .B1(n45), .B2(OldWriteAr[3]), .ZN(n155)
         );
  IAO21D1 U31 ( .A1(n73), .A2(n74), .B(n55), .ZN(n72) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n76), .B(n75), .Z(n81) );
  MOAI22D1 U88 ( .A1(n166), .A2(n40), .B1(n40), .B2(OldReadAr[0]), .ZN(n162)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n150), .CPN(StateClock), .CDN(n192), .Q(
        OldReadAr[3]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n148), .CPN(StateClock), .CDN(n192), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n162), .CPN(StateClock), .CDN(n191), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n155), .CPN(StateClock), .CDN(n191), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n154), .CPN(StateClock), .CDN(n192), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n153), .CPN(StateClock), .CDN(n192), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n152), .CPN(StateClock), .CDN(n192), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n149), .CPN(StateClock), .CDN(n192), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n159), .CPN(StateClock), .CDN(n191), .Q(
        NextState[0]), .QN(n144) );
  DFNCND1 \NextState_reg[1]  ( .D(n158), .CPN(StateClock), .CDN(n191), .Q(
        NextState[1]), .QN(n143) );
  DFNCND1 \NextState_reg[2]  ( .D(n156), .CPN(StateClock), .CDN(n191), .Q(
        NextState[2]), .QN(n141) );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n191), 
        .QN(n170) );
  DFNCND1 WriteCmdr_reg ( .D(n157), .CPN(StateClock), .CDN(n191), .Q(WriteCmd)
         );
  DFNCND1 ReadCmdr_reg ( .D(n160), .CPN(StateClock), .CDN(n191), .Q(ReadCmd)
         );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n191), 
        .QN(n171) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n191), 
        .Q(n52), .QN(n172) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N68), .E(N71), .CP(StateClock), .CDN(n193), 
        .Q(WriteAddr[1]), .QN(n46) );
  EDFCND1 \ReadAr_reg[3]  ( .D(N51), .E(N50), .CP(StateClock), .CDN(n193), .Q(
        ReadAddr[3]), .QN(n163) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N50), .CP(StateClock), .CDN(n193), .Q(
        ReadAddr[2]), .QN(n164) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N48), .E(N50), .CP(StateClock), .CDN(n193), .Q(
        ReadAddr[1]), .QN(n165) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N47), .E(N50), .CP(StateClock), .CDN(n193), .Q(
        ReadAddr[0]), .QN(n166) );
  EDFCND1 \WriteAr_reg[3]  ( .D(N70), .E(N71), .CP(StateClock), .CDN(n193), 
        .Q(WriteAddr[3]), .QN(n167) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N69), .E(N71), .CP(StateClock), .CDN(n193), 
        .Q(WriteAddr[2]), .QN(n168) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N67), .E(N71), .CP(StateClock), .CDN(n193), 
        .Q(WriteAddr[0]), .QN(n169) );
  INVD1 U3 ( .I(n195), .ZN(n192) );
  INVD1 U4 ( .I(n194), .ZN(n193) );
  BUFFD1 U5 ( .I(Reset), .Z(n194) );
  BUFFD1 U7 ( .I(Reset), .Z(n195) );
  INVD1 U8 ( .I(n196), .ZN(n191) );
  BUFFD1 U9 ( .I(Reset), .Z(n196) );
  INVD1 U10 ( .I(n48), .ZN(n49) );
  ND2D1 U16 ( .A1(n66), .A2(n42), .ZN(n119) );
  OAI211D1 U17 ( .A1(n35), .A2(n63), .B(n66), .C(n115), .ZN(n48) );
  INR2D1 U18 ( .A1(n71), .B1(n116), .ZN(n115) );
  AOI21D1 U19 ( .A1(n52), .A2(n117), .B(n190), .ZN(n116) );
  MAOI22D0 U20 ( .A1(n69), .A2(n190), .B1(n190), .B2(n71), .ZN(n66) );
  ND2D1 U21 ( .A1(n66), .A2(n35), .ZN(n47) );
  INVD1 U22 ( .I(n106), .ZN(n76) );
  OA211D0 U23 ( .A1(n75), .A2(n76), .B(n77), .C(n78), .Z(n55) );
  INVD1 U24 ( .I(n85), .ZN(n77) );
  NR3D0 U25 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n78) );
  NR3D0 U26 ( .A1(WriteAddr[2]), .A2(n46), .A3(ReadAddr[2]), .ZN(n80) );
  ND2D1 U27 ( .A1(n130), .A2(ReadAddr[2]), .ZN(n129) );
  INVD1 U28 ( .I(n40), .ZN(n38) );
  ND2D1 U29 ( .A1(n107), .A2(n108), .ZN(n85) );
  XNR2D1 U30 ( .A1(ReadAddr[1]), .A2(n46), .ZN(n107) );
  INVD1 U32 ( .I(n90), .ZN(n84) );
  INVD1 U33 ( .I(n97), .ZN(n108) );
  INVD1 U35 ( .I(n53), .ZN(n42) );
  OAI21D1 U36 ( .A1(n130), .A2(ReadAddr[2]), .B(n129), .ZN(n114) );
  ND3D1 U37 ( .A1(n42), .A2(n35), .A3(n56), .ZN(N71) );
  AOI21D1 U38 ( .A1(n76), .A2(n83), .B(ReadAddr[1]), .ZN(n105) );
  ND2D1 U39 ( .A1(n35), .A2(n118), .ZN(N50) );
  NR3D0 U40 ( .A1(n117), .A2(n124), .A3(n125), .ZN(n123) );
  XNR2D1 U41 ( .A1(ReadAddr[3]), .A2(n41), .ZN(n125) );
  XNR2D1 U42 ( .A1(ReadAddr[2]), .A2(n39), .ZN(n124) );
  XNR2D1 U43 ( .A1(n126), .A2(WriteAddr[3]), .ZN(n99) );
  XNR2D1 U44 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n104) );
  NR2D1 U45 ( .A1(n114), .A2(n118), .ZN(N49) );
  NR2D1 U46 ( .A1(n131), .A2(n118), .ZN(N48) );
  XNR2D1 U47 ( .A1(ReadAddr[1]), .A2(ReadAddr[0]), .ZN(n131) );
  NR2D1 U48 ( .A1(n112), .A2(n118), .ZN(N51) );
  NR2D1 U49 ( .A1(ReadAddr[0]), .A2(n118), .ZN(N47) );
  ND2D1 U50 ( .A1(WriteReq), .A2(n47), .ZN(n45) );
  OAI32D1 U51 ( .A1(n35), .A2(WriteReq), .A3(n194), .B1(n36), .B2(n132), .ZN(
        n147) );
  AOI21D1 U52 ( .A1(n37), .A2(n35), .B(n194), .ZN(n36) );
  OAI22D0 U53 ( .A1(n48), .A2(n141), .B1(n49), .B2(n50), .ZN(n156) );
  AOI21D1 U54 ( .A1(n51), .A2(n52), .B(n53), .ZN(n50) );
  OAI22D0 U55 ( .A1(n171), .A2(n54), .B1(n190), .B2(n55), .ZN(n51) );
  OAI22D0 U56 ( .A1(n48), .A2(n143), .B1(n49), .B2(n67), .ZN(n158) );
  AOI31D0 U57 ( .A1(n68), .A2(n69), .A3(n190), .B(n70), .ZN(n67) );
  IOA21D1 U58 ( .A1(n52), .A2(n54), .B(n86), .ZN(n68) );
  OAI31D0 U59 ( .A1(n71), .A2(n190), .A3(n72), .B(n35), .ZN(n70) );
  OAI22D0 U60 ( .A1(n48), .A2(n144), .B1(n49), .B2(n100), .ZN(n159) );
  AOI22D0 U61 ( .A1(n101), .A2(n52), .B1(n102), .B2(n103), .ZN(n100) );
  AOI211D1 U62 ( .A1(n164), .A2(n106), .B(n37), .C(n85), .ZN(n102) );
  AOI221D0 U63 ( .A1(n90), .A2(n76), .B1(n104), .B2(ReadAddr[1]), .C(n105), 
        .ZN(n103) );
  NR3D0 U64 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n60) );
  XNR2D1 U65 ( .A1(n167), .A2(OldWriteAr[3]), .ZN(n62) );
  XNR2D1 U66 ( .A1(n46), .A2(OldWriteAr[1]), .ZN(n61) );
  OAI21D1 U67 ( .A1(n56), .A2(n47), .B(n57), .ZN(n157) );
  ND4D1 U68 ( .A1(n58), .A2(n47), .A3(n59), .A4(n60), .ZN(n57) );
  XNR2D1 U69 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n58) );
  XNR2D1 U70 ( .A1(WriteAddr[2]), .A2(OldWriteAr[2]), .ZN(n59) );
  INVD1 U71 ( .I(WriteReq), .ZN(n63) );
  CKND2D0 U72 ( .A1(ReadReq), .A2(n119), .ZN(n40) );
  ND2D1 U73 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n128) );
  AOI21D1 U74 ( .A1(n128), .A2(n168), .B(n126), .ZN(n98) );
  ND2D1 U75 ( .A1(n171), .A2(n52), .ZN(n71) );
  OAI22D0 U76 ( .A1(n38), .A2(n39), .B1(n164), .B2(n40), .ZN(n148) );
  OAI22D0 U77 ( .A1(n38), .A2(n41), .B1(n163), .B2(n40), .ZN(n150) );
  AOI21D1 U78 ( .A1(n83), .A2(n84), .B(WriteAddr[1]), .ZN(n79) );
  NR2D1 U79 ( .A1(WriteAddr[2]), .A2(n164), .ZN(n90) );
  OAI21D1 U80 ( .A1(n171), .A2(n109), .B(n190), .ZN(n101) );
  NR4D0 U81 ( .A1(n108), .A2(n110), .A3(n95), .A4(n111), .ZN(n109) );
  XNR2D1 U82 ( .A1(WriteAddr[2]), .A2(n114), .ZN(n110) );
  XNR2D1 U83 ( .A1(WriteAddr[3]), .A2(n112), .ZN(n111) );
  ND4D1 U84 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(n54) );
  XNR2D1 U85 ( .A1(n99), .A2(n163), .ZN(n94) );
  XNR2D1 U86 ( .A1(ReadAddr[2]), .A2(n98), .ZN(n96) );
  NR2D1 U87 ( .A1(n128), .A2(n168), .ZN(n126) );
  NR2D1 U89 ( .A1(n46), .A2(n168), .ZN(n75) );
  XNR2D1 U90 ( .A1(ReadAddr[3]), .A2(n167), .ZN(n106) );
  XNR2D1 U91 ( .A1(WriteAddr[0]), .A2(n166), .ZN(n97) );
  XNR2D1 U92 ( .A1(n163), .A2(n129), .ZN(n112) );
  ND2D1 U93 ( .A1(ReadCmd), .A2(n35), .ZN(n118) );
  ND2D1 U94 ( .A1(WriteCmd), .A2(n42), .ZN(n56) );
  OAI211D1 U95 ( .A1(n46), .A2(ReadAddr[1]), .B(n83), .C(n92), .ZN(n74) );
  AOI22D0 U96 ( .A1(n163), .A2(WriteAddr[3]), .B1(n166), .B2(WriteAddr[0]), 
        .ZN(n92) );
  OAI21D1 U97 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n128), .ZN(n113) );
  ND3D1 U98 ( .A1(n171), .A2(n190), .A3(n172), .ZN(n35) );
  OAI211D1 U99 ( .A1(n165), .A2(WriteAddr[1]), .B(n84), .C(n87), .ZN(n73) );
  AOI22D0 U100 ( .A1(n167), .A2(ReadAddr[3]), .B1(n169), .B2(ReadAddr[0]), 
        .ZN(n87) );
  OAI22D0 U101 ( .A1(n165), .A2(n42), .B1(n113), .B2(n56), .ZN(N68) );
  OAI22D0 U102 ( .A1(n163), .A2(n42), .B1(n99), .B2(n56), .ZN(N70) );
  OAI22D0 U103 ( .A1(n164), .A2(n42), .B1(n127), .B2(n56), .ZN(N69) );
  INVD1 U104 ( .I(n98), .ZN(n127) );
  OAI22D0 U105 ( .A1(n166), .A2(n42), .B1(WriteAddr[0]), .B2(n56), .ZN(N67) );
  NR3D0 U106 ( .A1(n171), .A2(n172), .A3(n190), .ZN(n53) );
  ND2D1 U107 ( .A1(n164), .A2(WriteAddr[2]), .ZN(n83) );
  INVD1 U108 ( .I(n171), .ZN(n69) );
  ND3D1 U109 ( .A1(n190), .A2(n69), .A3(n172), .ZN(n37) );
  OAI21D1 U110 ( .A1(n118), .A2(n119), .B(n120), .ZN(n160) );
  ND4D1 U111 ( .A1(n121), .A2(n119), .A3(n122), .A4(n123), .ZN(n120) );
  XNR2D1 U112 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n121) );
  XNR2D1 U113 ( .A1(ReadAddr[1]), .A2(OldReadAr[1]), .ZN(n122) );
  OAI21D1 U114 ( .A1(n74), .A2(n73), .B(n172), .ZN(n86) );
  NR2D1 U115 ( .A1(n166), .A2(n165), .ZN(n130) );
  XNR2D1 U116 ( .A1(n113), .A2(n165), .ZN(n95) );
  OAI31D0 U117 ( .A1(n42), .A2(n195), .A3(ReadReq), .B(n43), .ZN(n151) );
  OAI21D1 U118 ( .A1(n44), .A2(n195), .B(FullFIFO), .ZN(n43) );
  BUFFD1 U119 ( .I(n170), .Z(n190) );
  INVD1 U120 ( .I(OldReadAr[2]), .ZN(n39) );
  INVD1 U121 ( .I(OldReadAr[3]), .ZN(n41) );
  ND2D1 U122 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U123 ( .I(ReadReq), .ZN(n117) );
endmodule


module DPMem1kx32_AWid4_DWid32_0 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, N133, N166, N199, N232, N265, N298, N331, N364, N397,
         N430, N463, N496, N529, N562, N595, N628, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n103, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n102,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  OR2D1 U3 ( .A1(n486), .A2(Dreadyr), .Z(n103) );
  XNR4D1 U13 ( .A1(n234), .A2(n233), .A3(n236), .A4(n235), .ZN(n76) );
  XOR4D1 U14 ( .A1(n238), .A2(n237), .A3(n240), .A4(n239), .Z(n75) );
  XOR4D1 U15 ( .A1(n230), .A2(n229), .A3(n232), .A4(n231), .Z(n72) );
  XOR4D1 U16 ( .A1(n223), .A2(n222), .A3(n225), .A4(n224), .Z(n69) );
  XNR4D1 U17 ( .A1(n216), .A2(n215), .A3(n218), .A4(n217), .ZN(n66) );
  XOR4D1 U21 ( .A1(n81), .A2(N71), .A3(n82), .A4(N74), .Z(n80) );
  XNR4D1 U22 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n82) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n88) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n87) );
  XNR4D1 U29 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .ZN(n84) );
  XNR4D1 U30 ( .A1(N79), .A2(N77), .A3(N81), .A4(N80), .ZN(n78) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N84), .E(n251), .CP(n379), .CDN(n540), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n240), .E(n251), .CP(n379), .CDN(n539), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n239), .E(n251), .CP(n379), .CDN(n539), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n238), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n233), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n232), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n231), .E(n252), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n230), .E(n252), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n229), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n228), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n227), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n226), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n225), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n224), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n223), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n222), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n221), .E(n253), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n220), .E(n253), .CP(n382), .CDN(n538), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n219), .E(n253), .CP(n382), .CDN(n538), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n218), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n217), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n216), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n215), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n214), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n213), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n212), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n211), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n210), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n209), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N84), .E(n259), .CP(n383), .CDN(n537), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n240), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n239), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n238), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n233), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n232), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n231), .E(n260), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n230), .E(n260), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n229), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n228), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n227), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n226), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n225), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n224), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n223), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n222), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n221), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n220), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n219), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n218), .E(n261), .CP(n385), .CDN(n534), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n217), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n216), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n215), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n214), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n213), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n212), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n211), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n210), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n209), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N84), .E(n283), .CP(n394), .CDN(n528), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n240), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n239), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n238), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n233), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n232), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n231), .E(n284), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n230), .E(n284), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n229), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n228), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n227), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n226), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n225), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n224), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n223), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n222), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n221), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n220), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n219), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n218), .E(n285), .CP(n396), .CDN(n525), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n217), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n216), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n215), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n214), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n213), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n212), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n211), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n210), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n209), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N84), .E(n291), .CP(n398), .CDN(n525), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n240), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n239), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n238), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n233), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n232), .E(n291), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n231), .E(n292), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n230), .E(n292), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n229), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n228), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n227), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n226), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n225), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n224), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n223), .E(n292), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n222), .E(n292), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n221), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n220), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n219), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n218), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n217), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n216), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n215), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n214), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n213), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n212), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n211), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n210), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n209), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N84), .E(n315), .CP(n409), .CDN(n516), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n240), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n239), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n238), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n233), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n232), .E(n315), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n231), .E(n316), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n230), .E(n316), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n229), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n228), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n227), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n226), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n225), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n224), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n223), .E(n316), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n222), .E(n316), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n221), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n220), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n219), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n218), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n217), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n216), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n215), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n214), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n213), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n212), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n211), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n210), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n209), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N84), .E(n323), .CP(n412), .CDN(n513), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n240), .E(n323), .CP(n412), .CDN(n512), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n239), .E(n323), .CP(n412), .CDN(n512), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n238), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n233), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n232), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n231), .E(n324), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n230), .E(n324), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n229), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n228), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n227), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n226), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n225), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n224), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n223), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n222), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n221), .E(n325), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n220), .E(n325), .CP(n415), .CDN(n511), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n219), .E(n325), .CP(n415), .CDN(n511), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n218), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n217), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n216), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n215), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n214), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n213), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n212), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n211), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n210), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n209), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N84), .E(n347), .CP(n423), .CDN(n504), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n240), .E(n347), .CP(n423), .CDN(n503), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n239), .E(n347), .CP(n423), .CDN(n503), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n238), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n233), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n232), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n231), .E(n348), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n230), .E(n348), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n229), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n228), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n227), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n226), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n225), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n224), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n223), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n222), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n221), .E(n349), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n220), .E(n349), .CP(n426), .CDN(n502), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n219), .E(n349), .CP(n426), .CDN(n502), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n218), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n217), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n216), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n215), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n214), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n213), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n212), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n211), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n210), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n209), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N84), .E(n355), .CP(n427), .CDN(n501), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n240), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n239), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n238), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n233), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n232), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n231), .E(n356), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n230), .E(n356), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n229), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n228), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n227), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n226), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n225), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n224), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n223), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n222), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n221), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n220), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n219), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n218), .E(n357), .CP(n429), .CDN(n498), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n217), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n216), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n215), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n214), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n213), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n212), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n211), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n210), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n209), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N84), .E(n243), .CP(n376), .CDN(n543), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n240), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n239), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n238), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n233), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n232), .E(n243), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n231), .E(n244), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n230), .E(n244), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n229), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n228), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n227), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n226), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n225), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n224), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n223), .E(n244), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n222), .E(n244), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n221), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n220), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n219), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n218), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n217), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n216), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n215), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n214), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n213), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n212), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n211), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n210), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n209), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N84), .E(n267), .CP(n387), .CDN(n534), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n240), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n239), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n238), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n233), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n232), .E(n267), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n231), .E(n268), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n230), .E(n268), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n229), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n228), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n227), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n226), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n225), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n224), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n223), .E(n268), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n222), .E(n268), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n221), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n220), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n219), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n218), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n217), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n216), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n215), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n214), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n213), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n212), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n211), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n210), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n209), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N84), .E(n275), .CP(n390), .CDN(n531), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n240), .E(n275), .CP(n390), .CDN(n530), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n239), .E(n275), .CP(n390), .CDN(n530), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n238), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n233), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n232), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n231), .E(n276), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n230), .E(n276), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n229), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n228), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n227), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n226), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n225), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n224), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n223), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n222), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n221), .E(n277), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n220), .E(n277), .CP(n393), .CDN(n529), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n219), .E(n277), .CP(n393), .CDN(n529), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n218), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n217), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n216), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n215), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n214), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n213), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n212), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n211), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n210), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n209), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N84), .E(n299), .CP(n401), .CDN(n522), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n240), .E(n299), .CP(n401), .CDN(n521), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n239), .E(n299), .CP(n401), .CDN(n521), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n238), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n233), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n232), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n231), .E(n300), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n230), .E(n300), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n229), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n228), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n227), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n226), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n225), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n224), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n223), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n222), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n221), .E(n301), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n220), .E(n301), .CP(n404), .CDN(n520), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n219), .E(n301), .CP(n404), .CDN(n520), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n218), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n217), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n216), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n215), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n214), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n213), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n212), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n211), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n210), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n209), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N84), .E(n307), .CP(n405), .CDN(n519), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n240), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n239), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n238), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n233), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n232), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n231), .E(n308), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n230), .E(n308), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n229), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n228), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n227), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n226), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n225), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n224), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n223), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n222), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n221), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n220), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n219), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n218), .E(n309), .CP(n407), .CDN(n516), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n217), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n216), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n215), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n214), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n213), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n212), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n211), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n210), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n209), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N84), .E(n331), .CP(n416), .CDN(n510), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n240), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n239), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n238), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n233), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n232), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n231), .E(n332), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n230), .E(n332), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n229), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n228), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n227), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n226), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n225), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n224), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n223), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n222), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n221), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n220), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n219), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n218), .E(n333), .CP(n418), .CDN(n507), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n217), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n216), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n215), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n214), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n213), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n212), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n211), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n210), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n209), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N84), .E(n339), .CP(n420), .CDN(n507), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n240), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n239), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n238), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n233), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n232), .E(n339), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n231), .E(n340), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n230), .E(n340), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n229), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n228), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n227), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n226), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n225), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n224), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n223), .E(n340), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n222), .E(n340), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n221), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n220), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n219), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n218), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n217), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n216), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n215), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n214), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n213), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n212), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n211), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n210), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n209), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N84), .E(n363), .CP(n431), .CDN(n498), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n240), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n239), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n238), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n233), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n232), .E(n363), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n231), .E(n364), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n230), .E(n364), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n229), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n228), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n227), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n226), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n225), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n224), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n223), .E(n364), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n222), .E(n364), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n221), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n220), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n219), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n218), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n217), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n216), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n215), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n214), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n213), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n212), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n211), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n210), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n209), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n103), .CP(n480), .CDN(n495), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n237), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n236), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n235), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n234), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n237), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n236), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n235), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n234), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n237), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n236), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n235), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n234), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n237), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n236), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n235), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n234), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n237), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n236), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n235), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n234), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n237), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n236), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n235), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n234), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n237), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n236), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n235), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n234), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n237), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n236), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n235), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n234), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n237), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n236), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n235), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n234), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n237), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n236), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n235), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n234), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n237), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n236), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n235), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n234), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n237), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n236), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n235), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n234), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n237), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n236), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n235), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n234), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n237), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n236), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n235), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n234), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n237), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n236), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n235), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n234), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n237), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n236), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n235), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n234), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N50), .E(n483), .CP(n477), .CDN(n546), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N51), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N52), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N53), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N54), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N55), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N56), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N57), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N58), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N59), .E(n483), .CP(n478), .CDN(n545), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N60), .E(n484), .CP(n478), .CDN(n545), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N61), .E(n484), .CP(n478), .CDN(n545), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N62), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N63), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N64), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N65), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N66), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N67), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N68), .E(n484), .CP(n479), .CDN(n544), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N69), .E(n484), .CP(n479), .CDN(n544), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N70), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N71), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N72), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N73), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N74), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N75), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N76), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N77), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N78), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N79), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N80), .E(n486), .CP(n480), .CDN(n543), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N81), .E(n486), .CP(n480), .CDN(n543), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N82), .E(n486), .CP(n480), .CDN(n543), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKAN2D0 U4 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  INVD1 U5 ( .I(n494), .ZN(n171) );
  INVD1 U6 ( .I(n493), .ZN(n175) );
  BUFFD1 U7 ( .I(n569), .Z(n501) );
  BUFFD1 U8 ( .I(n569), .Z(n502) );
  BUFFD1 U9 ( .I(n568), .Z(n503) );
  BUFFD1 U10 ( .I(n568), .Z(n504) );
  BUFFD1 U11 ( .I(n567), .Z(n505) );
  BUFFD1 U12 ( .I(n567), .Z(n506) );
  BUFFD1 U18 ( .I(n566), .Z(n507) );
  BUFFD1 U19 ( .I(n566), .Z(n508) );
  BUFFD1 U20 ( .I(n565), .Z(n509) );
  BUFFD1 U23 ( .I(n565), .Z(n510) );
  BUFFD1 U24 ( .I(n564), .Z(n511) );
  BUFFD1 U25 ( .I(n564), .Z(n512) );
  BUFFD1 U26 ( .I(n563), .Z(n513) );
  BUFFD1 U31 ( .I(n563), .Z(n514) );
  BUFFD1 U32 ( .I(n562), .Z(n515) );
  BUFFD1 U33 ( .I(n562), .Z(n516) );
  BUFFD1 U34 ( .I(n561), .Z(n517) );
  BUFFD1 U35 ( .I(n561), .Z(n518) );
  BUFFD1 U36 ( .I(n560), .Z(n519) );
  BUFFD1 U37 ( .I(n560), .Z(n520) );
  BUFFD1 U38 ( .I(n559), .Z(n521) );
  BUFFD1 U39 ( .I(n559), .Z(n522) );
  BUFFD1 U40 ( .I(n558), .Z(n523) );
  BUFFD1 U41 ( .I(n558), .Z(n524) );
  BUFFD1 U42 ( .I(n557), .Z(n525) );
  BUFFD1 U43 ( .I(n557), .Z(n526) );
  BUFFD1 U44 ( .I(n556), .Z(n527) );
  BUFFD1 U45 ( .I(n556), .Z(n528) );
  BUFFD1 U46 ( .I(n555), .Z(n529) );
  BUFFD1 U47 ( .I(n555), .Z(n530) );
  BUFFD1 U48 ( .I(n554), .Z(n531) );
  BUFFD1 U49 ( .I(n554), .Z(n532) );
  BUFFD1 U50 ( .I(n553), .Z(n533) );
  BUFFD1 U51 ( .I(n553), .Z(n534) );
  BUFFD1 U52 ( .I(n552), .Z(n535) );
  BUFFD1 U53 ( .I(n552), .Z(n536) );
  BUFFD1 U54 ( .I(n551), .Z(n537) );
  BUFFD1 U55 ( .I(n551), .Z(n538) );
  BUFFD1 U56 ( .I(n550), .Z(n539) );
  BUFFD1 U57 ( .I(n550), .Z(n540) );
  BUFFD1 U58 ( .I(n549), .Z(n541) );
  BUFFD1 U59 ( .I(n549), .Z(n542) );
  BUFFD1 U60 ( .I(n548), .Z(n543) );
  BUFFD1 U61 ( .I(n548), .Z(n544) );
  BUFFD1 U62 ( .I(n547), .Z(n545) );
  BUFFD1 U63 ( .I(n547), .Z(n546) );
  BUFFD1 U64 ( .I(n572), .Z(n495) );
  BUFFD1 U65 ( .I(n572), .Z(n496) );
  BUFFD1 U66 ( .I(n571), .Z(n497) );
  BUFFD1 U67 ( .I(n571), .Z(n498) );
  BUFFD1 U68 ( .I(n570), .Z(n499) );
  BUFFD1 U69 ( .I(n570), .Z(n500) );
  BUFFD1 U70 ( .I(n574), .Z(n569) );
  BUFFD1 U71 ( .I(n574), .Z(n568) );
  BUFFD1 U72 ( .I(n574), .Z(n567) );
  BUFFD1 U73 ( .I(n575), .Z(n566) );
  BUFFD1 U74 ( .I(n575), .Z(n565) );
  BUFFD1 U75 ( .I(n575), .Z(n564) );
  BUFFD1 U76 ( .I(n576), .Z(n563) );
  BUFFD1 U77 ( .I(n576), .Z(n562) );
  BUFFD1 U78 ( .I(n576), .Z(n561) );
  BUFFD1 U79 ( .I(n577), .Z(n560) );
  BUFFD1 U80 ( .I(n577), .Z(n559) );
  BUFFD1 U81 ( .I(n577), .Z(n558) );
  BUFFD1 U82 ( .I(n578), .Z(n557) );
  BUFFD1 U83 ( .I(n578), .Z(n556) );
  BUFFD1 U84 ( .I(n578), .Z(n555) );
  BUFFD1 U85 ( .I(n579), .Z(n554) );
  BUFFD1 U86 ( .I(n579), .Z(n553) );
  BUFFD1 U87 ( .I(n579), .Z(n552) );
  BUFFD1 U88 ( .I(n580), .Z(n551) );
  BUFFD1 U89 ( .I(n580), .Z(n550) );
  BUFFD1 U90 ( .I(n580), .Z(n549) );
  BUFFD1 U91 ( .I(n581), .Z(n548) );
  BUFFD1 U92 ( .I(n581), .Z(n547) );
  BUFFD1 U93 ( .I(n573), .Z(n571) );
  BUFFD1 U94 ( .I(n573), .Z(n570) );
  BUFFD1 U95 ( .I(n573), .Z(n572) );
  BUFFD1 U96 ( .I(n585), .Z(n574) );
  BUFFD1 U97 ( .I(n585), .Z(n575) );
  BUFFD1 U98 ( .I(n584), .Z(n576) );
  BUFFD1 U99 ( .I(n584), .Z(n577) );
  BUFFD1 U100 ( .I(n583), .Z(n578) );
  BUFFD1 U101 ( .I(n583), .Z(n579) );
  BUFFD1 U102 ( .I(n582), .Z(n580) );
  BUFFD1 U103 ( .I(n582), .Z(n581) );
  BUFFD1 U104 ( .I(n587), .Z(n585) );
  BUFFD1 U105 ( .I(n587), .Z(n584) );
  BUFFD1 U106 ( .I(n588), .Z(n583) );
  BUFFD1 U107 ( .I(n588), .Z(n582) );
  BUFFD1 U108 ( .I(n586), .Z(n573) );
  BUFFD1 U109 ( .I(n587), .Z(n586) );
  INVD1 U110 ( .I(n589), .ZN(n587) );
  INVD1 U111 ( .I(n589), .ZN(n588) );
  INVD1 U112 ( .I(n590), .ZN(n589) );
  INVD1 U113 ( .I(Reset), .ZN(n590) );
  BUFFD1 U114 ( .I(n435), .Z(n433) );
  BUFFD1 U115 ( .I(n436), .Z(n432) );
  BUFFD1 U116 ( .I(n436), .Z(n431) );
  BUFFD1 U117 ( .I(n437), .Z(n430) );
  BUFFD1 U118 ( .I(n437), .Z(n429) );
  BUFFD1 U119 ( .I(n438), .Z(n428) );
  BUFFD1 U120 ( .I(n438), .Z(n427) );
  BUFFD1 U121 ( .I(n439), .Z(n426) );
  BUFFD1 U122 ( .I(n439), .Z(n425) );
  BUFFD1 U123 ( .I(n440), .Z(n424) );
  BUFFD1 U124 ( .I(n440), .Z(n423) );
  BUFFD1 U125 ( .I(n441), .Z(n422) );
  BUFFD1 U126 ( .I(n441), .Z(n421) );
  BUFFD1 U127 ( .I(n442), .Z(n420) );
  BUFFD1 U128 ( .I(n442), .Z(n419) );
  BUFFD1 U129 ( .I(n443), .Z(n418) );
  BUFFD1 U130 ( .I(n443), .Z(n417) );
  BUFFD1 U131 ( .I(n444), .Z(n416) );
  BUFFD1 U132 ( .I(n444), .Z(n415) );
  BUFFD1 U133 ( .I(n445), .Z(n414) );
  BUFFD1 U134 ( .I(n445), .Z(n413) );
  BUFFD1 U135 ( .I(n446), .Z(n412) );
  BUFFD1 U136 ( .I(n446), .Z(n411) );
  BUFFD1 U137 ( .I(n447), .Z(n410) );
  BUFFD1 U138 ( .I(n447), .Z(n409) );
  BUFFD1 U139 ( .I(n448), .Z(n408) );
  BUFFD1 U140 ( .I(n448), .Z(n407) );
  BUFFD1 U141 ( .I(n449), .Z(n406) );
  BUFFD1 U142 ( .I(n449), .Z(n405) );
  BUFFD1 U143 ( .I(n450), .Z(n404) );
  BUFFD1 U144 ( .I(n450), .Z(n403) );
  BUFFD1 U145 ( .I(n451), .Z(n402) );
  BUFFD1 U146 ( .I(n451), .Z(n401) );
  BUFFD1 U147 ( .I(n452), .Z(n400) );
  BUFFD1 U148 ( .I(n452), .Z(n399) );
  BUFFD1 U149 ( .I(n453), .Z(n398) );
  BUFFD1 U150 ( .I(n453), .Z(n397) );
  BUFFD1 U151 ( .I(n454), .Z(n396) );
  BUFFD1 U152 ( .I(n454), .Z(n395) );
  BUFFD1 U153 ( .I(n455), .Z(n394) );
  BUFFD1 U154 ( .I(n455), .Z(n393) );
  BUFFD1 U155 ( .I(n456), .Z(n392) );
  BUFFD1 U156 ( .I(n456), .Z(n391) );
  BUFFD1 U157 ( .I(n457), .Z(n390) );
  BUFFD1 U158 ( .I(n457), .Z(n389) );
  BUFFD1 U159 ( .I(n458), .Z(n388) );
  BUFFD1 U160 ( .I(n458), .Z(n387) );
  BUFFD1 U161 ( .I(n459), .Z(n386) );
  BUFFD1 U162 ( .I(n459), .Z(n385) );
  BUFFD1 U163 ( .I(n460), .Z(n384) );
  BUFFD1 U164 ( .I(n460), .Z(n383) );
  BUFFD1 U165 ( .I(n461), .Z(n382) );
  BUFFD1 U166 ( .I(n461), .Z(n381) );
  BUFFD1 U167 ( .I(n462), .Z(n380) );
  BUFFD1 U168 ( .I(n462), .Z(n379) );
  BUFFD1 U169 ( .I(n463), .Z(n378) );
  BUFFD1 U170 ( .I(n463), .Z(n377) );
  BUFFD1 U171 ( .I(n435), .Z(n434) );
  INVD1 U172 ( .I(n367), .ZN(n365) );
  INVD1 U173 ( .I(n368), .ZN(n364) );
  INVD1 U174 ( .I(n368), .ZN(n363) );
  INVD1 U175 ( .I(n303), .ZN(n301) );
  INVD1 U176 ( .I(n304), .ZN(n300) );
  INVD1 U177 ( .I(n304), .ZN(n299) );
  INVD1 U178 ( .I(n367), .ZN(n366) );
  INVD1 U179 ( .I(n303), .ZN(n302) );
  BUFFD1 U180 ( .I(n464), .Z(n376) );
  BUFFD1 U181 ( .I(n465), .Z(n464) );
  BUFFD1 U182 ( .I(n474), .Z(n435) );
  BUFFD1 U183 ( .I(n474), .Z(n436) );
  BUFFD1 U184 ( .I(n474), .Z(n437) );
  BUFFD1 U185 ( .I(n473), .Z(n438) );
  BUFFD1 U186 ( .I(n473), .Z(n439) );
  BUFFD1 U187 ( .I(n473), .Z(n440) );
  BUFFD1 U188 ( .I(n472), .Z(n441) );
  BUFFD1 U189 ( .I(n472), .Z(n442) );
  BUFFD1 U190 ( .I(n472), .Z(n443) );
  BUFFD1 U191 ( .I(n471), .Z(n444) );
  BUFFD1 U192 ( .I(n471), .Z(n445) );
  BUFFD1 U193 ( .I(n471), .Z(n446) );
  BUFFD1 U194 ( .I(n470), .Z(n447) );
  BUFFD1 U195 ( .I(n470), .Z(n448) );
  BUFFD1 U196 ( .I(n470), .Z(n449) );
  BUFFD1 U197 ( .I(n469), .Z(n450) );
  BUFFD1 U198 ( .I(n469), .Z(n451) );
  BUFFD1 U199 ( .I(n469), .Z(n452) );
  BUFFD1 U200 ( .I(n468), .Z(n453) );
  BUFFD1 U201 ( .I(n468), .Z(n454) );
  BUFFD1 U202 ( .I(n468), .Z(n455) );
  BUFFD1 U203 ( .I(n467), .Z(n456) );
  BUFFD1 U204 ( .I(n467), .Z(n457) );
  BUFFD1 U205 ( .I(n467), .Z(n458) );
  BUFFD1 U206 ( .I(n466), .Z(n459) );
  BUFFD1 U207 ( .I(n466), .Z(n460) );
  BUFFD1 U208 ( .I(n466), .Z(n461) );
  BUFFD1 U209 ( .I(n465), .Z(n462) );
  BUFFD1 U210 ( .I(n465), .Z(n463) );
  INVD1 U211 ( .I(n361), .ZN(n367) );
  INVD1 U212 ( .I(n361), .ZN(n368) );
  INVD1 U213 ( .I(n297), .ZN(n303) );
  INVD1 U214 ( .I(n297), .ZN(n304) );
  INVD1 U215 ( .I(n359), .ZN(n357) );
  INVD1 U216 ( .I(n360), .ZN(n356) );
  INVD1 U217 ( .I(n360), .ZN(n355) );
  INVD1 U218 ( .I(n351), .ZN(n349) );
  INVD1 U219 ( .I(n352), .ZN(n348) );
  INVD1 U220 ( .I(n352), .ZN(n347) );
  INVD1 U221 ( .I(n343), .ZN(n341) );
  INVD1 U222 ( .I(n344), .ZN(n340) );
  INVD1 U223 ( .I(n344), .ZN(n339) );
  INVD1 U224 ( .I(n335), .ZN(n333) );
  INVD1 U225 ( .I(n336), .ZN(n332) );
  INVD1 U226 ( .I(n336), .ZN(n331) );
  INVD1 U227 ( .I(n327), .ZN(n325) );
  INVD1 U228 ( .I(n328), .ZN(n324) );
  INVD1 U229 ( .I(n328), .ZN(n323) );
  INVD1 U230 ( .I(n319), .ZN(n317) );
  INVD1 U231 ( .I(n320), .ZN(n316) );
  INVD1 U232 ( .I(n320), .ZN(n315) );
  INVD1 U233 ( .I(n311), .ZN(n309) );
  INVD1 U234 ( .I(n312), .ZN(n308) );
  INVD1 U235 ( .I(n312), .ZN(n307) );
  INVD1 U236 ( .I(n295), .ZN(n293) );
  INVD1 U237 ( .I(n296), .ZN(n292) );
  INVD1 U238 ( .I(n296), .ZN(n291) );
  INVD1 U239 ( .I(n287), .ZN(n285) );
  INVD1 U240 ( .I(n288), .ZN(n284) );
  INVD1 U241 ( .I(n288), .ZN(n283) );
  INVD1 U242 ( .I(n279), .ZN(n277) );
  INVD1 U243 ( .I(n280), .ZN(n276) );
  INVD1 U244 ( .I(n280), .ZN(n275) );
  INVD1 U245 ( .I(n271), .ZN(n269) );
  INVD1 U246 ( .I(n272), .ZN(n268) );
  INVD1 U247 ( .I(n272), .ZN(n267) );
  INVD1 U248 ( .I(n263), .ZN(n261) );
  INVD1 U249 ( .I(n264), .ZN(n260) );
  INVD1 U250 ( .I(n264), .ZN(n259) );
  INVD1 U251 ( .I(n255), .ZN(n253) );
  INVD1 U252 ( .I(n256), .ZN(n252) );
  INVD1 U253 ( .I(n256), .ZN(n251) );
  INVD1 U254 ( .I(n247), .ZN(n245) );
  INVD1 U255 ( .I(n248), .ZN(n244) );
  INVD1 U256 ( .I(n248), .ZN(n243) );
  INVD1 U257 ( .I(n351), .ZN(n350) );
  INVD1 U258 ( .I(n343), .ZN(n342) );
  INVD1 U259 ( .I(n359), .ZN(n358) );
  INVD1 U260 ( .I(n335), .ZN(n334) );
  INVD1 U261 ( .I(n327), .ZN(n326) );
  INVD1 U262 ( .I(n319), .ZN(n318) );
  INVD1 U263 ( .I(n311), .ZN(n310) );
  INVD1 U264 ( .I(n295), .ZN(n294) );
  INVD1 U265 ( .I(n287), .ZN(n286) );
  INVD1 U266 ( .I(n279), .ZN(n278) );
  INVD1 U267 ( .I(n271), .ZN(n270) );
  INVD1 U268 ( .I(n263), .ZN(n262) );
  INVD1 U269 ( .I(n255), .ZN(n254) );
  INVD1 U270 ( .I(n247), .ZN(n246) );
  BUFFD1 U271 ( .I(n373), .Z(n474) );
  BUFFD1 U272 ( .I(n373), .Z(n473) );
  BUFFD1 U273 ( .I(n372), .Z(n472) );
  BUFFD1 U274 ( .I(n372), .Z(n471) );
  BUFFD1 U275 ( .I(n371), .Z(n470) );
  BUFFD1 U276 ( .I(n371), .Z(n469) );
  BUFFD1 U277 ( .I(n370), .Z(n468) );
  BUFFD1 U278 ( .I(n370), .Z(n467) );
  BUFFD1 U279 ( .I(n369), .Z(n466) );
  BUFFD1 U280 ( .I(n369), .Z(n465) );
  BUFFD1 U281 ( .I(n197), .Z(n198) );
  BUFFD1 U282 ( .I(n197), .Z(n199) );
  BUFFD1 U283 ( .I(n197), .Z(n200) );
  BUFFD1 U284 ( .I(n196), .Z(n201) );
  BUFFD1 U285 ( .I(n196), .Z(n202) );
  BUFFD1 U286 ( .I(n196), .Z(n203) );
  BUFFD1 U287 ( .I(n195), .Z(n204) );
  BUFFD1 U288 ( .I(n195), .Z(n205) );
  BUFFD1 U289 ( .I(n195), .Z(n206) );
  BUFFD1 U290 ( .I(n194), .Z(n207) );
  BUFFD1 U291 ( .I(n194), .Z(n208) );
  BUFFD1 U292 ( .I(n182), .Z(n183) );
  BUFFD1 U293 ( .I(n182), .Z(n184) );
  BUFFD1 U294 ( .I(n182), .Z(n185) );
  BUFFD1 U295 ( .I(n181), .Z(n186) );
  BUFFD1 U296 ( .I(n181), .Z(n187) );
  BUFFD1 U297 ( .I(n181), .Z(n188) );
  BUFFD1 U298 ( .I(n180), .Z(n189) );
  BUFFD1 U299 ( .I(n180), .Z(n190) );
  BUFFD1 U300 ( .I(n180), .Z(n191) );
  BUFFD1 U301 ( .I(n179), .Z(n192) );
  BUFFD1 U302 ( .I(n179), .Z(n193) );
  INVD1 U303 ( .I(n353), .ZN(n359) );
  INVD1 U304 ( .I(n353), .ZN(n360) );
  INVD1 U305 ( .I(n345), .ZN(n351) );
  INVD1 U306 ( .I(n345), .ZN(n352) );
  INVD1 U307 ( .I(n337), .ZN(n343) );
  INVD1 U308 ( .I(n337), .ZN(n344) );
  INVD1 U309 ( .I(n329), .ZN(n335) );
  INVD1 U310 ( .I(n329), .ZN(n336) );
  INVD1 U311 ( .I(n321), .ZN(n327) );
  INVD1 U312 ( .I(n321), .ZN(n328) );
  INVD1 U313 ( .I(n313), .ZN(n319) );
  INVD1 U314 ( .I(n313), .ZN(n320) );
  INVD1 U315 ( .I(n305), .ZN(n311) );
  INVD1 U316 ( .I(n305), .ZN(n312) );
  INVD1 U317 ( .I(n289), .ZN(n295) );
  INVD1 U318 ( .I(n289), .ZN(n296) );
  INVD1 U319 ( .I(n281), .ZN(n287) );
  INVD1 U320 ( .I(n281), .ZN(n288) );
  INVD1 U321 ( .I(n273), .ZN(n279) );
  INVD1 U322 ( .I(n273), .ZN(n280) );
  INVD1 U323 ( .I(n265), .ZN(n271) );
  INVD1 U324 ( .I(n265), .ZN(n272) );
  INVD1 U325 ( .I(n257), .ZN(n263) );
  INVD1 U326 ( .I(n257), .ZN(n264) );
  INVD1 U327 ( .I(n249), .ZN(n255) );
  INVD1 U328 ( .I(n249), .ZN(n256) );
  INVD1 U329 ( .I(n241), .ZN(n247) );
  INVD1 U330 ( .I(n241), .ZN(n248) );
  INVD1 U331 ( .I(n362), .ZN(n361) );
  INVD1 U332 ( .I(N133), .ZN(n362) );
  NR2D1 U333 ( .A1(n94), .A2(n98), .ZN(N133) );
  INVD1 U334 ( .I(n298), .ZN(n297) );
  INVD1 U335 ( .I(N397), .ZN(n298) );
  NR2D1 U336 ( .A1(n91), .A2(n94), .ZN(N397) );
  INVD1 U337 ( .I(n487), .ZN(n485) );
  INVD1 U338 ( .I(n488), .ZN(n484) );
  INVD1 U339 ( .I(n488), .ZN(n483) );
  INVD1 U340 ( .I(n487), .ZN(n486) );
  BUFFD1 U341 ( .I(n374), .Z(n373) );
  BUFFD1 U342 ( .I(n374), .Z(n372) );
  BUFFD1 U343 ( .I(n374), .Z(n371) );
  BUFFD1 U344 ( .I(n375), .Z(n370) );
  BUFFD1 U345 ( .I(n375), .Z(n369) );
  INVD1 U346 ( .I(n481), .ZN(n479) );
  INVD1 U347 ( .I(n482), .ZN(n478) );
  INVD1 U348 ( .I(n482), .ZN(n477) );
  INVD1 U349 ( .I(n481), .ZN(n480) );
  XOR3D1 U350 ( .A1(n211), .A2(n210), .A3(n65), .Z(N84) );
  XOR3D1 U351 ( .A1(n209), .A2(n66), .A3(n67), .Z(n65) );
  XOR3D1 U352 ( .A1(n214), .A2(n213), .A3(n68), .Z(n67) );
  XOR3D1 U353 ( .A1(n228), .A2(n227), .A3(n74), .Z(n73) );
  XOR3D1 U354 ( .A1(n75), .A2(n226), .A3(n76), .Z(n74) );
  XOR3D1 U355 ( .A1(n69), .A2(n212), .A3(n70), .Z(n68) );
  XOR3D1 U356 ( .A1(n221), .A2(n220), .A3(n71), .Z(n70) );
  XOR3D1 U357 ( .A1(n72), .A2(n219), .A3(n73), .Z(n71) );
  XOR3D1 U358 ( .A1(N59), .A2(N58), .A3(n86), .Z(n85) );
  XOR3D1 U359 ( .A1(n87), .A2(N57), .A3(n88), .Z(n86) );
  XOR3D1 U360 ( .A1(N66), .A2(N65), .A3(n83), .Z(n81) );
  XOR3D1 U361 ( .A1(N64), .A2(n84), .A3(n85), .Z(n83) );
  XOR3D1 U362 ( .A1(N78), .A2(N73), .A3(n77), .Z(N82) );
  XOR3D1 U363 ( .A1(N72), .A2(n78), .A3(n79), .Z(n77) );
  XOR3D1 U364 ( .A1(N76), .A2(N75), .A3(n80), .Z(n79) );
  BUFFD1 U365 ( .I(n491), .Z(n197) );
  BUFFD1 U366 ( .I(n492), .Z(n182) );
  BUFFD1 U367 ( .I(n491), .Z(n196) );
  BUFFD1 U368 ( .I(n492), .Z(n181) );
  BUFFD1 U369 ( .I(n491), .Z(n195) );
  BUFFD1 U370 ( .I(n492), .Z(n180) );
  INVD1 U371 ( .I(n171), .ZN(n173) );
  INVD1 U372 ( .I(n171), .ZN(n174) );
  BUFFD1 U373 ( .I(n491), .Z(n194) );
  BUFFD1 U374 ( .I(n492), .Z(n179) );
  INVD1 U375 ( .I(n171), .ZN(n172) );
  INVD1 U376 ( .I(n175), .ZN(n177) );
  INVD1 U377 ( .I(n175), .ZN(n178) );
  INVD1 U378 ( .I(n175), .ZN(n176) );
  INVD1 U379 ( .I(n346), .ZN(n345) );
  INVD1 U380 ( .I(N199), .ZN(n346) );
  NR2D1 U381 ( .A1(n93), .A2(n98), .ZN(N199) );
  INVD1 U382 ( .I(n338), .ZN(n337) );
  INVD1 U383 ( .I(N232), .ZN(n338) );
  NR2D1 U384 ( .A1(n93), .A2(n97), .ZN(N232) );
  ND2D1 U385 ( .A1(n101), .A2(n96), .ZN(n98) );
  ND2D1 U386 ( .A1(n99), .A2(n100), .ZN(n94) );
  ND2D1 U387 ( .A1(n95), .A2(n96), .ZN(n91) );
  INVD1 U388 ( .I(n330), .ZN(n329) );
  INVD1 U389 ( .I(N265), .ZN(n330) );
  NR2D1 U390 ( .A1(n92), .A2(n98), .ZN(N265) );
  INVD1 U391 ( .I(n322), .ZN(n321) );
  INVD1 U392 ( .I(N298), .ZN(n322) );
  NR2D1 U393 ( .A1(n92), .A2(n97), .ZN(N298) );
  INVD1 U394 ( .I(n314), .ZN(n313) );
  INVD1 U395 ( .I(N331), .ZN(n314) );
  NR2D1 U396 ( .A1(n90), .A2(n98), .ZN(N331) );
  INVD1 U397 ( .I(n306), .ZN(n305) );
  INVD1 U398 ( .I(N364), .ZN(n306) );
  NR2D1 U399 ( .A1(n90), .A2(n97), .ZN(N364) );
  INVD1 U400 ( .I(n250), .ZN(n249) );
  INVD1 U401 ( .I(N595), .ZN(n250) );
  NR2D1 U402 ( .A1(n90), .A2(n91), .ZN(N595) );
  INVD1 U403 ( .I(n354), .ZN(n353) );
  INVD1 U404 ( .I(N166), .ZN(n354) );
  NR2D1 U405 ( .A1(n94), .A2(n97), .ZN(N166) );
  INVD1 U406 ( .I(n290), .ZN(n289) );
  INVD1 U407 ( .I(N430), .ZN(n290) );
  NR2D1 U408 ( .A1(n89), .A2(n94), .ZN(N430) );
  INVD1 U409 ( .I(n282), .ZN(n281) );
  INVD1 U410 ( .I(N463), .ZN(n282) );
  NR2D1 U411 ( .A1(n91), .A2(n93), .ZN(N463) );
  INVD1 U412 ( .I(n274), .ZN(n273) );
  INVD1 U413 ( .I(N496), .ZN(n274) );
  NR2D1 U414 ( .A1(n89), .A2(n93), .ZN(N496) );
  INVD1 U415 ( .I(n266), .ZN(n265) );
  INVD1 U416 ( .I(N529), .ZN(n266) );
  NR2D1 U417 ( .A1(n91), .A2(n92), .ZN(N529) );
  INVD1 U418 ( .I(n258), .ZN(n257) );
  INVD1 U419 ( .I(N562), .ZN(n258) );
  NR2D1 U420 ( .A1(n89), .A2(n92), .ZN(N562) );
  INVD1 U421 ( .I(n242), .ZN(n241) );
  INVD1 U422 ( .I(N628), .ZN(n242) );
  NR2D1 U423 ( .A1(n89), .A2(n90), .ZN(N628) );
  INVD1 U424 ( .I(n489), .ZN(n487) );
  INVD1 U425 ( .I(n489), .ZN(n488) );
  INVD1 U426 ( .I(n475), .ZN(n482) );
  INVD1 U427 ( .I(n475), .ZN(n481) );
  BUFFD1 U428 ( .I(ClockW), .Z(n374) );
  BUFFD1 U429 ( .I(ClockW), .Z(n375) );
  BUFFD1 U430 ( .I(DataI[14]), .Z(n223) );
  BUFFD1 U431 ( .I(DataI[15]), .Z(n224) );
  BUFFD1 U432 ( .I(DataI[21]), .Z(n230) );
  BUFFD1 U433 ( .I(DataI[22]), .Z(n231) );
  BUFFD1 U434 ( .I(DataI[25]), .Z(n234) );
  BUFFD1 U435 ( .I(DataI[26]), .Z(n235) );
  BUFFD1 U436 ( .I(DataI[29]), .Z(n238) );
  BUFFD1 U437 ( .I(DataI[30]), .Z(n239) );
  BUFFD1 U438 ( .I(DataI[10]), .Z(n219) );
  BUFFD1 U439 ( .I(DataI[11]), .Z(n220) );
  BUFFD1 U440 ( .I(DataI[17]), .Z(n226) );
  BUFFD1 U441 ( .I(DataI[18]), .Z(n227) );
  BUFFD1 U442 ( .I(DataI[13]), .Z(n222) );
  BUFFD1 U443 ( .I(DataI[16]), .Z(n225) );
  BUFFD1 U444 ( .I(DataI[20]), .Z(n229) );
  BUFFD1 U445 ( .I(DataI[23]), .Z(n232) );
  BUFFD1 U446 ( .I(DataI[24]), .Z(n233) );
  BUFFD1 U447 ( .I(DataI[27]), .Z(n236) );
  BUFFD1 U448 ( .I(DataI[28]), .Z(n237) );
  BUFFD1 U449 ( .I(DataI[31]), .Z(n240) );
  BUFFD1 U450 ( .I(DataI[12]), .Z(n221) );
  BUFFD1 U451 ( .I(DataI[19]), .Z(n228) );
  BUFFD1 U452 ( .I(DataI[2]), .Z(n211) );
  BUFFD1 U453 ( .I(DataI[1]), .Z(n210) );
  BUFFD1 U454 ( .I(DataI[7]), .Z(n216) );
  BUFFD1 U455 ( .I(DataI[8]), .Z(n217) );
  BUFFD1 U456 ( .I(DataI[3]), .Z(n212) );
  BUFFD1 U457 ( .I(DataI[4]), .Z(n213) );
  BUFFD1 U458 ( .I(DataI[6]), .Z(n215) );
  BUFFD1 U459 ( .I(DataI[9]), .Z(n218) );
  BUFFD1 U460 ( .I(DataI[0]), .Z(n209) );
  BUFFD1 U461 ( .I(DataI[5]), .Z(n214) );
  MUX4D0 U462 ( .I0(n8), .I1(n6), .I2(n7), .I3(n5), .S0(n172), .S1(n176), .Z(
        N80) );
  MUX4D0 U463 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n198), .S1(n183), .Z(n7)
         );
  MUX4D0 U464 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n198), .S1(n183), .Z(n6)
         );
  MUX4D0 U465 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n198), .S1(n183), .Z(n8)
         );
  MUX4D0 U466 ( .I0(n12), .I1(n10), .I2(n11), .I3(n9), .S0(n172), .S1(n176), 
        .Z(N79) );
  MUX4D0 U467 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n198), .S1(n183), .Z(n11)
         );
  MUX4D0 U468 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n198), .S1(n183), .Z(n10) );
  MUX4D0 U469 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n198), .S1(n183), .Z(n12)
         );
  MUX4D0 U470 ( .I0(n32), .I1(n30), .I2(n31), .I3(n29), .S0(n172), .S1(n176), 
        .Z(N74) );
  MUX4D0 U471 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n200), .S1(n185), .Z(n31)
         );
  MUX4D0 U472 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n200), .S1(n185), .Z(n30) );
  MUX4D0 U473 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n200), .S1(n185), .Z(n32)
         );
  MUX4D0 U474 ( .I0(n52), .I1(n50), .I2(n51), .I3(n49), .S0(n173), .S1(n177), 
        .Z(N69) );
  MUX4D0 U475 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n202), .S1(n187), .Z(n51) );
  MUX4D0 U476 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n202), .S1(n187), .Z(
        n50) );
  MUX4D0 U477 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n202), .S1(n187), .Z(n52) );
  MUX4D0 U478 ( .I0(n56), .I1(n54), .I2(n55), .I3(n53), .S0(n173), .S1(n177), 
        .Z(N68) );
  MUX4D0 U479 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n202), .S1(n187), .Z(n55) );
  MUX4D0 U480 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n202), .S1(n187), .Z(
        n54) );
  MUX4D0 U481 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n202), .S1(n187), .Z(n56) );
  MUX4D0 U482 ( .I0(n118), .I1(n116), .I2(n117), .I3(n115), .S0(n173), .S1(
        n177), .Z(N62) );
  MUX4D0 U483 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n204), .S1(n189), .Z(
        n117) );
  MUX4D0 U484 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n204), .S1(n189), .Z(
        n116) );
  MUX4D0 U485 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n204), .S1(n189), .Z(
        n118) );
  MUX4D0 U486 ( .I0(n122), .I1(n120), .I2(n121), .I3(n119), .S0(n173), .S1(
        n177), .Z(N61) );
  MUX4D0 U487 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n204), .S1(n189), .Z(
        n121) );
  MUX4D0 U488 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n204), .S1(n189), .Z(
        n120) );
  MUX4D0 U489 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n204), .S1(n189), .Z(
        n122) );
  MUX4D0 U490 ( .I0(n146), .I1(n144), .I2(n145), .I3(n143), .S0(n174), .S1(
        n178), .Z(N55) );
  MUX4D0 U491 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n206), .S1(n191), .Z(
        n145) );
  MUX4D0 U492 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n206), .S1(n191), .Z(
        n144) );
  MUX4D0 U493 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n206), .S1(n191), .Z(
        n146) );
  MUX4D0 U494 ( .I0(n150), .I1(n148), .I2(n149), .I3(n147), .S0(n174), .S1(
        n178), .Z(N54) );
  MUX4D0 U495 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n207), .S1(n192), .Z(
        n149) );
  MUX4D0 U496 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n207), .S1(n192), .Z(
        n148) );
  MUX4D0 U497 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n207), .S1(n192), .Z(
        n150) );
  MUX4D0 U498 ( .I0(n162), .I1(n160), .I2(n161), .I3(n159), .S0(n174), .S1(
        n178), .Z(N51) );
  MUX4D0 U499 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n208), .S1(n193), .Z(
        n161) );
  MUX4D0 U500 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n208), .S1(n193), .Z(
        n160) );
  MUX4D0 U501 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n208), .S1(n193), .Z(
        n162) );
  MUX4D0 U502 ( .I0(n166), .I1(n164), .I2(n165), .I3(n163), .S0(n174), .S1(
        n178), .Z(N50) );
  MUX4D0 U503 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n208), .S1(n193), .Z(
        n165) );
  MUX4D0 U504 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n208), .S1(n193), .Z(
        n164) );
  MUX4D0 U505 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n208), .S1(n193), .Z(
        n166) );
  MUX4D0 U506 ( .I0(n28), .I1(n26), .I2(n27), .I3(n25), .S0(n172), .S1(n176), 
        .Z(N75) );
  MUX4D0 U507 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n200), .S1(n185), .Z(n27)
         );
  MUX4D0 U508 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n200), .S1(n185), .Z(n26) );
  MUX4D0 U509 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n200), .S1(n185), .Z(n28)
         );
  MUX4D0 U510 ( .I0(n106), .I1(n104), .I2(n105), .I3(n102), .S0(n173), .S1(
        n177), .Z(N65) );
  MUX4D0 U511 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n203), .S1(n188), .Z(
        n105) );
  MUX4D0 U512 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n203), .S1(n188), .Z(
        n104) );
  MUX4D0 U513 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n203), .S1(n188), .Z(
        n106) );
  MUX4D0 U514 ( .I0(n134), .I1(n132), .I2(n133), .I3(n131), .S0(n174), .S1(
        n178), .Z(N58) );
  MUX4D0 U515 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n205), .S1(n190), .Z(
        n133) );
  MUX4D0 U516 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n205), .S1(n190), .Z(
        n132) );
  MUX4D0 U517 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n205), .S1(n190), .Z(
        n134) );
  MUX4D0 U518 ( .I0(n138), .I1(n136), .I2(n137), .I3(n135), .S0(n174), .S1(
        n178), .Z(N57) );
  MUX4D0 U519 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n206), .S1(n191), .Z(
        n137) );
  MUX4D0 U520 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n206), .S1(n191), .Z(
        n136) );
  MUX4D0 U521 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n206), .S1(n191), .Z(
        n138) );
  MUX4D0 U522 ( .I0(n4), .I1(n2), .I2(n3), .I3(n1), .S0(n172), .S1(n176), .Z(
        N81) );
  MUX4D0 U523 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n198), .S1(n183), .Z(n3)
         );
  MUX4D0 U524 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n198), .S1(n183), .Z(n2)
         );
  MUX4D0 U525 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n198), .S1(n183), .Z(n4)
         );
  MUX4D0 U526 ( .I0(n20), .I1(n18), .I2(n19), .I3(n17), .S0(n172), .S1(n176), 
        .Z(N77) );
  MUX4D0 U527 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n199), .S1(n184), .Z(n19)
         );
  MUX4D0 U528 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n199), .S1(n184), .Z(n18) );
  MUX4D0 U529 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n199), .S1(n184), .Z(n20)
         );
  MUX4D0 U530 ( .I0(n44), .I1(n42), .I2(n43), .I3(n41), .S0(n173), .S1(n177), 
        .Z(N71) );
  MUX4D0 U531 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n201), .S1(n186), .Z(n43) );
  MUX4D0 U532 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n201), .S1(n186), .Z(
        n42) );
  MUX4D0 U533 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n201), .S1(n186), .Z(n44) );
  MUX4D0 U534 ( .I0(n48), .I1(n46), .I2(n47), .I3(n45), .S0(n173), .S1(n177), 
        .Z(N70) );
  MUX4D0 U535 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n201), .S1(n186), .Z(n47) );
  MUX4D0 U536 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n201), .S1(n186), .Z(
        n46) );
  MUX4D0 U537 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n201), .S1(n186), .Z(n48) );
  MUX4D0 U538 ( .I0(n60), .I1(n58), .I2(n59), .I3(n57), .S0(n173), .S1(n177), 
        .Z(N67) );
  MUX4D0 U539 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n202), .S1(n187), .Z(n59) );
  MUX4D0 U540 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n202), .S1(n187), .Z(
        n58) );
  MUX4D0 U541 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n202), .S1(n187), .Z(n60) );
  MUX4D0 U542 ( .I0(n114), .I1(n112), .I2(n113), .I3(n111), .S0(n173), .S1(
        n177), .Z(N63) );
  MUX4D0 U543 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n204), .S1(n189), .Z(
        n113) );
  MUX4D0 U544 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n204), .S1(n189), .Z(
        n112) );
  MUX4D0 U545 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n204), .S1(n189), .Z(
        n114) );
  MUX4D0 U546 ( .I0(n126), .I1(n124), .I2(n125), .I3(n123), .S0(n174), .S1(
        n178), .Z(N60) );
  MUX4D0 U547 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n205), .S1(n190), .Z(
        n125) );
  MUX4D0 U548 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n205), .S1(n190), .Z(
        n124) );
  MUX4D0 U549 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n205), .S1(n190), .Z(
        n126) );
  MUX4D0 U550 ( .I0(n142), .I1(n140), .I2(n141), .I3(n139), .S0(n174), .S1(
        n178), .Z(N56) );
  MUX4D0 U551 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n206), .S1(n191), .Z(
        n141) );
  MUX4D0 U552 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n206), .S1(n191), .Z(
        n140) );
  MUX4D0 U553 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n206), .S1(n191), .Z(
        n142) );
  MUX4D0 U554 ( .I0(n154), .I1(n152), .I2(n153), .I3(n151), .S0(n174), .S1(
        n178), .Z(N53) );
  MUX4D0 U555 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n207), .S1(n192), .Z(
        n153) );
  MUX4D0 U556 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n207), .S1(n192), .Z(
        n152) );
  MUX4D0 U557 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n207), .S1(n192), .Z(
        n154) );
  MUX4D0 U558 ( .I0(n158), .I1(n156), .I2(n157), .I3(n155), .S0(n174), .S1(
        n178), .Z(N52) );
  MUX4D0 U559 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n207), .S1(n192), .Z(
        n157) );
  MUX4D0 U560 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n207), .S1(n192), .Z(
        n156) );
  MUX4D0 U561 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n207), .S1(n192), .Z(
        n158) );
  MUX4D0 U562 ( .I0(n24), .I1(n22), .I2(n23), .I3(n21), .S0(n172), .S1(n176), 
        .Z(N76) );
  MUX4D0 U563 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n199), .S1(n184), .Z(n23)
         );
  MUX4D0 U564 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n199), .S1(n184), .Z(n22) );
  MUX4D0 U565 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n199), .S1(n184), .Z(n24)
         );
  MUX4D0 U566 ( .I0(n40), .I1(n38), .I2(n39), .I3(n37), .S0(n173), .S1(n177), 
        .Z(N72) );
  MUX4D0 U567 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n201), .S1(n186), .Z(n39)
         );
  MUX4D0 U568 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n201), .S1(n186), .Z(n38) );
  MUX4D0 U569 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n201), .S1(n186), .Z(n40)
         );
  MUX4D0 U570 ( .I0(n64), .I1(n62), .I2(n63), .I3(n61), .S0(n173), .S1(n177), 
        .Z(N66) );
  MUX4D0 U571 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n203), .S1(n188), .Z(n63) );
  MUX4D0 U572 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n203), .S1(n188), .Z(
        n62) );
  MUX4D0 U573 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n203), .S1(n188), .Z(n64) );
  MUX4D0 U574 ( .I0(n110), .I1(n108), .I2(n109), .I3(n107), .S0(n173), .S1(
        n177), .Z(N64) );
  MUX4D0 U575 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n203), .S1(n188), .Z(
        n109) );
  MUX4D0 U576 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n203), .S1(n188), .Z(
        n108) );
  MUX4D0 U577 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n203), .S1(n188), .Z(
        n110) );
  MUX4D0 U578 ( .I0(n130), .I1(n128), .I2(n129), .I3(n127), .S0(n174), .S1(
        n178), .Z(N59) );
  MUX4D0 U579 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n205), .S1(n190), .Z(
        n129) );
  MUX4D0 U580 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n205), .S1(n190), .Z(
        n128) );
  MUX4D0 U581 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n205), .S1(n190), .Z(
        n130) );
  MUX4D0 U582 ( .I0(n170), .I1(n168), .I2(n169), .I3(n167), .S0(n174), .S1(
        n178), .Z(N49) );
  MUX4D0 U583 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n208), .S1(n193), .Z(
        n169) );
  MUX4D0 U584 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n208), .S1(n193), .Z(
        n168) );
  MUX4D0 U585 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n208), .S1(n193), .Z(
        n170) );
  MUX4D0 U586 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n208), .S1(n193), .Z(
        n167) );
  MUX4D0 U587 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n198), .S1(n183), .Z(n1)
         );
  MUX4D0 U588 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n198), .S1(n183), .Z(n5)
         );
  MUX4D0 U589 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n198), .S1(n183), .Z(n9)
         );
  MUX4D0 U590 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n199), .S1(n184), .Z(n17) );
  MUX4D0 U591 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n199), .S1(n184), .Z(n21) );
  MUX4D0 U592 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n200), .S1(n185), .Z(n25) );
  MUX4D0 U593 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n200), .S1(n185), .Z(n29) );
  MUX4D0 U594 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n201), .S1(n186), .Z(n37) );
  MUX4D0 U595 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n201), .S1(n186), .Z(
        n41) );
  MUX4D0 U596 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n201), .S1(n186), .Z(
        n45) );
  MUX4D0 U597 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n202), .S1(n187), .Z(
        n49) );
  MUX4D0 U598 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n202), .S1(n187), .Z(
        n53) );
  MUX4D0 U599 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n202), .S1(n187), .Z(
        n57) );
  MUX4D0 U600 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n203), .S1(n188), .Z(
        n61) );
  MUX4D0 U601 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n203), .S1(n188), .Z(
        n102) );
  MUX4D0 U602 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n203), .S1(n188), .Z(
        n107) );
  MUX4D0 U603 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n204), .S1(n189), .Z(
        n111) );
  MUX4D0 U604 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n204), .S1(n189), .Z(
        n115) );
  MUX4D0 U605 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n204), .S1(n189), .Z(
        n119) );
  MUX4D0 U606 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n205), .S1(n190), .Z(
        n123) );
  MUX4D0 U607 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n205), .S1(n190), .Z(
        n127) );
  MUX4D0 U608 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n205), .S1(n190), .Z(
        n131) );
  MUX4D0 U609 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n206), .S1(n191), .Z(
        n135) );
  MUX4D0 U610 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n206), .S1(n191), .Z(
        n139) );
  MUX4D0 U611 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n206), .S1(n191), .Z(
        n143) );
  MUX4D0 U612 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n207), .S1(n192), .Z(
        n147) );
  MUX4D0 U613 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n207), .S1(n192), .Z(
        n151) );
  MUX4D0 U614 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n207), .S1(n192), .Z(
        n155) );
  MUX4D0 U615 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n208), .S1(n193), .Z(
        n159) );
  MUX4D0 U616 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n208), .S1(n193), .Z(
        n163) );
  BUFFD1 U617 ( .I(N47), .Z(n494) );
  BUFFD1 U618 ( .I(N46), .Z(n493) );
  BUFFD1 U619 ( .I(N44), .Z(n491) );
  BUFFD1 U620 ( .I(N45), .Z(n492) );
  MUX4D0 U621 ( .I0(n36), .I1(n34), .I2(n35), .I3(n33), .S0(n172), .S1(n176), 
        .Z(N73) );
  MUX4D0 U622 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n200), .S1(n185), .Z(n35)
         );
  MUX4D0 U623 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n200), .S1(n185), .Z(n34) );
  MUX4D0 U624 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n200), .S1(n185), .Z(n36)
         );
  MUX4D0 U625 ( .I0(n16), .I1(n14), .I2(n15), .I3(n13), .S0(n172), .S1(n176), 
        .Z(N78) );
  MUX4D0 U626 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n199), .S1(n184), .Z(n15)
         );
  MUX4D0 U627 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n199), .S1(n184), .Z(n14) );
  MUX4D0 U628 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n199), .S1(n184), .Z(n16)
         );
  MUX4D0 U629 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n199), .S1(n184), .Z(n13) );
  MUX4D0 U630 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n200), .S1(n185), .Z(n33) );
  ND2D1 U631 ( .A1(AddrW[1]), .A2(n100), .ZN(n93) );
  ND2D1 U632 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n90) );
  ND2D1 U633 ( .A1(n101), .A2(AddrW[0]), .ZN(n97) );
  ND2D1 U634 ( .A1(AddrW[2]), .A2(n99), .ZN(n92) );
  ND2D1 U635 ( .A1(AddrW[0]), .A2(n95), .ZN(n89) );
  INR2D1 U636 ( .A1(Write), .B1(AddrW[3]), .ZN(n101) );
  INVD1 U637 ( .I(AddrW[1]), .ZN(n99) );
  INVD1 U638 ( .I(AddrW[0]), .ZN(n96) );
  INVD1 U639 ( .I(AddrW[2]), .ZN(n100) );
  AN2D1 U640 ( .A1(Write), .A2(AddrW[3]), .Z(n95) );
  INVD1 U641 ( .I(n490), .ZN(n489) );
  INVD1 U642 ( .I(Read), .ZN(n490) );
  INR2D1 U643 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INVD1 U644 ( .I(n476), .ZN(n475) );
  INVD1 U645 ( .I(ClockR), .ZN(n476) );
  INR2D1 U646 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U647 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_0 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n5,
         n7, n8, n9, n12;

  AO211D1 U8 ( .A1(n7), .A2(n8), .B(N8), .C(N5), .Z(n9) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n5), .QN(N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n5), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n12), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n12), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n5), .Q(\ClockInN[0] ), 
        .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n5), .QN(n7) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n12), .QN(n5) );
  INVD1 U3 ( .I(Reset), .ZN(n12) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n7), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n8), .A2(n7), .B(n9), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n8) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_0 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n17, n18, n19, n21, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_0_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_0_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_0_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n26), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n17), .CP(FastClock), .CDN(n26), .Q(ClockOut)
         );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n26), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n26), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n19), .CP(Sample), .SDN(n29), .Q(
        DivideFactor[4]), .QN(n41) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n18), .CP(Sample), .SDN(n29), .Q(
        DivideFactor[1]), .QN(n53) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n21), .CP(Sample), .SDN(n29), .Q(
        DivideFactor[0]), .QN(n51) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n29), 
        .Q(DivideFactor[3]), .QN(n46) );
  INVD1 U3 ( .I(n28), .ZN(n26) );
  INVD1 U4 ( .I(n28), .ZN(n27) );
  INVD1 U5 ( .I(n29), .ZN(n28) );
  INVD1 U6 ( .I(Reset), .ZN(n29) );
  AO222D0 U7 ( .A1(N27), .A2(n30), .B1(N35), .B2(n31), .C1(DivideFactor[0]), 
        .C2(n32), .Z(n21) );
  AO222D0 U8 ( .A1(N31), .A2(n30), .B1(N39), .B2(n31), .C1(DivideFactor[4]), 
        .C2(n32), .Z(n19) );
  AO222D0 U9 ( .A1(N28), .A2(n30), .B1(N36), .B2(n31), .C1(DivideFactor[1]), 
        .C2(n32), .Z(n18) );
  CKND0 U10 ( .CLK(N54), .CN(n32) );
  AN2D0 U11 ( .A1(n33), .A2(n34), .Z(n31) );
  AN3D0 U12 ( .A1(n35), .A2(n36), .A3(n37), .Z(n30) );
  CKXOR2D0 U13 ( .A1(ClockOut), .A2(n38), .Z(n17) );
  AO22D0 U14 ( .A1(N32), .A2(n37), .B1(N40), .B2(n33), .Z(N55) );
  MUX2ND0 U15 ( .I0(n39), .I1(n40), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U16 ( .A1(AdjustFreq[1]), .A2(n34), .ZN(n40) );
  ND3D0 U17 ( .A1(n41), .A2(n36), .A3(n42), .ZN(n34) );
  ND4D0 U18 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n42) );
  IND3D0 U19 ( .A1(AdjustFreq[1]), .B1(n36), .B2(n35), .ZN(n39) );
  CKND2D0 U20 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n35) );
  AO22D0 U21 ( .A1(N30), .A2(n37), .B1(N38), .B2(n33), .Z(N51) );
  AO22D0 U22 ( .A1(N29), .A2(n37), .B1(N37), .B2(n33), .Z(N49) );
  AN2D0 U23 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n33) );
  NR2D0 U24 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n37) );
  INR2D0 U25 ( .A1(N14), .B1(n38), .ZN(N21) );
  INR2D0 U26 ( .A1(N13), .B1(n38), .ZN(N20) );
  INR2D0 U27 ( .A1(N12), .B1(n38), .ZN(N19) );
  INR2D0 U28 ( .A1(N11), .B1(n38), .ZN(N18) );
  INR2D0 U29 ( .A1(N10), .B1(n38), .ZN(N17) );
  INR2D0 U30 ( .A1(N9), .B1(n38), .ZN(N16) );
  OA21D0 U31 ( .A1(FastDivvy[5]), .A2(n36), .B(n43), .Z(n38) );
  IOA22D0 U32 ( .B1(n44), .B2(n45), .A1(n36), .A2(FastDivvy[5]), .ZN(n43) );
  AOI221D0 U33 ( .A1(FastDivvy[4]), .A2(n41), .B1(FastDivvy[3]), .B2(n46), .C(
        n47), .ZN(n45) );
  AOI221D0 U34 ( .A1(DivideFactor[3]), .A2(n48), .B1(DivideFactor[2]), .B2(n49), .C(n50), .ZN(n47) );
  IAO21D0 U35 ( .A1(n49), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n50) );
  OAI32D0 U36 ( .A1(n51), .A2(FastDivvy[0]), .A3(n52), .B1(FastDivvy[1]), .B2(
        n53), .ZN(n49) );
  AN2D0 U37 ( .A1(FastDivvy[1]), .A2(n53), .Z(n52) );
  CKND0 U38 ( .CLK(FastDivvy[3]), .CN(n48) );
  NR2D0 U39 ( .A1(FastDivvy[4]), .A2(n41), .ZN(n44) );
  CKND0 U40 ( .CLK(DivideFactor[5]), .CN(n36) );
  CKND0 U41 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U42 ( .A1(WireD[5]), .A2(n27), .ZN(WireD[0]) );
endmodule


module MultiCounter_0 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_0_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module FIFOTop_AWid3_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [2:0] SM_ReadAddr;
  wire   [2:0] SM_WriteAddr;

  FIFOStateM_AWid3_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid3_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD1 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module SerEncoder_DWid32_1 ( SerOut, SerValid, FIFO_ReadReq, ParIn, F_Empty, 
        ParClk, SerClk, ParValid, Reset );
  input [31:0] ParIn;
  input F_Empty, ParClk, SerClk, ParValid, Reset;
  output SerOut, SerValid, FIFO_ReadReq;
  wire   N2, N3, N4, N5, N6, HalfParClkr, \Sh_N[5] , N8, N9, N10, N11, N12,
         N13, N23, N24, N25, N26, N27, N28, N29, N31, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80;
  wire   [31:0] InBuf;

  SerEncoder_DWid32_1_DW01_dec_0 \ShifterBlock/sub_132  ( .A({n3, n8, n2, n7, 
        n5, n4}), .SUM({N13, N12, N11, N10, N9, N8}) );
  DFCNQD1 SerValidr_reg ( .D(n35), .CP(n45), .CDN(n57), .Q(SerValid) );
  DFCNQD1 HalfParClkr_reg ( .D(n49), .CP(ParClk), .CDN(n54), .Q(HalfParClkr)
         );
  DFCNQD1 \InBuf_reg[30]  ( .D(N83), .CP(n48), .CDN(n54), .Q(InBuf[30]) );
  DFCNQD1 \InBuf_reg[29]  ( .D(N82), .CP(n48), .CDN(n54), .Q(InBuf[29]) );
  DFCNQD1 \InBuf_reg[26]  ( .D(N79), .CP(n48), .CDN(n55), .Q(InBuf[26]) );
  DFCNQD1 \InBuf_reg[25]  ( .D(N78), .CP(n47), .CDN(n55), .Q(InBuf[25]) );
  DFCNQD1 \InBuf_reg[22]  ( .D(N75), .CP(n47), .CDN(n55), .Q(InBuf[22]) );
  DFCNQD1 \InBuf_reg[21]  ( .D(N74), .CP(n47), .CDN(n55), .Q(InBuf[21]) );
  DFCNQD1 \InBuf_reg[18]  ( .D(N71), .CP(n47), .CDN(n56), .Q(InBuf[18]) );
  DFCNQD1 \InBuf_reg[17]  ( .D(N70), .CP(n47), .CDN(n56), .Q(InBuf[17]) );
  DFCNQD1 \InBuf_reg[14]  ( .D(N67), .CP(n46), .CDN(n56), .Q(InBuf[14]) );
  DFCNQD1 \InBuf_reg[13]  ( .D(N66), .CP(n46), .CDN(n56), .Q(InBuf[13]) );
  DFCNQD1 \InBuf_reg[10]  ( .D(N63), .CP(n46), .CDN(n56), .Q(InBuf[10]) );
  DFCNQD1 \InBuf_reg[9]  ( .D(N62), .CP(n46), .CDN(n56), .Q(InBuf[9]) );
  DFCNQD1 \InBuf_reg[6]  ( .D(N59), .CP(n45), .CDN(n57), .Q(InBuf[6]) );
  DFCNQD1 \InBuf_reg[5]  ( .D(N58), .CP(n45), .CDN(n57), .Q(InBuf[5]) );
  DFCNQD1 \InBuf_reg[2]  ( .D(N55), .CP(n45), .CDN(n57), .Q(InBuf[2]) );
  DFCNQD1 \InBuf_reg[1]  ( .D(N54), .CP(n45), .CDN(n57), .Q(InBuf[1]) );
  DFCNQD1 \InBuf_reg[31]  ( .D(N84), .CP(n48), .CDN(n54), .Q(InBuf[31]) );
  DFCNQD1 \InBuf_reg[28]  ( .D(N81), .CP(n48), .CDN(n55), .Q(InBuf[28]) );
  DFCNQD1 \InBuf_reg[27]  ( .D(N80), .CP(n48), .CDN(n55), .Q(InBuf[27]) );
  DFCNQD1 \InBuf_reg[24]  ( .D(N77), .CP(n47), .CDN(n55), .Q(InBuf[24]) );
  DFCNQD1 \InBuf_reg[23]  ( .D(N76), .CP(n47), .CDN(n55), .Q(InBuf[23]) );
  DFCNQD1 \InBuf_reg[20]  ( .D(N73), .CP(n47), .CDN(n55), .Q(InBuf[20]) );
  DFCNQD1 \InBuf_reg[19]  ( .D(N72), .CP(n47), .CDN(n55), .Q(InBuf[19]) );
  DFCNQD1 \InBuf_reg[16]  ( .D(N69), .CP(n46), .CDN(n56), .Q(InBuf[16]) );
  DFCNQD1 \InBuf_reg[15]  ( .D(N68), .CP(n46), .CDN(n56), .Q(InBuf[15]) );
  DFCNQD1 \InBuf_reg[12]  ( .D(N65), .CP(n46), .CDN(n56), .Q(InBuf[12]) );
  DFCNQD1 \InBuf_reg[11]  ( .D(N64), .CP(n46), .CDN(n56), .Q(InBuf[11]) );
  DFCNQD1 \InBuf_reg[8]  ( .D(N61), .CP(n46), .CDN(n57), .Q(InBuf[8]) );
  DFCNQD1 \InBuf_reg[7]  ( .D(N60), .CP(n45), .CDN(n57), .Q(InBuf[7]) );
  DFCNQD1 \InBuf_reg[4]  ( .D(N57), .CP(n45), .CDN(n57), .Q(InBuf[4]) );
  DFCNQD1 \InBuf_reg[3]  ( .D(N56), .CP(n45), .CDN(n57), .Q(InBuf[3]) );
  DFCNQD1 \InBuf_reg[0]  ( .D(N53), .CP(n45), .CDN(n57), .Q(InBuf[0]) );
  DFCNQD1 \Sh_N_reg[5]  ( .D(N13), .CP(SerClk), .CDN(n54), .Q(\Sh_N[5] ) );
  DFCNQD1 \Sh_N_reg[4]  ( .D(N12), .CP(SerClk), .CDN(n54), .Q(N6) );
  DFCNQD1 \Sh_N_reg[2]  ( .D(N10), .CP(SerClk), .CDN(n54), .Q(N4) );
  DFCNQD1 \Sh_N_reg[3]  ( .D(N11), .CP(SerClk), .CDN(n54), .Q(N5) );
  DFCNQD1 \Sh_N_reg[1]  ( .D(N9), .CP(SerClk), .CDN(n54), .Q(N3) );
  DFCNQD1 \Sh_N_reg[0]  ( .D(N8), .CP(SerClk), .CDN(n54), .Q(N2) );
  DFCNQD1 SerOutr_reg ( .D(n1), .CP(SerClk), .CDN(n56), .Q(SerOut) );
  BUFFD0 U3 ( .I(N31), .Z(n1) );
  CKBD0 U4 ( .CLK(N3), .C(n5) );
  BUFFD0 U5 ( .I(n9), .Z(n2) );
  CKBD0 U6 ( .CLK(n6), .C(n3) );
  CKBXD0 U7 ( .I(\Sh_N[5] ), .Z(n6) );
  CKBD0 U8 ( .CLK(N2), .C(n4) );
  OR2D0 U9 ( .A1(n4), .A2(n5), .Z(n64) );
  CKND2D0 U10 ( .A1(n5), .A2(n4), .ZN(n65) );
  BUFFD0 U11 ( .I(N4), .Z(n7) );
  CKBXD0 U12 ( .I(N6), .Z(n8) );
  BUFFD0 U13 ( .I(N5), .Z(n9) );
  BUFFD1 U14 ( .I(n51), .Z(n58) );
  INVD1 U15 ( .I(n59), .ZN(n57) );
  BUFFD1 U16 ( .I(n51), .Z(n59) );
  INVD1 U17 ( .I(n60), .ZN(n56) );
  BUFFD1 U18 ( .I(n52), .Z(n60) );
  INVD1 U19 ( .I(n61), .ZN(n55) );
  BUFFD1 U20 ( .I(n52), .Z(n61) );
  BUFFD1 U21 ( .I(Reset), .Z(n51) );
  BUFFD1 U22 ( .I(Reset), .Z(n52) );
  INVD1 U23 ( .I(n62), .ZN(n54) );
  BUFFD1 U24 ( .I(n53), .Z(n62) );
  BUFFD1 U25 ( .I(Reset), .Z(n53) );
  INVD1 U26 ( .I(n40), .ZN(n35) );
  INVD1 U27 ( .I(n40), .ZN(n36) );
  INVD1 U28 ( .I(n39), .ZN(n37) );
  INVD1 U29 ( .I(n49), .ZN(n45) );
  INVD1 U30 ( .I(n49), .ZN(n46) );
  INVD1 U31 ( .I(n50), .ZN(n47) );
  INVD1 U32 ( .I(n50), .ZN(n48) );
  INVD1 U33 ( .I(n39), .ZN(n38) );
  INVD1 U34 ( .I(n64), .ZN(n63) );
  INVD1 U35 ( .I(n42), .ZN(n40) );
  INVD1 U36 ( .I(n43), .ZN(n49) );
  INVD1 U37 ( .I(n42), .ZN(n39) );
  INVD1 U38 ( .I(n43), .ZN(n50) );
  AN2D1 U39 ( .A1(n7), .A2(n63), .Z(N26) );
  MUX2D0 U40 ( .I0(n15), .I1(n16), .S(n7), .Z(n31) );
  MUX4ND0 U41 ( .I0(InBuf[8]), .I1(InBuf[9]), .I2(InBuf[10]), .I3(InBuf[11]), 
        .S0(N2), .S1(N3), .ZN(n15) );
  MUX4ND0 U42 ( .I0(InBuf[12]), .I1(InBuf[13]), .I2(InBuf[14]), .I3(InBuf[15]), 
        .S0(N2), .S1(N3), .ZN(n16) );
  MUX2D0 U43 ( .I0(n17), .I1(n18), .S(n7), .Z(n29) );
  MUX4ND0 U44 ( .I0(InBuf[16]), .I1(InBuf[17]), .I2(InBuf[18]), .I3(InBuf[19]), 
        .S0(N2), .S1(N3), .ZN(n17) );
  MUX4ND0 U45 ( .I0(InBuf[20]), .I1(InBuf[21]), .I2(InBuf[22]), .I3(InBuf[23]), 
        .S0(N2), .S1(N3), .ZN(n18) );
  MUX2D0 U46 ( .I0(n19), .I1(n20), .S(n7), .Z(n27) );
  MUX4ND0 U47 ( .I0(InBuf[24]), .I1(InBuf[25]), .I2(InBuf[26]), .I3(InBuf[27]), 
        .S0(N2), .S1(N3), .ZN(n19) );
  MUX4ND0 U48 ( .I0(InBuf[28]), .I1(InBuf[29]), .I2(InBuf[30]), .I3(InBuf[31]), 
        .S0(N2), .S1(N3), .ZN(n20) );
  MUX2D0 U49 ( .I0(n21), .I1(n22), .S(n7), .Z(n33) );
  MUX4ND0 U50 ( .I0(InBuf[0]), .I1(InBuf[1]), .I2(InBuf[2]), .I3(InBuf[3]), 
        .S0(N2), .S1(N3), .ZN(n21) );
  MUX4ND0 U51 ( .I0(InBuf[4]), .I1(InBuf[5]), .I2(InBuf[6]), .I3(InBuf[7]), 
        .S0(N2), .S1(N3), .ZN(n22) );
  NR2D1 U52 ( .A1(n65), .A2(n7), .ZN(N24) );
  INVD1 U53 ( .I(n41), .ZN(n42) );
  INVD1 U54 ( .I(N85), .ZN(n41) );
  INVD1 U55 ( .I(n44), .ZN(n43) );
  INVD1 U56 ( .I(HalfParClkr), .ZN(n44) );
  MUX2ND0 U57 ( .I0(n23), .I1(n24), .S(n8), .ZN(N29) );
  MUX2ND0 U58 ( .I0(n25), .I1(n26), .S(n8), .ZN(N27) );
  MUX2ND0 U59 ( .I0(n24), .I1(n23), .S(n8), .ZN(N25) );
  MUX2ND0 U60 ( .I0(n26), .I1(n25), .S(n8), .ZN(N23) );
  CKND1 U61 ( .CLK(n27), .CN(n28) );
  CKND1 U62 ( .CLK(n29), .CN(n30) );
  MUX2ND0 U63 ( .I0(n30), .I1(n28), .S(n9), .ZN(n24) );
  CKND1 U64 ( .CLK(n31), .CN(n32) );
  CKND1 U65 ( .CLK(n33), .CN(n34) );
  MUX2ND0 U66 ( .I0(n34), .I1(n32), .S(n9), .ZN(n23) );
  MUX2ND0 U67 ( .I0(n28), .I1(n34), .S(n9), .ZN(n26) );
  MUX2ND0 U68 ( .I0(n32), .I1(n30), .S(n9), .ZN(n25) );
  MUX2ND0 U69 ( .I0(n65), .I1(n64), .S(n7), .ZN(N28) );
  AN2D0 U70 ( .A1(ParIn[31]), .A2(n38), .Z(N84) );
  AN2D0 U71 ( .A1(ParIn[30]), .A2(n38), .Z(N83) );
  AN2D0 U72 ( .A1(ParIn[29]), .A2(n38), .Z(N82) );
  AN2D0 U73 ( .A1(ParIn[28]), .A2(n38), .Z(N81) );
  AN2D0 U74 ( .A1(ParIn[27]), .A2(n37), .Z(N80) );
  AN2D0 U75 ( .A1(ParIn[26]), .A2(n37), .Z(N79) );
  AN2D0 U76 ( .A1(ParIn[25]), .A2(n37), .Z(N78) );
  AN2D0 U77 ( .A1(ParIn[24]), .A2(n37), .Z(N77) );
  AN2D0 U78 ( .A1(ParIn[23]), .A2(n37), .Z(N76) );
  AN2D0 U79 ( .A1(ParIn[22]), .A2(n37), .Z(N75) );
  AN2D0 U80 ( .A1(ParIn[21]), .A2(n37), .Z(N74) );
  AN2D0 U81 ( .A1(ParIn[20]), .A2(n37), .Z(N73) );
  AN2D0 U82 ( .A1(ParIn[19]), .A2(n37), .Z(N72) );
  AN2D0 U83 ( .A1(ParIn[18]), .A2(n37), .Z(N71) );
  AN2D0 U84 ( .A1(ParIn[17]), .A2(n36), .Z(N70) );
  AN2D0 U85 ( .A1(ParIn[16]), .A2(n36), .Z(N69) );
  AN2D0 U86 ( .A1(ParIn[15]), .A2(n36), .Z(N68) );
  AN2D0 U87 ( .A1(ParIn[14]), .A2(n36), .Z(N67) );
  AN2D0 U88 ( .A1(ParIn[13]), .A2(n36), .Z(N66) );
  AN2D0 U89 ( .A1(ParIn[12]), .A2(n36), .Z(N65) );
  AN2D0 U90 ( .A1(ParIn[11]), .A2(n36), .Z(N64) );
  AN2D0 U91 ( .A1(ParIn[10]), .A2(n36), .Z(N63) );
  AN2D0 U92 ( .A1(ParIn[9]), .A2(n36), .Z(N62) );
  AN2D0 U93 ( .A1(ParIn[8]), .A2(n36), .Z(N61) );
  AN2D0 U94 ( .A1(ParIn[7]), .A2(n35), .Z(N60) );
  AN2D0 U95 ( .A1(ParIn[6]), .A2(n35), .Z(N59) );
  AN2D0 U96 ( .A1(ParIn[5]), .A2(n35), .Z(N58) );
  AN2D0 U97 ( .A1(ParIn[4]), .A2(n35), .Z(N57) );
  AN2D0 U98 ( .A1(ParIn[3]), .A2(n35), .Z(N56) );
  AN2D0 U99 ( .A1(ParIn[2]), .A2(n35), .Z(N55) );
  AN2D0 U100 ( .A1(ParIn[1]), .A2(n35), .Z(N54) );
  AN2D0 U101 ( .A1(ParIn[0]), .A2(n35), .Z(N53) );
  IND2D0 U102 ( .A1(n66), .B1(n67), .ZN(N31) );
  OAI21D0 U103 ( .A1(N23), .A2(n68), .B(n69), .ZN(n67) );
  MUX2ND0 U104 ( .I0(n70), .I1(n71), .S(n68), .ZN(n69) );
  MUX3ND0 U105 ( .I0(N25), .I1(n72), .I2(N24), .S0(n3), .S1(n73), .ZN(n71) );
  NR2D0 U106 ( .A1(n3), .A2(n9), .ZN(n73) );
  MUX2D0 U107 ( .I0(n74), .I1(N26), .S(n75), .Z(n72) );
  NR2D0 U108 ( .A1(n8), .A2(n9), .ZN(n75) );
  INR2D0 U109 ( .A1(N27), .B1(n8), .ZN(n74) );
  CKND0 U110 ( .CLK(n2), .CN(n70) );
  CKND2D0 U111 ( .A1(n76), .A2(n77), .ZN(n68) );
  MUX2ND0 U112 ( .I0(n78), .I1(n79), .S(n2), .ZN(n66) );
  CKND2D0 U113 ( .A1(N29), .A2(n80), .ZN(n79) );
  CKND2D0 U114 ( .A1(N28), .A2(n80), .ZN(n78) );
  NR2D0 U115 ( .A1(n77), .A2(n76), .ZN(n80) );
  CKND0 U116 ( .CLK(n8), .CN(n76) );
  CKND0 U117 ( .CLK(n3), .CN(n77) );
  INR3D0 U118 ( .A1(n35), .B1(n58), .B2(n49), .ZN(FIFO_ReadReq) );
  INR2D0 U119 ( .A1(ParValid), .B1(F_Empty), .ZN(N85) );
endmodule


module SerialTx_1 ( SerOut, SerClk, SerIn, ParClk, Reset );
  input SerIn, ParClk, Reset;
  output SerOut, SerClk;
  wire   n2;

  PLLTop_2 PLL_TxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerIn), .Z(SerOut) );
endmodule


module FIFOTop_AWid4_DWid32_1 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3;
  wire   [3:0] SM_ReadAddr;
  wire   [3:0] SM_WriteAddr;

  FIFOStateM_AWid4_1 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(
        SM_WriteAddr), .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(
        SM_MemReadCmd), .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), 
        .WriteReq(WriteIn), .ClkR(ClkR), .ClkW(ClkW), .Reset(n2) );
  DPMem1kx32_AWid4_DWid32_1 FIFO_Mem1 ( .DataO(Dout), .DataI(Din), .AddrR(
        SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(n2) );
  INVD1 U2 ( .I(n3), .ZN(n2) );
  INVD1 U3 ( .I(Reseter), .ZN(n3) );
  BUFFD1 U4 ( .I(SM_MemReadCmd), .Z(n1) );
  TIEH U5 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32_1 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   SerClock, N30, N31, N32, N33, N34, N37, N38, N39, N40, N41, N42, N43,
         N47, n84, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453;
  wire   [3:0] ParValidTimer;
  wire   [31:0] Decoder;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  MOAI22D1 U17 ( .A1(n266), .A2(n426), .B1(n268), .B2(Decoder[31]), .ZN(n389)
         );
  MOAI22D1 U18 ( .A1(n266), .A2(n425), .B1(n268), .B2(Decoder[30]), .ZN(n388)
         );
  MOAI22D1 U19 ( .A1(n266), .A2(n424), .B1(n268), .B2(Decoder[29]), .ZN(n387)
         );
  MOAI22D1 U20 ( .A1(n266), .A2(n423), .B1(n268), .B2(Decoder[28]), .ZN(n386)
         );
  MOAI22D1 U21 ( .A1(n266), .A2(n422), .B1(n267), .B2(Decoder[27]), .ZN(n385)
         );
  MOAI22D1 U22 ( .A1(n266), .A2(n421), .B1(n267), .B2(Decoder[26]), .ZN(n384)
         );
  MOAI22D1 U23 ( .A1(n266), .A2(n420), .B1(n267), .B2(Decoder[25]), .ZN(n383)
         );
  MOAI22D1 U24 ( .A1(n266), .A2(n419), .B1(n267), .B2(Decoder[24]), .ZN(n382)
         );
  MOAI22D1 U25 ( .A1(n266), .A2(n418), .B1(n267), .B2(Decoder[23]), .ZN(n381)
         );
  MOAI22D1 U26 ( .A1(n266), .A2(n417), .B1(n267), .B2(Decoder[22]), .ZN(n380)
         );
  MOAI22D1 U27 ( .A1(n266), .A2(n416), .B1(n267), .B2(Decoder[21]), .ZN(n379)
         );
  MOAI22D1 U28 ( .A1(n266), .A2(n415), .B1(n266), .B2(Decoder[20]), .ZN(n378)
         );
  MOAI22D1 U29 ( .A1(n266), .A2(n414), .B1(n267), .B2(Decoder[19]), .ZN(n377)
         );
  MOAI22D1 U30 ( .A1(n266), .A2(n413), .B1(n267), .B2(Decoder[18]), .ZN(n376)
         );
  MOAI22D1 U31 ( .A1(n266), .A2(n412), .B1(n267), .B2(Decoder[17]), .ZN(n375)
         );
  MOAI22D1 U32 ( .A1(n266), .A2(n411), .B1(n267), .B2(Decoder[16]), .ZN(n374)
         );
  MOAI22D1 U33 ( .A1(n266), .A2(n410), .B1(n267), .B2(Decoder[15]), .ZN(n373)
         );
  MOAI22D1 U34 ( .A1(n266), .A2(n409), .B1(n267), .B2(Decoder[14]), .ZN(n372)
         );
  MOAI22D1 U35 ( .A1(n265), .A2(n408), .B1(n267), .B2(Decoder[13]), .ZN(n371)
         );
  MOAI22D1 U36 ( .A1(n265), .A2(n407), .B1(n267), .B2(Decoder[12]), .ZN(n370)
         );
  MOAI22D1 U37 ( .A1(n265), .A2(n406), .B1(n267), .B2(Decoder[11]), .ZN(n369)
         );
  MOAI22D1 U38 ( .A1(n265), .A2(n405), .B1(n267), .B2(Decoder[10]), .ZN(n368)
         );
  MOAI22D1 U39 ( .A1(n265), .A2(n404), .B1(n267), .B2(Decoder[9]), .ZN(n367)
         );
  MOAI22D1 U40 ( .A1(n265), .A2(n403), .B1(n267), .B2(Decoder[8]), .ZN(n366)
         );
  MOAI22D1 U41 ( .A1(n265), .A2(n402), .B1(n268), .B2(Decoder[7]), .ZN(n365)
         );
  MOAI22D1 U42 ( .A1(n265), .A2(n401), .B1(n267), .B2(Decoder[6]), .ZN(n364)
         );
  MOAI22D1 U43 ( .A1(n265), .A2(n400), .B1(n268), .B2(Decoder[5]), .ZN(n363)
         );
  MOAI22D1 U44 ( .A1(n265), .A2(n399), .B1(n268), .B2(Decoder[4]), .ZN(n362)
         );
  MOAI22D1 U45 ( .A1(n265), .A2(n398), .B1(n268), .B2(Decoder[3]), .ZN(n361)
         );
  MOAI22D1 U46 ( .A1(n265), .A2(n397), .B1(n268), .B2(Decoder[2]), .ZN(n360)
         );
  MOAI22D1 U47 ( .A1(n265), .A2(n396), .B1(n268), .B2(Decoder[1]), .ZN(n359)
         );
  MOAI22D1 U48 ( .A1(n266), .A2(n395), .B1(n268), .B2(Decoder[0]), .ZN(n358)
         );
  OR3D1 U92 ( .A1(FrameSR[55]), .A2(FrameSR[54]), .A3(FrameSR[53]), .Z(n434)
         );
  OR3D1 U94 ( .A1(FrameSR[39]), .A2(FrameSR[38]), .A3(FrameSR[37]), .Z(n433)
         );
  OR3D1 U96 ( .A1(FrameSR[32]), .A2(FrameSR[23]), .A3(FrameSR[22]), .Z(n432)
         );
  OA21D1 U99 ( .A1(n430), .A2(n429), .B(SerValid), .Z(N43) );
  OR2D1 U101 ( .A1(Count32[1]), .A2(Count32[0]), .Z(n428) );
  DesDecoder_DWid32_1_DW01_inc_0 \ClkGen/add_206  ( .A(Count32), .SUM({N34, 
        N33, N32, N31, N30}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(FrameSR[62]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[63]) );
  DFNCND1 \FrameSR_reg[22]  ( .D(FrameSR[21]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[22]) );
  DFNCND1 \FrameSR_reg[23]  ( .D(FrameSR[22]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[23]) );
  DFNCND1 \FrameSR_reg[37]  ( .D(FrameSR[36]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[37]) );
  DFNCND1 \FrameSR_reg[38]  ( .D(FrameSR[37]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[38]) );
  DFNCND1 \FrameSR_reg[53]  ( .D(FrameSR[52]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[53]) );
  DFNCND1 \FrameSR_reg[54]  ( .D(FrameSR[53]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[54]) );
  DFNCND1 \FrameSR_reg[32]  ( .D(FrameSR[31]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[32]) );
  DFNCND1 \FrameSR_reg[39]  ( .D(FrameSR[38]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[39]) );
  DFNCND1 \FrameSR_reg[55]  ( .D(FrameSR[54]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[55]) );
  DFNCND1 \FrameSR_reg[8]  ( .D(FrameSR[7]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[8]) );
  DFNCND1 \FrameSR_reg[9]  ( .D(FrameSR[8]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[9]) );
  DFNCND1 \FrameSR_reg[10]  ( .D(FrameSR[9]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[10]) );
  DFNCND1 \FrameSR_reg[11]  ( .D(FrameSR[10]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[11]) );
  DFNCND1 \FrameSR_reg[12]  ( .D(FrameSR[11]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[12]) );
  DFNCND1 \FrameSR_reg[13]  ( .D(FrameSR[12]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[13]) );
  DFNCND1 \FrameSR_reg[14]  ( .D(FrameSR[13]), .CPN(n296), .CDN(n299), .Q(
        FrameSR[14]) );
  DFNCND1 \FrameSR_reg[15]  ( .D(FrameSR[14]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[15]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(FrameSR[18]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[19]) );
  DFNCND1 \FrameSR_reg[24]  ( .D(FrameSR[23]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[24]) );
  DFNCND1 \FrameSR_reg[25]  ( .D(FrameSR[24]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[25]) );
  DFNCND1 \FrameSR_reg[26]  ( .D(FrameSR[25]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[26]) );
  DFNCND1 \FrameSR_reg[27]  ( .D(FrameSR[26]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[27]) );
  DFNCND1 \FrameSR_reg[28]  ( .D(FrameSR[27]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[28]) );
  DFNCND1 \FrameSR_reg[29]  ( .D(FrameSR[28]), .CPN(n294), .CDN(n300), .Q(
        FrameSR[29]) );
  DFNCND1 \FrameSR_reg[30]  ( .D(FrameSR[29]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[30]) );
  DFNCND1 \FrameSR_reg[31]  ( .D(FrameSR[30]), .CPN(n294), .CDN(n301), .Q(
        FrameSR[31]) );
  DFNCND1 \FrameSR_reg[40]  ( .D(FrameSR[39]), .CPN(n293), .CDN(n302), .Q(
        FrameSR[40]) );
  DFNCND1 \FrameSR_reg[41]  ( .D(FrameSR[40]), .CPN(n293), .CDN(n302), .Q(
        FrameSR[41]) );
  DFNCND1 \FrameSR_reg[42]  ( .D(FrameSR[41]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[42]) );
  DFNCND1 \FrameSR_reg[43]  ( .D(FrameSR[42]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[43]) );
  DFNCND1 \FrameSR_reg[44]  ( .D(FrameSR[43]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[44]) );
  DFNCND1 \FrameSR_reg[45]  ( .D(FrameSR[44]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[45]) );
  DFNCND1 \FrameSR_reg[46]  ( .D(FrameSR[45]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[46]) );
  DFNCND1 \FrameSR_reg[47]  ( .D(FrameSR[46]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[47]) );
  DFNCND1 \FrameSR_reg[56]  ( .D(FrameSR[55]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[56]) );
  DFNCND1 \FrameSR_reg[57]  ( .D(FrameSR[56]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[57]) );
  DFNCND1 \FrameSR_reg[58]  ( .D(FrameSR[57]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[58]) );
  DFNCND1 \FrameSR_reg[59]  ( .D(FrameSR[58]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[59]) );
  DFNCND1 \FrameSR_reg[60]  ( .D(FrameSR[59]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[60]) );
  DFNCND1 \FrameSR_reg[61]  ( .D(FrameSR[60]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[61]) );
  DFNCND1 \FrameSR_reg[62]  ( .D(FrameSR[61]), .CPN(n290), .CDN(n304), .Q(
        FrameSR[62]) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n297), .CDN(n298), .Q(FrameSR[0])
         );
  DFNCND1 \FrameSR_reg[4]  ( .D(FrameSR[3]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(FrameSR[19]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(FrameSR[33]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(FrameSR[48]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(FrameSR[1]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(FrameSR[5]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(FrameSR[17]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(FrameSR[32]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(FrameSR[47]), .CPN(n292), .CDN(n302), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(FrameSR[0]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(FrameSR[2]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(FrameSR[4]), .CPN(n297), .CDN(n298), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(FrameSR[6]), .CPN(n296), .CDN(n298), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(FrameSR[20]), .CPN(n295), .CDN(n300), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(FrameSR[34]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(FrameSR[49]), .CPN(n292), .CDN(n303), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[51]  ( .D(FrameSR[50]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[51]) );
  DFNCND1 \FrameSR_reg[36]  ( .D(FrameSR[35]), .CPN(n293), .CDN(n301), .Q(
        FrameSR[36]) );
  DFNCND1 \FrameSR_reg[52]  ( .D(FrameSR[51]), .CPN(n291), .CDN(n303), .Q(
        FrameSR[52]) );
  DFNCND1 \FrameSR_reg[17]  ( .D(FrameSR[16]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[17]) );
  DFNCND1 \FrameSR_reg[16]  ( .D(FrameSR[15]), .CPN(n295), .CDN(n299), .Q(
        FrameSR[16]) );
  EDFCNQD1 \Count32_reg[4]  ( .D(N42), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[4]) );
  DFNCND1 \Decoder_reg[31]  ( .D(n326), .CPN(n290), .CDN(n304), .Q(Decoder[31]) );
  DFNCND1 \Decoder_reg[30]  ( .D(n327), .CPN(n290), .CDN(n304), .Q(Decoder[30]) );
  DFNCND1 \Decoder_reg[29]  ( .D(n328), .CPN(n290), .CDN(n304), .Q(Decoder[29]) );
  DFNCND1 \Decoder_reg[28]  ( .D(n329), .CPN(n290), .CDN(n304), .Q(Decoder[28]) );
  DFNCND1 \Decoder_reg[27]  ( .D(n330), .CPN(n290), .CDN(n304), .Q(Decoder[27]) );
  DFNCND1 \Decoder_reg[26]  ( .D(n331), .CPN(n289), .CDN(n304), .Q(Decoder[26]) );
  DFNCND1 \Decoder_reg[25]  ( .D(n332), .CPN(n289), .CDN(n305), .Q(Decoder[25]) );
  DFNCND1 \Decoder_reg[24]  ( .D(n333), .CPN(n289), .CDN(n305), .Q(Decoder[24]) );
  DFNCND1 \Decoder_reg[23]  ( .D(n334), .CPN(n289), .CDN(n305), .Q(Decoder[23]) );
  DFNCND1 \Decoder_reg[22]  ( .D(n335), .CPN(n289), .CDN(n305), .Q(Decoder[22]) );
  DFNCND1 \Decoder_reg[21]  ( .D(n336), .CPN(n289), .CDN(n305), .Q(Decoder[21]) );
  DFNCND1 \Decoder_reg[20]  ( .D(n337), .CPN(n289), .CDN(n305), .Q(Decoder[20]) );
  DFNCND1 \Decoder_reg[19]  ( .D(n338), .CPN(n289), .CDN(n305), .Q(Decoder[19]) );
  DFNCND1 \Decoder_reg[18]  ( .D(n339), .CPN(n289), .CDN(n305), .Q(Decoder[18]) );
  DFNCND1 \Decoder_reg[17]  ( .D(n340), .CPN(n288), .CDN(n305), .Q(Decoder[17]) );
  DFNCND1 \Decoder_reg[16]  ( .D(n341), .CPN(n288), .CDN(n305), .Q(Decoder[16]) );
  DFNCND1 \Decoder_reg[15]  ( .D(n342), .CPN(n288), .CDN(n306), .Q(Decoder[15]) );
  DFNCND1 \Decoder_reg[14]  ( .D(n343), .CPN(n288), .CDN(n306), .Q(Decoder[14]) );
  DFNCND1 \Decoder_reg[13]  ( .D(n344), .CPN(n288), .CDN(n306), .Q(Decoder[13]) );
  DFNCND1 \Decoder_reg[12]  ( .D(n345), .CPN(n288), .CDN(n306), .Q(Decoder[12]) );
  DFNCND1 \Decoder_reg[11]  ( .D(n346), .CPN(n288), .CDN(n306), .Q(Decoder[11]) );
  DFNCND1 \Decoder_reg[10]  ( .D(n347), .CPN(n288), .CDN(n306), .Q(Decoder[10]) );
  DFNCND1 \Decoder_reg[9]  ( .D(n348), .CPN(n288), .CDN(n306), .Q(Decoder[9])
         );
  DFNCND1 \Decoder_reg[8]  ( .D(n349), .CPN(n287), .CDN(n306), .Q(Decoder[8])
         );
  DFNCND1 \Decoder_reg[7]  ( .D(n350), .CPN(n287), .CDN(n306), .Q(Decoder[7])
         );
  DFNCND1 \Decoder_reg[6]  ( .D(n351), .CPN(n287), .CDN(n306), .Q(Decoder[6])
         );
  DFNCND1 \Decoder_reg[5]  ( .D(n352), .CPN(n287), .CDN(n307), .Q(Decoder[5])
         );
  DFNCND1 \Decoder_reg[4]  ( .D(n353), .CPN(n287), .CDN(n307), .Q(Decoder[4])
         );
  DFNCND1 \Decoder_reg[3]  ( .D(n354), .CPN(n287), .CDN(n307), .Q(Decoder[3])
         );
  DFNCND1 \Decoder_reg[2]  ( .D(n355), .CPN(n287), .CDN(n307), .Q(Decoder[2])
         );
  DFNCND1 \Decoder_reg[1]  ( .D(n356), .CPN(n287), .CDN(n307), .Q(Decoder[1])
         );
  DFNCND1 \Decoder_reg[0]  ( .D(n357), .CPN(n287), .CDN(n307), .Q(Decoder[0])
         );
  DFNCND1 \ParValidTimer_reg[1]  ( .D(n391), .CPN(n283), .CDN(n311), .Q(
        ParValidTimer[1]) );
  EDFCNQD1 \Count32_reg[1]  ( .D(N39), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[1]) );
  DFNCND1 \ParValidTimer_reg[0]  ( .D(n390), .CPN(n283), .CDN(n311), .Q(
        ParValidTimer[0]) );
  EDFCNQD1 \Count32_reg[3]  ( .D(N41), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[3]) );
  EDFCNQD1 \Count32_reg[2]  ( .D(N40), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[2]) );
  EDFCNQD1 \Count32_reg[0]  ( .D(N38), .E(SerValid), .CP(n282), .CDN(n311), 
        .Q(Count32[0]) );
  DFNCND1 \ParOutr_reg[2]  ( .D(n360), .CPN(n286), .CDN(n308), .Q(ParOut[2]), 
        .QN(n397) );
  DFNCND1 \ParOutr_reg[1]  ( .D(n359), .CPN(n286), .CDN(n307), .Q(ParOut[1]), 
        .QN(n396) );
  EDFCNQD1 ParClkr_reg ( .D(N37), .E(N43), .CP(n282), .CDN(n311), .Q(ParClk)
         );
  DFNCND1 \ParOutr_reg[0]  ( .D(n358), .CPN(n286), .CDN(n307), .Q(ParOut[0]), 
        .QN(n395) );
  DFNCND1 \ParOutr_reg[5]  ( .D(n363), .CPN(n286), .CDN(n308), .Q(ParOut[5]), 
        .QN(n400) );
  DFNCND1 \ParOutr_reg[12]  ( .D(n370), .CPN(n285), .CDN(n309), .Q(ParOut[12]), 
        .QN(n407) );
  DFNCND1 \ParOutr_reg[19]  ( .D(n377), .CPN(n284), .CDN(n309), .Q(ParOut[19]), 
        .QN(n414) );
  DFNCND1 \ParOutr_reg[6]  ( .D(n364), .CPN(n286), .CDN(n308), .Q(ParOut[6]), 
        .QN(n401) );
  DFNCND1 \ParOutr_reg[9]  ( .D(n367), .CPN(n285), .CDN(n308), .Q(ParOut[9]), 
        .QN(n404) );
  DFNCND1 \ParOutr_reg[13]  ( .D(n371), .CPN(n285), .CDN(n309), .Q(ParOut[13]), 
        .QN(n408) );
  DFNCND1 \ParOutr_reg[16]  ( .D(n374), .CPN(n284), .CDN(n309), .Q(ParOut[16]), 
        .QN(n411) );
  DFNCND1 \ParOutr_reg[20]  ( .D(n378), .CPN(n284), .CDN(n309), .Q(ParOut[20]), 
        .QN(n415) );
  DFNCND1 \ParOutr_reg[23]  ( .D(n381), .CPN(n284), .CDN(n310), .Q(ParOut[23]), 
        .QN(n418) );
  DFNCND1 \ParOutr_reg[24]  ( .D(n382), .CPN(n284), .CDN(n310), .Q(ParOut[24]), 
        .QN(n419) );
  DFNCND1 \ParOutr_reg[27]  ( .D(n385), .CPN(n283), .CDN(n310), .Q(ParOut[27]), 
        .QN(n422) );
  DFNCND1 \ParOutr_reg[28]  ( .D(n386), .CPN(n283), .CDN(n310), .Q(ParOut[28]), 
        .QN(n423) );
  DFNCND1 \ParOutr_reg[31]  ( .D(n389), .CPN(n283), .CDN(n310), .Q(ParOut[31]), 
        .QN(n426) );
  DFNCND1 \ParOutr_reg[3]  ( .D(n361), .CPN(n286), .CDN(n308), .Q(ParOut[3]), 
        .QN(n398) );
  DFNCND1 \ParOutr_reg[4]  ( .D(n362), .CPN(n286), .CDN(n308), .Q(ParOut[4]), 
        .QN(n399) );
  DFNCND1 \ParOutr_reg[10]  ( .D(n368), .CPN(n285), .CDN(n308), .Q(ParOut[10]), 
        .QN(n405) );
  DFNCND1 \ParOutr_reg[11]  ( .D(n369), .CPN(n285), .CDN(n308), .Q(ParOut[11]), 
        .QN(n406) );
  DFNCND1 \ParOutr_reg[17]  ( .D(n375), .CPN(n284), .CDN(n309), .Q(ParOut[17]), 
        .QN(n412) );
  DFNCND1 \ParOutr_reg[18]  ( .D(n376), .CPN(n284), .CDN(n309), .Q(ParOut[18]), 
        .QN(n413) );
  DFNCND1 \ParOutr_reg[7]  ( .D(n365), .CPN(n285), .CDN(n308), .Q(ParOut[7]), 
        .QN(n402) );
  DFNCND1 \ParOutr_reg[8]  ( .D(n366), .CPN(n285), .CDN(n308), .Q(ParOut[8]), 
        .QN(n403) );
  DFNCND1 \ParOutr_reg[14]  ( .D(n372), .CPN(n285), .CDN(n309), .Q(ParOut[14]), 
        .QN(n409) );
  DFNCND1 \ParOutr_reg[15]  ( .D(n373), .CPN(n285), .CDN(n309), .Q(ParOut[15]), 
        .QN(n410) );
  DFNCND1 \ParOutr_reg[21]  ( .D(n379), .CPN(n284), .CDN(n309), .Q(ParOut[21]), 
        .QN(n416) );
  DFNCND1 \ParOutr_reg[22]  ( .D(n380), .CPN(n284), .CDN(n310), .Q(ParOut[22]), 
        .QN(n417) );
  DFNCND1 \ParOutr_reg[25]  ( .D(n383), .CPN(n283), .CDN(n310), .Q(ParOut[25]), 
        .QN(n420) );
  DFNCND1 \ParOutr_reg[26]  ( .D(n384), .CPN(n283), .CDN(n310), .Q(ParOut[26]), 
        .QN(n421) );
  DFNCND1 \ParOutr_reg[29]  ( .D(n387), .CPN(n283), .CDN(n310), .Q(ParOut[29]), 
        .QN(n424) );
  DFNCND1 \ParOutr_reg[30]  ( .D(n388), .CPN(n283), .CDN(n310), .Q(ParOut[30]), 
        .QN(n425) );
  DFNCND1 ParValidr_reg ( .D(n394), .CPN(n282), .CDN(n311), .Q(ParValid), .QN(
        n427) );
  DFNCND1 doParSync_reg ( .D(N47), .CPN(n286), .CDN(n322), .Q(n429), .QN(n453)
         );
  DFNCND1 UnLoad_reg ( .D(n258), .CPN(n286), .CDN(n322), .Q(n451), .QN(n324)
         );
  DFNCND1 \ParValidTimer_reg[3]  ( .D(n393), .CPN(n282), .CDN(n322), .QN(n323)
         );
  DFNCND1 \ParValidTimer_reg[2]  ( .D(n392), .CPN(n282), .CDN(n322), .QN(n325)
         );
  BUFFD1 U3 ( .I(n313), .Z(n309) );
  BUFFD1 U4 ( .I(n313), .Z(n308) );
  BUFFD1 U5 ( .I(n314), .Z(n307) );
  BUFFD1 U6 ( .I(n314), .Z(n306) );
  BUFFD1 U7 ( .I(n315), .Z(n305) );
  BUFFD1 U8 ( .I(n315), .Z(n304) );
  BUFFD1 U9 ( .I(n316), .Z(n303) );
  BUFFD1 U10 ( .I(n316), .Z(n302) );
  BUFFD1 U11 ( .I(n317), .Z(n301) );
  BUFFD1 U12 ( .I(n317), .Z(n300) );
  BUFFD1 U13 ( .I(n318), .Z(n299) );
  BUFFD1 U14 ( .I(n318), .Z(n298) );
  BUFFD1 U15 ( .I(n312), .Z(n311) );
  BUFFD1 U16 ( .I(n312), .Z(n310) );
  BUFFD1 U49 ( .I(n320), .Z(n313) );
  BUFFD1 U50 ( .I(n320), .Z(n314) );
  BUFFD1 U51 ( .I(n320), .Z(n315) );
  BUFFD1 U52 ( .I(n319), .Z(n316) );
  BUFFD1 U53 ( .I(n319), .Z(n317) );
  BUFFD1 U54 ( .I(n319), .Z(n318) );
  BUFFD1 U55 ( .I(n321), .Z(n312) );
  BUFFD1 U56 ( .I(n322), .Z(n321) );
  BUFFD1 U57 ( .I(n322), .Z(n320) );
  BUFFD1 U58 ( .I(n322), .Z(n319) );
  INVD1 U59 ( .I(Reset), .ZN(n322) );
  INVD1 U60 ( .I(n260), .ZN(n257) );
  INVD1 U61 ( .I(n261), .ZN(n256) );
  INVD1 U62 ( .I(n262), .ZN(n255) );
  INVD1 U63 ( .I(n259), .ZN(n258) );
  BUFFD1 U64 ( .I(n271), .Z(n282) );
  BUFFD1 U65 ( .I(n271), .Z(n283) );
  BUFFD1 U66 ( .I(n272), .Z(n284) );
  BUFFD1 U67 ( .I(n272), .Z(n285) );
  BUFFD1 U68 ( .I(n273), .Z(n286) );
  BUFFD1 U69 ( .I(n273), .Z(n287) );
  BUFFD1 U70 ( .I(n274), .Z(n288) );
  BUFFD1 U71 ( .I(n274), .Z(n289) );
  BUFFD1 U72 ( .I(n275), .Z(n290) );
  BUFFD1 U73 ( .I(n275), .Z(n291) );
  BUFFD1 U74 ( .I(n276), .Z(n292) );
  BUFFD1 U75 ( .I(n276), .Z(n293) );
  BUFFD1 U76 ( .I(n277), .Z(n294) );
  BUFFD1 U77 ( .I(n277), .Z(n295) );
  BUFFD1 U78 ( .I(n278), .Z(n296) );
  BUFFD1 U79 ( .I(n278), .Z(n297) );
  INVD1 U80 ( .I(n270), .ZN(n265) );
  INVD1 U81 ( .I(n270), .ZN(n266) );
  INVD1 U82 ( .I(n269), .ZN(n267) );
  INVD1 U83 ( .I(n269), .ZN(n268) );
  BUFFD1 U84 ( .I(n443), .Z(n259) );
  BUFFD1 U85 ( .I(n443), .Z(n260) );
  BUFFD1 U86 ( .I(n443), .Z(n261) );
  BUFFD1 U87 ( .I(n443), .Z(n262) );
  BUFFD1 U88 ( .I(n280), .Z(n273) );
  BUFFD1 U89 ( .I(n280), .Z(n274) );
  BUFFD1 U90 ( .I(n280), .Z(n275) );
  BUFFD1 U91 ( .I(n279), .Z(n276) );
  BUFFD1 U93 ( .I(n279), .Z(n277) );
  BUFFD1 U95 ( .I(n279), .Z(n278) );
  BUFFD1 U97 ( .I(n281), .Z(n271) );
  BUFFD1 U98 ( .I(n281), .Z(n272) );
  INVD1 U100 ( .I(n263), .ZN(n270) );
  INVD1 U102 ( .I(n263), .ZN(n269) );
  IND2D1 U103 ( .A1(n442), .B1(n441), .ZN(n443) );
  NR2D1 U104 ( .A1(n441), .A2(n442), .ZN(N47) );
  BUFFD1 U105 ( .I(SerClock), .Z(n280) );
  BUFFD1 U106 ( .I(SerClock), .Z(n279) );
  BUFFD1 U107 ( .I(SerClock), .Z(n281) );
  OAI21D1 U108 ( .A1(n452), .A2(n427), .B(n324), .ZN(n394) );
  NR2D1 U109 ( .A1(ParClk), .A2(n323), .ZN(n452) );
  NR2D1 U110 ( .A1(ParClk), .A2(n429), .ZN(N37) );
  NR4D0 U111 ( .A1(n428), .A2(Count32[2]), .A3(Count32[4]), .A4(Count32[3]), 
        .ZN(n430) );
  AN2D1 U112 ( .A1(N34), .A2(n453), .Z(N42) );
  AN2D1 U113 ( .A1(N33), .A2(n453), .Z(N41) );
  AN2D1 U114 ( .A1(N32), .A2(n453), .Z(N40) );
  AN2D1 U115 ( .A1(N31), .A2(n453), .Z(N39) );
  AN2D1 U116 ( .A1(N30), .A2(n453), .Z(N38) );
  ND2D1 U117 ( .A1(n323), .A2(ParValidTimer[0]), .ZN(n446) );
  INVD1 U118 ( .I(ParValidTimer[1]), .ZN(n449) );
  AO22D0 U119 ( .A1(FrameSR[8]), .A2(n257), .B1(Decoder[0]), .B2(n259), .Z(
        n357) );
  AO22D0 U120 ( .A1(FrameSR[9]), .A2(n257), .B1(Decoder[1]), .B2(n259), .Z(
        n356) );
  AO22D0 U121 ( .A1(FrameSR[10]), .A2(n257), .B1(Decoder[2]), .B2(n259), .Z(
        n355) );
  AO22D0 U122 ( .A1(FrameSR[11]), .A2(n258), .B1(Decoder[3]), .B2(n259), .Z(
        n354) );
  AO22D0 U123 ( .A1(FrameSR[12]), .A2(n258), .B1(Decoder[4]), .B2(n259), .Z(
        n353) );
  AO22D0 U124 ( .A1(FrameSR[13]), .A2(n258), .B1(Decoder[5]), .B2(n259), .Z(
        n352) );
  AO22D0 U125 ( .A1(FrameSR[14]), .A2(n258), .B1(Decoder[6]), .B2(n259), .Z(
        n351) );
  AO22D0 U126 ( .A1(FrameSR[15]), .A2(n258), .B1(Decoder[7]), .B2(n259), .Z(
        n350) );
  AO22D0 U127 ( .A1(FrameSR[24]), .A2(n255), .B1(Decoder[8]), .B2(n260), .Z(
        n349) );
  AO22D0 U128 ( .A1(FrameSR[25]), .A2(n256), .B1(Decoder[9]), .B2(n260), .Z(
        n348) );
  AO22D0 U129 ( .A1(FrameSR[26]), .A2(n256), .B1(Decoder[10]), .B2(n260), .Z(
        n347) );
  AO22D0 U130 ( .A1(FrameSR[27]), .A2(n256), .B1(Decoder[11]), .B2(n260), .Z(
        n346) );
  AO22D0 U131 ( .A1(FrameSR[28]), .A2(n257), .B1(Decoder[12]), .B2(n260), .Z(
        n345) );
  AO22D0 U132 ( .A1(FrameSR[29]), .A2(n257), .B1(Decoder[13]), .B2(n260), .Z(
        n344) );
  AO22D0 U133 ( .A1(FrameSR[30]), .A2(n257), .B1(Decoder[14]), .B2(n260), .Z(
        n343) );
  AO22D0 U134 ( .A1(FrameSR[31]), .A2(n257), .B1(Decoder[15]), .B2(n260), .Z(
        n342) );
  AO22D0 U135 ( .A1(FrameSR[40]), .A2(n257), .B1(Decoder[16]), .B2(n261), .Z(
        n341) );
  AO22D0 U136 ( .A1(FrameSR[41]), .A2(n257), .B1(Decoder[17]), .B2(n261), .Z(
        n340) );
  AO22D0 U137 ( .A1(FrameSR[42]), .A2(n255), .B1(Decoder[18]), .B2(n261), .Z(
        n339) );
  AO22D0 U138 ( .A1(FrameSR[43]), .A2(n255), .B1(Decoder[19]), .B2(n261), .Z(
        n338) );
  AO22D0 U139 ( .A1(FrameSR[44]), .A2(n255), .B1(Decoder[20]), .B2(n261), .Z(
        n337) );
  AO22D0 U140 ( .A1(FrameSR[45]), .A2(n255), .B1(Decoder[21]), .B2(n261), .Z(
        n336) );
  AO22D0 U141 ( .A1(FrameSR[46]), .A2(n256), .B1(Decoder[22]), .B2(n261), .Z(
        n335) );
  AO22D0 U142 ( .A1(FrameSR[47]), .A2(n256), .B1(Decoder[23]), .B2(n261), .Z(
        n334) );
  AO22D0 U143 ( .A1(FrameSR[56]), .A2(n256), .B1(Decoder[24]), .B2(n262), .Z(
        n333) );
  AO22D0 U144 ( .A1(FrameSR[57]), .A2(n256), .B1(Decoder[25]), .B2(n262), .Z(
        n332) );
  AO22D0 U145 ( .A1(FrameSR[58]), .A2(n256), .B1(Decoder[26]), .B2(n262), .Z(
        n331) );
  AO22D0 U146 ( .A1(FrameSR[59]), .A2(n256), .B1(Decoder[27]), .B2(n262), .Z(
        n330) );
  AO22D0 U147 ( .A1(FrameSR[60]), .A2(n255), .B1(Decoder[28]), .B2(n262), .Z(
        n329) );
  AO22D0 U148 ( .A1(FrameSR[61]), .A2(n255), .B1(Decoder[29]), .B2(n262), .Z(
        n328) );
  AO22D0 U149 ( .A1(FrameSR[62]), .A2(n255), .B1(Decoder[30]), .B2(n262), .Z(
        n327) );
  AO22D0 U150 ( .A1(FrameSR[63]), .A2(n255), .B1(Decoder[31]), .B2(n262), .Z(
        n326) );
  INVD1 U151 ( .I(ParValidTimer[0]), .ZN(n450) );
  INR2D1 U152 ( .A1(n84), .B1(n265), .ZN(n393) );
  OAI31D0 U153 ( .A1(n450), .A2(n325), .A3(n449), .B(n323), .ZN(n84) );
  NR2D1 U154 ( .A1(n445), .A2(n265), .ZN(n391) );
  XOR2D1 U155 ( .A1(ParValidTimer[1]), .A2(n446), .Z(n445) );
  NR2D1 U156 ( .A1(n444), .A2(n265), .ZN(n390) );
  XOR2D1 U157 ( .A1(n323), .A2(n450), .Z(n444) );
  INVD1 U158 ( .I(n264), .ZN(n263) );
  INVD1 U159 ( .I(n451), .ZN(n264) );
  NR2D1 U160 ( .A1(n265), .A2(n448), .ZN(n392) );
  XOR2D1 U161 ( .A1(n325), .A2(n447), .Z(n448) );
  NR2D1 U162 ( .A1(n449), .A2(n446), .ZN(n447) );
  NR4D0 U163 ( .A1(n434), .A2(FrameSR[48]), .A3(FrameSR[50]), .A4(FrameSR[49]), 
        .ZN(n435) );
  ND2D1 U164 ( .A1(n440), .A2(n439), .ZN(n442) );
  NR4D0 U165 ( .A1(FrameSR[3]), .A2(FrameSR[2]), .A3(FrameSR[1]), .A4(
        FrameSR[0]), .ZN(n440) );
  NR4D0 U166 ( .A1(FrameSR[7]), .A2(FrameSR[6]), .A3(FrameSR[5]), .A4(
        FrameSR[4]), .ZN(n439) );
  AN4D1 U167 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .Z(n441) );
  INR4D0 U168 ( .A1(FrameSR[19]), .B1(n431), .B2(FrameSR[17]), .B3(FrameSR[16]), .ZN(n438) );
  NR4D0 U169 ( .A1(n432), .A2(FrameSR[18]), .A3(FrameSR[21]), .A4(FrameSR[20]), 
        .ZN(n437) );
  NR4D0 U170 ( .A1(n433), .A2(FrameSR[33]), .A3(FrameSR[35]), .A4(FrameSR[34]), 
        .ZN(n436) );
  ND3D1 U171 ( .A1(FrameSR[51]), .A2(FrameSR[36]), .A3(FrameSR[52]), .ZN(n431)
         );
  AN2D1 U172 ( .A1(SerClk), .A2(SerValid), .Z(SerClock) );
endmodule


module SerialRx_1 ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n2;

  PLLTop_1 PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(ParClk), .Reset(n2) );
  BUFFD1 U1 ( .I(Reset), .Z(n2) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid3_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [2:0] ReadAddr;
  output [2:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n278, StateClockRaw, StateClock, N46, N47, N48, N49, N63, N64, N65,
         N66, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  wire   [2:0] OldReadAr;
  wire   [2:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n197), .CPN(StateClock), .Q(FullFIFO), .QN(n202) );
  DFND1 EmptyFIFOr_reg ( .D(n198), .CPN(StateClock), .Q(EmptyFIFO) );
  IAO21D1 U6 ( .A1(n273), .A2(n272), .B(n180), .ZN(n274) );
  MOAI22D1 U7 ( .A1(n184), .A2(n271), .B1(n271), .B2(OldReadAr[1]), .ZN(n196)
         );
  MOAI22D1 U8 ( .A1(n185), .A2(n271), .B1(n271), .B2(OldReadAr[2]), .ZN(n195)
         );
  MOAI22D1 U9 ( .A1(n270), .A2(n269), .B1(n270), .B2(OldWriteAr[1]), .ZN(n194)
         );
  MOAI22D1 U10 ( .A1(n270), .A2(n268), .B1(n270), .B2(OldWriteAr[2]), .ZN(n193) );
  MOAI22D1 U11 ( .A1(n182), .A2(n270), .B1(n270), .B2(OldWriteAr[0]), .ZN(n192) );
  MOAI22D1 U70 ( .A1(n183), .A2(n271), .B1(n271), .B2(OldReadAr[0]), .ZN(n186)
         );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n186), .CPN(StateClock), .CDN(n179), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n192), .CPN(StateClock), .CDN(n179), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n193), .CPN(StateClock), .CDN(n179), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n194), .CPN(StateClock), .CDN(n179), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n195), .CPN(StateClock), .CDN(n179), .Q(
        OldReadAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n196), .CPN(StateClock), .CDN(n179), .Q(
        OldReadAr[1]) );
  DFNCND1 ReadCmdr_reg ( .D(n187), .CPN(StateClock), .CDN(n179), .Q(ReadCmd)
         );
  DFNCND1 WriteCmdr_reg ( .D(n189), .CPN(StateClock), .CDN(n179), .Q(WriteCmd)
         );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n181), 
        .Q(CurState[2]), .QN(n245) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n181), 
        .Q(CurState[1]), .QN(n261) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n181), 
        .Q(CurState[0]), .QN(n236) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N65), .E(N66), .CP(StateClock), .CDN(n181), 
        .Q(WriteAddr[2]), .QN(n268) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N64), .E(N66), .CP(StateClock), .CDN(n181), 
        .Q(WriteAddr[1]), .QN(n269) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N49), .E(N48), .CP(StateClock), .CDN(n181), .Q(
        ReadAddr[2]), .QN(n185) );
  EDFCND1 \ReadAr_reg[1]  ( .D(N47), .E(N48), .CP(StateClock), .CDN(n181), .Q(
        ReadAddr[1]), .QN(n184) );
  EDFCND1 \ReadAr_reg[0]  ( .D(N46), .E(N48), .CP(StateClock), .CDN(n181), .Q(
        ReadAddr[0]), .QN(n183) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N63), .E(N66), .CP(StateClock), .CDN(n181), 
        .Q(n278), .QN(n182) );
  DFNCND1 \NextState_reg[1]  ( .D(n190), .CPN(StateClock), .CDN(n181), .Q(
        NextState[1]), .QN(n200) );
  DFNCND1 \NextState_reg[0]  ( .D(n188), .CPN(StateClock), .CDN(n181), .Q(
        NextState[0]), .QN(n199) );
  DFNCND1 \NextState_reg[2]  ( .D(n191), .CPN(StateClock), .CDN(n181), .Q(
        NextState[2]), .QN(n201) );
  INVD1 U3 ( .I(n180), .ZN(n179) );
  INVD1 U4 ( .I(n181), .ZN(n180) );
  INVD1 U5 ( .I(Reset), .ZN(n181) );
  INVD1 U12 ( .I(n238), .ZN(n231) );
  INVD1 U13 ( .I(n266), .ZN(n260) );
  MAOI22D0 U14 ( .A1(ReadAddr[0]), .A2(n240), .B1(n269), .B2(n218), .ZN(n215)
         );
  XNR2D1 U15 ( .A1(n268), .A2(n240), .ZN(n238) );
  INVD1 U16 ( .I(n240), .ZN(n234) );
  XNR2D1 U17 ( .A1(n231), .A2(ReadAddr[2]), .ZN(n257) );
  INVD1 U18 ( .I(n272), .ZN(n277) );
  ND2D1 U19 ( .A1(n232), .A2(n275), .ZN(n229) );
  ND3D1 U20 ( .A1(n275), .A2(n277), .A3(n204), .ZN(N66) );
  NR2D1 U21 ( .A1(n245), .A2(n236), .ZN(n273) );
  ND2D1 U22 ( .A1(n232), .A2(n277), .ZN(n267) );
  NR2D1 U23 ( .A1(ReadAddr[0]), .A2(n207), .ZN(N46) );
  NR2D1 U24 ( .A1(n217), .A2(n207), .ZN(N49) );
  NR2D1 U25 ( .A1(n203), .A2(n207), .ZN(N47) );
  XNR2D1 U26 ( .A1(ReadAddr[0]), .A2(ReadAddr[1]), .ZN(n203) );
  OAI211D1 U27 ( .A1(CurState[1]), .A2(n236), .B(n232), .C(n212), .ZN(n266) );
  AOI21D1 U28 ( .A1(WriteReq), .A2(n272), .B(n211), .ZN(n212) );
  AOI21D1 U29 ( .A1(CurState[0]), .A2(n210), .B(n245), .ZN(n211) );
  OAI33D1 U30 ( .A1(n230), .A2(n272), .A3(n229), .B1(n228), .B2(n227), .B3(
        n226), .ZN(n189) );
  INVD1 U31 ( .I(WriteCmd), .ZN(n230) );
  XNR2D1 U32 ( .A1(n268), .A2(OldWriteAr[2]), .ZN(n226) );
  XNR2D1 U33 ( .A1(n269), .A2(OldWriteAr[1]), .ZN(n227) );
  ND2D1 U34 ( .A1(WriteReq), .A2(n267), .ZN(n270) );
  OAI22D0 U35 ( .A1(n266), .A2(n200), .B1(n260), .B2(n254), .ZN(n190) );
  AOI31D0 U36 ( .A1(n253), .A2(n252), .A3(n251), .B(n272), .ZN(n254) );
  IIND4D1 U37 ( .A1(n244), .A2(n242), .B1(n237), .B2(n236), .ZN(n252) );
  AOI31D0 U38 ( .A1(n183), .A2(CurState[0]), .A3(n250), .B(n249), .ZN(n251) );
  OAI22D0 U39 ( .A1(n266), .A2(n199), .B1(n260), .B2(n224), .ZN(n188) );
  AOI21D1 U40 ( .A1(CurState[1]), .A2(n223), .B(n273), .ZN(n224) );
  OAI21D1 U41 ( .A1(CurState[2]), .A2(n222), .B(n221), .ZN(n223) );
  AOI22D0 U42 ( .A1(n258), .A2(ReadAddr[2]), .B1(n185), .B2(n259), .ZN(n222)
         );
  OAI31D0 U43 ( .A1(n277), .A2(WriteReq), .A3(n180), .B(n276), .ZN(n198) );
  OAI31D0 U44 ( .A1(CurState[0]), .A2(n180), .A3(CurState[2]), .B(EmptyFIFO), 
        .ZN(n276) );
  OAI21D1 U45 ( .A1(n266), .A2(n201), .B(n265), .ZN(n191) );
  OAI211D1 U46 ( .A1(CurState[2]), .A2(n264), .B(CurState[0]), .C(n263), .ZN(
        n265) );
  NR4D0 U47 ( .A1(n257), .A2(n256), .A3(n261), .A4(n255), .ZN(n264) );
  AOI21D1 U48 ( .A1(n262), .A2(n261), .B(n260), .ZN(n263) );
  ND3D1 U49 ( .A1(n225), .A2(n267), .A3(WriteReq), .ZN(n228) );
  XNR2D1 U50 ( .A1(n278), .A2(OldWriteAr[0]), .ZN(n225) );
  MAOI22D0 U51 ( .A1(n278), .A2(n213), .B1(n184), .B2(n218), .ZN(n214) );
  OAI33D1 U52 ( .A1(ReadAddr[1]), .A2(WriteAddr[2]), .A3(n215), .B1(n268), 
        .B2(WriteAddr[1]), .B3(n214), .ZN(n259) );
  OAI33D1 U53 ( .A1(ReadAddr[1]), .A2(n215), .A3(n268), .B1(n214), .B2(
        WriteAddr[2]), .B3(WriteAddr[1]), .ZN(n258) );
  NR2D1 U54 ( .A1(n269), .A2(n182), .ZN(n240) );
  OAI21D1 U55 ( .A1(WriteAddr[1]), .A2(n278), .B(n234), .ZN(n216) );
  XOR2D1 U56 ( .A1(n216), .A2(n184), .Z(n256) );
  AOI31D0 U57 ( .A1(n182), .A2(CurState[0]), .A3(n233), .B(n232), .ZN(n253) );
  NR3D0 U58 ( .A1(n256), .A2(n183), .A3(n257), .ZN(n233) );
  OAI31D0 U59 ( .A1(n220), .A2(n219), .A3(n255), .B(CurState[0]), .ZN(n221) );
  XNR2D1 U60 ( .A1(WriteAddr[2]), .A2(n217), .ZN(n219) );
  INVD1 U61 ( .I(n256), .ZN(n220) );
  NR3D0 U62 ( .A1(n256), .A2(n182), .A3(n241), .ZN(n250) );
  AOI21D1 U63 ( .A1(n244), .A2(n240), .B(n239), .ZN(n241) );
  OAI32D1 U64 ( .A1(n268), .A2(n185), .A3(n240), .B1(ReadAddr[2]), .B2(n238), 
        .ZN(n239) );
  AO22D0 U65 ( .A1(ReadAddr[2]), .A2(n259), .B1(n258), .B2(n185), .Z(n262) );
  OAI222D0 U66 ( .A1(n268), .A2(ReadAddr[2]), .B1(n269), .B2(ReadAddr[1]), 
        .C1(n182), .C2(ReadAddr[0]), .ZN(n242) );
  AOI22D0 U67 ( .A1(n245), .A2(CurState[1]), .B1(n261), .B2(n273), .ZN(n232)
         );
  NR3D0 U68 ( .A1(CurState[1]), .A2(CurState[2]), .A3(CurState[0]), .ZN(n272)
         );
  ND2D1 U69 ( .A1(CurState[1]), .A2(n273), .ZN(n275) );
  ND2D1 U71 ( .A1(ReadCmd), .A2(n277), .ZN(n207) );
  OAI21D1 U72 ( .A1(n182), .A2(n183), .B(n218), .ZN(n255) );
  OAI32D0 U73 ( .A1(n275), .A2(n180), .A3(ReadReq), .B1(n274), .B2(n202), .ZN(
        n197) );
  ND2D1 U74 ( .A1(WriteCmd), .A2(n275), .ZN(n204) );
  OAI211D1 U75 ( .A1(n182), .A2(ReadAddr[1]), .B(n235), .C(n234), .ZN(n237) );
  OAI21D1 U76 ( .A1(WriteAddr[1]), .A2(n184), .B(n183), .ZN(n235) );
  CKND2D0 U77 ( .A1(ReadReq), .A2(n229), .ZN(n271) );
  NR2D1 U78 ( .A1(WriteAddr[2]), .A2(n185), .ZN(n244) );
  ND2D1 U79 ( .A1(n182), .A2(n183), .ZN(n218) );
  OAI22D0 U80 ( .A1(n183), .A2(n275), .B1(n278), .B2(n204), .ZN(N63) );
  OAI22D0 U81 ( .A1(n185), .A2(n275), .B1(n231), .B2(n204), .ZN(N65) );
  OAI22D0 U82 ( .A1(n184), .A2(n275), .B1(n216), .B2(n204), .ZN(N64) );
  AOI31D0 U83 ( .A1(n248), .A2(n247), .A3(n246), .B(n245), .ZN(n249) );
  AOI22D0 U84 ( .A1(n244), .A2(ReadAddr[1]), .B1(n182), .B2(ReadAddr[0]), .ZN(
        n246) );
  OAI21D1 U85 ( .A1(n244), .A2(n242), .B(n269), .ZN(n248) );
  OAI21D1 U86 ( .A1(ReadAddr[1]), .A2(n243), .B(n242), .ZN(n247) );
  OAI32D1 U87 ( .A1(n209), .A2(n208), .A3(n210), .B1(n229), .B2(n207), .ZN(
        n187) );
  XNR2D1 U88 ( .A1(n184), .A2(OldReadAr[1]), .ZN(n208) );
  ND3D1 U89 ( .A1(n206), .A2(n229), .A3(n205), .ZN(n209) );
  XNR2D1 U90 ( .A1(ReadAddr[2]), .A2(OldReadAr[2]), .ZN(n206) );
  IND2D1 U91 ( .A1(ReadCmd), .B1(n277), .ZN(N48) );
  NR2D1 U92 ( .A1(n183), .A2(n184), .ZN(n213) );
  XOR2D1 U93 ( .A1(n213), .A2(n185), .Z(n217) );
  XNR2D1 U94 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n243) );
  XNR2D1 U95 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n205) );
  BUFFD1 U96 ( .I(n278), .Z(WriteAddr[0]) );
  ND2D1 U97 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  INVD0 U98 ( .I(ReadReq), .ZN(n210) );
endmodule


module DPMem1kx32_AWid3_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [2:0] AddrR;
  input [2:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N48, N49, N50, ClockR, ClockW, Dreadyr, \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N87, N99, N161, N194, N227, N260, N293, N326, N359, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361;
  wire   [31:0] DataOr;
  assign N48 = AddrR[0];
  assign N49 = AddrR[1];
  assign N50 = AddrR[2];

  XNR4D1 U13 ( .A1(DataI[25]), .A2(DataI[24]), .A3(DataI[27]), .A4(DataI[26]), 
        .ZN(n349) );
  XOR4D1 U14 ( .A1(DataI[29]), .A2(DataI[28]), .A3(DataI[31]), .A4(DataI[30]), 
        .Z(n350) );
  XOR4D1 U15 ( .A1(DataI[21]), .A2(DataI[20]), .A3(DataI[23]), .A4(DataI[22]), 
        .Z(n353) );
  XOR4D1 U16 ( .A1(DataI[14]), .A2(DataI[13]), .A3(DataI[16]), .A4(DataI[15]), 
        .Z(n356) );
  XNR4D1 U17 ( .A1(DataI[7]), .A2(DataI[6]), .A3(DataI[9]), .A4(DataI[8]), 
        .ZN(n359) );
  XOR4D1 U21 ( .A1(n344), .A2(N74), .A3(n343), .A4(N77), .Z(n345) );
  XNR4D1 U22 ( .A1(N71), .A2(N70), .A3(N73), .A4(N72), .ZN(n343) );
  XNR4D1 U27 ( .A1(N53), .A2(N52), .A3(N55), .A4(N54), .ZN(n337) );
  XOR4D1 U28 ( .A1(N57), .A2(N56), .A3(N59), .A4(N58), .Z(n338) );
  XNR4D1 U29 ( .A1(N64), .A2(N63), .A3(N66), .A4(N65), .ZN(n341) );
  XNR4D1 U30 ( .A1(N82), .A2(N80), .A3(N84), .A4(N83), .ZN(n347) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(DataI[23]), .E(n193), .CP(n242), .CDN(
        n290), .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(DataI[22]), .E(n194), .CP(n242), .CDN(
        n290), .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(DataI[17]), .E(n194), .CP(n243), .CDN(
        n289), .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(DataI[16]), .E(n194), .CP(n243), .CDN(
        n289), .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(DataI[15]), .E(n194), .CP(n243), .CDN(
        n289), .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(DataI[14]), .E(n194), .CP(n243), .CDN(
        n289), .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(DataI[13]), .E(n194), .CP(n243), .CDN(
        n289), .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(DataI[12]), .E(n195), .CP(n243), .CDN(
        n289), .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(DataI[11]), .E(n195), .CP(n243), .CDN(
        n289), .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(DataI[10]), .E(n195), .CP(n243), .CDN(
        n289), .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(DataI[9]), .E(n195), .CP(n243), .CDN(n288), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(DataI[8]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(DataI[7]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(DataI[6]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(DataI[5]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(DataI[4]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(DataI[3]), .E(n195), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(DataI[2]), .E(n196), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(DataI[1]), .E(n196), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(DataI[0]), .E(n196), .CP(n244), .CDN(n288), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(DataI[23]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(DataI[22]), .E(n210), .CP(n249), .CDN(
        n284), .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(DataI[17]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(DataI[16]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(DataI[15]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(DataI[14]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(DataI[13]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(DataI[12]), .E(n211), .CP(n250), .CDN(
        n283), .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(DataI[11]), .E(n211), .CP(n251), .CDN(
        n283), .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(DataI[10]), .E(n211), .CP(n251), .CDN(
        n283), .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(DataI[9]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(DataI[8]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(DataI[7]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(DataI[6]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(DataI[5]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(DataI[4]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(DataI[3]), .E(n211), .CP(n251), .CDN(n282), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(DataI[2]), .E(n212), .CP(n252), .CDN(n282), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(DataI[1]), .E(n212), .CP(n252), .CDN(n282), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(DataI[0]), .E(n212), .CP(n252), .CDN(n282), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(DataI[23]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(DataI[22]), .E(n162), .CP(n227), .CDN(
        n302), .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(DataI[17]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(DataI[16]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(DataI[15]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(DataI[14]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(DataI[13]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(DataI[12]), .E(n163), .CP(n228), .CDN(
        n301), .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(DataI[11]), .E(n163), .CP(n229), .CDN(
        n301), .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(DataI[10]), .E(n163), .CP(n229), .CDN(
        n301), .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(DataI[9]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(DataI[8]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(DataI[7]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(DataI[6]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(DataI[5]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(DataI[4]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(DataI[3]), .E(n163), .CP(n229), .CDN(n300), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(DataI[2]), .E(n164), .CP(n230), .CDN(n300), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(DataI[1]), .E(n164), .CP(n230), .CDN(n300), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(DataI[0]), .E(n164), .CP(n230), .CDN(n300), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(DataI[23]), .E(n169), .CP(n231), .CDN(
        n299), .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(DataI[22]), .E(n170), .CP(n231), .CDN(
        n299), .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(DataI[17]), .E(n170), .CP(n232), .CDN(
        n298), .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(DataI[16]), .E(n170), .CP(n232), .CDN(
        n298), .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(DataI[15]), .E(n170), .CP(n232), .CDN(
        n298), .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(DataI[14]), .E(n170), .CP(n232), .CDN(
        n298), .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(DataI[13]), .E(n170), .CP(n232), .CDN(
        n298), .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(DataI[12]), .E(n171), .CP(n232), .CDN(
        n298), .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(DataI[11]), .E(n171), .CP(n232), .CDN(
        n298), .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(DataI[10]), .E(n171), .CP(n232), .CDN(
        n298), .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(DataI[9]), .E(n171), .CP(n232), .CDN(n297), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(DataI[8]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(DataI[7]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(DataI[6]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(DataI[5]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(DataI[4]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(DataI[3]), .E(n171), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(DataI[2]), .E(n172), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(DataI[1]), .E(n172), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(DataI[0]), .E(n172), .CP(n233), .CDN(n297), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(DataI[23]), .E(n177), .CP(n235), .CDN(
        n296), .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(DataI[22]), .E(n178), .CP(n235), .CDN(
        n296), .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(DataI[17]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(DataI[16]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(DataI[15]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(DataI[14]), .E(n178), .CP(n236), .CDN(
        n295), .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(DataI[13]), .E(n178), .CP(n236), .CDN(
        n295), .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(DataI[12]), .E(n179), .CP(n236), .CDN(
        n295), .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(DataI[11]), .E(n179), .CP(n236), .CDN(
        n295), .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(DataI[10]), .E(n179), .CP(n236), .CDN(
        n295), .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(DataI[9]), .E(n179), .CP(n236), .CDN(n294), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(DataI[8]), .E(n179), .CP(n236), .CDN(n294), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(DataI[7]), .E(n179), .CP(n236), .CDN(n294), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(DataI[6]), .E(n179), .CP(n236), .CDN(n294), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(DataI[5]), .E(n179), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(DataI[4]), .E(n179), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(DataI[3]), .E(n179), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(DataI[2]), .E(n180), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(DataI[1]), .E(n180), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(DataI[0]), .E(n180), .CP(n237), .CDN(n294), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(DataI[23]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(DataI[22]), .E(n186), .CP(n238), .CDN(
        n293), .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(DataI[17]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(DataI[16]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(DataI[15]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(DataI[14]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(DataI[13]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(DataI[12]), .E(n187), .CP(n239), .CDN(
        n292), .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(DataI[11]), .E(n187), .CP(n240), .CDN(
        n292), .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(DataI[10]), .E(n187), .CP(n240), .CDN(
        n292), .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(DataI[9]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(DataI[8]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(DataI[7]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(DataI[6]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(DataI[5]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(DataI[4]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(DataI[3]), .E(n187), .CP(n240), .CDN(n291), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(DataI[2]), .E(n188), .CP(n241), .CDN(n291), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(DataI[1]), .E(n188), .CP(n241), .CDN(n291), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(DataI[0]), .E(n188), .CP(n241), .CDN(n291), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(DataI[23]), .E(n201), .CP(n246), .CDN(
        n287), .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(DataI[22]), .E(n202), .CP(n246), .CDN(
        n287), .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(DataI[17]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(DataI[16]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(DataI[15]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(DataI[14]), .E(n202), .CP(n247), .CDN(
        n286), .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(DataI[13]), .E(n202), .CP(n247), .CDN(
        n286), .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(DataI[12]), .E(n203), .CP(n247), .CDN(
        n286), .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(DataI[11]), .E(n203), .CP(n247), .CDN(
        n286), .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(DataI[10]), .E(n203), .CP(n247), .CDN(
        n286), .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(DataI[9]), .E(n203), .CP(n247), .CDN(n285), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(DataI[8]), .E(n203), .CP(n247), .CDN(n285), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(DataI[7]), .E(n203), .CP(n247), .CDN(n285), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(DataI[6]), .E(n203), .CP(n247), .CDN(n285), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(DataI[5]), .E(n203), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(DataI[4]), .E(n203), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(DataI[3]), .E(n203), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(DataI[2]), .E(n204), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(DataI[1]), .E(n204), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(DataI[0]), .E(n204), .CP(n248), .CDN(n285), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(DataI[23]), .E(n153), .CP(n224), .CDN(
        n305), .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(DataI[22]), .E(n154), .CP(n224), .CDN(
        n305), .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(DataI[17]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(DataI[16]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(DataI[15]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(DataI[14]), .E(n154), .CP(n225), .CDN(
        n304), .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(DataI[13]), .E(n154), .CP(n225), .CDN(
        n304), .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(DataI[12]), .E(n155), .CP(n225), .CDN(
        n304), .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(DataI[11]), .E(n155), .CP(n225), .CDN(
        n304), .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(DataI[10]), .E(n155), .CP(n225), .CDN(
        n304), .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(DataI[9]), .E(n155), .CP(n225), .CDN(n303), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(DataI[8]), .E(n155), .CP(n225), .CDN(n303), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(DataI[7]), .E(n155), .CP(n225), .CDN(n303), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(DataI[6]), .E(n155), .CP(n225), .CDN(n303), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(DataI[5]), .E(n155), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(DataI[4]), .E(n155), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(DataI[3]), .E(n155), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(DataI[2]), .E(n156), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(DataI[1]), .E(n156), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(DataI[0]), .E(n156), .CP(n226), .CDN(n303), 
        .Q(\Storage[7][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n1), .CP(n273), .CDN(n282), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N87), .E(n193), .CP(n241), .CDN(n291), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(DataI[31]), .E(n193), .CP(n241), .CDN(
        n290), .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(DataI[30]), .E(n193), .CP(n241), .CDN(
        n290), .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(DataI[29]), .E(n193), .CP(n241), .CDN(
        n290), .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(DataI[28]), .E(n193), .CP(n241), .CDN(
        n290), .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(DataI[27]), .E(n193), .CP(n241), .CDN(
        n290), .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(DataI[26]), .E(n193), .CP(n242), .CDN(
        n290), .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(DataI[25]), .E(n193), .CP(n242), .CDN(
        n290), .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(DataI[24]), .E(n193), .CP(n242), .CDN(
        n290), .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(DataI[21]), .E(n194), .CP(n242), .CDN(
        n290), .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(DataI[20]), .E(n194), .CP(n242), .CDN(
        n289), .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(DataI[19]), .E(n194), .CP(n242), .CDN(
        n289), .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(DataI[18]), .E(n194), .CP(n242), .CDN(
        n289), .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N87), .E(n209), .CP(n248), .CDN(n285), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(DataI[31]), .E(n209), .CP(n248), .CDN(
        n284), .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(DataI[30]), .E(n209), .CP(n248), .CDN(
        n284), .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(DataI[29]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(DataI[28]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(DataI[27]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(DataI[26]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(DataI[25]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(DataI[24]), .E(n209), .CP(n249), .CDN(
        n284), .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(DataI[21]), .E(n210), .CP(n249), .CDN(
        n284), .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(DataI[20]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(DataI[19]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(DataI[18]), .E(n210), .CP(n250), .CDN(
        n283), .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N87), .E(n161), .CP(n226), .CDN(n303), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(DataI[31]), .E(n161), .CP(n226), .CDN(
        n302), .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(DataI[30]), .E(n161), .CP(n226), .CDN(
        n302), .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(DataI[29]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(DataI[28]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(DataI[27]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(DataI[26]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(DataI[25]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(DataI[24]), .E(n161), .CP(n227), .CDN(
        n302), .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(DataI[21]), .E(n162), .CP(n227), .CDN(
        n302), .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(DataI[20]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(DataI[19]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(DataI[18]), .E(n162), .CP(n228), .CDN(
        n301), .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N87), .E(n169), .CP(n230), .CDN(n300), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(DataI[31]), .E(n169), .CP(n230), .CDN(
        n299), .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(DataI[30]), .E(n169), .CP(n230), .CDN(
        n299), .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(DataI[29]), .E(n169), .CP(n230), .CDN(
        n299), .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(DataI[28]), .E(n169), .CP(n230), .CDN(
        n299), .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(DataI[27]), .E(n169), .CP(n230), .CDN(
        n299), .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(DataI[26]), .E(n169), .CP(n231), .CDN(
        n299), .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(DataI[25]), .E(n169), .CP(n231), .CDN(
        n299), .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(DataI[24]), .E(n169), .CP(n231), .CDN(
        n299), .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(DataI[21]), .E(n170), .CP(n231), .CDN(
        n299), .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(DataI[20]), .E(n170), .CP(n231), .CDN(
        n298), .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(DataI[19]), .E(n170), .CP(n231), .CDN(
        n298), .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(DataI[18]), .E(n170), .CP(n231), .CDN(
        n298), .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N87), .E(n177), .CP(n234), .CDN(n297), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(DataI[31]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(DataI[30]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(DataI[29]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(DataI[28]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(DataI[27]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(DataI[26]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(DataI[25]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(DataI[24]), .E(n177), .CP(n234), .CDN(
        n296), .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(DataI[21]), .E(n178), .CP(n235), .CDN(
        n296), .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(DataI[20]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(DataI[19]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(DataI[18]), .E(n178), .CP(n235), .CDN(
        n295), .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N87), .E(n185), .CP(n237), .CDN(n294), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(DataI[31]), .E(n185), .CP(n237), .CDN(
        n293), .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(DataI[30]), .E(n185), .CP(n237), .CDN(
        n293), .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(DataI[29]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(DataI[28]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(DataI[27]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(DataI[26]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(DataI[25]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(DataI[24]), .E(n185), .CP(n238), .CDN(
        n293), .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(DataI[21]), .E(n186), .CP(n238), .CDN(
        n293), .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(DataI[20]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(DataI[19]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(DataI[18]), .E(n186), .CP(n239), .CDN(
        n292), .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N87), .E(n201), .CP(n245), .CDN(n288), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(DataI[31]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(DataI[30]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(DataI[29]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(DataI[28]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(DataI[27]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(DataI[26]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(DataI[25]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(DataI[24]), .E(n201), .CP(n245), .CDN(
        n287), .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(DataI[21]), .E(n202), .CP(n246), .CDN(
        n287), .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(DataI[20]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(DataI[19]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(DataI[18]), .E(n202), .CP(n246), .CDN(
        n286), .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N87), .E(n153), .CP(n223), .CDN(n306), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(DataI[31]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(DataI[30]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(DataI[29]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(DataI[28]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(DataI[27]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(DataI[26]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(DataI[25]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(DataI[24]), .E(n153), .CP(n223), .CDN(
        n305), .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(DataI[21]), .E(n154), .CP(n224), .CDN(
        n305), .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(DataI[20]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(DataI[19]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(DataI[18]), .E(n154), .CP(n224), .CDN(
        n304), .Q(\Storage[7][18] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N53), .E(n277), .CP(n270), .CDN(n309), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N54), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N55), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N56), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N57), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N58), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N59), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N60), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N61), .E(n277), .CP(n270), .CDN(n308), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N62), .E(n277), .CP(n271), .CDN(n308), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N63), .E(n277), .CP(n271), .CDN(n308), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N64), .E(n277), .CP(n271), .CDN(n308), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N65), .E(n277), .CP(n271), .CDN(n307), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N66), .E(n277), .CP(n271), .CDN(n307), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N67), .E(n277), .CP(n271), .CDN(n307), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N68), .E(n277), .CP(n271), .CDN(n307), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N69), .E(n277), .CP(n271), .CDN(n307), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N70), .E(n276), .CP(n271), .CDN(n307), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N71), .E(n276), .CP(n272), .CDN(n307), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N72), .E(n276), .CP(n272), .CDN(n307), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N73), .E(n276), .CP(n272), .CDN(n307), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N74), .E(n276), .CP(n272), .CDN(n307), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N75), .E(n276), .CP(n272), .CDN(n307), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N76), .E(n276), .CP(n272), .CDN(n306), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N77), .E(n276), .CP(n272), .CDN(n306), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N78), .E(n276), .CP(n272), .CDN(n306), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N79), .E(n276), .CP(n272), .CDN(n306), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N80), .E(n276), .CP(n273), .CDN(n306), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N81), .E(n276), .CP(n273), .CDN(n306), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N82), .E(n276), .CP(n273), .CDN(n306), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N83), .E(n276), .CP(n273), .CDN(n306), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N84), .E(n276), .CP(n273), .CDN(n306), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N85), .E(n276), .CP(n273), .CDN(n306), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKAN2D0 U3 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  INVD1 U4 ( .I(n281), .ZN(n129) );
  BUFFD1 U5 ( .I(n320), .Z(n288) );
  BUFFD1 U6 ( .I(n320), .Z(n289) );
  BUFFD1 U7 ( .I(n319), .Z(n290) );
  BUFFD1 U8 ( .I(n319), .Z(n291) );
  BUFFD1 U9 ( .I(n318), .Z(n292) );
  BUFFD1 U10 ( .I(n318), .Z(n293) );
  BUFFD1 U11 ( .I(n317), .Z(n294) );
  BUFFD1 U12 ( .I(n317), .Z(n295) );
  BUFFD1 U18 ( .I(n316), .Z(n296) );
  BUFFD1 U19 ( .I(n316), .Z(n297) );
  BUFFD1 U20 ( .I(n315), .Z(n298) );
  BUFFD1 U23 ( .I(n315), .Z(n299) );
  BUFFD1 U24 ( .I(n314), .Z(n300) );
  BUFFD1 U25 ( .I(n314), .Z(n301) );
  BUFFD1 U26 ( .I(n313), .Z(n302) );
  BUFFD1 U31 ( .I(n313), .Z(n303) );
  BUFFD1 U32 ( .I(n312), .Z(n304) );
  BUFFD1 U33 ( .I(n312), .Z(n305) );
  BUFFD1 U34 ( .I(n311), .Z(n306) );
  BUFFD1 U35 ( .I(n311), .Z(n307) );
  BUFFD1 U36 ( .I(n310), .Z(n308) );
  BUFFD1 U37 ( .I(n310), .Z(n309) );
  BUFFD1 U38 ( .I(n323), .Z(n282) );
  BUFFD1 U39 ( .I(n323), .Z(n283) );
  BUFFD1 U40 ( .I(n322), .Z(n284) );
  BUFFD1 U41 ( .I(n322), .Z(n285) );
  BUFFD1 U42 ( .I(n321), .Z(n286) );
  BUFFD1 U43 ( .I(n321), .Z(n287) );
  BUFFD1 U44 ( .I(n325), .Z(n320) );
  BUFFD1 U45 ( .I(n325), .Z(n319) );
  BUFFD1 U46 ( .I(n325), .Z(n318) );
  BUFFD1 U47 ( .I(n326), .Z(n317) );
  BUFFD1 U48 ( .I(n326), .Z(n316) );
  BUFFD1 U49 ( .I(n326), .Z(n315) );
  BUFFD1 U50 ( .I(n327), .Z(n314) );
  BUFFD1 U51 ( .I(n327), .Z(n313) );
  BUFFD1 U52 ( .I(n327), .Z(n312) );
  BUFFD1 U53 ( .I(n328), .Z(n311) );
  BUFFD1 U54 ( .I(n328), .Z(n310) );
  BUFFD1 U55 ( .I(n324), .Z(n322) );
  BUFFD1 U56 ( .I(n324), .Z(n321) );
  BUFFD1 U57 ( .I(n324), .Z(n323) );
  BUFFD1 U58 ( .I(n330), .Z(n325) );
  BUFFD1 U59 ( .I(n330), .Z(n326) );
  BUFFD1 U60 ( .I(n329), .Z(n327) );
  BUFFD1 U61 ( .I(n329), .Z(n328) );
  BUFFD1 U62 ( .I(n331), .Z(n324) );
  INVD1 U63 ( .I(n332), .ZN(n331) );
  INVD1 U64 ( .I(n332), .ZN(n330) );
  INVD1 U65 ( .I(n332), .ZN(n329) );
  INVD1 U66 ( .I(n333), .ZN(n332) );
  INVD1 U67 ( .I(Reset), .ZN(n333) );
  BUFFD1 U68 ( .I(n256), .Z(n246) );
  BUFFD1 U69 ( .I(n256), .Z(n245) );
  BUFFD1 U70 ( .I(n257), .Z(n244) );
  BUFFD1 U71 ( .I(n257), .Z(n243) );
  BUFFD1 U72 ( .I(n258), .Z(n242) );
  BUFFD1 U73 ( .I(n258), .Z(n241) );
  BUFFD1 U74 ( .I(n259), .Z(n240) );
  BUFFD1 U75 ( .I(n259), .Z(n239) );
  BUFFD1 U76 ( .I(n260), .Z(n238) );
  BUFFD1 U77 ( .I(n260), .Z(n237) );
  BUFFD1 U78 ( .I(n261), .Z(n236) );
  BUFFD1 U79 ( .I(n261), .Z(n235) );
  BUFFD1 U80 ( .I(n262), .Z(n234) );
  BUFFD1 U81 ( .I(n262), .Z(n233) );
  BUFFD1 U82 ( .I(n263), .Z(n232) );
  BUFFD1 U83 ( .I(n263), .Z(n231) );
  BUFFD1 U84 ( .I(n264), .Z(n230) );
  BUFFD1 U85 ( .I(n264), .Z(n229) );
  BUFFD1 U86 ( .I(n265), .Z(n228) );
  BUFFD1 U87 ( .I(n265), .Z(n227) );
  BUFFD1 U88 ( .I(n266), .Z(n226) );
  BUFFD1 U89 ( .I(n266), .Z(n225) );
  BUFFD1 U90 ( .I(n267), .Z(n224) );
  BUFFD1 U91 ( .I(n267), .Z(n223) );
  INVD1 U92 ( .I(n197), .ZN(n195) );
  INVD1 U93 ( .I(n198), .ZN(n194) );
  INVD1 U94 ( .I(n198), .ZN(n193) );
  INVD1 U95 ( .I(n189), .ZN(n187) );
  INVD1 U96 ( .I(n190), .ZN(n186) );
  INVD1 U97 ( .I(n190), .ZN(n185) );
  INVD1 U98 ( .I(n165), .ZN(n163) );
  INVD1 U99 ( .I(n166), .ZN(n162) );
  INVD1 U100 ( .I(n166), .ZN(n161) );
  INVD1 U101 ( .I(n157), .ZN(n155) );
  INVD1 U102 ( .I(n158), .ZN(n154) );
  INVD1 U103 ( .I(n158), .ZN(n153) );
  INVD1 U104 ( .I(n197), .ZN(n196) );
  INVD1 U105 ( .I(n189), .ZN(n188) );
  INVD1 U106 ( .I(n165), .ZN(n164) );
  INVD1 U107 ( .I(n157), .ZN(n156) );
  BUFFD1 U108 ( .I(n253), .Z(n251) );
  BUFFD1 U109 ( .I(n254), .Z(n250) );
  BUFFD1 U110 ( .I(n254), .Z(n249) );
  BUFFD1 U111 ( .I(n255), .Z(n248) );
  BUFFD1 U112 ( .I(n255), .Z(n247) );
  BUFFD1 U113 ( .I(n216), .Z(n256) );
  BUFFD1 U114 ( .I(n216), .Z(n257) );
  BUFFD1 U115 ( .I(n216), .Z(n258) );
  BUFFD1 U116 ( .I(n217), .Z(n259) );
  BUFFD1 U117 ( .I(n217), .Z(n260) );
  BUFFD1 U118 ( .I(n217), .Z(n261) );
  BUFFD1 U119 ( .I(n218), .Z(n262) );
  BUFFD1 U120 ( .I(n218), .Z(n263) );
  BUFFD1 U121 ( .I(n218), .Z(n264) );
  BUFFD1 U122 ( .I(n219), .Z(n265) );
  BUFFD1 U123 ( .I(n219), .Z(n266) );
  BUFFD1 U124 ( .I(n219), .Z(n267) );
  BUFFD1 U125 ( .I(n253), .Z(n252) );
  BUFFD1 U126 ( .I(n143), .Z(n145) );
  BUFFD1 U127 ( .I(n142), .Z(n149) );
  BUFFD1 U128 ( .I(n142), .Z(n147) );
  BUFFD1 U129 ( .I(n143), .Z(n146) );
  BUFFD1 U130 ( .I(n142), .Z(n148) );
  BUFFD1 U131 ( .I(n140), .Z(n138) );
  BUFFD1 U132 ( .I(n140), .Z(n137) );
  BUFFD1 U133 ( .I(n140), .Z(n136) );
  BUFFD1 U134 ( .I(n139), .Z(n135) );
  BUFFD1 U135 ( .I(n139), .Z(n134) );
  BUFFD1 U136 ( .I(n143), .Z(n144) );
  BUFFD1 U137 ( .I(n139), .Z(n133) );
  INVD1 U138 ( .I(n183), .ZN(n189) );
  INVD1 U139 ( .I(n183), .ZN(n190) );
  INVD1 U140 ( .I(n159), .ZN(n165) );
  INVD1 U141 ( .I(n159), .ZN(n166) );
  INVD1 U142 ( .I(n151), .ZN(n157) );
  INVD1 U143 ( .I(n151), .ZN(n158) );
  INVD1 U144 ( .I(n191), .ZN(n197) );
  INVD1 U145 ( .I(n191), .ZN(n198) );
  INVD1 U146 ( .I(n213), .ZN(n211) );
  INVD1 U147 ( .I(n214), .ZN(n210) );
  INVD1 U148 ( .I(n214), .ZN(n209) );
  INVD1 U149 ( .I(n205), .ZN(n203) );
  INVD1 U150 ( .I(n206), .ZN(n202) );
  INVD1 U151 ( .I(n206), .ZN(n201) );
  INVD1 U152 ( .I(n181), .ZN(n179) );
  INVD1 U153 ( .I(n182), .ZN(n178) );
  INVD1 U154 ( .I(n182), .ZN(n177) );
  INVD1 U155 ( .I(n173), .ZN(n171) );
  INVD1 U156 ( .I(n174), .ZN(n170) );
  INVD1 U157 ( .I(n174), .ZN(n169) );
  INVD1 U158 ( .I(n213), .ZN(n212) );
  INVD1 U159 ( .I(n205), .ZN(n204) );
  INVD1 U160 ( .I(n181), .ZN(n180) );
  INVD1 U161 ( .I(n173), .ZN(n172) );
  BUFFD1 U162 ( .I(n215), .Z(n253) );
  BUFFD1 U163 ( .I(n215), .Z(n254) );
  BUFFD1 U164 ( .I(n215), .Z(n255) );
  BUFFD1 U165 ( .I(n221), .Z(n216) );
  BUFFD1 U166 ( .I(n221), .Z(n217) );
  BUFFD1 U167 ( .I(n220), .Z(n218) );
  BUFFD1 U168 ( .I(n220), .Z(n219) );
  INVD1 U169 ( .I(n274), .ZN(n272) );
  INVD1 U170 ( .I(n275), .ZN(n271) );
  INVD1 U171 ( .I(n275), .ZN(n270) );
  INVD1 U172 ( .I(n274), .ZN(n273) );
  XOR3D1 U173 ( .A1(N69), .A2(N68), .A3(n342), .Z(n344) );
  XOR3D1 U174 ( .A1(N67), .A2(n341), .A3(n340), .Z(n342) );
  XOR3D1 U175 ( .A1(N62), .A2(N61), .A3(n339), .Z(n340) );
  XOR3D1 U176 ( .A1(n338), .A2(N60), .A3(n337), .Z(n339) );
  XOR3D1 U177 ( .A1(N81), .A2(N76), .A3(n348), .Z(N85) );
  XOR3D1 U178 ( .A1(N75), .A2(n347), .A3(n346), .Z(n348) );
  XOR3D1 U179 ( .A1(N79), .A2(N78), .A3(n345), .Z(n346) );
  BUFFD1 U180 ( .I(n279), .Z(n142) );
  BUFFD1 U181 ( .I(n279), .Z(n143) );
  BUFFD1 U182 ( .I(n141), .Z(n150) );
  BUFFD1 U183 ( .I(n279), .Z(n141) );
  BUFFD1 U184 ( .I(n280), .Z(n140) );
  BUFFD1 U185 ( .I(n280), .Z(n139) );
  INVD1 U186 ( .I(n129), .ZN(n131) );
  INVD1 U187 ( .I(n129), .ZN(n132) );
  INVD1 U188 ( .I(n129), .ZN(n130) );
  INVD1 U189 ( .I(AddrW[0]), .ZN(n334) );
  INVD1 U190 ( .I(n207), .ZN(n213) );
  INVD1 U191 ( .I(n207), .ZN(n214) );
  INVD1 U192 ( .I(n199), .ZN(n205) );
  INVD1 U193 ( .I(n199), .ZN(n206) );
  INVD1 U194 ( .I(n175), .ZN(n181) );
  INVD1 U195 ( .I(n175), .ZN(n182) );
  INVD1 U196 ( .I(n167), .ZN(n173) );
  INVD1 U197 ( .I(n167), .ZN(n174) );
  INVD1 U198 ( .I(n192), .ZN(n191) );
  INVD1 U199 ( .I(N194), .ZN(n192) );
  NR3D0 U200 ( .A1(n336), .A2(AddrW[0]), .A3(n361), .ZN(N194) );
  INVD1 U201 ( .I(n184), .ZN(n183) );
  INVD1 U202 ( .I(N227), .ZN(n184) );
  NR3D0 U203 ( .A1(n336), .A2(n361), .A3(n334), .ZN(N227) );
  INVD1 U204 ( .I(n160), .ZN(n159) );
  INVD1 U205 ( .I(N326), .ZN(n160) );
  NR3D0 U206 ( .A1(n336), .A2(AddrW[0]), .A3(n335), .ZN(N326) );
  INVD1 U207 ( .I(n152), .ZN(n151) );
  INVD1 U208 ( .I(N359), .ZN(n152) );
  NR3D0 U209 ( .A1(n336), .A2(n335), .A3(n334), .ZN(N359) );
  INVD1 U210 ( .I(n278), .ZN(n276) );
  INVD1 U211 ( .I(n278), .ZN(n277) );
  INVD1 U212 ( .I(n268), .ZN(n275) );
  INVD1 U213 ( .I(n268), .ZN(n274) );
  BUFFD1 U214 ( .I(ClockW), .Z(n221) );
  BUFFD1 U215 ( .I(ClockW), .Z(n220) );
  BUFFD1 U216 ( .I(n222), .Z(n215) );
  BUFFD1 U217 ( .I(ClockW), .Z(n222) );
  XOR3D1 U218 ( .A1(DataI[2]), .A2(DataI[1]), .A3(n360), .Z(N87) );
  XOR3D1 U219 ( .A1(DataI[0]), .A2(n359), .A3(n358), .Z(n360) );
  XOR3D1 U220 ( .A1(DataI[5]), .A2(DataI[4]), .A3(n357), .Z(n358) );
  XOR3D1 U221 ( .A1(DataI[19]), .A2(DataI[18]), .A3(n351), .Z(n352) );
  XOR3D1 U222 ( .A1(n350), .A2(DataI[17]), .A3(n349), .Z(n351) );
  XOR3D1 U223 ( .A1(n356), .A2(DataI[3]), .A3(n355), .Z(n357) );
  XOR3D1 U224 ( .A1(DataI[12]), .A2(DataI[11]), .A3(n354), .Z(n355) );
  XOR3D1 U225 ( .A1(n353), .A2(DataI[10]), .A3(n352), .Z(n354) );
  MUX4ND0 U226 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n149), .S1(n134), .ZN(
        n110) );
  MUX4ND0 U227 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n150), .S1(n134), .ZN(
        n113) );
  MUX4ND0 U228 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n149), .S1(n134), .ZN(
        n107) );
  MUX4ND0 U229 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n150), .S1(n134), .ZN(
        n116) );
  BUFFD1 U230 ( .I(N48), .Z(n279) );
  MUX4ND0 U231 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n150), .S1(n136), .ZN(n7)
         );
  MUX4ND0 U232 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n150), .S1(n136), .ZN(n10)
         );
  MUX4ND0 U233 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n150), .S1(n135), .ZN(n25)
         );
  MUX4ND0 U234 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n148), .S1(n135), .ZN(
        n40) );
  MUX4ND0 U235 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n149), .S1(n135), .ZN(
        n43) );
  MUX4ND0 U236 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n149), .S1(n134), .ZN(
        n61) );
  MUX4ND0 U237 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n148), .S1(n134), .ZN(
        n64) );
  MUX4ND0 U238 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n150), .S1(n134), .ZN(
        n122) );
  MUX4ND0 U239 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n150), .S1(n134), .ZN(
        n125) );
  MUX4ND0 U240 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n148), .S1(n135), .ZN(n22)
         );
  MUX4ND0 U241 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n149), .S1(n135), .ZN(n28)
         );
  MUX4ND0 U242 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n148), .S1(n135), .ZN(
        n52) );
  MUX4ND0 U243 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n149), .S1(n134), .ZN(
        n101) );
  MUX4ND0 U244 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n150), .S1(n134), .ZN(
        n104) );
  MUX4ND0 U245 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n150), .S1(n136), .ZN(n4)
         );
  MUX4ND0 U246 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n149), .S1(n136), .ZN(n16)
         );
  MUX4ND0 U247 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n148), .S1(n135), .ZN(
        n34) );
  MUX4ND0 U248 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n149), .S1(n135), .ZN(
        n37) );
  MUX4ND0 U249 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n148), .S1(n135), .ZN(
        n46) );
  MUX4ND0 U250 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n149), .S1(n135), .ZN(
        n58) );
  MUX4ND0 U251 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n149), .S1(n134), .ZN(
        n95) );
  MUX4ND0 U252 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n150), .S1(n134), .ZN(
        n119) );
  MUX4ND0 U253 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n150), .S1(n136), .ZN(n13)
         );
  MUX4ND0 U254 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n149), .S1(n136), .ZN(n19)
         );
  MUX4ND0 U255 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n148), .S1(n135), .ZN(n31)
         );
  MUX4ND0 U256 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n148), .S1(n135), .ZN(
        n49) );
  MUX4ND0 U257 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n149), .S1(n135), .ZN(
        n55) );
  MUX4ND0 U258 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n148), .S1(n134), .ZN(
        n98) );
  MUX4ND0 U259 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n150), .S1(n133), .ZN(
        n128) );
  BUFFD1 U260 ( .I(N50), .Z(n281) );
  BUFFD1 U261 ( .I(N49), .Z(n280) );
  INVD1 U262 ( .I(n176), .ZN(n175) );
  INVD1 U263 ( .I(N260), .ZN(n176) );
  NR3D0 U264 ( .A1(n335), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N260) );
  INVD1 U265 ( .I(n208), .ZN(n207) );
  INVD1 U266 ( .I(N99), .ZN(n208) );
  NR3D0 U267 ( .A1(n361), .A2(AddrW[1]), .A3(AddrW[0]), .ZN(N99) );
  INVD1 U268 ( .I(n168), .ZN(n167) );
  INVD1 U269 ( .I(N293), .ZN(n168) );
  NR3D0 U270 ( .A1(n334), .A2(AddrW[1]), .A3(n335), .ZN(N293) );
  INVD1 U271 ( .I(AddrW[1]), .ZN(n336) );
  ND2D1 U272 ( .A1(AddrW[2]), .A2(Write), .ZN(n335) );
  IND2D1 U273 ( .A1(AddrW[2]), .B1(Write), .ZN(n361) );
  INVD1 U274 ( .I(n200), .ZN(n199) );
  INVD1 U275 ( .I(N161), .ZN(n200) );
  NR3D0 U276 ( .A1(n334), .A2(AddrW[1]), .A3(n361), .ZN(N161) );
  INVD1 U277 ( .I(Read), .ZN(n278) );
  OR2D1 U278 ( .A1(n276), .A2(Dreadyr), .Z(n1) );
  CKAN2D0 U279 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  INVD1 U280 ( .I(n269), .ZN(n268) );
  INVD1 U281 ( .I(ClockR), .ZN(n269) );
  CKAN2D0 U282 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U283 ( .I0(n2), .I1(n3), .I2(n4), .S0(n138), .S1(n130), .ZN(N84) );
  MUX3ND0 U284 ( .I0(n5), .I1(n6), .I2(n7), .S0(n138), .S1(n130), .ZN(N83) );
  MUX3ND0 U285 ( .I0(n8), .I1(n9), .I2(n10), .S0(n138), .S1(n130), .ZN(N82) );
  MUX3ND0 U286 ( .I0(n11), .I1(n12), .I2(n13), .S0(n138), .S1(n130), .ZN(N81)
         );
  MUX3ND0 U287 ( .I0(n14), .I1(n15), .I2(n16), .S0(n138), .S1(n130), .ZN(N80)
         );
  MUX3ND0 U288 ( .I0(n17), .I1(n18), .I2(n19), .S0(n138), .S1(n130), .ZN(N79)
         );
  MUX3ND0 U289 ( .I0(n20), .I1(n21), .I2(n22), .S0(n138), .S1(n130), .ZN(N78)
         );
  MUX3ND0 U290 ( .I0(n23), .I1(n24), .I2(n25), .S0(n138), .S1(n131), .ZN(N77)
         );
  MUX3ND0 U291 ( .I0(n26), .I1(n27), .I2(n28), .S0(n138), .S1(n131), .ZN(N76)
         );
  MUX3ND0 U292 ( .I0(n29), .I1(n30), .I2(n31), .S0(n138), .S1(n131), .ZN(N75)
         );
  MUX3ND0 U293 ( .I0(n32), .I1(n33), .I2(n34), .S0(n138), .S1(n131), .ZN(N74)
         );
  MUX3ND0 U294 ( .I0(n35), .I1(n36), .I2(n37), .S0(n138), .S1(n131), .ZN(N73)
         );
  MUX3ND0 U295 ( .I0(n38), .I1(n39), .I2(n40), .S0(n138), .S1(n131), .ZN(N72)
         );
  MUX3ND0 U296 ( .I0(n41), .I1(n42), .I2(n43), .S0(n137), .S1(n131), .ZN(N71)
         );
  MUX3ND0 U297 ( .I0(n44), .I1(n45), .I2(n46), .S0(n137), .S1(n131), .ZN(N70)
         );
  MUX3ND0 U298 ( .I0(n47), .I1(n48), .I2(n49), .S0(n137), .S1(n131), .ZN(N69)
         );
  MUX3ND0 U299 ( .I0(n50), .I1(n51), .I2(n52), .S0(n137), .S1(n131), .ZN(N68)
         );
  MUX3ND0 U300 ( .I0(n53), .I1(n54), .I2(n55), .S0(n137), .S1(n131), .ZN(N67)
         );
  MUX3ND0 U301 ( .I0(n56), .I1(n57), .I2(n58), .S0(n137), .S1(n131), .ZN(N66)
         );
  MUX3ND0 U302 ( .I0(n59), .I1(n60), .I2(n61), .S0(n137), .S1(n131), .ZN(N65)
         );
  MUX3ND0 U303 ( .I0(n62), .I1(n63), .I2(n64), .S0(n137), .S1(n132), .ZN(N64)
         );
  MUX3ND0 U304 ( .I0(n65), .I1(n94), .I2(n95), .S0(n137), .S1(n132), .ZN(N63)
         );
  MUX3ND0 U305 ( .I0(n96), .I1(n97), .I2(n98), .S0(n137), .S1(n132), .ZN(N62)
         );
  MUX3ND0 U306 ( .I0(n99), .I1(n100), .I2(n101), .S0(n137), .S1(n132), .ZN(N61) );
  MUX3ND0 U307 ( .I0(n102), .I1(n103), .I2(n104), .S0(n137), .S1(n132), .ZN(
        N60) );
  MUX3ND0 U308 ( .I0(n105), .I1(n106), .I2(n107), .S0(n137), .S1(n132), .ZN(
        N59) );
  MUX3ND0 U309 ( .I0(n108), .I1(n109), .I2(n110), .S0(n136), .S1(n132), .ZN(
        N58) );
  MUX3ND0 U310 ( .I0(n111), .I1(n112), .I2(n113), .S0(n136), .S1(n132), .ZN(
        N57) );
  MUX3ND0 U311 ( .I0(n114), .I1(n115), .I2(n116), .S0(n136), .S1(n132), .ZN(
        N56) );
  MUX3ND0 U312 ( .I0(n117), .I1(n118), .I2(n119), .S0(n136), .S1(n132), .ZN(
        N55) );
  MUX3ND0 U313 ( .I0(n120), .I1(n121), .I2(n122), .S0(n136), .S1(n132), .ZN(
        N54) );
  MUX3ND0 U314 ( .I0(n123), .I1(n124), .I2(n125), .S0(n136), .S1(n132), .ZN(
        N53) );
  MUX3ND0 U315 ( .I0(n126), .I1(n127), .I2(n128), .S0(n136), .S1(n132), .ZN(
        N52) );
  MUX2ND0 U316 ( .I0(\Storage[2][0] ), .I1(\Storage[3][0] ), .S(n147), .ZN(n3)
         );
  MUX2ND0 U317 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .S(n147), .ZN(n2)
         );
  MUX2ND0 U318 ( .I0(\Storage[2][1] ), .I1(\Storage[3][1] ), .S(n146), .ZN(n6)
         );
  MUX2ND0 U319 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .S(n147), .ZN(n5)
         );
  MUX2ND0 U320 ( .I0(\Storage[2][2] ), .I1(\Storage[3][2] ), .S(n148), .ZN(n9)
         );
  MUX2ND0 U321 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .S(n147), .ZN(n8)
         );
  MUX2ND0 U322 ( .I0(\Storage[2][3] ), .I1(\Storage[3][3] ), .S(n148), .ZN(n12) );
  MUX2ND0 U323 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .S(n148), .ZN(n11) );
  MUX2ND0 U324 ( .I0(\Storage[2][4] ), .I1(\Storage[3][4] ), .S(n147), .ZN(n15) );
  MUX2ND0 U325 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .S(n148), .ZN(n14) );
  MUX2ND0 U326 ( .I0(\Storage[2][5] ), .I1(\Storage[3][5] ), .S(n147), .ZN(n18) );
  MUX2ND0 U327 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .S(n147), .ZN(n17) );
  MUX2ND0 U328 ( .I0(\Storage[2][6] ), .I1(\Storage[3][6] ), .S(n148), .ZN(n21) );
  MUX2ND0 U329 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .S(n147), .ZN(n20) );
  MUX2ND0 U330 ( .I0(\Storage[2][7] ), .I1(\Storage[3][7] ), .S(n147), .ZN(n24) );
  MUX2ND0 U331 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .S(n147), .ZN(n23) );
  MUX2ND0 U332 ( .I0(\Storage[2][8] ), .I1(\Storage[3][8] ), .S(n147), .ZN(n27) );
  MUX2ND0 U333 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .S(n147), .ZN(n26) );
  MUX2ND0 U334 ( .I0(\Storage[2][9] ), .I1(\Storage[3][9] ), .S(n147), .ZN(n30) );
  MUX2ND0 U335 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .S(n147), .ZN(n29) );
  MUX2ND0 U336 ( .I0(\Storage[2][10] ), .I1(\Storage[3][10] ), .S(n147), .ZN(
        n33) );
  MUX2ND0 U337 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .S(n147), .ZN(
        n32) );
  MUX2ND0 U338 ( .I0(\Storage[2][11] ), .I1(\Storage[3][11] ), .S(n147), .ZN(
        n36) );
  MUX2ND0 U339 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .S(n147), .ZN(
        n35) );
  MUX2ND0 U340 ( .I0(\Storage[2][12] ), .I1(\Storage[3][12] ), .S(n147), .ZN(
        n39) );
  MUX2ND0 U341 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .S(n146), .ZN(
        n38) );
  MUX2ND0 U342 ( .I0(\Storage[2][13] ), .I1(\Storage[3][13] ), .S(n146), .ZN(
        n42) );
  MUX2ND0 U343 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .S(n146), .ZN(
        n41) );
  MUX2ND0 U344 ( .I0(\Storage[2][14] ), .I1(\Storage[3][14] ), .S(n146), .ZN(
        n45) );
  MUX2ND0 U345 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .S(n146), .ZN(
        n44) );
  MUX2ND0 U346 ( .I0(\Storage[2][15] ), .I1(\Storage[3][15] ), .S(n146), .ZN(
        n48) );
  MUX2ND0 U347 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .S(n146), .ZN(
        n47) );
  MUX2ND0 U348 ( .I0(\Storage[2][16] ), .I1(\Storage[3][16] ), .S(n146), .ZN(
        n51) );
  MUX2ND0 U349 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .S(n146), .ZN(
        n50) );
  MUX2ND0 U350 ( .I0(\Storage[2][17] ), .I1(\Storage[3][17] ), .S(n146), .ZN(
        n54) );
  MUX2ND0 U351 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .S(n146), .ZN(
        n53) );
  MUX2ND0 U352 ( .I0(\Storage[2][18] ), .I1(\Storage[3][18] ), .S(n146), .ZN(
        n57) );
  MUX2ND0 U353 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .S(n146), .ZN(
        n56) );
  MUX2ND0 U354 ( .I0(\Storage[2][19] ), .I1(\Storage[3][19] ), .S(n146), .ZN(
        n60) );
  MUX2ND0 U355 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .S(n146), .ZN(
        n59) );
  MUX2ND0 U356 ( .I0(\Storage[2][20] ), .I1(\Storage[3][20] ), .S(n146), .ZN(
        n63) );
  MUX2ND0 U357 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .S(n146), .ZN(
        n62) );
  MUX2ND0 U358 ( .I0(\Storage[2][21] ), .I1(\Storage[3][21] ), .S(n146), .ZN(
        n94) );
  MUX2ND0 U359 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .S(n145), .ZN(
        n65) );
  MUX2ND0 U360 ( .I0(\Storage[2][22] ), .I1(\Storage[3][22] ), .S(n145), .ZN(
        n97) );
  MUX2ND0 U361 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .S(n145), .ZN(
        n96) );
  MUX2ND0 U362 ( .I0(\Storage[2][23] ), .I1(\Storage[3][23] ), .S(n145), .ZN(
        n100) );
  MUX2ND0 U363 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .S(n145), .ZN(
        n99) );
  MUX2ND0 U364 ( .I0(\Storage[2][24] ), .I1(\Storage[3][24] ), .S(n145), .ZN(
        n103) );
  MUX2ND0 U365 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .S(n145), .ZN(
        n102) );
  MUX2ND0 U366 ( .I0(\Storage[2][25] ), .I1(\Storage[3][25] ), .S(n145), .ZN(
        n106) );
  MUX2ND0 U367 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .S(n145), .ZN(
        n105) );
  MUX2ND0 U368 ( .I0(\Storage[2][26] ), .I1(\Storage[3][26] ), .S(n145), .ZN(
        n109) );
  MUX2ND0 U369 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .S(n145), .ZN(
        n108) );
  MUX2ND0 U370 ( .I0(\Storage[2][27] ), .I1(\Storage[3][27] ), .S(n145), .ZN(
        n112) );
  MUX2ND0 U371 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .S(n145), .ZN(
        n111) );
  MUX2ND0 U372 ( .I0(\Storage[2][28] ), .I1(\Storage[3][28] ), .S(n145), .ZN(
        n115) );
  MUX2ND0 U373 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .S(n145), .ZN(
        n114) );
  MUX2ND0 U374 ( .I0(\Storage[2][29] ), .I1(\Storage[3][29] ), .S(n145), .ZN(
        n118) );
  MUX2ND0 U375 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .S(n145), .ZN(
        n117) );
  MUX2ND0 U376 ( .I0(\Storage[2][30] ), .I1(\Storage[3][30] ), .S(n145), .ZN(
        n121) );
  MUX2ND0 U377 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .S(n145), .ZN(
        n120) );
  MUX2ND0 U378 ( .I0(\Storage[2][31] ), .I1(\Storage[3][31] ), .S(n145), .ZN(
        n124) );
  MUX2ND0 U379 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .S(n144), .ZN(
        n123) );
  MUX2ND0 U380 ( .I0(\Storage[2][32] ), .I1(\Storage[3][32] ), .S(n147), .ZN(
        n127) );
  MUX2ND0 U381 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .S(n146), .ZN(
        n126) );
endmodule


module PLLTop_1 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_1 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_1 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_1 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_2 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_2 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_2 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_2 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module PLLTop_3 ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry, n1, n2;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator_3 Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(n1) );
  VFO_3 VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(n1) );
  MultiCounter_3 MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(n1) );
  INVD1 U1 ( .I(n2), .ZN(n1) );
  INVD1 U2 ( .I(Reset), .ZN(n2) );
endmodule


module FIFOStateM_AWid4_1 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [3:0] ReadAddr;
  output [3:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   StateClockRaw, StateClock, N47, N48, N49, N50, N51, N67, N68, N69,
         N70, N71, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n88, n89, n93, n133, n134, n135, n136,
         n137, n138, n139, n140, n142, n145, n146, n161, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n767, n768, n769, n770, n771, n772, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820;
  wire   [2:0] NextState;
  wire   [3:0] OldReadAr;
  wire   [3:0] OldWriteAr;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n718), .CPN(StateClock), .Q(FullFIFO) );
  DFND1 EmptyFIFOr_reg ( .D(n722), .CPN(StateClock), .Q(EmptyFIFO), .QN(n726)
         );
  MOAI22D1 U6 ( .A1(n705), .A2(n815), .B1(n815), .B2(OldReadAr[1]), .ZN(n720)
         );
  OA21D1 U11 ( .A1(n698), .A2(n691), .B(n820), .Z(n811) );
  MOAI22D1 U12 ( .A1(n702), .A2(n810), .B1(n810), .B2(OldWriteAr[2]), .ZN(n717) );
  MOAI22D1 U13 ( .A1(n701), .A2(n810), .B1(n810), .B2(OldWriteAr[0]), .ZN(n716) );
  MOAI22D1 U14 ( .A1(n810), .A2(n809), .B1(n810), .B2(OldWriteAr[1]), .ZN(n715) );
  MOAI22D1 U15 ( .A1(n703), .A2(n810), .B1(n810), .B2(OldWriteAr[3]), .ZN(n714) );
  IAO21D1 U31 ( .A1(n782), .A2(n781), .B(n800), .ZN(n783) );
  OA21D1 U34 ( .A1(ReadAddr[2]), .A2(n779), .B(n780), .Z(n774) );
  MOAI22D1 U88 ( .A1(n704), .A2(n815), .B1(n815), .B2(OldReadAr[0]), .ZN(n708)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n719), .CPN(StateClock), .CDN(n693), .Q(
        OldReadAr[3]), .QN(n814) );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n721), .CPN(StateClock), .CDN(n693), .Q(
        OldReadAr[2]), .QN(n816) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n708), .CPN(StateClock), .CDN(n692), .Q(
        OldReadAr[0]) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n714), .CPN(StateClock), .CDN(n692), .Q(
        OldWriteAr[3]) );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n715), .CPN(StateClock), .CDN(n693), .Q(
        OldWriteAr[1]) );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n716), .CPN(StateClock), .CDN(n693), .Q(
        OldWriteAr[0]) );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n717), .CPN(StateClock), .CDN(n693), .Q(
        OldWriteAr[2]) );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n720), .CPN(StateClock), .CDN(n693), .Q(
        OldReadAr[1]) );
  DFNCND1 \NextState_reg[0]  ( .D(n710), .CPN(StateClock), .CDN(n692), .Q(
        NextState[0]), .QN(n723) );
  DFNCND1 \NextState_reg[1]  ( .D(n711), .CPN(StateClock), .CDN(n692), .Q(
        NextState[1]), .QN(n724) );
  DFNCND1 \NextState_reg[2]  ( .D(n713), .CPN(StateClock), .CDN(n692), .Q(
        NextState[2]), .QN(n725) );
  DFNCND1 WriteCmdr_reg ( .D(n712), .CPN(StateClock), .CDN(n692), .Q(WriteCmd)
         );
  DFNCND1 ReadCmdr_reg ( .D(n709), .CPN(StateClock), .CDN(n692), .Q(ReadCmd)
         );
  DFCND1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n692), 
        .QN(n700) );
  DFCND1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n692), 
        .Q(n803), .QN(n698) );
  DFCND1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n692), 
        .QN(n699) );
  EDFCNQD1 \WriteAr_reg[1]  ( .D(N68), .E(n582), .CP(StateClock), .CDN(n693), 
        .Q(WriteAddr[1]) );
  EDFCND1 \ReadAr_reg[3]  ( .D(n1), .E(n352), .CP(StateClock), .CDN(n694), .Q(
        ReadAddr[3]), .QN(n707) );
  EDFCND1 \ReadAr_reg[2]  ( .D(n178), .E(n352), .CP(StateClock), .CDN(n694), 
        .Q(ReadAddr[2]), .QN(n706) );
  EDFCND1 \ReadAr_reg[1]  ( .D(n236), .E(n352), .CP(StateClock), .CDN(n694), 
        .Q(ReadAddr[1]), .QN(n705) );
  EDFCND1 \ReadAr_reg[0]  ( .D(n293), .E(n352), .CP(StateClock), .CDN(n694), 
        .Q(ReadAddr[0]), .QN(n704) );
  EDFCND1 \WriteAr_reg[3]  ( .D(n399), .E(n582), .CP(StateClock), .CDN(n694), 
        .Q(WriteAddr[3]), .QN(n703) );
  EDFCND1 \WriteAr_reg[2]  ( .D(n459), .E(n582), .CP(StateClock), .CDN(n694), 
        .Q(WriteAddr[2]), .QN(n702) );
  EDFCND1 \WriteAr_reg[0]  ( .D(n519), .E(n582), .CP(StateClock), .CDN(n694), 
        .Q(WriteAddr[0]), .QN(n701) );
  CKBD0 U3 ( .CLK(n746), .C(n177) );
  BUFFD0 U4 ( .I(n3), .Z(n1) );
  BUFFD0 U5 ( .I(n4), .Z(n2) );
  BUFFD0 U7 ( .I(n5), .Z(n3) );
  BUFFD0 U8 ( .I(n6), .Z(n4) );
  BUFFD0 U9 ( .I(n7), .Z(n5) );
  BUFFD0 U10 ( .I(n8), .Z(n6) );
  BUFFD0 U16 ( .I(n9), .Z(n7) );
  BUFFD0 U17 ( .I(n10), .Z(n8) );
  BUFFD0 U18 ( .I(n11), .Z(n9) );
  BUFFD0 U19 ( .I(n12), .Z(n10) );
  BUFFD0 U20 ( .I(n13), .Z(n11) );
  BUFFD0 U21 ( .I(n14), .Z(n12) );
  BUFFD0 U22 ( .I(n15), .Z(n13) );
  BUFFD0 U23 ( .I(n16), .Z(n14) );
  BUFFD0 U24 ( .I(n17), .Z(n15) );
  BUFFD0 U25 ( .I(n18), .Z(n16) );
  BUFFD0 U26 ( .I(n19), .Z(n17) );
  BUFFD0 U27 ( .I(n20), .Z(n18) );
  BUFFD0 U28 ( .I(n21), .Z(n19) );
  BUFFD0 U29 ( .I(n22), .Z(n20) );
  BUFFD0 U30 ( .I(n23), .Z(n21) );
  BUFFD0 U32 ( .I(n24), .Z(n22) );
  BUFFD0 U33 ( .I(n25), .Z(n23) );
  BUFFD0 U35 ( .I(n26), .Z(n24) );
  BUFFD0 U36 ( .I(n32), .Z(n25) );
  BUFFD0 U37 ( .I(n27), .Z(n26) );
  BUFFD0 U38 ( .I(n28), .Z(n27) );
  BUFFD0 U39 ( .I(n29), .Z(n28) );
  BUFFD0 U40 ( .I(n30), .Z(n29) );
  BUFFD0 U41 ( .I(n31), .Z(n30) );
  CKBD0 U42 ( .CLK(n707), .C(n458) );
  BUFFD0 U43 ( .I(n33), .Z(n31) );
  BUFFD0 U44 ( .I(N51), .Z(n32) );
  BUFFD0 U45 ( .I(n34), .Z(n33) );
  BUFFD0 U46 ( .I(n88), .Z(n34) );
  BUFFD0 U47 ( .I(n89), .Z(n88) );
  BUFFD0 U48 ( .I(n93), .Z(n89) );
  BUFFD0 U49 ( .I(n133), .Z(n93) );
  BUFFD0 U50 ( .I(n134), .Z(n133) );
  BUFFD0 U51 ( .I(n135), .Z(n134) );
  BUFFD0 U52 ( .I(n136), .Z(n135) );
  BUFFD0 U53 ( .I(n137), .Z(n136) );
  BUFFD0 U54 ( .I(n138), .Z(n137) );
  BUFFD0 U55 ( .I(n139), .Z(n138) );
  BUFFD0 U56 ( .I(n140), .Z(n139) );
  BUFFD0 U57 ( .I(n142), .Z(n140) );
  BUFFD0 U58 ( .I(n145), .Z(n142) );
  BUFFD0 U59 ( .I(n146), .Z(n145) );
  BUFFD0 U60 ( .I(n161), .Z(n146) );
  BUFFD0 U61 ( .I(n173), .Z(n161) );
  BUFFD0 U62 ( .I(n174), .Z(n173) );
  BUFFD0 U63 ( .I(n175), .Z(n174) );
  BUFFD0 U64 ( .I(n176), .Z(n175) );
  BUFFD0 U65 ( .I(n177), .Z(n176) );
  XNR2D0 U66 ( .A1(n458), .A2(n729), .ZN(n746) );
  BUFFD0 U67 ( .I(n179), .Z(n178) );
  BUFFD0 U68 ( .I(n180), .Z(n179) );
  BUFFD0 U69 ( .I(n181), .Z(n180) );
  BUFFD0 U70 ( .I(n182), .Z(n181) );
  BUFFD0 U71 ( .I(n183), .Z(n182) );
  BUFFD0 U72 ( .I(n184), .Z(n183) );
  BUFFD0 U73 ( .I(n185), .Z(n184) );
  BUFFD0 U74 ( .I(n186), .Z(n185) );
  BUFFD0 U75 ( .I(n187), .Z(n186) );
  BUFFD0 U76 ( .I(n188), .Z(n187) );
  BUFFD0 U77 ( .I(n189), .Z(n188) );
  BUFFD0 U78 ( .I(n190), .Z(n189) );
  BUFFD0 U79 ( .I(n191), .Z(n190) );
  BUFFD0 U80 ( .I(n192), .Z(n191) );
  BUFFD0 U81 ( .I(n193), .Z(n192) );
  BUFFD0 U82 ( .I(n194), .Z(n193) );
  BUFFD0 U83 ( .I(n195), .Z(n194) );
  BUFFD0 U84 ( .I(n196), .Z(n195) );
  BUFFD0 U85 ( .I(n197), .Z(n196) );
  BUFFD0 U86 ( .I(n198), .Z(n197) );
  BUFFD0 U87 ( .I(n199), .Z(n198) );
  BUFFD0 U89 ( .I(n200), .Z(n199) );
  BUFFD0 U90 ( .I(n201), .Z(n200) );
  BUFFD0 U91 ( .I(n202), .Z(n201) );
  BUFFD0 U92 ( .I(n203), .Z(n202) );
  BUFFD0 U93 ( .I(n204), .Z(n203) );
  BUFFD0 U94 ( .I(n205), .Z(n204) );
  BUFFD0 U95 ( .I(n206), .Z(n205) );
  BUFFD0 U96 ( .I(n207), .Z(n206) );
  BUFFD0 U97 ( .I(n208), .Z(n207) );
  BUFFD0 U98 ( .I(n209), .Z(n208) );
  BUFFD0 U99 ( .I(n210), .Z(n209) );
  BUFFD0 U100 ( .I(n211), .Z(n210) );
  BUFFD0 U101 ( .I(n212), .Z(n211) );
  BUFFD0 U102 ( .I(n213), .Z(n212) );
  BUFFD0 U103 ( .I(n214), .Z(n213) );
  BUFFD0 U104 ( .I(n215), .Z(n214) );
  BUFFD0 U105 ( .I(n216), .Z(n215) );
  BUFFD0 U106 ( .I(n217), .Z(n216) );
  BUFFD0 U107 ( .I(n218), .Z(n217) );
  BUFFD0 U108 ( .I(n219), .Z(n218) );
  BUFFD0 U109 ( .I(n220), .Z(n219) );
  BUFFD0 U110 ( .I(n221), .Z(n220) );
  BUFFD0 U111 ( .I(n222), .Z(n221) );
  BUFFD0 U112 ( .I(n223), .Z(n222) );
  BUFFD0 U113 ( .I(n224), .Z(n223) );
  BUFFD0 U114 ( .I(n225), .Z(n224) );
  BUFFD0 U115 ( .I(n226), .Z(n225) );
  BUFFD0 U116 ( .I(n227), .Z(n226) );
  BUFFD0 U117 ( .I(n228), .Z(n227) );
  BUFFD0 U118 ( .I(n229), .Z(n228) );
  BUFFD0 U119 ( .I(n230), .Z(n229) );
  BUFFD0 U120 ( .I(n231), .Z(n230) );
  BUFFD0 U121 ( .I(n232), .Z(n231) );
  BUFFD0 U122 ( .I(n233), .Z(n232) );
  BUFFD0 U123 ( .I(n234), .Z(n233) );
  BUFFD0 U124 ( .I(N49), .Z(n234) );
  CKBD0 U125 ( .CLK(ReadAddr[2]), .C(n235) );
  OAI21D0 U126 ( .A1(n728), .A2(n235), .B(n729), .ZN(n744) );
  BUFFD0 U127 ( .I(n237), .Z(n236) );
  BUFFD0 U128 ( .I(n239), .Z(n237) );
  BUFFD0 U129 ( .I(n240), .Z(n238) );
  BUFFD0 U130 ( .I(n241), .Z(n239) );
  BUFFD0 U131 ( .I(n242), .Z(n240) );
  BUFFD0 U132 ( .I(n243), .Z(n241) );
  BUFFD0 U133 ( .I(n244), .Z(n242) );
  BUFFD0 U134 ( .I(n245), .Z(n243) );
  BUFFD0 U135 ( .I(n246), .Z(n244) );
  BUFFD0 U136 ( .I(n247), .Z(n245) );
  BUFFD0 U137 ( .I(n248), .Z(n246) );
  BUFFD0 U138 ( .I(n249), .Z(n247) );
  BUFFD0 U139 ( .I(n250), .Z(n248) );
  BUFFD0 U140 ( .I(n251), .Z(n249) );
  BUFFD0 U141 ( .I(n252), .Z(n250) );
  BUFFD0 U142 ( .I(n253), .Z(n251) );
  BUFFD0 U143 ( .I(n254), .Z(n252) );
  BUFFD0 U144 ( .I(n255), .Z(n253) );
  BUFFD0 U145 ( .I(n256), .Z(n254) );
  BUFFD0 U146 ( .I(n257), .Z(n255) );
  BUFFD0 U147 ( .I(n258), .Z(n256) );
  BUFFD0 U148 ( .I(n259), .Z(n257) );
  BUFFD0 U149 ( .I(n260), .Z(n258) );
  BUFFD0 U150 ( .I(n261), .Z(n259) );
  BUFFD0 U151 ( .I(n262), .Z(n260) );
  BUFFD0 U152 ( .I(n263), .Z(n261) );
  BUFFD0 U153 ( .I(n264), .Z(n262) );
  BUFFD0 U154 ( .I(n265), .Z(n263) );
  BUFFD0 U155 ( .I(n266), .Z(n264) );
  BUFFD0 U156 ( .I(N48), .Z(n265) );
  BUFFD0 U157 ( .I(n267), .Z(n266) );
  BUFFD0 U158 ( .I(n268), .Z(n267) );
  BUFFD0 U159 ( .I(n269), .Z(n268) );
  BUFFD0 U160 ( .I(n270), .Z(n269) );
  BUFFD0 U161 ( .I(n271), .Z(n270) );
  BUFFD0 U162 ( .I(n272), .Z(n271) );
  BUFFD0 U163 ( .I(n273), .Z(n272) );
  BUFFD0 U164 ( .I(n274), .Z(n273) );
  BUFFD0 U165 ( .I(n275), .Z(n274) );
  BUFFD0 U166 ( .I(n276), .Z(n275) );
  BUFFD0 U167 ( .I(n277), .Z(n276) );
  BUFFD0 U168 ( .I(n278), .Z(n277) );
  BUFFD0 U169 ( .I(n279), .Z(n278) );
  BUFFD0 U170 ( .I(n280), .Z(n279) );
  BUFFD0 U171 ( .I(n281), .Z(n280) );
  BUFFD0 U172 ( .I(n282), .Z(n281) );
  BUFFD0 U173 ( .I(n283), .Z(n282) );
  BUFFD0 U174 ( .I(n284), .Z(n283) );
  BUFFD0 U175 ( .I(n285), .Z(n284) );
  BUFFD0 U176 ( .I(n286), .Z(n285) );
  BUFFD0 U177 ( .I(n287), .Z(n286) );
  BUFFD0 U178 ( .I(n288), .Z(n287) );
  BUFFD0 U179 ( .I(n289), .Z(n288) );
  BUFFD0 U180 ( .I(n290), .Z(n289) );
  BUFFD0 U181 ( .I(n727), .Z(n290) );
  BUFFD0 U182 ( .I(n292), .Z(n291) );
  BUFFD0 U183 ( .I(ReadAddr[1]), .Z(n292) );
  XNR2D0 U184 ( .A1(n291), .A2(n294), .ZN(n727) );
  BUFFD0 U185 ( .I(n295), .Z(n293) );
  BUFFD0 U186 ( .I(n296), .Z(n294) );
  BUFFD0 U187 ( .I(n297), .Z(n295) );
  BUFFD0 U188 ( .I(n298), .Z(n296) );
  BUFFD0 U189 ( .I(n299), .Z(n297) );
  BUFFD0 U190 ( .I(n300), .Z(n298) );
  BUFFD0 U191 ( .I(n301), .Z(n299) );
  BUFFD0 U192 ( .I(n302), .Z(n300) );
  BUFFD0 U193 ( .I(n303), .Z(n301) );
  BUFFD0 U194 ( .I(n304), .Z(n302) );
  BUFFD0 U195 ( .I(n305), .Z(n303) );
  BUFFD0 U196 ( .I(n306), .Z(n304) );
  BUFFD0 U197 ( .I(n307), .Z(n305) );
  BUFFD0 U198 ( .I(n308), .Z(n306) );
  BUFFD0 U199 ( .I(n309), .Z(n307) );
  BUFFD0 U200 ( .I(n310), .Z(n308) );
  BUFFD0 U201 ( .I(n311), .Z(n309) );
  BUFFD0 U202 ( .I(n312), .Z(n310) );
  BUFFD0 U203 ( .I(n313), .Z(n311) );
  BUFFD0 U204 ( .I(n314), .Z(n312) );
  BUFFD0 U205 ( .I(n315), .Z(n313) );
  BUFFD0 U206 ( .I(n316), .Z(n314) );
  BUFFD0 U207 ( .I(n317), .Z(n315) );
  BUFFD0 U208 ( .I(n318), .Z(n316) );
  BUFFD0 U209 ( .I(n319), .Z(n317) );
  BUFFD0 U210 ( .I(n320), .Z(n318) );
  BUFFD0 U211 ( .I(n321), .Z(n319) );
  BUFFD0 U212 ( .I(n322), .Z(n320) );
  BUFFD0 U213 ( .I(n323), .Z(n321) );
  BUFFD0 U214 ( .I(n324), .Z(n322) );
  BUFFD0 U215 ( .I(n325), .Z(n323) );
  BUFFD0 U216 ( .I(n326), .Z(n324) );
  BUFFD0 U217 ( .I(n327), .Z(n325) );
  BUFFD0 U218 ( .I(n328), .Z(n326) );
  BUFFD0 U219 ( .I(n329), .Z(n327) );
  BUFFD0 U220 ( .I(n330), .Z(n328) );
  BUFFD0 U221 ( .I(N47), .Z(n329) );
  BUFFD0 U222 ( .I(n331), .Z(n330) );
  BUFFD0 U223 ( .I(n332), .Z(n331) );
  BUFFD0 U224 ( .I(n333), .Z(n332) );
  BUFFD0 U225 ( .I(n334), .Z(n333) );
  BUFFD0 U226 ( .I(n335), .Z(n334) );
  BUFFD0 U227 ( .I(n336), .Z(n335) );
  BUFFD0 U228 ( .I(n337), .Z(n336) );
  BUFFD0 U229 ( .I(n338), .Z(n337) );
  BUFFD0 U230 ( .I(n339), .Z(n338) );
  BUFFD0 U231 ( .I(n340), .Z(n339) );
  BUFFD0 U232 ( .I(n341), .Z(n340) );
  BUFFD0 U233 ( .I(n342), .Z(n341) );
  BUFFD0 U234 ( .I(n343), .Z(n342) );
  BUFFD0 U235 ( .I(n344), .Z(n343) );
  BUFFD0 U236 ( .I(n345), .Z(n344) );
  BUFFD0 U237 ( .I(n346), .Z(n345) );
  BUFFD0 U238 ( .I(n347), .Z(n346) );
  BUFFD0 U239 ( .I(n348), .Z(n347) );
  BUFFD0 U240 ( .I(n349), .Z(n348) );
  BUFFD0 U241 ( .I(n350), .Z(n349) );
  BUFFD0 U242 ( .I(n351), .Z(n350) );
  BUFFD0 U243 ( .I(ReadAddr[0]), .Z(n351) );
  BUFFD0 U244 ( .I(n354), .Z(n352) );
  BUFFD0 U245 ( .I(n355), .Z(n353) );
  BUFFD0 U246 ( .I(n356), .Z(n354) );
  BUFFD0 U247 ( .I(n357), .Z(n355) );
  BUFFD0 U248 ( .I(n358), .Z(n356) );
  BUFFD0 U249 ( .I(n359), .Z(n357) );
  BUFFD0 U250 ( .I(n360), .Z(n358) );
  BUFFD0 U251 ( .I(n361), .Z(n359) );
  BUFFD0 U252 ( .I(n362), .Z(n360) );
  BUFFD0 U253 ( .I(n363), .Z(n361) );
  BUFFD0 U254 ( .I(n380), .Z(n362) );
  BUFFD0 U255 ( .I(n364), .Z(n363) );
  BUFFD0 U256 ( .I(n365), .Z(n364) );
  BUFFD0 U257 ( .I(n366), .Z(n365) );
  BUFFD0 U258 ( .I(n367), .Z(n366) );
  BUFFD0 U259 ( .I(n368), .Z(n367) );
  BUFFD0 U260 ( .I(n369), .Z(n368) );
  BUFFD0 U261 ( .I(n370), .Z(n369) );
  BUFFD0 U262 ( .I(n371), .Z(n370) );
  BUFFD0 U263 ( .I(n372), .Z(n371) );
  BUFFD0 U264 ( .I(n373), .Z(n372) );
  BUFFD0 U265 ( .I(n374), .Z(n373) );
  BUFFD0 U266 ( .I(n375), .Z(n374) );
  BUFFD0 U267 ( .I(n376), .Z(n375) );
  BUFFD0 U268 ( .I(n377), .Z(n376) );
  BUFFD0 U269 ( .I(n378), .Z(n377) );
  BUFFD0 U270 ( .I(n379), .Z(n378) );
  BUFFD0 U271 ( .I(n631), .Z(n379) );
  BUFFD0 U272 ( .I(N50), .Z(n380) );
  BUFFD0 U273 ( .I(n820), .Z(n381) );
  BUFFD0 U274 ( .I(n381), .Z(n382) );
  BUFFD0 U275 ( .I(n382), .Z(n383) );
  BUFFD0 U276 ( .I(n383), .Z(n384) );
  BUFFD0 U277 ( .I(n384), .Z(n385) );
  BUFFD0 U278 ( .I(n385), .Z(n386) );
  BUFFD0 U279 ( .I(n386), .Z(n387) );
  BUFFD0 U280 ( .I(n387), .Z(n388) );
  BUFFD0 U281 ( .I(n388), .Z(n389) );
  BUFFD0 U282 ( .I(n389), .Z(n390) );
  BUFFD0 U283 ( .I(n390), .Z(n391) );
  BUFFD0 U284 ( .I(n391), .Z(n392) );
  BUFFD0 U285 ( .I(n392), .Z(n393) );
  BUFFD0 U286 ( .I(n393), .Z(n394) );
  BUFFD0 U287 ( .I(n394), .Z(n395) );
  BUFFD0 U288 ( .I(n395), .Z(n396) );
  BUFFD0 U289 ( .I(n396), .Z(n397) );
  BUFFD0 U290 ( .I(n397), .Z(n398) );
  BUFFD0 U291 ( .I(n404), .Z(n399) );
  BUFFD0 U292 ( .I(N70), .Z(n400) );
  BUFFD0 U293 ( .I(n400), .Z(n401) );
  BUFFD0 U294 ( .I(n401), .Z(n402) );
  BUFFD0 U295 ( .I(n402), .Z(n403) );
  BUFFD0 U296 ( .I(n405), .Z(n404) );
  BUFFD0 U297 ( .I(n406), .Z(n405) );
  BUFFD0 U298 ( .I(n407), .Z(n406) );
  BUFFD0 U299 ( .I(n408), .Z(n407) );
  BUFFD0 U300 ( .I(n409), .Z(n408) );
  BUFFD0 U301 ( .I(n410), .Z(n409) );
  BUFFD0 U302 ( .I(n411), .Z(n410) );
  BUFFD0 U303 ( .I(n412), .Z(n411) );
  BUFFD0 U304 ( .I(n413), .Z(n412) );
  BUFFD0 U305 ( .I(n414), .Z(n413) );
  BUFFD0 U306 ( .I(n415), .Z(n414) );
  BUFFD0 U307 ( .I(n416), .Z(n415) );
  BUFFD0 U308 ( .I(n417), .Z(n416) );
  BUFFD0 U309 ( .I(n418), .Z(n417) );
  BUFFD0 U310 ( .I(n419), .Z(n418) );
  BUFFD0 U311 ( .I(n420), .Z(n419) );
  BUFFD0 U312 ( .I(n421), .Z(n420) );
  BUFFD0 U313 ( .I(n422), .Z(n421) );
  BUFFD0 U314 ( .I(n423), .Z(n422) );
  BUFFD0 U315 ( .I(n424), .Z(n423) );
  BUFFD0 U316 ( .I(n425), .Z(n424) );
  BUFFD0 U317 ( .I(n426), .Z(n425) );
  BUFFD0 U318 ( .I(n427), .Z(n426) );
  BUFFD0 U319 ( .I(n428), .Z(n427) );
  BUFFD0 U320 ( .I(n429), .Z(n428) );
  BUFFD0 U321 ( .I(n430), .Z(n429) );
  BUFFD0 U322 ( .I(n431), .Z(n430) );
  BUFFD0 U323 ( .I(n432), .Z(n431) );
  BUFFD0 U324 ( .I(n433), .Z(n432) );
  BUFFD0 U325 ( .I(n434), .Z(n433) );
  BUFFD0 U326 ( .I(n435), .Z(n434) );
  BUFFD0 U327 ( .I(n436), .Z(n435) );
  BUFFD0 U328 ( .I(n437), .Z(n436) );
  BUFFD0 U329 ( .I(n438), .Z(n437) );
  BUFFD0 U330 ( .I(n439), .Z(n438) );
  BUFFD0 U331 ( .I(n440), .Z(n439) );
  BUFFD0 U332 ( .I(n441), .Z(n440) );
  BUFFD0 U333 ( .I(n442), .Z(n441) );
  BUFFD0 U334 ( .I(n443), .Z(n442) );
  BUFFD0 U335 ( .I(n444), .Z(n443) );
  BUFFD0 U336 ( .I(n445), .Z(n444) );
  BUFFD0 U337 ( .I(n446), .Z(n445) );
  BUFFD0 U338 ( .I(n447), .Z(n446) );
  BUFFD0 U339 ( .I(n448), .Z(n447) );
  BUFFD0 U340 ( .I(n449), .Z(n448) );
  BUFFD0 U341 ( .I(n450), .Z(n449) );
  BUFFD0 U342 ( .I(n451), .Z(n450) );
  BUFFD0 U343 ( .I(n452), .Z(n451) );
  BUFFD0 U344 ( .I(n453), .Z(n452) );
  BUFFD0 U345 ( .I(n454), .Z(n453) );
  BUFFD0 U346 ( .I(n455), .Z(n454) );
  BUFFD0 U347 ( .I(n456), .Z(n455) );
  BUFFD0 U348 ( .I(n457), .Z(n456) );
  BUFFD0 U349 ( .I(n403), .Z(n457) );
  XNR2D0 U350 ( .A1(n732), .A2(WriteAddr[3]), .ZN(n759) );
  BUFFD0 U351 ( .I(n464), .Z(n459) );
  BUFFD0 U352 ( .I(N69), .Z(n460) );
  BUFFD0 U353 ( .I(n460), .Z(n461) );
  BUFFD0 U354 ( .I(n461), .Z(n462) );
  BUFFD0 U355 ( .I(n462), .Z(n463) );
  BUFFD0 U356 ( .I(n465), .Z(n464) );
  BUFFD0 U357 ( .I(n466), .Z(n465) );
  BUFFD0 U358 ( .I(n467), .Z(n466) );
  BUFFD0 U359 ( .I(n468), .Z(n467) );
  BUFFD0 U360 ( .I(n469), .Z(n468) );
  BUFFD0 U361 ( .I(n470), .Z(n469) );
  BUFFD0 U362 ( .I(n471), .Z(n470) );
  BUFFD0 U363 ( .I(n472), .Z(n471) );
  BUFFD0 U364 ( .I(n473), .Z(n472) );
  BUFFD0 U365 ( .I(n474), .Z(n473) );
  BUFFD0 U366 ( .I(n475), .Z(n474) );
  BUFFD0 U367 ( .I(n476), .Z(n475) );
  BUFFD0 U368 ( .I(n477), .Z(n476) );
  BUFFD0 U369 ( .I(n478), .Z(n477) );
  BUFFD0 U370 ( .I(n479), .Z(n478) );
  BUFFD0 U371 ( .I(n480), .Z(n479) );
  BUFFD0 U372 ( .I(n481), .Z(n480) );
  BUFFD0 U373 ( .I(n482), .Z(n481) );
  BUFFD0 U374 ( .I(n483), .Z(n482) );
  BUFFD0 U375 ( .I(n484), .Z(n483) );
  BUFFD0 U376 ( .I(n485), .Z(n484) );
  BUFFD0 U377 ( .I(n486), .Z(n485) );
  BUFFD0 U378 ( .I(n487), .Z(n486) );
  BUFFD0 U379 ( .I(n488), .Z(n487) );
  BUFFD0 U380 ( .I(n489), .Z(n488) );
  BUFFD0 U381 ( .I(n490), .Z(n489) );
  BUFFD0 U382 ( .I(n491), .Z(n490) );
  BUFFD0 U383 ( .I(n492), .Z(n491) );
  BUFFD0 U384 ( .I(n493), .Z(n492) );
  BUFFD0 U385 ( .I(n494), .Z(n493) );
  BUFFD0 U386 ( .I(n495), .Z(n494) );
  BUFFD0 U387 ( .I(n496), .Z(n495) );
  BUFFD0 U388 ( .I(n497), .Z(n496) );
  BUFFD0 U389 ( .I(n498), .Z(n497) );
  BUFFD0 U390 ( .I(n499), .Z(n498) );
  BUFFD0 U391 ( .I(n500), .Z(n499) );
  BUFFD0 U392 ( .I(n501), .Z(n500) );
  BUFFD0 U393 ( .I(n502), .Z(n501) );
  BUFFD0 U394 ( .I(n503), .Z(n502) );
  BUFFD0 U395 ( .I(n504), .Z(n503) );
  BUFFD0 U396 ( .I(n505), .Z(n504) );
  BUFFD0 U397 ( .I(n506), .Z(n505) );
  BUFFD0 U398 ( .I(n507), .Z(n506) );
  BUFFD0 U399 ( .I(n508), .Z(n507) );
  BUFFD0 U400 ( .I(n509), .Z(n508) );
  BUFFD0 U401 ( .I(n510), .Z(n509) );
  BUFFD0 U402 ( .I(n511), .Z(n510) );
  BUFFD0 U403 ( .I(n512), .Z(n511) );
  BUFFD0 U404 ( .I(n513), .Z(n512) );
  BUFFD0 U405 ( .I(n514), .Z(n513) );
  BUFFD0 U406 ( .I(n515), .Z(n514) );
  BUFFD0 U407 ( .I(n516), .Z(n515) );
  BUFFD0 U408 ( .I(n517), .Z(n516) );
  BUFFD0 U409 ( .I(n518), .Z(n517) );
  BUFFD0 U410 ( .I(n463), .Z(n518) );
  BUFFD0 U411 ( .I(n524), .Z(n519) );
  BUFFD0 U412 ( .I(N67), .Z(n520) );
  BUFFD0 U413 ( .I(n520), .Z(n521) );
  BUFFD0 U414 ( .I(n521), .Z(n522) );
  BUFFD0 U415 ( .I(n522), .Z(n523) );
  BUFFD0 U416 ( .I(n525), .Z(n524) );
  BUFFD0 U417 ( .I(n526), .Z(n525) );
  BUFFD0 U418 ( .I(n527), .Z(n526) );
  BUFFD0 U419 ( .I(n528), .Z(n527) );
  BUFFD0 U420 ( .I(n529), .Z(n528) );
  BUFFD0 U421 ( .I(n530), .Z(n529) );
  BUFFD0 U422 ( .I(n531), .Z(n530) );
  BUFFD0 U423 ( .I(n532), .Z(n531) );
  BUFFD0 U424 ( .I(n533), .Z(n532) );
  BUFFD0 U425 ( .I(n534), .Z(n533) );
  BUFFD0 U426 ( .I(n535), .Z(n534) );
  BUFFD0 U427 ( .I(n536), .Z(n535) );
  BUFFD0 U428 ( .I(n537), .Z(n536) );
  BUFFD0 U429 ( .I(n538), .Z(n537) );
  BUFFD0 U430 ( .I(n539), .Z(n538) );
  BUFFD0 U431 ( .I(n540), .Z(n539) );
  BUFFD0 U432 ( .I(n541), .Z(n540) );
  BUFFD0 U433 ( .I(n542), .Z(n541) );
  BUFFD0 U434 ( .I(n543), .Z(n542) );
  BUFFD0 U435 ( .I(n544), .Z(n543) );
  BUFFD0 U436 ( .I(n545), .Z(n544) );
  BUFFD0 U437 ( .I(n546), .Z(n545) );
  BUFFD0 U438 ( .I(n547), .Z(n546) );
  BUFFD0 U439 ( .I(n548), .Z(n547) );
  BUFFD0 U440 ( .I(n549), .Z(n548) );
  BUFFD0 U441 ( .I(n550), .Z(n549) );
  BUFFD0 U442 ( .I(n551), .Z(n550) );
  BUFFD0 U443 ( .I(n552), .Z(n551) );
  BUFFD0 U444 ( .I(n553), .Z(n552) );
  BUFFD0 U445 ( .I(n554), .Z(n553) );
  BUFFD0 U446 ( .I(n555), .Z(n554) );
  BUFFD0 U447 ( .I(n556), .Z(n555) );
  BUFFD0 U448 ( .I(n557), .Z(n556) );
  BUFFD0 U449 ( .I(n558), .Z(n557) );
  BUFFD0 U450 ( .I(n559), .Z(n558) );
  BUFFD0 U451 ( .I(n560), .Z(n559) );
  BUFFD0 U452 ( .I(n561), .Z(n560) );
  BUFFD0 U453 ( .I(n562), .Z(n561) );
  BUFFD0 U454 ( .I(n563), .Z(n562) );
  BUFFD0 U455 ( .I(n564), .Z(n563) );
  BUFFD0 U456 ( .I(n565), .Z(n564) );
  BUFFD0 U457 ( .I(n566), .Z(n565) );
  BUFFD0 U458 ( .I(n567), .Z(n566) );
  BUFFD0 U459 ( .I(n568), .Z(n567) );
  BUFFD0 U460 ( .I(n569), .Z(n568) );
  BUFFD0 U461 ( .I(n570), .Z(n569) );
  BUFFD0 U462 ( .I(n571), .Z(n570) );
  BUFFD0 U463 ( .I(n572), .Z(n571) );
  BUFFD0 U464 ( .I(n573), .Z(n572) );
  BUFFD0 U465 ( .I(n574), .Z(n573) );
  BUFFD0 U466 ( .I(n575), .Z(n574) );
  BUFFD0 U467 ( .I(n576), .Z(n575) );
  BUFFD0 U468 ( .I(n577), .Z(n576) );
  BUFFD0 U469 ( .I(n578), .Z(n577) );
  BUFFD0 U470 ( .I(n523), .Z(n578) );
  ND3D8 U471 ( .A1(n813), .A2(n631), .A3(n799), .ZN(N71) );
  BUFFD0 U472 ( .I(N71), .Z(n579) );
  BUFFD0 U473 ( .I(n579), .Z(n580) );
  BUFFD0 U474 ( .I(n580), .Z(n581) );
  BUFFD0 U475 ( .I(n583), .Z(n582) );
  BUFFD0 U476 ( .I(n584), .Z(n583) );
  BUFFD0 U477 ( .I(n585), .Z(n584) );
  BUFFD0 U478 ( .I(n586), .Z(n585) );
  BUFFD0 U479 ( .I(n587), .Z(n586) );
  BUFFD0 U480 ( .I(n588), .Z(n587) );
  BUFFD0 U481 ( .I(n589), .Z(n588) );
  BUFFD0 U482 ( .I(n590), .Z(n589) );
  BUFFD0 U483 ( .I(n591), .Z(n590) );
  BUFFD0 U484 ( .I(n592), .Z(n591) );
  BUFFD0 U485 ( .I(n593), .Z(n592) );
  BUFFD0 U486 ( .I(n594), .Z(n593) );
  BUFFD0 U487 ( .I(n595), .Z(n594) );
  BUFFD0 U488 ( .I(n596), .Z(n595) );
  BUFFD0 U489 ( .I(n597), .Z(n596) );
  BUFFD0 U490 ( .I(n598), .Z(n597) );
  BUFFD0 U491 ( .I(n599), .Z(n598) );
  BUFFD0 U492 ( .I(n600), .Z(n599) );
  BUFFD0 U493 ( .I(n601), .Z(n600) );
  BUFFD0 U494 ( .I(n602), .Z(n601) );
  BUFFD0 U495 ( .I(n603), .Z(n602) );
  BUFFD0 U496 ( .I(n604), .Z(n603) );
  BUFFD0 U497 ( .I(n605), .Z(n604) );
  BUFFD0 U498 ( .I(n606), .Z(n605) );
  BUFFD0 U499 ( .I(n607), .Z(n606) );
  BUFFD0 U500 ( .I(n608), .Z(n607) );
  BUFFD0 U501 ( .I(n609), .Z(n608) );
  BUFFD0 U502 ( .I(n610), .Z(n609) );
  BUFFD0 U503 ( .I(n611), .Z(n610) );
  BUFFD0 U504 ( .I(n612), .Z(n611) );
  BUFFD0 U505 ( .I(n613), .Z(n612) );
  BUFFD0 U506 ( .I(n614), .Z(n613) );
  BUFFD0 U507 ( .I(n615), .Z(n614) );
  BUFFD0 U508 ( .I(n616), .Z(n615) );
  BUFFD0 U509 ( .I(n617), .Z(n616) );
  BUFFD0 U510 ( .I(n618), .Z(n617) );
  BUFFD0 U511 ( .I(n619), .Z(n618) );
  BUFFD0 U512 ( .I(n620), .Z(n619) );
  BUFFD0 U513 ( .I(n621), .Z(n620) );
  BUFFD0 U514 ( .I(n622), .Z(n621) );
  BUFFD0 U515 ( .I(n623), .Z(n622) );
  BUFFD0 U516 ( .I(n624), .Z(n623) );
  BUFFD0 U517 ( .I(n625), .Z(n624) );
  BUFFD0 U518 ( .I(n626), .Z(n625) );
  BUFFD0 U519 ( .I(n627), .Z(n626) );
  BUFFD0 U520 ( .I(n628), .Z(n627) );
  BUFFD0 U521 ( .I(n629), .Z(n628) );
  BUFFD0 U522 ( .I(n630), .Z(n629) );
  BUFFD0 U523 ( .I(n581), .Z(n630) );
  ND3D0 U524 ( .A1(n699), .A2(n691), .A3(n698), .ZN(n820) );
  INVD0 U525 ( .I(n802), .ZN(n813) );
  BUFFD0 U526 ( .I(n398), .Z(n631) );
  INVD1 U527 ( .I(n696), .ZN(n693) );
  INVD1 U528 ( .I(n695), .ZN(n694) );
  BUFFD1 U529 ( .I(Reset), .Z(n695) );
  BUFFD1 U530 ( .I(Reset), .Z(n696) );
  INVD1 U531 ( .I(n697), .ZN(n692) );
  BUFFD1 U532 ( .I(Reset), .Z(n697) );
  ND2D1 U533 ( .A1(n789), .A2(n813), .ZN(n739) );
  INVD1 U534 ( .I(n807), .ZN(n806) );
  INVD1 U535 ( .I(n815), .ZN(n817) );
  MAOI22D0 U536 ( .A1(n786), .A2(n691), .B1(n691), .B2(n784), .ZN(n789) );
  OAI211D1 U537 ( .A1(n820), .A2(n792), .B(n789), .C(n743), .ZN(n807) );
  INR2D1 U538 ( .A1(n784), .B1(n742), .ZN(n743) );
  AOI21D1 U539 ( .A1(n803), .A2(n741), .B(n691), .ZN(n742) );
  ND2D1 U540 ( .A1(WriteReq), .A2(n808), .ZN(n810) );
  ND2D1 U541 ( .A1(ReadReq), .A2(n739), .ZN(n815) );
  ND2D1 U542 ( .A1(n789), .A2(n820), .ZN(n808) );
  AOI21D1 U543 ( .A1(n779), .A2(n772), .B(ReadAddr[1]), .ZN(n753) );
  INVD1 U544 ( .I(n752), .ZN(n779) );
  OA211D0 U545 ( .A1(n780), .A2(n779), .B(n778), .C(n777), .Z(n800) );
  INVD1 U546 ( .I(n770), .ZN(n778) );
  NR3D0 U547 ( .A1(n776), .A2(n775), .A3(n774), .ZN(n777) );
  NR3D0 U548 ( .A1(WriteAddr[2]), .A2(n809), .A3(ReadAddr[2]), .ZN(n775) );
  ND2D1 U549 ( .A1(n728), .A2(n235), .ZN(n729) );
  ND2D1 U550 ( .A1(n751), .A2(n750), .ZN(n770) );
  XNR2D1 U551 ( .A1(ReadAddr[1]), .A2(n809), .ZN(n751) );
  INVD1 U552 ( .I(n767), .ZN(n771) );
  INVD1 U553 ( .I(n761), .ZN(n750) );
  ND2D1 U554 ( .A1(n353), .A2(n740), .ZN(N50) );
  NR3D0 U555 ( .A1(n741), .A2(n734), .A3(n733), .ZN(n735) );
  XNR2D1 U556 ( .A1(ReadAddr[3]), .A2(n814), .ZN(n733) );
  XNR2D1 U557 ( .A1(ReadAddr[2]), .A2(n816), .ZN(n734) );
  XNR2D1 U558 ( .A1(ReadAddr[2]), .A2(WriteAddr[2]), .ZN(n754) );
  NR2D1 U559 ( .A1(n744), .A2(n740), .ZN(N49) );
  NR2D1 U560 ( .A1(n238), .A2(n740), .ZN(N48) );
  NR2D1 U561 ( .A1(n2), .A2(n740), .ZN(N51) );
  NR2D1 U562 ( .A1(n294), .A2(n740), .ZN(N47) );
  INVD1 U563 ( .I(ReadReq), .ZN(n741) );
  INVD1 U564 ( .I(WriteReq), .ZN(n792) );
  INVD1 U565 ( .I(WriteAddr[1]), .ZN(n809) );
  OAI211D1 U566 ( .A1(n809), .A2(ReadAddr[1]), .B(n772), .C(n765), .ZN(n781)
         );
  AOI22D0 U567 ( .A1(n707), .A2(WriteAddr[3]), .B1(n704), .B2(WriteAddr[0]), 
        .ZN(n765) );
  ND2D1 U568 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .ZN(n730) );
  OAI21D1 U569 ( .A1(WriteAddr[1]), .A2(WriteAddr[0]), .B(n730), .ZN(n745) );
  AOI21D1 U570 ( .A1(n730), .A2(n702), .B(n732), .ZN(n760) );
  OAI211D1 U571 ( .A1(n705), .A2(WriteAddr[1]), .B(n771), .C(n768), .ZN(n782)
         );
  AOI22D0 U572 ( .A1(n703), .A2(ReadAddr[3]), .B1(n701), .B2(ReadAddr[0]), 
        .ZN(n768) );
  ND2D1 U573 ( .A1(n699), .A2(n803), .ZN(n784) );
  OAI22D0 U574 ( .A1(n817), .A2(n816), .B1(n706), .B2(n815), .ZN(n721) );
  OAI22D0 U575 ( .A1(n817), .A2(n814), .B1(n707), .B2(n815), .ZN(n719) );
  NR3D0 U576 ( .A1(n699), .A2(n698), .A3(n691), .ZN(n802) );
  ND2D1 U577 ( .A1(n706), .A2(WriteAddr[2]), .ZN(n772) );
  OAI22D0 U578 ( .A1(n807), .A2(n725), .B1(n806), .B2(n805), .ZN(n713) );
  AOI21D1 U579 ( .A1(n804), .A2(n803), .B(n802), .ZN(n805) );
  OAI22D0 U580 ( .A1(n699), .A2(n801), .B1(n691), .B2(n800), .ZN(n804) );
  OAI22D0 U581 ( .A1(n807), .A2(n724), .B1(n806), .B2(n788), .ZN(n711) );
  AOI31D0 U582 ( .A1(n787), .A2(n786), .A3(n691), .B(n785), .ZN(n788) );
  IOA21D1 U583 ( .A1(n803), .A2(n801), .B(n769), .ZN(n787) );
  OAI31D0 U584 ( .A1(n784), .A2(n691), .A3(n783), .B(n820), .ZN(n785) );
  OAI22D0 U585 ( .A1(n807), .A2(n723), .B1(n806), .B2(n758), .ZN(n710) );
  AOI22D0 U586 ( .A1(n757), .A2(n803), .B1(n756), .B2(n755), .ZN(n758) );
  AOI211D1 U587 ( .A1(n706), .A2(n752), .B(n818), .C(n770), .ZN(n756) );
  AOI221D0 U588 ( .A1(n767), .A2(n779), .B1(n754), .B2(ReadAddr[1]), .C(n753), 
        .ZN(n755) );
  AOI21D1 U589 ( .A1(n772), .A2(n771), .B(WriteAddr[1]), .ZN(n776) );
  INVD1 U590 ( .I(n699), .ZN(n786) );
  NR2D1 U591 ( .A1(WriteAddr[2]), .A2(n706), .ZN(n767) );
  OAI21D1 U592 ( .A1(n740), .A2(n739), .B(n738), .ZN(n709) );
  ND4D1 U593 ( .A1(n737), .A2(n739), .A3(n736), .A4(n735), .ZN(n738) );
  XNR2D1 U594 ( .A1(ReadAddr[0]), .A2(OldReadAr[0]), .ZN(n737) );
  XNR2D1 U595 ( .A1(ReadAddr[1]), .A2(OldReadAr[1]), .ZN(n736) );
  OAI21D1 U596 ( .A1(n699), .A2(n749), .B(n691), .ZN(n757) );
  NR4D0 U597 ( .A1(n750), .A2(n748), .A3(n763), .A4(n747), .ZN(n749) );
  XNR2D1 U598 ( .A1(WriteAddr[2]), .A2(n744), .ZN(n748) );
  XNR2D1 U599 ( .A1(WriteAddr[3]), .A2(n746), .ZN(n747) );
  OAI21D1 U600 ( .A1(n799), .A2(n808), .B(n798), .ZN(n712) );
  ND4D1 U601 ( .A1(n797), .A2(n808), .A3(n796), .A4(n795), .ZN(n798) );
  XNR2D1 U602 ( .A1(WriteAddr[0]), .A2(OldWriteAr[0]), .ZN(n797) );
  XNR2D1 U603 ( .A1(WriteAddr[2]), .A2(OldWriteAr[2]), .ZN(n796) );
  ND4D1 U604 ( .A1(n764), .A2(n763), .A3(n762), .A4(n761), .ZN(n801) );
  XNR2D1 U605 ( .A1(n759), .A2(n707), .ZN(n764) );
  XNR2D1 U606 ( .A1(ReadAddr[2]), .A2(n760), .ZN(n762) );
  NR2D1 U607 ( .A1(n730), .A2(n702), .ZN(n732) );
  NR2D1 U608 ( .A1(n809), .A2(n702), .ZN(n780) );
  XNR2D1 U609 ( .A1(ReadAddr[3]), .A2(n703), .ZN(n752) );
  XNR2D1 U610 ( .A1(WriteAddr[0]), .A2(n704), .ZN(n761) );
  NR2D1 U611 ( .A1(n704), .A2(n705), .ZN(n728) );
  XNR2D1 U612 ( .A1(n745), .A2(n705), .ZN(n763) );
  BUFFD1 U613 ( .I(n700), .Z(n691) );
  ND2D1 U614 ( .A1(ReadCmd), .A2(n353), .ZN(n740) );
  ND2D1 U615 ( .A1(WriteCmd), .A2(n813), .ZN(n799) );
  OAI32D1 U616 ( .A1(n820), .A2(WriteReq), .A3(n695), .B1(n819), .B2(n726), 
        .ZN(n722) );
  AOI21D1 U617 ( .A1(n818), .A2(n820), .B(n695), .ZN(n819) );
  OAI22D0 U618 ( .A1(n705), .A2(n813), .B1(n745), .B2(n799), .ZN(N68) );
  OAI22D0 U619 ( .A1(n458), .A2(n813), .B1(n759), .B2(n799), .ZN(N70) );
  OAI22D0 U620 ( .A1(n706), .A2(n813), .B1(n731), .B2(n799), .ZN(N69) );
  INVD1 U621 ( .I(n760), .ZN(n731) );
  OAI22D0 U622 ( .A1(n704), .A2(n813), .B1(WriteAddr[0]), .B2(n799), .ZN(N67)
         );
  ND3D1 U623 ( .A1(n691), .A2(n786), .A3(n698), .ZN(n818) );
  NR3D0 U624 ( .A1(n794), .A2(n793), .A3(n792), .ZN(n795) );
  XNR2D1 U625 ( .A1(n703), .A2(OldWriteAr[3]), .ZN(n793) );
  XNR2D1 U626 ( .A1(n809), .A2(OldWriteAr[1]), .ZN(n794) );
  OAI21D1 U627 ( .A1(n781), .A2(n782), .B(n698), .ZN(n769) );
  OAI31D0 U628 ( .A1(n813), .A2(n696), .A3(ReadReq), .B(n812), .ZN(n718) );
  OAI21D1 U629 ( .A1(n811), .A2(n696), .B(FullFIFO), .ZN(n812) );
  ND2D1 U630 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
endmodule


module DPMem1kx32_AWid4_DWid32_1 ( Dready, ParityErr, DataO, DataI, AddrR, 
        AddrW, ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [3:0] AddrR;
  input [3:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N9, N44, N45, N46, N47, ClockR, ClockW, Dreadyr, \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N84, N133, N166, N199, N232, N265, N298, N331, N364, N397,
         N430, N463, N496, N529, N562, N595, N628, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];

  OR2D1 U3 ( .A1(n486), .A2(Dreadyr), .Z(n591) );
  XNR4D1 U13 ( .A1(n234), .A2(n233), .A3(n236), .A4(n235), .ZN(n617) );
  XOR4D1 U14 ( .A1(n238), .A2(n237), .A3(n240), .A4(n239), .Z(n618) );
  XOR4D1 U15 ( .A1(n230), .A2(n229), .A3(n232), .A4(n231), .Z(n621) );
  XOR4D1 U16 ( .A1(n223), .A2(n222), .A3(n225), .A4(n224), .Z(n624) );
  XNR4D1 U17 ( .A1(n216), .A2(n215), .A3(n218), .A4(n217), .ZN(n627) );
  XOR4D1 U21 ( .A1(n612), .A2(N71), .A3(n611), .A4(N74), .Z(n613) );
  XNR4D1 U22 ( .A1(N68), .A2(N67), .A3(N70), .A4(N69), .ZN(n611) );
  XNR4D1 U27 ( .A1(N50), .A2(N49), .A3(N52), .A4(N51), .ZN(n605) );
  XOR4D1 U28 ( .A1(N54), .A2(N53), .A3(N56), .A4(N55), .Z(n606) );
  XNR4D1 U29 ( .A1(N61), .A2(N60), .A3(N63), .A4(N62), .ZN(n609) );
  XNR4D1 U30 ( .A1(N79), .A2(N77), .A3(N81), .A4(N80), .ZN(n615) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(N84), .E(n251), .CP(n379), .CDN(n540), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n240), .E(n251), .CP(n379), .CDN(n539), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n239), .E(n251), .CP(n379), .CDN(n539), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n238), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n233), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n232), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n231), .E(n252), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n230), .E(n252), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n229), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n228), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n227), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n226), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n225), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n224), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n223), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n222), .E(n252), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n221), .E(n253), .CP(n381), .CDN(n538), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n220), .E(n253), .CP(n382), .CDN(n538), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n219), .E(n253), .CP(n382), .CDN(n538), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n218), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n217), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n216), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n215), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n214), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n213), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n212), .E(n253), .CP(n382), .CDN(n537), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n211), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n210), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n209), .E(n254), .CP(n383), .CDN(n537), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(N84), .E(n259), .CP(n383), .CDN(n537), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n240), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n239), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n238), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n233), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n232), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n231), .E(n260), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n230), .E(n260), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n229), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n228), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n227), .E(n260), .CP(n384), .CDN(n535), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n226), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n225), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n224), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n223), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n222), .E(n260), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n221), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n220), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n219), .E(n261), .CP(n385), .CDN(n535), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n218), .E(n261), .CP(n385), .CDN(n534), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n217), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n216), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n215), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n214), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n213), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n212), .E(n261), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n211), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n210), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n209), .E(n262), .CP(n386), .CDN(n534), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(N84), .E(n283), .CP(n394), .CDN(n528), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n240), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n239), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n238), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n233), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n232), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n231), .E(n284), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n230), .E(n284), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n229), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n228), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n227), .E(n284), .CP(n395), .CDN(n526), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n226), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n225), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n224), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n223), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n222), .E(n284), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n221), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n220), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n219), .E(n285), .CP(n396), .CDN(n526), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n218), .E(n285), .CP(n396), .CDN(n525), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n217), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n216), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n215), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n214), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n213), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n212), .E(n285), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n211), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n210), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n209), .E(n286), .CP(n397), .CDN(n525), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(N84), .E(n291), .CP(n398), .CDN(n525), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n240), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n239), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n238), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n233), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n232), .E(n291), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n231), .E(n292), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n230), .E(n292), .CP(n399), .CDN(n524), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n229), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n228), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n227), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n226), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n225), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n224), .E(n292), .CP(n399), .CDN(n523), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n223), .E(n292), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n222), .E(n292), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n221), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n220), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n219), .E(n293), .CP(n400), .CDN(n523), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n218), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n217), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n216), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n215), .E(n293), .CP(n400), .CDN(n522), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n214), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n213), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n212), .E(n293), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n211), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n210), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n209), .E(n294), .CP(n401), .CDN(n522), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(N84), .E(n315), .CP(n409), .CDN(n516), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n240), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n239), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n238), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n233), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n232), .E(n315), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n231), .E(n316), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n230), .E(n316), .CP(n410), .CDN(n515), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n229), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n228), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n227), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n226), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n225), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n224), .E(n316), .CP(n410), .CDN(n514), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n223), .E(n316), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n222), .E(n316), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n221), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n220), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n219), .E(n317), .CP(n411), .CDN(n514), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n218), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n217), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n216), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n215), .E(n317), .CP(n411), .CDN(n513), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n214), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n213), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n212), .E(n317), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n211), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n210), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n209), .E(n318), .CP(n412), .CDN(n513), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(N84), .E(n323), .CP(n412), .CDN(n513), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n240), .E(n323), .CP(n412), .CDN(n512), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n239), .E(n323), .CP(n412), .CDN(n512), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n238), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n233), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n232), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n231), .E(n324), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n230), .E(n324), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n229), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n228), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n227), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n226), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n225), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n224), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n223), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n222), .E(n324), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n221), .E(n325), .CP(n414), .CDN(n511), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n220), .E(n325), .CP(n415), .CDN(n511), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n219), .E(n325), .CP(n415), .CDN(n511), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n218), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n217), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n216), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n215), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n214), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n213), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n212), .E(n325), .CP(n415), .CDN(n510), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n211), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n210), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n209), .E(n326), .CP(n416), .CDN(n510), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(N84), .E(n347), .CP(n423), .CDN(n504), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n240), .E(n347), .CP(n423), .CDN(n503), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n239), .E(n347), .CP(n423), .CDN(n503), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n238), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n233), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n232), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n231), .E(n348), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n230), .E(n348), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n229), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n228), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n227), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n226), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n225), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n224), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n223), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n222), .E(n348), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n221), .E(n349), .CP(n425), .CDN(n502), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n220), .E(n349), .CP(n426), .CDN(n502), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n219), .E(n349), .CP(n426), .CDN(n502), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n218), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n217), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n216), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n215), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n214), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n213), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n212), .E(n349), .CP(n426), .CDN(n501), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n211), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n210), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n209), .E(n350), .CP(n427), .CDN(n501), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N84), .E(n355), .CP(n427), .CDN(n501), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n240), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n239), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n238), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n233), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n232), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n231), .E(n356), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n230), .E(n356), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n229), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n228), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n227), .E(n356), .CP(n428), .CDN(n499), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n226), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n225), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n224), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n223), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n222), .E(n356), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n221), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n220), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n219), .E(n357), .CP(n429), .CDN(n499), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n218), .E(n357), .CP(n429), .CDN(n498), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n217), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n216), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n215), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n214), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n213), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n212), .E(n357), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n211), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n210), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n209), .E(n358), .CP(n430), .CDN(n498), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(N84), .E(n243), .CP(n376), .CDN(n543), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n240), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n239), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n238), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n233), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n232), .E(n243), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n231), .E(n244), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n230), .E(n244), .CP(n377), .CDN(n542), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n229), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n228), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n227), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n226), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n225), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n224), .E(n244), .CP(n377), .CDN(n541), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n223), .E(n244), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n222), .E(n244), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n221), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n220), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n219), .E(n245), .CP(n378), .CDN(n541), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n218), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n217), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n216), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n215), .E(n245), .CP(n378), .CDN(n540), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n214), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n213), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n212), .E(n245), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n211), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n210), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n209), .E(n246), .CP(n379), .CDN(n540), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(N84), .E(n267), .CP(n387), .CDN(n534), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n240), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n239), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n238), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n233), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n232), .E(n267), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n231), .E(n268), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n230), .E(n268), .CP(n388), .CDN(n533), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n229), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n228), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n227), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n226), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n225), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n224), .E(n268), .CP(n388), .CDN(n532), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n223), .E(n268), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n222), .E(n268), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n221), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n220), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n219), .E(n269), .CP(n389), .CDN(n532), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n218), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n217), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n216), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n215), .E(n269), .CP(n389), .CDN(n531), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n214), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n213), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n212), .E(n269), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n211), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n210), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n209), .E(n270), .CP(n390), .CDN(n531), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(N84), .E(n275), .CP(n390), .CDN(n531), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n240), .E(n275), .CP(n390), .CDN(n530), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n239), .E(n275), .CP(n390), .CDN(n530), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n238), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n233), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n232), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n231), .E(n276), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n230), .E(n276), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n229), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n228), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n227), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n226), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n225), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n224), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n223), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n222), .E(n276), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n221), .E(n277), .CP(n392), .CDN(n529), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n220), .E(n277), .CP(n393), .CDN(n529), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n219), .E(n277), .CP(n393), .CDN(n529), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n218), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n217), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n216), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n215), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n214), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n213), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n212), .E(n277), .CP(n393), .CDN(n528), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n211), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n210), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n209), .E(n278), .CP(n394), .CDN(n528), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(N84), .E(n299), .CP(n401), .CDN(n522), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n240), .E(n299), .CP(n401), .CDN(n521), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n239), .E(n299), .CP(n401), .CDN(n521), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n238), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n233), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n232), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n231), .E(n300), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n230), .E(n300), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n229), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n228), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n227), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n226), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n225), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n224), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n223), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n222), .E(n300), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n221), .E(n301), .CP(n403), .CDN(n520), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n220), .E(n301), .CP(n404), .CDN(n520), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n219), .E(n301), .CP(n404), .CDN(n520), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n218), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n217), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n216), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n215), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n214), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n213), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n212), .E(n301), .CP(n404), .CDN(n519), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n211), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n210), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n209), .E(n302), .CP(n405), .CDN(n519), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(N84), .E(n307), .CP(n405), .CDN(n519), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n240), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n239), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n238), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n233), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n232), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n231), .E(n308), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n230), .E(n308), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n229), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n228), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n227), .E(n308), .CP(n406), .CDN(n517), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n226), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n225), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n224), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n223), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n222), .E(n308), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n221), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n220), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n219), .E(n309), .CP(n407), .CDN(n517), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n218), .E(n309), .CP(n407), .CDN(n516), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n217), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n216), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n215), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n214), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n213), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n212), .E(n309), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n211), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n210), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n209), .E(n310), .CP(n408), .CDN(n516), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(N84), .E(n331), .CP(n416), .CDN(n510), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n240), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n239), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n238), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n233), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n232), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n231), .E(n332), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n230), .E(n332), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n229), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n228), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n227), .E(n332), .CP(n417), .CDN(n508), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n226), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n225), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n224), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n223), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n222), .E(n332), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n221), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n220), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n219), .E(n333), .CP(n418), .CDN(n508), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n218), .E(n333), .CP(n418), .CDN(n507), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n217), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n216), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n215), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n214), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n213), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n212), .E(n333), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n211), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n210), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n209), .E(n334), .CP(n419), .CDN(n507), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(N84), .E(n339), .CP(n420), .CDN(n507), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n240), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n239), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n238), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n233), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n232), .E(n339), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n231), .E(n340), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n230), .E(n340), .CP(n421), .CDN(n506), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n229), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n228), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n227), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n226), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n225), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n224), .E(n340), .CP(n421), .CDN(n505), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n223), .E(n340), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n222), .E(n340), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n221), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n220), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n219), .E(n341), .CP(n422), .CDN(n505), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n218), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n217), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n216), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n215), .E(n341), .CP(n422), .CDN(n504), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n214), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n213), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n212), .E(n341), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n211), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n210), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n209), .E(n342), .CP(n423), .CDN(n504), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N84), .E(n363), .CP(n431), .CDN(n498), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n240), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n239), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n238), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n233), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n232), .E(n363), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n231), .E(n364), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n230), .E(n364), .CP(n432), .CDN(n497), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n229), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n228), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n227), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n226), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n225), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n224), .E(n364), .CP(n432), .CDN(n496), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n223), .E(n364), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n222), .E(n364), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n221), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n220), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n219), .E(n365), .CP(n433), .CDN(n496), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n218), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n217), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n216), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n215), .E(n365), .CP(n433), .CDN(n495), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n214), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n213), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n212), .E(n365), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n211), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n210), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n209), .E(n366), .CP(n434), .CDN(n495), 
        .Q(\Storage[0][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n591), .CP(n480), .CDN(n495), .Q(Dreadyr) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n237), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n236), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n235), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n234), .E(n251), .CP(n380), .CDN(n539), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n237), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n236), .E(n259), .CP(n383), .CDN(n536), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n235), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n234), .E(n259), .CP(n384), .CDN(n536), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n237), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n236), .E(n283), .CP(n394), .CDN(n527), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n235), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n234), .E(n283), .CP(n395), .CDN(n527), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n237), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n236), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n235), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n234), .E(n291), .CP(n398), .CDN(n524), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n237), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n236), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n235), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n234), .E(n315), .CP(n409), .CDN(n515), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n237), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n236), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n235), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n234), .E(n323), .CP(n413), .CDN(n512), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n237), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n236), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n235), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n234), .E(n347), .CP(n424), .CDN(n503), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n237), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n236), .E(n355), .CP(n427), .CDN(n500), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n235), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n234), .E(n355), .CP(n428), .CDN(n500), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n237), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n236), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n235), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n234), .E(n243), .CP(n376), .CDN(n542), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n237), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n236), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n235), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n234), .E(n267), .CP(n387), .CDN(n533), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n237), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n236), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n235), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n234), .E(n275), .CP(n391), .CDN(n530), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n237), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n236), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n235), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n234), .E(n299), .CP(n402), .CDN(n521), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n237), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n236), .E(n307), .CP(n405), .CDN(n518), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n235), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n234), .E(n307), .CP(n406), .CDN(n518), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n237), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n236), .E(n331), .CP(n416), .CDN(n509), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n235), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n234), .E(n331), .CP(n417), .CDN(n509), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n237), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n236), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n235), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n234), .E(n339), .CP(n420), .CDN(n506), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n237), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n236), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n235), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n234), .E(n363), .CP(n431), .CDN(n497), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \DataOr_reg[31]  ( .D(N50), .E(n483), .CP(n477), .CDN(n546), .Q(
        DataOr[31]) );
  EDFCNQD1 \DataOr_reg[30]  ( .D(N51), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[30]) );
  EDFCNQD1 \DataOr_reg[29]  ( .D(N52), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[29]) );
  EDFCNQD1 \DataOr_reg[28]  ( .D(N53), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[28]) );
  EDFCNQD1 \DataOr_reg[27]  ( .D(N54), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[27]) );
  EDFCNQD1 \DataOr_reg[26]  ( .D(N55), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[26]) );
  EDFCNQD1 \DataOr_reg[25]  ( .D(N56), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[25]) );
  EDFCNQD1 \DataOr_reg[24]  ( .D(N57), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[24]) );
  EDFCNQD1 \DataOr_reg[23]  ( .D(N58), .E(n483), .CP(n477), .CDN(n545), .Q(
        DataOr[23]) );
  EDFCNQD1 \DataOr_reg[22]  ( .D(N59), .E(n483), .CP(n478), .CDN(n545), .Q(
        DataOr[22]) );
  EDFCNQD1 \DataOr_reg[21]  ( .D(N60), .E(n484), .CP(n478), .CDN(n545), .Q(
        DataOr[21]) );
  EDFCNQD1 \DataOr_reg[20]  ( .D(N61), .E(n484), .CP(n478), .CDN(n545), .Q(
        DataOr[20]) );
  EDFCNQD1 \DataOr_reg[19]  ( .D(N62), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[19]) );
  EDFCNQD1 \DataOr_reg[18]  ( .D(N63), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[18]) );
  EDFCNQD1 \DataOr_reg[17]  ( .D(N64), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[17]) );
  EDFCNQD1 \DataOr_reg[16]  ( .D(N65), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[16]) );
  EDFCNQD1 \DataOr_reg[15]  ( .D(N66), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[15]) );
  EDFCNQD1 \DataOr_reg[14]  ( .D(N67), .E(n484), .CP(n478), .CDN(n544), .Q(
        DataOr[14]) );
  EDFCNQD1 \DataOr_reg[13]  ( .D(N68), .E(n484), .CP(n479), .CDN(n544), .Q(
        DataOr[13]) );
  EDFCNQD1 \DataOr_reg[12]  ( .D(N69), .E(n484), .CP(n479), .CDN(n544), .Q(
        DataOr[12]) );
  EDFCNQD1 \DataOr_reg[11]  ( .D(N70), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[11]) );
  EDFCNQD1 \DataOr_reg[10]  ( .D(N71), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[10]) );
  EDFCNQD1 \DataOr_reg[9]  ( .D(N72), .E(n485), .CP(n479), .CDN(n544), .Q(
        DataOr[9]) );
  EDFCNQD1 \DataOr_reg[8]  ( .D(N73), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[8]) );
  EDFCNQD1 \DataOr_reg[7]  ( .D(N74), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[7]) );
  EDFCNQD1 \DataOr_reg[6]  ( .D(N75), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[6]) );
  EDFCNQD1 \DataOr_reg[5]  ( .D(N76), .E(n485), .CP(n479), .CDN(n543), .Q(
        DataOr[5]) );
  EDFCNQD1 \DataOr_reg[4]  ( .D(N77), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[4]) );
  EDFCNQD1 \DataOr_reg[3]  ( .D(N78), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[3]) );
  EDFCNQD1 \DataOr_reg[2]  ( .D(N79), .E(n485), .CP(n480), .CDN(n543), .Q(
        DataOr[2]) );
  EDFCNQD1 \DataOr_reg[1]  ( .D(N80), .E(n486), .CP(n480), .CDN(n543), .Q(
        DataOr[1]) );
  EDFCNQD1 \DataOr_reg[0]  ( .D(N81), .E(n486), .CP(n480), .CDN(n543), .Q(
        DataOr[0]) );
  EDFCNQD1 Parityr_reg ( .D(N82), .E(n486), .CP(n480), .CDN(n543), .Q(
        ParityErr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  CKAN2D0 U4 ( .A1(Dreadyr), .A2(ChipEna), .Z(Dready) );
  INVD1 U5 ( .I(n494), .ZN(n171) );
  INVD1 U6 ( .I(n493), .ZN(n175) );
  BUFFD1 U7 ( .I(n569), .Z(n501) );
  BUFFD1 U8 ( .I(n569), .Z(n502) );
  BUFFD1 U9 ( .I(n568), .Z(n503) );
  BUFFD1 U10 ( .I(n568), .Z(n504) );
  BUFFD1 U11 ( .I(n567), .Z(n505) );
  BUFFD1 U12 ( .I(n567), .Z(n506) );
  BUFFD1 U18 ( .I(n566), .Z(n507) );
  BUFFD1 U19 ( .I(n566), .Z(n508) );
  BUFFD1 U20 ( .I(n565), .Z(n509) );
  BUFFD1 U23 ( .I(n565), .Z(n510) );
  BUFFD1 U24 ( .I(n564), .Z(n511) );
  BUFFD1 U25 ( .I(n564), .Z(n512) );
  BUFFD1 U26 ( .I(n563), .Z(n513) );
  BUFFD1 U31 ( .I(n563), .Z(n514) );
  BUFFD1 U32 ( .I(n562), .Z(n515) );
  BUFFD1 U33 ( .I(n562), .Z(n516) );
  BUFFD1 U34 ( .I(n561), .Z(n517) );
  BUFFD1 U35 ( .I(n561), .Z(n518) );
  BUFFD1 U36 ( .I(n560), .Z(n519) );
  BUFFD1 U37 ( .I(n560), .Z(n520) );
  BUFFD1 U38 ( .I(n559), .Z(n521) );
  BUFFD1 U39 ( .I(n559), .Z(n522) );
  BUFFD1 U40 ( .I(n558), .Z(n523) );
  BUFFD1 U41 ( .I(n558), .Z(n524) );
  BUFFD1 U42 ( .I(n557), .Z(n525) );
  BUFFD1 U43 ( .I(n557), .Z(n526) );
  BUFFD1 U44 ( .I(n556), .Z(n527) );
  BUFFD1 U45 ( .I(n556), .Z(n528) );
  BUFFD1 U46 ( .I(n555), .Z(n529) );
  BUFFD1 U47 ( .I(n555), .Z(n530) );
  BUFFD1 U48 ( .I(n554), .Z(n531) );
  BUFFD1 U49 ( .I(n554), .Z(n532) );
  BUFFD1 U50 ( .I(n553), .Z(n533) );
  BUFFD1 U51 ( .I(n553), .Z(n534) );
  BUFFD1 U52 ( .I(n552), .Z(n535) );
  BUFFD1 U53 ( .I(n552), .Z(n536) );
  BUFFD1 U54 ( .I(n551), .Z(n537) );
  BUFFD1 U55 ( .I(n551), .Z(n538) );
  BUFFD1 U56 ( .I(n550), .Z(n539) );
  BUFFD1 U57 ( .I(n550), .Z(n540) );
  BUFFD1 U58 ( .I(n549), .Z(n541) );
  BUFFD1 U59 ( .I(n549), .Z(n542) );
  BUFFD1 U60 ( .I(n548), .Z(n543) );
  BUFFD1 U61 ( .I(n548), .Z(n544) );
  BUFFD1 U62 ( .I(n547), .Z(n545) );
  BUFFD1 U63 ( .I(n547), .Z(n546) );
  BUFFD1 U64 ( .I(n572), .Z(n495) );
  BUFFD1 U65 ( .I(n572), .Z(n496) );
  BUFFD1 U66 ( .I(n571), .Z(n497) );
  BUFFD1 U67 ( .I(n571), .Z(n498) );
  BUFFD1 U68 ( .I(n570), .Z(n499) );
  BUFFD1 U69 ( .I(n570), .Z(n500) );
  BUFFD1 U70 ( .I(n574), .Z(n569) );
  BUFFD1 U71 ( .I(n574), .Z(n568) );
  BUFFD1 U72 ( .I(n574), .Z(n567) );
  BUFFD1 U73 ( .I(n575), .Z(n566) );
  BUFFD1 U74 ( .I(n575), .Z(n565) );
  BUFFD1 U75 ( .I(n575), .Z(n564) );
  BUFFD1 U76 ( .I(n576), .Z(n563) );
  BUFFD1 U77 ( .I(n576), .Z(n562) );
  BUFFD1 U78 ( .I(n576), .Z(n561) );
  BUFFD1 U79 ( .I(n577), .Z(n560) );
  BUFFD1 U80 ( .I(n577), .Z(n559) );
  BUFFD1 U81 ( .I(n577), .Z(n558) );
  BUFFD1 U82 ( .I(n578), .Z(n557) );
  BUFFD1 U83 ( .I(n578), .Z(n556) );
  BUFFD1 U84 ( .I(n578), .Z(n555) );
  BUFFD1 U85 ( .I(n579), .Z(n554) );
  BUFFD1 U86 ( .I(n579), .Z(n553) );
  BUFFD1 U87 ( .I(n579), .Z(n552) );
  BUFFD1 U88 ( .I(n580), .Z(n551) );
  BUFFD1 U89 ( .I(n580), .Z(n550) );
  BUFFD1 U90 ( .I(n580), .Z(n549) );
  BUFFD1 U91 ( .I(n581), .Z(n548) );
  BUFFD1 U92 ( .I(n581), .Z(n547) );
  BUFFD1 U93 ( .I(n573), .Z(n571) );
  BUFFD1 U94 ( .I(n573), .Z(n570) );
  BUFFD1 U95 ( .I(n573), .Z(n572) );
  BUFFD1 U96 ( .I(n585), .Z(n574) );
  BUFFD1 U97 ( .I(n585), .Z(n575) );
  BUFFD1 U98 ( .I(n584), .Z(n576) );
  BUFFD1 U99 ( .I(n584), .Z(n577) );
  BUFFD1 U100 ( .I(n583), .Z(n578) );
  BUFFD1 U101 ( .I(n583), .Z(n579) );
  BUFFD1 U102 ( .I(n582), .Z(n580) );
  BUFFD1 U103 ( .I(n582), .Z(n581) );
  BUFFD1 U104 ( .I(n587), .Z(n585) );
  BUFFD1 U105 ( .I(n587), .Z(n584) );
  BUFFD1 U106 ( .I(n588), .Z(n583) );
  BUFFD1 U107 ( .I(n588), .Z(n582) );
  BUFFD1 U108 ( .I(n586), .Z(n573) );
  BUFFD1 U109 ( .I(n587), .Z(n586) );
  INVD1 U110 ( .I(n589), .ZN(n587) );
  INVD1 U111 ( .I(n589), .ZN(n588) );
  BUFFD1 U112 ( .I(n435), .Z(n433) );
  BUFFD1 U113 ( .I(n436), .Z(n432) );
  BUFFD1 U114 ( .I(n436), .Z(n431) );
  BUFFD1 U115 ( .I(n437), .Z(n430) );
  BUFFD1 U116 ( .I(n437), .Z(n429) );
  BUFFD1 U117 ( .I(n438), .Z(n428) );
  BUFFD1 U118 ( .I(n438), .Z(n427) );
  BUFFD1 U119 ( .I(n439), .Z(n426) );
  BUFFD1 U120 ( .I(n439), .Z(n425) );
  BUFFD1 U121 ( .I(n440), .Z(n424) );
  BUFFD1 U122 ( .I(n440), .Z(n423) );
  BUFFD1 U123 ( .I(n441), .Z(n422) );
  BUFFD1 U124 ( .I(n441), .Z(n421) );
  BUFFD1 U125 ( .I(n442), .Z(n420) );
  BUFFD1 U126 ( .I(n442), .Z(n419) );
  BUFFD1 U127 ( .I(n443), .Z(n418) );
  BUFFD1 U128 ( .I(n443), .Z(n417) );
  BUFFD1 U129 ( .I(n444), .Z(n416) );
  BUFFD1 U130 ( .I(n444), .Z(n415) );
  BUFFD1 U131 ( .I(n445), .Z(n414) );
  BUFFD1 U132 ( .I(n445), .Z(n413) );
  BUFFD1 U133 ( .I(n446), .Z(n412) );
  BUFFD1 U134 ( .I(n446), .Z(n411) );
  BUFFD1 U135 ( .I(n447), .Z(n410) );
  BUFFD1 U136 ( .I(n447), .Z(n409) );
  BUFFD1 U137 ( .I(n448), .Z(n408) );
  BUFFD1 U138 ( .I(n448), .Z(n407) );
  BUFFD1 U139 ( .I(n449), .Z(n406) );
  BUFFD1 U140 ( .I(n449), .Z(n405) );
  BUFFD1 U141 ( .I(n450), .Z(n404) );
  BUFFD1 U142 ( .I(n450), .Z(n403) );
  BUFFD1 U143 ( .I(n451), .Z(n402) );
  BUFFD1 U144 ( .I(n451), .Z(n401) );
  BUFFD1 U145 ( .I(n452), .Z(n400) );
  BUFFD1 U146 ( .I(n452), .Z(n399) );
  BUFFD1 U147 ( .I(n453), .Z(n398) );
  BUFFD1 U148 ( .I(n453), .Z(n397) );
  BUFFD1 U149 ( .I(n454), .Z(n396) );
  BUFFD1 U150 ( .I(n454), .Z(n395) );
  BUFFD1 U151 ( .I(n455), .Z(n394) );
  BUFFD1 U152 ( .I(n455), .Z(n393) );
  BUFFD1 U153 ( .I(n456), .Z(n392) );
  BUFFD1 U154 ( .I(n456), .Z(n391) );
  BUFFD1 U155 ( .I(n457), .Z(n390) );
  BUFFD1 U156 ( .I(n457), .Z(n389) );
  BUFFD1 U157 ( .I(n458), .Z(n388) );
  BUFFD1 U158 ( .I(n458), .Z(n387) );
  BUFFD1 U159 ( .I(n459), .Z(n386) );
  BUFFD1 U160 ( .I(n459), .Z(n385) );
  BUFFD1 U161 ( .I(n460), .Z(n384) );
  BUFFD1 U162 ( .I(n460), .Z(n383) );
  BUFFD1 U163 ( .I(n461), .Z(n382) );
  BUFFD1 U164 ( .I(n461), .Z(n381) );
  BUFFD1 U165 ( .I(n462), .Z(n380) );
  BUFFD1 U166 ( .I(n462), .Z(n379) );
  BUFFD1 U167 ( .I(n463), .Z(n378) );
  BUFFD1 U168 ( .I(n463), .Z(n377) );
  BUFFD1 U169 ( .I(n435), .Z(n434) );
  INVD1 U170 ( .I(n590), .ZN(n589) );
  INVD1 U171 ( .I(Reset), .ZN(n590) );
  INVD1 U172 ( .I(n367), .ZN(n365) );
  INVD1 U173 ( .I(n368), .ZN(n364) );
  INVD1 U174 ( .I(n368), .ZN(n363) );
  INVD1 U175 ( .I(n303), .ZN(n301) );
  INVD1 U176 ( .I(n304), .ZN(n300) );
  INVD1 U177 ( .I(n304), .ZN(n299) );
  INVD1 U178 ( .I(n367), .ZN(n366) );
  INVD1 U179 ( .I(n303), .ZN(n302) );
  BUFFD1 U180 ( .I(n464), .Z(n376) );
  BUFFD1 U181 ( .I(n465), .Z(n464) );
  BUFFD1 U182 ( .I(n474), .Z(n435) );
  BUFFD1 U183 ( .I(n474), .Z(n436) );
  BUFFD1 U184 ( .I(n474), .Z(n437) );
  BUFFD1 U185 ( .I(n473), .Z(n438) );
  BUFFD1 U186 ( .I(n473), .Z(n439) );
  BUFFD1 U187 ( .I(n473), .Z(n440) );
  BUFFD1 U188 ( .I(n472), .Z(n441) );
  BUFFD1 U189 ( .I(n472), .Z(n442) );
  BUFFD1 U190 ( .I(n472), .Z(n443) );
  BUFFD1 U191 ( .I(n471), .Z(n444) );
  BUFFD1 U192 ( .I(n471), .Z(n445) );
  BUFFD1 U193 ( .I(n471), .Z(n446) );
  BUFFD1 U194 ( .I(n470), .Z(n447) );
  BUFFD1 U195 ( .I(n470), .Z(n448) );
  BUFFD1 U196 ( .I(n470), .Z(n449) );
  BUFFD1 U197 ( .I(n469), .Z(n450) );
  BUFFD1 U198 ( .I(n469), .Z(n451) );
  BUFFD1 U199 ( .I(n469), .Z(n452) );
  BUFFD1 U200 ( .I(n468), .Z(n453) );
  BUFFD1 U201 ( .I(n468), .Z(n454) );
  BUFFD1 U202 ( .I(n468), .Z(n455) );
  BUFFD1 U203 ( .I(n467), .Z(n456) );
  BUFFD1 U204 ( .I(n467), .Z(n457) );
  BUFFD1 U205 ( .I(n467), .Z(n458) );
  BUFFD1 U206 ( .I(n466), .Z(n459) );
  BUFFD1 U207 ( .I(n466), .Z(n460) );
  BUFFD1 U208 ( .I(n466), .Z(n461) );
  BUFFD1 U209 ( .I(n465), .Z(n462) );
  BUFFD1 U210 ( .I(n465), .Z(n463) );
  INVD1 U211 ( .I(n361), .ZN(n367) );
  INVD1 U212 ( .I(n361), .ZN(n368) );
  INVD1 U213 ( .I(n297), .ZN(n303) );
  INVD1 U214 ( .I(n297), .ZN(n304) );
  INVD1 U215 ( .I(n359), .ZN(n357) );
  INVD1 U216 ( .I(n360), .ZN(n356) );
  INVD1 U217 ( .I(n360), .ZN(n355) );
  INVD1 U218 ( .I(n351), .ZN(n349) );
  INVD1 U219 ( .I(n352), .ZN(n348) );
  INVD1 U220 ( .I(n352), .ZN(n347) );
  INVD1 U221 ( .I(n343), .ZN(n341) );
  INVD1 U222 ( .I(n344), .ZN(n340) );
  INVD1 U223 ( .I(n344), .ZN(n339) );
  INVD1 U224 ( .I(n335), .ZN(n333) );
  INVD1 U225 ( .I(n336), .ZN(n332) );
  INVD1 U226 ( .I(n336), .ZN(n331) );
  INVD1 U227 ( .I(n327), .ZN(n325) );
  INVD1 U228 ( .I(n328), .ZN(n324) );
  INVD1 U229 ( .I(n328), .ZN(n323) );
  INVD1 U230 ( .I(n319), .ZN(n317) );
  INVD1 U231 ( .I(n320), .ZN(n316) );
  INVD1 U232 ( .I(n320), .ZN(n315) );
  INVD1 U233 ( .I(n311), .ZN(n309) );
  INVD1 U234 ( .I(n312), .ZN(n308) );
  INVD1 U235 ( .I(n312), .ZN(n307) );
  INVD1 U236 ( .I(n295), .ZN(n293) );
  INVD1 U237 ( .I(n296), .ZN(n292) );
  INVD1 U238 ( .I(n296), .ZN(n291) );
  INVD1 U239 ( .I(n287), .ZN(n285) );
  INVD1 U240 ( .I(n288), .ZN(n284) );
  INVD1 U241 ( .I(n288), .ZN(n283) );
  INVD1 U242 ( .I(n279), .ZN(n277) );
  INVD1 U243 ( .I(n280), .ZN(n276) );
  INVD1 U244 ( .I(n280), .ZN(n275) );
  INVD1 U245 ( .I(n271), .ZN(n269) );
  INVD1 U246 ( .I(n272), .ZN(n268) );
  INVD1 U247 ( .I(n272), .ZN(n267) );
  INVD1 U248 ( .I(n263), .ZN(n261) );
  INVD1 U249 ( .I(n264), .ZN(n260) );
  INVD1 U250 ( .I(n264), .ZN(n259) );
  INVD1 U251 ( .I(n255), .ZN(n253) );
  INVD1 U252 ( .I(n256), .ZN(n252) );
  INVD1 U253 ( .I(n256), .ZN(n251) );
  INVD1 U254 ( .I(n247), .ZN(n245) );
  INVD1 U255 ( .I(n248), .ZN(n244) );
  INVD1 U256 ( .I(n248), .ZN(n243) );
  INVD1 U257 ( .I(n351), .ZN(n350) );
  INVD1 U258 ( .I(n343), .ZN(n342) );
  INVD1 U259 ( .I(n359), .ZN(n358) );
  INVD1 U260 ( .I(n335), .ZN(n334) );
  INVD1 U261 ( .I(n327), .ZN(n326) );
  INVD1 U262 ( .I(n319), .ZN(n318) );
  INVD1 U263 ( .I(n311), .ZN(n310) );
  INVD1 U264 ( .I(n295), .ZN(n294) );
  INVD1 U265 ( .I(n287), .ZN(n286) );
  INVD1 U266 ( .I(n279), .ZN(n278) );
  INVD1 U267 ( .I(n271), .ZN(n270) );
  INVD1 U268 ( .I(n263), .ZN(n262) );
  INVD1 U269 ( .I(n255), .ZN(n254) );
  INVD1 U270 ( .I(n247), .ZN(n246) );
  BUFFD1 U271 ( .I(n373), .Z(n474) );
  BUFFD1 U272 ( .I(n373), .Z(n473) );
  BUFFD1 U273 ( .I(n372), .Z(n472) );
  BUFFD1 U274 ( .I(n372), .Z(n471) );
  BUFFD1 U275 ( .I(n371), .Z(n470) );
  BUFFD1 U276 ( .I(n371), .Z(n469) );
  BUFFD1 U277 ( .I(n370), .Z(n468) );
  BUFFD1 U278 ( .I(n370), .Z(n467) );
  BUFFD1 U279 ( .I(n369), .Z(n466) );
  BUFFD1 U280 ( .I(n369), .Z(n465) );
  BUFFD1 U281 ( .I(n197), .Z(n198) );
  BUFFD1 U282 ( .I(n197), .Z(n199) );
  BUFFD1 U283 ( .I(n197), .Z(n200) );
  BUFFD1 U284 ( .I(n196), .Z(n201) );
  BUFFD1 U285 ( .I(n196), .Z(n202) );
  BUFFD1 U286 ( .I(n196), .Z(n203) );
  BUFFD1 U287 ( .I(n195), .Z(n204) );
  BUFFD1 U288 ( .I(n195), .Z(n205) );
  BUFFD1 U289 ( .I(n195), .Z(n206) );
  BUFFD1 U290 ( .I(n194), .Z(n207) );
  BUFFD1 U291 ( .I(n194), .Z(n208) );
  BUFFD1 U292 ( .I(n182), .Z(n183) );
  BUFFD1 U293 ( .I(n182), .Z(n184) );
  BUFFD1 U294 ( .I(n182), .Z(n185) );
  BUFFD1 U295 ( .I(n181), .Z(n186) );
  BUFFD1 U296 ( .I(n181), .Z(n187) );
  BUFFD1 U297 ( .I(n181), .Z(n188) );
  BUFFD1 U298 ( .I(n180), .Z(n189) );
  BUFFD1 U299 ( .I(n180), .Z(n190) );
  BUFFD1 U300 ( .I(n180), .Z(n191) );
  BUFFD1 U301 ( .I(n179), .Z(n192) );
  BUFFD1 U302 ( .I(n179), .Z(n193) );
  INVD1 U303 ( .I(n353), .ZN(n359) );
  INVD1 U304 ( .I(n353), .ZN(n360) );
  INVD1 U305 ( .I(n345), .ZN(n351) );
  INVD1 U306 ( .I(n345), .ZN(n352) );
  INVD1 U307 ( .I(n337), .ZN(n343) );
  INVD1 U308 ( .I(n337), .ZN(n344) );
  INVD1 U309 ( .I(n329), .ZN(n335) );
  INVD1 U310 ( .I(n329), .ZN(n336) );
  INVD1 U311 ( .I(n321), .ZN(n327) );
  INVD1 U312 ( .I(n321), .ZN(n328) );
  INVD1 U313 ( .I(n313), .ZN(n319) );
  INVD1 U314 ( .I(n313), .ZN(n320) );
  INVD1 U315 ( .I(n305), .ZN(n311) );
  INVD1 U316 ( .I(n305), .ZN(n312) );
  INVD1 U317 ( .I(n289), .ZN(n295) );
  INVD1 U318 ( .I(n289), .ZN(n296) );
  INVD1 U319 ( .I(n281), .ZN(n287) );
  INVD1 U320 ( .I(n281), .ZN(n288) );
  INVD1 U321 ( .I(n273), .ZN(n279) );
  INVD1 U322 ( .I(n273), .ZN(n280) );
  INVD1 U323 ( .I(n265), .ZN(n271) );
  INVD1 U324 ( .I(n265), .ZN(n272) );
  INVD1 U325 ( .I(n257), .ZN(n263) );
  INVD1 U326 ( .I(n257), .ZN(n264) );
  INVD1 U327 ( .I(n249), .ZN(n255) );
  INVD1 U328 ( .I(n249), .ZN(n256) );
  INVD1 U329 ( .I(n241), .ZN(n247) );
  INVD1 U330 ( .I(n241), .ZN(n248) );
  INVD1 U331 ( .I(n362), .ZN(n361) );
  INVD1 U332 ( .I(N133), .ZN(n362) );
  NR2D1 U333 ( .A1(n599), .A2(n595), .ZN(N133) );
  INVD1 U334 ( .I(n298), .ZN(n297) );
  INVD1 U335 ( .I(N397), .ZN(n298) );
  NR2D1 U336 ( .A1(n602), .A2(n599), .ZN(N397) );
  INVD1 U337 ( .I(n487), .ZN(n485) );
  INVD1 U338 ( .I(n488), .ZN(n484) );
  INVD1 U339 ( .I(n488), .ZN(n483) );
  INVD1 U340 ( .I(n487), .ZN(n486) );
  BUFFD1 U341 ( .I(n374), .Z(n373) );
  BUFFD1 U342 ( .I(n374), .Z(n372) );
  BUFFD1 U343 ( .I(n374), .Z(n371) );
  BUFFD1 U344 ( .I(n375), .Z(n370) );
  BUFFD1 U345 ( .I(n375), .Z(n369) );
  INVD1 U346 ( .I(n481), .ZN(n479) );
  INVD1 U347 ( .I(n482), .ZN(n478) );
  INVD1 U348 ( .I(n482), .ZN(n477) );
  INVD1 U349 ( .I(n481), .ZN(n480) );
  XOR3D1 U350 ( .A1(n211), .A2(n210), .A3(n628), .Z(N84) );
  XOR3D1 U351 ( .A1(n209), .A2(n627), .A3(n626), .Z(n628) );
  XOR3D1 U352 ( .A1(n214), .A2(n213), .A3(n625), .Z(n626) );
  XOR3D1 U353 ( .A1(n228), .A2(n227), .A3(n619), .Z(n620) );
  XOR3D1 U354 ( .A1(n618), .A2(n226), .A3(n617), .Z(n619) );
  XOR3D1 U355 ( .A1(n624), .A2(n212), .A3(n623), .Z(n625) );
  XOR3D1 U356 ( .A1(n221), .A2(n220), .A3(n622), .Z(n623) );
  XOR3D1 U357 ( .A1(n621), .A2(n219), .A3(n620), .Z(n622) );
  XOR3D1 U358 ( .A1(N66), .A2(N65), .A3(n610), .Z(n612) );
  XOR3D1 U359 ( .A1(N64), .A2(n609), .A3(n608), .Z(n610) );
  XOR3D1 U360 ( .A1(N59), .A2(N58), .A3(n607), .Z(n608) );
  XOR3D1 U361 ( .A1(n606), .A2(N57), .A3(n605), .Z(n607) );
  XOR3D1 U362 ( .A1(N78), .A2(N73), .A3(n616), .Z(N82) );
  XOR3D1 U363 ( .A1(N72), .A2(n615), .A3(n614), .Z(n616) );
  XOR3D1 U364 ( .A1(N76), .A2(N75), .A3(n613), .Z(n614) );
  BUFFD1 U365 ( .I(n491), .Z(n197) );
  BUFFD1 U366 ( .I(n492), .Z(n182) );
  BUFFD1 U367 ( .I(n491), .Z(n196) );
  BUFFD1 U368 ( .I(n492), .Z(n181) );
  BUFFD1 U369 ( .I(n491), .Z(n195) );
  BUFFD1 U370 ( .I(n492), .Z(n180) );
  INVD1 U371 ( .I(n171), .ZN(n173) );
  INVD1 U372 ( .I(n171), .ZN(n174) );
  BUFFD1 U373 ( .I(n491), .Z(n194) );
  BUFFD1 U374 ( .I(n492), .Z(n179) );
  INVD1 U375 ( .I(n171), .ZN(n172) );
  INVD1 U376 ( .I(n175), .ZN(n177) );
  INVD1 U377 ( .I(n175), .ZN(n178) );
  INVD1 U378 ( .I(n175), .ZN(n176) );
  ND2D1 U379 ( .A1(n592), .A2(n597), .ZN(n595) );
  ND2D1 U380 ( .A1(n594), .A2(n593), .ZN(n599) );
  ND2D1 U381 ( .A1(n598), .A2(n597), .ZN(n602) );
  INVD1 U382 ( .I(n346), .ZN(n345) );
  INVD1 U383 ( .I(N199), .ZN(n346) );
  NR2D1 U384 ( .A1(n600), .A2(n595), .ZN(N199) );
  INVD1 U385 ( .I(n338), .ZN(n337) );
  INVD1 U386 ( .I(N232), .ZN(n338) );
  NR2D1 U387 ( .A1(n600), .A2(n596), .ZN(N232) );
  INVD1 U388 ( .I(n330), .ZN(n329) );
  INVD1 U389 ( .I(N265), .ZN(n330) );
  NR2D1 U390 ( .A1(n601), .A2(n595), .ZN(N265) );
  INVD1 U391 ( .I(n322), .ZN(n321) );
  INVD1 U392 ( .I(N298), .ZN(n322) );
  NR2D1 U393 ( .A1(n601), .A2(n596), .ZN(N298) );
  INVD1 U394 ( .I(n314), .ZN(n313) );
  INVD1 U395 ( .I(N331), .ZN(n314) );
  NR2D1 U396 ( .A1(n603), .A2(n595), .ZN(N331) );
  INVD1 U397 ( .I(n306), .ZN(n305) );
  INVD1 U398 ( .I(N364), .ZN(n306) );
  NR2D1 U399 ( .A1(n603), .A2(n596), .ZN(N364) );
  INVD1 U400 ( .I(n250), .ZN(n249) );
  INVD1 U401 ( .I(N595), .ZN(n250) );
  NR2D1 U402 ( .A1(n603), .A2(n602), .ZN(N595) );
  INVD1 U403 ( .I(n354), .ZN(n353) );
  INVD1 U404 ( .I(N166), .ZN(n354) );
  NR2D1 U405 ( .A1(n599), .A2(n596), .ZN(N166) );
  INVD1 U406 ( .I(n290), .ZN(n289) );
  INVD1 U407 ( .I(N430), .ZN(n290) );
  NR2D1 U408 ( .A1(n604), .A2(n599), .ZN(N430) );
  INVD1 U409 ( .I(n282), .ZN(n281) );
  INVD1 U410 ( .I(N463), .ZN(n282) );
  NR2D1 U411 ( .A1(n602), .A2(n600), .ZN(N463) );
  INVD1 U412 ( .I(n274), .ZN(n273) );
  INVD1 U413 ( .I(N496), .ZN(n274) );
  NR2D1 U414 ( .A1(n604), .A2(n600), .ZN(N496) );
  INVD1 U415 ( .I(n266), .ZN(n265) );
  INVD1 U416 ( .I(N529), .ZN(n266) );
  NR2D1 U417 ( .A1(n602), .A2(n601), .ZN(N529) );
  INVD1 U418 ( .I(n258), .ZN(n257) );
  INVD1 U419 ( .I(N562), .ZN(n258) );
  NR2D1 U420 ( .A1(n604), .A2(n601), .ZN(N562) );
  INVD1 U421 ( .I(n242), .ZN(n241) );
  INVD1 U422 ( .I(N628), .ZN(n242) );
  NR2D1 U423 ( .A1(n604), .A2(n603), .ZN(N628) );
  INVD1 U424 ( .I(n489), .ZN(n487) );
  INVD1 U425 ( .I(n489), .ZN(n488) );
  INVD1 U426 ( .I(n475), .ZN(n482) );
  INVD1 U427 ( .I(n475), .ZN(n481) );
  BUFFD1 U428 ( .I(ClockW), .Z(n374) );
  BUFFD1 U429 ( .I(ClockW), .Z(n375) );
  BUFFD1 U430 ( .I(DataI[14]), .Z(n223) );
  BUFFD1 U431 ( .I(DataI[15]), .Z(n224) );
  BUFFD1 U432 ( .I(DataI[21]), .Z(n230) );
  BUFFD1 U433 ( .I(DataI[22]), .Z(n231) );
  BUFFD1 U434 ( .I(DataI[25]), .Z(n234) );
  BUFFD1 U435 ( .I(DataI[26]), .Z(n235) );
  BUFFD1 U436 ( .I(DataI[29]), .Z(n238) );
  BUFFD1 U437 ( .I(DataI[30]), .Z(n239) );
  BUFFD1 U438 ( .I(DataI[10]), .Z(n219) );
  BUFFD1 U439 ( .I(DataI[17]), .Z(n226) );
  BUFFD1 U440 ( .I(DataI[18]), .Z(n227) );
  BUFFD1 U441 ( .I(DataI[13]), .Z(n222) );
  BUFFD1 U442 ( .I(DataI[16]), .Z(n225) );
  BUFFD1 U443 ( .I(DataI[20]), .Z(n229) );
  BUFFD1 U444 ( .I(DataI[23]), .Z(n232) );
  BUFFD1 U445 ( .I(DataI[24]), .Z(n233) );
  BUFFD1 U446 ( .I(DataI[27]), .Z(n236) );
  BUFFD1 U447 ( .I(DataI[28]), .Z(n237) );
  BUFFD1 U448 ( .I(DataI[31]), .Z(n240) );
  BUFFD1 U449 ( .I(DataI[19]), .Z(n228) );
  BUFFD1 U450 ( .I(DataI[2]), .Z(n211) );
  BUFFD1 U451 ( .I(DataI[1]), .Z(n210) );
  BUFFD1 U452 ( .I(DataI[7]), .Z(n216) );
  BUFFD1 U453 ( .I(DataI[8]), .Z(n217) );
  BUFFD1 U454 ( .I(DataI[3]), .Z(n212) );
  BUFFD1 U455 ( .I(DataI[4]), .Z(n213) );
  BUFFD1 U456 ( .I(DataI[11]), .Z(n220) );
  BUFFD1 U457 ( .I(DataI[6]), .Z(n215) );
  BUFFD1 U458 ( .I(DataI[9]), .Z(n218) );
  BUFFD1 U459 ( .I(DataI[0]), .Z(n209) );
  BUFFD1 U460 ( .I(DataI[5]), .Z(n214) );
  BUFFD1 U461 ( .I(DataI[12]), .Z(n221) );
  MUX4D0 U462 ( .I0(n8), .I1(n6), .I2(n7), .I3(n5), .S0(n172), .S1(n176), .Z(
        N80) );
  MUX4D0 U463 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n198), .S1(n183), .Z(n7)
         );
  MUX4D0 U464 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n198), .S1(n183), .Z(n6)
         );
  MUX4D0 U465 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n198), .S1(n183), .Z(n8)
         );
  MUX4D0 U466 ( .I0(n12), .I1(n10), .I2(n11), .I3(n9), .S0(n172), .S1(n176), 
        .Z(N79) );
  MUX4D0 U467 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n198), .S1(n183), .Z(n11)
         );
  MUX4D0 U468 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n198), .S1(n183), .Z(n10) );
  MUX4D0 U469 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n198), .S1(n183), .Z(n12)
         );
  MUX4D0 U470 ( .I0(n32), .I1(n30), .I2(n31), .I3(n29), .S0(n172), .S1(n176), 
        .Z(N74) );
  MUX4D0 U471 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n200), .S1(n185), .Z(n31)
         );
  MUX4D0 U472 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n200), .S1(n185), .Z(n30) );
  MUX4D0 U473 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n200), .S1(n185), .Z(n32)
         );
  MUX4D0 U474 ( .I0(n52), .I1(n50), .I2(n51), .I3(n49), .S0(n173), .S1(n177), 
        .Z(N69) );
  MUX4D0 U475 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n202), .S1(n187), .Z(n51) );
  MUX4D0 U476 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n202), .S1(n187), .Z(
        n50) );
  MUX4D0 U477 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n202), .S1(n187), .Z(n52) );
  MUX4D0 U478 ( .I0(n56), .I1(n54), .I2(n55), .I3(n53), .S0(n173), .S1(n177), 
        .Z(N68) );
  MUX4D0 U479 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n202), .S1(n187), .Z(n55) );
  MUX4D0 U480 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n202), .S1(n187), .Z(
        n54) );
  MUX4D0 U481 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n202), .S1(n187), .Z(n56) );
  MUX4D0 U482 ( .I0(n118), .I1(n116), .I2(n117), .I3(n115), .S0(n173), .S1(
        n177), .Z(N62) );
  MUX4D0 U483 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n204), .S1(n189), .Z(
        n117) );
  MUX4D0 U484 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n204), .S1(n189), .Z(
        n116) );
  MUX4D0 U485 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n204), .S1(n189), .Z(
        n118) );
  MUX4D0 U486 ( .I0(n122), .I1(n120), .I2(n121), .I3(n119), .S0(n173), .S1(
        n177), .Z(N61) );
  MUX4D0 U487 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n204), .S1(n189), .Z(
        n121) );
  MUX4D0 U488 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n204), .S1(n189), .Z(
        n120) );
  MUX4D0 U489 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n204), .S1(n189), .Z(
        n122) );
  MUX4D0 U490 ( .I0(n146), .I1(n144), .I2(n145), .I3(n143), .S0(n174), .S1(
        n178), .Z(N55) );
  MUX4D0 U491 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n206), .S1(n191), .Z(
        n145) );
  MUX4D0 U492 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n206), .S1(n191), .Z(
        n144) );
  MUX4D0 U493 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n206), .S1(n191), .Z(
        n146) );
  MUX4D0 U494 ( .I0(n150), .I1(n148), .I2(n149), .I3(n147), .S0(n174), .S1(
        n178), .Z(N54) );
  MUX4D0 U495 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n207), .S1(n192), .Z(
        n149) );
  MUX4D0 U496 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n207), .S1(n192), .Z(
        n148) );
  MUX4D0 U497 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n207), .S1(n192), .Z(
        n150) );
  MUX4D0 U498 ( .I0(n162), .I1(n160), .I2(n161), .I3(n159), .S0(n174), .S1(
        n178), .Z(N51) );
  MUX4D0 U499 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n208), .S1(n193), .Z(
        n161) );
  MUX4D0 U500 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n208), .S1(n193), .Z(
        n160) );
  MUX4D0 U501 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n208), .S1(n193), .Z(
        n162) );
  MUX4D0 U502 ( .I0(n166), .I1(n164), .I2(n165), .I3(n163), .S0(n174), .S1(
        n178), .Z(N50) );
  MUX4D0 U503 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n208), .S1(n193), .Z(
        n165) );
  MUX4D0 U504 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n208), .S1(n193), .Z(
        n164) );
  MUX4D0 U505 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n208), .S1(n193), .Z(
        n166) );
  MUX4D0 U506 ( .I0(n28), .I1(n26), .I2(n27), .I3(n25), .S0(n172), .S1(n176), 
        .Z(N75) );
  MUX4D0 U507 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n200), .S1(n185), .Z(n27)
         );
  MUX4D0 U508 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n200), .S1(n185), .Z(n26) );
  MUX4D0 U509 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n200), .S1(n185), .Z(n28)
         );
  MUX4D0 U510 ( .I0(n106), .I1(n104), .I2(n105), .I3(n102), .S0(n173), .S1(
        n177), .Z(N65) );
  MUX4D0 U511 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n203), .S1(n188), .Z(
        n105) );
  MUX4D0 U512 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n203), .S1(n188), .Z(
        n104) );
  MUX4D0 U513 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n203), .S1(n188), .Z(
        n106) );
  MUX4D0 U514 ( .I0(n134), .I1(n132), .I2(n133), .I3(n131), .S0(n174), .S1(
        n178), .Z(N58) );
  MUX4D0 U515 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n205), .S1(n190), .Z(
        n133) );
  MUX4D0 U516 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n205), .S1(n190), .Z(
        n132) );
  MUX4D0 U517 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n205), .S1(n190), .Z(
        n134) );
  MUX4D0 U518 ( .I0(n138), .I1(n136), .I2(n137), .I3(n135), .S0(n174), .S1(
        n178), .Z(N57) );
  MUX4D0 U519 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n206), .S1(n191), .Z(
        n137) );
  MUX4D0 U520 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n206), .S1(n191), .Z(
        n136) );
  MUX4D0 U521 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n206), .S1(n191), .Z(
        n138) );
  MUX4D0 U522 ( .I0(n4), .I1(n2), .I2(n3), .I3(n1), .S0(n172), .S1(n176), .Z(
        N81) );
  MUX4D0 U523 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n198), .S1(n183), .Z(n3)
         );
  MUX4D0 U524 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n198), .S1(n183), .Z(n2)
         );
  MUX4D0 U525 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n198), .S1(n183), .Z(n4)
         );
  MUX4D0 U526 ( .I0(n20), .I1(n18), .I2(n19), .I3(n17), .S0(n172), .S1(n176), 
        .Z(N77) );
  MUX4D0 U527 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n199), .S1(n184), .Z(n19)
         );
  MUX4D0 U528 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n199), .S1(n184), .Z(n18) );
  MUX4D0 U529 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n199), .S1(n184), .Z(n20)
         );
  MUX4D0 U530 ( .I0(n44), .I1(n42), .I2(n43), .I3(n41), .S0(n173), .S1(n177), 
        .Z(N71) );
  MUX4D0 U531 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n201), .S1(n186), .Z(n43) );
  MUX4D0 U532 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n201), .S1(n186), .Z(
        n42) );
  MUX4D0 U533 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n201), .S1(n186), .Z(n44) );
  MUX4D0 U534 ( .I0(n48), .I1(n46), .I2(n47), .I3(n45), .S0(n173), .S1(n177), 
        .Z(N70) );
  MUX4D0 U535 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n201), .S1(n186), .Z(n47) );
  MUX4D0 U536 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n201), .S1(n186), .Z(
        n46) );
  MUX4D0 U537 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n201), .S1(n186), .Z(n48) );
  MUX4D0 U538 ( .I0(n60), .I1(n58), .I2(n59), .I3(n57), .S0(n173), .S1(n177), 
        .Z(N67) );
  MUX4D0 U539 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n202), .S1(n187), .Z(n59) );
  MUX4D0 U540 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n202), .S1(n187), .Z(
        n58) );
  MUX4D0 U541 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n202), .S1(n187), .Z(n60) );
  MUX4D0 U542 ( .I0(n114), .I1(n112), .I2(n113), .I3(n111), .S0(n173), .S1(
        n177), .Z(N63) );
  MUX4D0 U543 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n204), .S1(n189), .Z(
        n113) );
  MUX4D0 U544 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n204), .S1(n189), .Z(
        n112) );
  MUX4D0 U545 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n204), .S1(n189), .Z(
        n114) );
  MUX4D0 U546 ( .I0(n126), .I1(n124), .I2(n125), .I3(n123), .S0(n174), .S1(
        n178), .Z(N60) );
  MUX4D0 U547 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n205), .S1(n190), .Z(
        n125) );
  MUX4D0 U548 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n205), .S1(n190), .Z(
        n124) );
  MUX4D0 U549 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n205), .S1(n190), .Z(
        n126) );
  MUX4D0 U550 ( .I0(n142), .I1(n140), .I2(n141), .I3(n139), .S0(n174), .S1(
        n178), .Z(N56) );
  MUX4D0 U551 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n206), .S1(n191), .Z(
        n141) );
  MUX4D0 U552 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n206), .S1(n191), .Z(
        n140) );
  MUX4D0 U553 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n206), .S1(n191), .Z(
        n142) );
  MUX4D0 U554 ( .I0(n154), .I1(n152), .I2(n153), .I3(n151), .S0(n174), .S1(
        n178), .Z(N53) );
  MUX4D0 U555 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n207), .S1(n192), .Z(
        n153) );
  MUX4D0 U556 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n207), .S1(n192), .Z(
        n152) );
  MUX4D0 U557 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n207), .S1(n192), .Z(
        n154) );
  MUX4D0 U558 ( .I0(n158), .I1(n156), .I2(n157), .I3(n155), .S0(n174), .S1(
        n178), .Z(N52) );
  MUX4D0 U559 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n207), .S1(n192), .Z(
        n157) );
  MUX4D0 U560 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n207), .S1(n192), .Z(
        n156) );
  MUX4D0 U561 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n207), .S1(n192), .Z(
        n158) );
  MUX4D0 U562 ( .I0(n24), .I1(n22), .I2(n23), .I3(n21), .S0(n172), .S1(n176), 
        .Z(N76) );
  MUX4D0 U563 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n199), .S1(n184), .Z(n23)
         );
  MUX4D0 U564 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n199), .S1(n184), .Z(n22) );
  MUX4D0 U565 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n199), .S1(n184), .Z(n24)
         );
  MUX4D0 U566 ( .I0(n40), .I1(n38), .I2(n39), .I3(n37), .S0(n173), .S1(n177), 
        .Z(N72) );
  MUX4D0 U567 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n201), .S1(n186), .Z(n39)
         );
  MUX4D0 U568 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n201), .S1(n186), .Z(n38) );
  MUX4D0 U569 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n201), .S1(n186), .Z(n40)
         );
  MUX4D0 U570 ( .I0(n64), .I1(n62), .I2(n63), .I3(n61), .S0(n173), .S1(n177), 
        .Z(N66) );
  MUX4D0 U571 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n203), .S1(n188), .Z(n63) );
  MUX4D0 U572 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n203), .S1(n188), .Z(
        n62) );
  MUX4D0 U573 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n203), .S1(n188), .Z(n64) );
  MUX4D0 U574 ( .I0(n110), .I1(n108), .I2(n109), .I3(n107), .S0(n173), .S1(
        n177), .Z(N64) );
  MUX4D0 U575 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n203), .S1(n188), .Z(
        n109) );
  MUX4D0 U576 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n203), .S1(n188), .Z(
        n108) );
  MUX4D0 U577 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n203), .S1(n188), .Z(
        n110) );
  MUX4D0 U578 ( .I0(n130), .I1(n128), .I2(n129), .I3(n127), .S0(n174), .S1(
        n178), .Z(N59) );
  MUX4D0 U579 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n205), .S1(n190), .Z(
        n129) );
  MUX4D0 U580 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n205), .S1(n190), .Z(
        n128) );
  MUX4D0 U581 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n205), .S1(n190), .Z(
        n130) );
  MUX4D0 U582 ( .I0(n170), .I1(n168), .I2(n169), .I3(n167), .S0(n174), .S1(
        n178), .Z(N49) );
  MUX4D0 U583 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n208), .S1(n193), .Z(
        n169) );
  MUX4D0 U584 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n208), .S1(n193), .Z(
        n168) );
  MUX4D0 U585 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n208), .S1(n193), .Z(
        n170) );
  MUX4D0 U586 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n208), .S1(n193), .Z(
        n167) );
  MUX4D0 U587 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n198), .S1(n183), .Z(n1)
         );
  MUX4D0 U588 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n198), .S1(n183), .Z(n5)
         );
  MUX4D0 U589 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n198), .S1(n183), .Z(n9)
         );
  MUX4D0 U590 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n199), .S1(n184), .Z(n17) );
  MUX4D0 U591 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n199), .S1(n184), .Z(n21) );
  MUX4D0 U592 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n200), .S1(n185), .Z(n25) );
  MUX4D0 U593 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n200), .S1(n185), .Z(n29) );
  MUX4D0 U594 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n201), .S1(n186), .Z(n37) );
  MUX4D0 U595 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n201), .S1(n186), .Z(
        n41) );
  MUX4D0 U596 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n201), .S1(n186), .Z(
        n45) );
  MUX4D0 U597 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n202), .S1(n187), .Z(
        n49) );
  MUX4D0 U598 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n202), .S1(n187), .Z(
        n53) );
  MUX4D0 U599 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n202), .S1(n187), .Z(
        n57) );
  MUX4D0 U600 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n203), .S1(n188), .Z(
        n61) );
  MUX4D0 U601 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n203), .S1(n188), .Z(
        n102) );
  MUX4D0 U602 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n203), .S1(n188), .Z(
        n107) );
  MUX4D0 U603 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n204), .S1(n189), .Z(
        n111) );
  MUX4D0 U604 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n204), .S1(n189), .Z(
        n115) );
  MUX4D0 U605 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n204), .S1(n189), .Z(
        n119) );
  MUX4D0 U606 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n205), .S1(n190), .Z(
        n123) );
  MUX4D0 U607 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n205), .S1(n190), .Z(
        n127) );
  MUX4D0 U608 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n205), .S1(n190), .Z(
        n131) );
  MUX4D0 U609 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n206), .S1(n191), .Z(
        n135) );
  MUX4D0 U610 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n206), .S1(n191), .Z(
        n139) );
  MUX4D0 U611 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n206), .S1(n191), .Z(
        n143) );
  MUX4D0 U612 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n207), .S1(n192), .Z(
        n147) );
  MUX4D0 U613 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n207), .S1(n192), .Z(
        n151) );
  MUX4D0 U614 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n207), .S1(n192), .Z(
        n155) );
  MUX4D0 U615 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n208), .S1(n193), .Z(
        n159) );
  MUX4D0 U616 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n208), .S1(n193), .Z(
        n163) );
  BUFFD1 U617 ( .I(N47), .Z(n494) );
  BUFFD1 U618 ( .I(N46), .Z(n493) );
  BUFFD1 U619 ( .I(N44), .Z(n491) );
  BUFFD1 U620 ( .I(N45), .Z(n492) );
  MUX4D0 U621 ( .I0(n36), .I1(n34), .I2(n35), .I3(n33), .S0(n172), .S1(n176), 
        .Z(N73) );
  MUX4D0 U622 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n200), .S1(n185), .Z(n35)
         );
  MUX4D0 U623 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n200), .S1(n185), .Z(n34) );
  MUX4D0 U624 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n200), .S1(n185), .Z(n36)
         );
  MUX4D0 U625 ( .I0(n16), .I1(n14), .I2(n15), .I3(n13), .S0(n172), .S1(n176), 
        .Z(N78) );
  MUX4D0 U626 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n199), .S1(n184), .Z(n15)
         );
  MUX4D0 U627 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n199), .S1(n184), .Z(n14) );
  MUX4D0 U628 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n199), .S1(n184), .Z(n16)
         );
  MUX4D0 U629 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n199), .S1(n184), .Z(n13) );
  MUX4D0 U630 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n200), .S1(n185), .Z(n33) );
  ND2D1 U631 ( .A1(AddrW[1]), .A2(n593), .ZN(n600) );
  ND2D1 U632 ( .A1(AddrW[2]), .A2(AddrW[1]), .ZN(n603) );
  ND2D1 U633 ( .A1(n592), .A2(AddrW[0]), .ZN(n596) );
  ND2D1 U634 ( .A1(AddrW[2]), .A2(n594), .ZN(n601) );
  ND2D1 U635 ( .A1(AddrW[0]), .A2(n598), .ZN(n604) );
  INR2D1 U636 ( .A1(Write), .B1(AddrW[3]), .ZN(n592) );
  INVD1 U637 ( .I(AddrW[1]), .ZN(n594) );
  INVD1 U638 ( .I(AddrW[0]), .ZN(n597) );
  INVD1 U639 ( .I(AddrW[2]), .ZN(n593) );
  AN2D1 U640 ( .A1(Write), .A2(AddrW[3]), .Z(n598) );
  INVD1 U641 ( .I(n490), .ZN(n489) );
  INVD1 U642 ( .I(Read), .ZN(n490) );
  INR2D1 U643 ( .A1(ClkW), .B1(N9), .ZN(ClockW) );
  INVD1 U644 ( .I(n476), .ZN(n475) );
  INVD1 U645 ( .I(ClockR), .ZN(n476) );
  INR2D1 U646 ( .A1(ClkR), .B1(N9), .ZN(ClockR) );
  INVD0 U647 ( .I(ChipEna), .ZN(N9) );
endmodule


module ClockComparator_1 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n12,
         n13, n14, n15, n16;

  AO211D1 U8 ( .A1(n15), .A2(n14), .B(N8), .C(N5), .Z(n13) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n16), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n16), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n12), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n12), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n16), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n16), .QN(n15) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n12), .QN(n16) );
  INVD1 U3 ( .I(Reset), .ZN(n12) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n15), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n14), .A2(n15), .B(n13), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n14) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_2 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n12,
         n13, n14, n15, n16;

  AO211D1 U8 ( .A1(n15), .A2(n14), .B(N8), .C(N5), .Z(n13) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n16), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n16), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n12), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n12), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n16), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n16), .QN(n15) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n12), .QN(n16) );
  INVD1 U3 ( .I(Reset), .ZN(n12) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n15), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n14), .A2(n15), .B(n13), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n14) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module ClockComparator_3 ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   \ClockInN[0] , N5, N6, \CounterClockN[0] , N7, N8, N9, N19, N20, n12,
         n13, n14, n15, n16;

  AO211D1 U8 ( .A1(n15), .A2(n14), .B(N8), .C(N5), .Z(n13) );
  DFCND1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n16), .QN(
        N19) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n16), .Q(
        \CounterClockN[0] ), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n12), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n12), .Q(
        AdjustFreq[1]) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n16), .Q(\ClockInN[0] ), .QN(N5) );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n16), .QN(n15) );
  DFSND1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n12), .QN(n16) );
  INVD1 U3 ( .I(Reset), .ZN(n12) );
  XNR2D1 U4 ( .A1(\ClockInN[0] ), .A2(n15), .ZN(N6) );
  NR2D1 U5 ( .A1(N6), .A2(N5), .ZN(N9) );
  OAI21D1 U6 ( .A1(n14), .A2(n15), .B(n13), .ZN(N20) );
  NR2D1 U7 ( .A1(N19), .A2(N7), .ZN(n14) );
  XNR2D1 U9 ( .A1(N19), .A2(\CounterClockN[0] ), .ZN(N8) );
endmodule


module VFO_1 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_1_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_1_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_1_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n69), .CP(FastClock), .CDN(n38), .Q(ClockOut)
         );
  DFSND1 \DivideFactor_reg[4]  ( .D(n67), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[4]), .QN(n53) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n68), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[1]), .QN(n65) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n66), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[0]), .QN(n63) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[3]), .QN(n58) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[5]), .QN(n48) );
  INVD1 U3 ( .I(n40), .ZN(n38) );
  INVD1 U4 ( .I(n40), .ZN(n39) );
  INVD1 U5 ( .I(n41), .ZN(n40) );
  INVD1 U6 ( .I(Reset), .ZN(n41) );
  AO222D0 U7 ( .A1(N27), .A2(n42), .B1(N35), .B2(n43), .C1(DivideFactor[0]), 
        .C2(n44), .Z(n66) );
  AO222D0 U8 ( .A1(N31), .A2(n42), .B1(N39), .B2(n43), .C1(DivideFactor[4]), 
        .C2(n44), .Z(n67) );
  AO222D0 U9 ( .A1(N28), .A2(n42), .B1(N36), .B2(n43), .C1(DivideFactor[1]), 
        .C2(n44), .Z(n68) );
  CKND0 U10 ( .CLK(N54), .CN(n44) );
  AN2D0 U11 ( .A1(n45), .A2(n46), .Z(n43) );
  AN3D0 U12 ( .A1(n47), .A2(n48), .A3(n49), .Z(n42) );
  CKXOR2D0 U13 ( .A1(ClockOut), .A2(n50), .Z(n69) );
  AO22D0 U14 ( .A1(N32), .A2(n49), .B1(N40), .B2(n45), .Z(N55) );
  MUX2ND0 U15 ( .I0(n51), .I1(n52), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U16 ( .A1(AdjustFreq[1]), .A2(n46), .ZN(n52) );
  ND3D0 U17 ( .A1(n53), .A2(n48), .A3(n54), .ZN(n46) );
  ND4D0 U18 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n54) );
  IND3D0 U19 ( .A1(AdjustFreq[1]), .B1(n48), .B2(n47), .ZN(n51) );
  CKND2D0 U20 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n47) );
  AO22D0 U21 ( .A1(N30), .A2(n49), .B1(N38), .B2(n45), .Z(N51) );
  AO22D0 U22 ( .A1(N29), .A2(n49), .B1(N37), .B2(n45), .Z(N49) );
  AN2D0 U23 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n45) );
  NR2D0 U24 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n49) );
  INR2D0 U25 ( .A1(N14), .B1(n50), .ZN(N21) );
  INR2D0 U26 ( .A1(N13), .B1(n50), .ZN(N20) );
  INR2D0 U27 ( .A1(N12), .B1(n50), .ZN(N19) );
  INR2D0 U28 ( .A1(N11), .B1(n50), .ZN(N18) );
  INR2D0 U29 ( .A1(N10), .B1(n50), .ZN(N17) );
  INR2D0 U30 ( .A1(N9), .B1(n50), .ZN(N16) );
  OA21D0 U31 ( .A1(FastDivvy[5]), .A2(n48), .B(n55), .Z(n50) );
  IOA22D0 U32 ( .B1(n56), .B2(n57), .A1(n48), .A2(FastDivvy[5]), .ZN(n55) );
  AOI221D0 U33 ( .A1(FastDivvy[4]), .A2(n53), .B1(FastDivvy[3]), .B2(n58), .C(
        n59), .ZN(n57) );
  AOI221D0 U34 ( .A1(DivideFactor[3]), .A2(n60), .B1(DivideFactor[2]), .B2(n61), .C(n62), .ZN(n59) );
  IAO21D0 U35 ( .A1(n61), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n62) );
  OAI32D0 U36 ( .A1(n63), .A2(FastDivvy[0]), .A3(n64), .B1(FastDivvy[1]), .B2(
        n65), .ZN(n61) );
  AN2D0 U37 ( .A1(FastDivvy[1]), .A2(n65), .Z(n64) );
  CKND0 U38 ( .CLK(FastDivvy[3]), .CN(n60) );
  NR2D0 U39 ( .A1(FastDivvy[4]), .A2(n53), .ZN(n56) );
  CKND0 U40 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U41 ( .A1(WireD[5]), .A2(n39), .ZN(WireD[0]) );
endmodule


module VFO_2 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_2_DW01_dec_0 \Sampler/sub_193  ( .A({DivideFactor[5:2], n16, n80}), 
        .SUM({N40, N39, N38, N37, N36, N35}) );
  VFO_2_DW01_inc_0 \Sampler/add_190  ( .A({DivideFactor[5:2], n16, n80}), 
        .SUM({N32, N31, N30, N29, N28, N27}) );
  VFO_2_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n218), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n249), .CP(FastClock), .CDN(n218), .Q(ClockOut)
         );
  EDFCNQD1 \DivideFactor_reg[5]  ( .D(N55), .E(n142), .CP(Sample), .CDN(n218), 
        .Q(DivideFactor[5]) );
  EDFCNQD1 \DivideFactor_reg[2]  ( .D(N49), .E(n142), .CP(Sample), .CDN(n218), 
        .Q(DivideFactor[2]) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n247), .CP(Sample), .SDN(n221), .Q(
        DivideFactor[4]), .QN(n233) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n1), .CP(Sample), .SDN(n221), .Q(
        DivideFactor[1]), .QN(n245) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n22), .CP(Sample), .SDN(n221), .Q(
        DivideFactor[0]), .QN(n243) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(n81), .E(n142), .CP(Sample), .CDN(n221), 
        .Q(DivideFactor[3]), .QN(n238) );
  BUFFD0 U3 ( .I(n2), .Z(n1) );
  BUFFD0 U4 ( .I(n3), .Z(n2) );
  BUFFD0 U5 ( .I(n4), .Z(n3) );
  BUFFD0 U6 ( .I(n5), .Z(n4) );
  BUFFD0 U7 ( .I(n6), .Z(n5) );
  BUFFD0 U8 ( .I(n7), .Z(n6) );
  BUFFD0 U9 ( .I(n8), .Z(n7) );
  BUFFD0 U10 ( .I(n9), .Z(n8) );
  BUFFD0 U11 ( .I(n10), .Z(n9) );
  BUFFD0 U12 ( .I(n11), .Z(n10) );
  BUFFD0 U13 ( .I(n12), .Z(n11) );
  BUFFD0 U14 ( .I(n13), .Z(n12) );
  BUFFD0 U15 ( .I(n14), .Z(n13) );
  BUFFD0 U16 ( .I(n15), .Z(n14) );
  BUFFD0 U17 ( .I(n248), .Z(n15) );
  BUFFD0 U18 ( .I(n20), .Z(n16) );
  BUFFD0 U19 ( .I(DivideFactor[1]), .Z(n20) );
  BUFFD0 U20 ( .I(n25), .Z(n22) );
  BUFFD0 U21 ( .I(n246), .Z(n23) );
  BUFFD0 U22 ( .I(n23), .Z(n24) );
  BUFFD0 U23 ( .I(n26), .Z(n25) );
  BUFFD0 U24 ( .I(n27), .Z(n26) );
  BUFFD0 U25 ( .I(n28), .Z(n27) );
  BUFFD0 U26 ( .I(n29), .Z(n28) );
  BUFFD0 U27 ( .I(n30), .Z(n29) );
  BUFFD0 U28 ( .I(n31), .Z(n30) );
  BUFFD0 U29 ( .I(n32), .Z(n31) );
  BUFFD0 U30 ( .I(n33), .Z(n32) );
  BUFFD0 U31 ( .I(n34), .Z(n33) );
  BUFFD0 U32 ( .I(n35), .Z(n34) );
  BUFFD0 U33 ( .I(n36), .Z(n35) );
  BUFFD0 U34 ( .I(n37), .Z(n36) );
  BUFFD0 U35 ( .I(n38), .Z(n37) );
  BUFFD0 U36 ( .I(n39), .Z(n38) );
  BUFFD0 U37 ( .I(n40), .Z(n39) );
  BUFFD0 U38 ( .I(n41), .Z(n40) );
  BUFFD0 U39 ( .I(n42), .Z(n41) );
  BUFFD0 U40 ( .I(n43), .Z(n42) );
  BUFFD0 U41 ( .I(n44), .Z(n43) );
  BUFFD0 U42 ( .I(n45), .Z(n44) );
  BUFFD0 U43 ( .I(n46), .Z(n45) );
  BUFFD0 U44 ( .I(n47), .Z(n46) );
  BUFFD0 U45 ( .I(n48), .Z(n47) );
  BUFFD0 U46 ( .I(n49), .Z(n48) );
  BUFFD0 U47 ( .I(n50), .Z(n49) );
  BUFFD0 U48 ( .I(n51), .Z(n50) );
  BUFFD0 U49 ( .I(n52), .Z(n51) );
  BUFFD0 U50 ( .I(n53), .Z(n52) );
  BUFFD0 U51 ( .I(n54), .Z(n53) );
  BUFFD0 U52 ( .I(n55), .Z(n54) );
  BUFFD0 U53 ( .I(n56), .Z(n55) );
  BUFFD0 U54 ( .I(n57), .Z(n56) );
  BUFFD0 U55 ( .I(n58), .Z(n57) );
  BUFFD0 U56 ( .I(n59), .Z(n58) );
  BUFFD0 U57 ( .I(n60), .Z(n59) );
  BUFFD0 U58 ( .I(n61), .Z(n60) );
  BUFFD0 U59 ( .I(n62), .Z(n61) );
  BUFFD0 U60 ( .I(n63), .Z(n62) );
  BUFFD0 U61 ( .I(n64), .Z(n63) );
  BUFFD0 U62 ( .I(n65), .Z(n64) );
  BUFFD0 U63 ( .I(n66), .Z(n65) );
  BUFFD0 U64 ( .I(n67), .Z(n66) );
  BUFFD0 U65 ( .I(n68), .Z(n67) );
  BUFFD0 U66 ( .I(n69), .Z(n68) );
  BUFFD0 U67 ( .I(n70), .Z(n69) );
  BUFFD0 U68 ( .I(n71), .Z(n70) );
  BUFFD0 U69 ( .I(n72), .Z(n71) );
  BUFFD0 U70 ( .I(n73), .Z(n72) );
  BUFFD0 U71 ( .I(n74), .Z(n73) );
  BUFFD0 U72 ( .I(n75), .Z(n74) );
  BUFFD0 U73 ( .I(n76), .Z(n75) );
  BUFFD0 U74 ( .I(n77), .Z(n76) );
  BUFFD0 U75 ( .I(n78), .Z(n77) );
  BUFFD0 U76 ( .I(n24), .Z(n78) );
  BUFFD0 U77 ( .I(DivideFactor[0]), .Z(n79) );
  CKBXD0 U78 ( .I(n79), .Z(n80) );
  BUFFD0 U79 ( .I(n85), .Z(n81) );
  BUFFD0 U80 ( .I(N51), .Z(n82) );
  BUFFD0 U81 ( .I(n82), .Z(n83) );
  BUFFD0 U82 ( .I(n83), .Z(n84) );
  BUFFD0 U83 ( .I(n86), .Z(n85) );
  BUFFD0 U84 ( .I(n87), .Z(n86) );
  BUFFD0 U85 ( .I(n88), .Z(n87) );
  BUFFD0 U86 ( .I(n89), .Z(n88) );
  BUFFD0 U87 ( .I(n90), .Z(n89) );
  BUFFD0 U88 ( .I(n91), .Z(n90) );
  BUFFD0 U89 ( .I(n92), .Z(n91) );
  BUFFD0 U90 ( .I(n93), .Z(n92) );
  BUFFD0 U91 ( .I(n94), .Z(n93) );
  BUFFD0 U92 ( .I(n95), .Z(n94) );
  BUFFD0 U93 ( .I(n96), .Z(n95) );
  BUFFD0 U94 ( .I(n97), .Z(n96) );
  BUFFD0 U95 ( .I(n98), .Z(n97) );
  BUFFD0 U96 ( .I(n99), .Z(n98) );
  BUFFD0 U97 ( .I(n100), .Z(n99) );
  BUFFD0 U98 ( .I(n101), .Z(n100) );
  BUFFD0 U99 ( .I(n102), .Z(n101) );
  BUFFD0 U100 ( .I(n103), .Z(n102) );
  BUFFD0 U101 ( .I(n104), .Z(n103) );
  BUFFD0 U102 ( .I(n105), .Z(n104) );
  BUFFD0 U103 ( .I(n106), .Z(n105) );
  BUFFD0 U104 ( .I(n107), .Z(n106) );
  BUFFD0 U105 ( .I(n108), .Z(n107) );
  BUFFD0 U106 ( .I(n109), .Z(n108) );
  BUFFD0 U107 ( .I(n110), .Z(n109) );
  BUFFD0 U108 ( .I(n111), .Z(n110) );
  BUFFD0 U109 ( .I(n112), .Z(n111) );
  BUFFD0 U110 ( .I(n113), .Z(n112) );
  BUFFD0 U111 ( .I(n114), .Z(n113) );
  BUFFD0 U112 ( .I(n115), .Z(n114) );
  BUFFD0 U113 ( .I(n116), .Z(n115) );
  BUFFD0 U114 ( .I(n117), .Z(n116) );
  BUFFD0 U115 ( .I(n118), .Z(n117) );
  BUFFD0 U116 ( .I(n119), .Z(n118) );
  BUFFD0 U117 ( .I(n120), .Z(n119) );
  BUFFD0 U118 ( .I(n121), .Z(n120) );
  BUFFD0 U119 ( .I(n122), .Z(n121) );
  BUFFD0 U120 ( .I(n123), .Z(n122) );
  BUFFD0 U121 ( .I(n124), .Z(n123) );
  BUFFD0 U122 ( .I(n125), .Z(n124) );
  BUFFD0 U123 ( .I(n126), .Z(n125) );
  BUFFD0 U124 ( .I(n127), .Z(n126) );
  BUFFD0 U125 ( .I(n128), .Z(n127) );
  BUFFD0 U126 ( .I(n129), .Z(n128) );
  BUFFD0 U127 ( .I(n130), .Z(n129) );
  BUFFD0 U128 ( .I(n131), .Z(n130) );
  BUFFD0 U129 ( .I(n132), .Z(n131) );
  BUFFD0 U130 ( .I(n133), .Z(n132) );
  BUFFD0 U131 ( .I(n134), .Z(n133) );
  BUFFD0 U132 ( .I(n135), .Z(n134) );
  BUFFD0 U133 ( .I(n136), .Z(n135) );
  BUFFD0 U134 ( .I(n137), .Z(n136) );
  BUFFD0 U135 ( .I(n138), .Z(n137) );
  BUFFD0 U136 ( .I(n139), .Z(n138) );
  BUFFD0 U137 ( .I(n84), .Z(n139) );
  MUX2ND1 U138 ( .I0(n196), .I1(n232), .S(AdjustFreq[0]), .ZN(N54) );
  BUFFD0 U139 ( .I(N54), .Z(n140) );
  BUFFD0 U140 ( .I(n143), .Z(n141) );
  BUFFD0 U141 ( .I(n141), .Z(n142) );
  BUFFD0 U142 ( .I(n144), .Z(n143) );
  BUFFD0 U143 ( .I(n145), .Z(n144) );
  BUFFD0 U144 ( .I(n146), .Z(n145) );
  BUFFD0 U145 ( .I(n147), .Z(n146) );
  BUFFD0 U146 ( .I(n148), .Z(n147) );
  BUFFD0 U147 ( .I(n149), .Z(n148) );
  BUFFD0 U148 ( .I(n150), .Z(n149) );
  BUFFD0 U149 ( .I(n151), .Z(n150) );
  BUFFD0 U150 ( .I(n152), .Z(n151) );
  BUFFD0 U151 ( .I(n153), .Z(n152) );
  BUFFD0 U152 ( .I(n154), .Z(n153) );
  BUFFD0 U153 ( .I(n155), .Z(n154) );
  BUFFD0 U154 ( .I(n156), .Z(n155) );
  BUFFD0 U155 ( .I(n157), .Z(n156) );
  BUFFD0 U156 ( .I(n158), .Z(n157) );
  BUFFD0 U157 ( .I(n159), .Z(n158) );
  BUFFD0 U158 ( .I(n160), .Z(n159) );
  BUFFD0 U159 ( .I(n161), .Z(n160) );
  BUFFD0 U160 ( .I(n162), .Z(n161) );
  BUFFD0 U161 ( .I(n163), .Z(n162) );
  BUFFD0 U162 ( .I(n164), .Z(n163) );
  BUFFD0 U163 ( .I(n165), .Z(n164) );
  BUFFD0 U164 ( .I(n166), .Z(n165) );
  BUFFD0 U165 ( .I(n167), .Z(n166) );
  BUFFD0 U166 ( .I(n168), .Z(n167) );
  BUFFD0 U167 ( .I(n169), .Z(n168) );
  BUFFD0 U168 ( .I(n170), .Z(n169) );
  BUFFD0 U169 ( .I(n171), .Z(n170) );
  BUFFD0 U170 ( .I(n172), .Z(n171) );
  BUFFD0 U171 ( .I(n173), .Z(n172) );
  BUFFD0 U172 ( .I(n174), .Z(n173) );
  BUFFD0 U173 ( .I(n175), .Z(n174) );
  BUFFD0 U174 ( .I(n176), .Z(n175) );
  BUFFD0 U175 ( .I(n177), .Z(n176) );
  BUFFD0 U176 ( .I(n178), .Z(n177) );
  BUFFD0 U177 ( .I(n179), .Z(n178) );
  BUFFD0 U178 ( .I(n180), .Z(n179) );
  BUFFD0 U179 ( .I(n181), .Z(n180) );
  BUFFD0 U180 ( .I(n182), .Z(n181) );
  BUFFD0 U181 ( .I(n183), .Z(n182) );
  BUFFD0 U182 ( .I(n184), .Z(n183) );
  BUFFD0 U183 ( .I(n185), .Z(n184) );
  BUFFD0 U184 ( .I(n186), .Z(n185) );
  BUFFD0 U185 ( .I(n187), .Z(n186) );
  BUFFD0 U186 ( .I(n188), .Z(n187) );
  BUFFD0 U187 ( .I(n189), .Z(n188) );
  BUFFD0 U188 ( .I(n190), .Z(n189) );
  BUFFD0 U189 ( .I(n191), .Z(n190) );
  BUFFD0 U190 ( .I(n192), .Z(n191) );
  BUFFD0 U191 ( .I(n193), .Z(n192) );
  BUFFD0 U192 ( .I(n194), .Z(n193) );
  BUFFD0 U193 ( .I(n195), .Z(n194) );
  BUFFD0 U194 ( .I(n140), .Z(n195) );
  BUFFD0 U195 ( .I(n231), .Z(n196) );
  INVD1 U196 ( .I(n220), .ZN(n218) );
  INVD1 U197 ( .I(n220), .ZN(n219) );
  INVD1 U198 ( .I(n221), .ZN(n220) );
  INVD1 U199 ( .I(Reset), .ZN(n221) );
  AO222D0 U200 ( .A1(N27), .A2(n222), .B1(N35), .B2(n223), .C1(n80), .C2(n224), 
        .Z(n246) );
  AO222D0 U201 ( .A1(N31), .A2(n222), .B1(N39), .B2(n223), .C1(DivideFactor[4]), .C2(n224), .Z(n247) );
  AO222D0 U202 ( .A1(N28), .A2(n222), .B1(N36), .B2(n223), .C1(n16), .C2(n224), 
        .Z(n248) );
  CKND0 U203 ( .CLK(n141), .CN(n224) );
  AN2D0 U204 ( .A1(n225), .A2(n226), .Z(n223) );
  AN3D0 U205 ( .A1(n227), .A2(n228), .A3(n229), .Z(n222) );
  CKXOR2D0 U206 ( .A1(ClockOut), .A2(n230), .Z(n249) );
  AO22D0 U207 ( .A1(N32), .A2(n229), .B1(N40), .B2(n225), .Z(N55) );
  CKND2D0 U208 ( .A1(AdjustFreq[1]), .A2(n226), .ZN(n232) );
  ND3D0 U209 ( .A1(n233), .A2(n228), .A3(n234), .ZN(n226) );
  ND4D0 U210 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(n16), .A4(n80), 
        .ZN(n234) );
  IND3D0 U211 ( .A1(AdjustFreq[1]), .B1(n228), .B2(n227), .ZN(n231) );
  CKND2D0 U212 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n227) );
  AO22D0 U213 ( .A1(N30), .A2(n229), .B1(N38), .B2(n225), .Z(N51) );
  AO22D0 U214 ( .A1(N29), .A2(n229), .B1(N37), .B2(n225), .Z(N49) );
  AN2D0 U215 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n225) );
  NR2D0 U216 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n229) );
  INR2D0 U217 ( .A1(N14), .B1(n230), .ZN(N21) );
  INR2D0 U218 ( .A1(N13), .B1(n230), .ZN(N20) );
  INR2D0 U219 ( .A1(N12), .B1(n230), .ZN(N19) );
  INR2D0 U220 ( .A1(N11), .B1(n230), .ZN(N18) );
  INR2D0 U221 ( .A1(N10), .B1(n230), .ZN(N17) );
  INR2D0 U222 ( .A1(N9), .B1(n230), .ZN(N16) );
  OA21D0 U223 ( .A1(FastDivvy[5]), .A2(n228), .B(n235), .Z(n230) );
  IOA22D0 U224 ( .B1(n236), .B2(n237), .A1(n228), .A2(FastDivvy[5]), .ZN(n235)
         );
  AOI221D0 U225 ( .A1(FastDivvy[4]), .A2(n233), .B1(FastDivvy[3]), .B2(n238), 
        .C(n239), .ZN(n237) );
  AOI221D0 U226 ( .A1(DivideFactor[3]), .A2(n240), .B1(DivideFactor[2]), .B2(
        n241), .C(n242), .ZN(n239) );
  IAO21D0 U227 ( .A1(n241), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n242)
         );
  OAI32D0 U228 ( .A1(n243), .A2(FastDivvy[0]), .A3(n244), .B1(FastDivvy[1]), 
        .B2(n245), .ZN(n241) );
  AN2D0 U229 ( .A1(FastDivvy[1]), .A2(n245), .Z(n244) );
  CKND0 U230 ( .CLK(FastDivvy[3]), .CN(n240) );
  NR2D0 U231 ( .A1(FastDivvy[4]), .A2(n233), .ZN(n236) );
  CKND0 U232 ( .CLK(DivideFactor[5]), .CN(n228) );
  CKND0 U233 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U234 ( .A1(WireD[5]), .A2(n219), .ZN(WireD[0]) );
endmodule


module VFO_3 ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay85ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay85ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay85ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay85ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay85ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_3_DW01_dec_0 \Sampler/sub_193  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_3_DW01_inc_0 \Sampler/add_190  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_3_DW01_inc_1 \ClockOutGen/add_171  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n38), .Q(
        FastDivvy[3]) );
  DFCNQD1 ClockOutReg_reg ( .D(n69), .CP(FastClock), .CDN(n38), .Q(ClockOut)
         );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[3]), .QN(n58) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n41), 
        .Q(DivideFactor[5]), .QN(n48) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n67), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[4]), .QN(n53) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n68), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[1]), .QN(n65) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n66), .CP(Sample), .SDN(n41), .Q(
        DivideFactor[0]), .QN(n63) );
  INVD1 U3 ( .I(n40), .ZN(n38) );
  INVD1 U4 ( .I(n40), .ZN(n39) );
  INVD1 U5 ( .I(n41), .ZN(n40) );
  INVD1 U6 ( .I(Reset), .ZN(n41) );
  AO222D0 U7 ( .A1(N27), .A2(n42), .B1(N35), .B2(n43), .C1(DivideFactor[0]), 
        .C2(n44), .Z(n66) );
  AO222D0 U8 ( .A1(N31), .A2(n42), .B1(N39), .B2(n43), .C1(DivideFactor[4]), 
        .C2(n44), .Z(n67) );
  AO222D0 U9 ( .A1(N28), .A2(n42), .B1(N36), .B2(n43), .C1(DivideFactor[1]), 
        .C2(n44), .Z(n68) );
  CKND0 U10 ( .CLK(N54), .CN(n44) );
  AN2D0 U11 ( .A1(n45), .A2(n46), .Z(n43) );
  AN3D0 U12 ( .A1(n47), .A2(n48), .A3(n49), .Z(n42) );
  CKXOR2D0 U13 ( .A1(ClockOut), .A2(n50), .Z(n69) );
  AO22D0 U14 ( .A1(N32), .A2(n49), .B1(N40), .B2(n45), .Z(N55) );
  MUX2ND0 U15 ( .I0(n51), .I1(n52), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U16 ( .A1(AdjustFreq[1]), .A2(n46), .ZN(n52) );
  ND3D0 U17 ( .A1(n53), .A2(n48), .A3(n54), .ZN(n46) );
  ND4D0 U18 ( .A1(DivideFactor[3]), .A2(DivideFactor[2]), .A3(DivideFactor[1]), 
        .A4(DivideFactor[0]), .ZN(n54) );
  IND3D0 U19 ( .A1(AdjustFreq[1]), .B1(n48), .B2(n47), .ZN(n51) );
  CKND2D0 U20 ( .A1(DivideFactor[4]), .A2(DivideFactor[3]), .ZN(n47) );
  AO22D0 U21 ( .A1(N30), .A2(n49), .B1(N38), .B2(n45), .Z(N51) );
  AO22D0 U22 ( .A1(N29), .A2(n49), .B1(N37), .B2(n45), .Z(N49) );
  AN2D0 U23 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n45) );
  NR2D0 U24 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n49) );
  INR2D0 U25 ( .A1(N14), .B1(n50), .ZN(N21) );
  INR2D0 U26 ( .A1(N13), .B1(n50), .ZN(N20) );
  INR2D0 U27 ( .A1(N12), .B1(n50), .ZN(N19) );
  INR2D0 U28 ( .A1(N11), .B1(n50), .ZN(N18) );
  INR2D0 U29 ( .A1(N10), .B1(n50), .ZN(N17) );
  INR2D0 U30 ( .A1(N9), .B1(n50), .ZN(N16) );
  OA21D0 U31 ( .A1(FastDivvy[5]), .A2(n48), .B(n55), .Z(n50) );
  IOA22D0 U32 ( .B1(n56), .B2(n57), .A1(n48), .A2(FastDivvy[5]), .ZN(n55) );
  AOI221D0 U33 ( .A1(FastDivvy[4]), .A2(n53), .B1(FastDivvy[3]), .B2(n58), .C(
        n59), .ZN(n57) );
  AOI221D0 U34 ( .A1(DivideFactor[3]), .A2(n60), .B1(DivideFactor[2]), .B2(n61), .C(n62), .ZN(n59) );
  IAO21D0 U35 ( .A1(n61), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n62) );
  OAI32D0 U36 ( .A1(n63), .A2(FastDivvy[0]), .A3(n64), .B1(FastDivvy[1]), .B2(
        n65), .ZN(n61) );
  AN2D0 U37 ( .A1(FastDivvy[1]), .A2(n65), .Z(n64) );
  CKND0 U38 ( .CLK(FastDivvy[3]), .CN(n60) );
  NR2D0 U39 ( .A1(FastDivvy[4]), .A2(n53), .ZN(n56) );
  CKND0 U40 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U41 ( .A1(WireD[5]), .A2(n39), .ZN(WireD[0]) );
endmodule


module MultiCounter_1 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_1_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_2 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_2_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_3 ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_3_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_1_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_1_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_2_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_2_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_1_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_3_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_3_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module MultiCounter_0_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_0_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module SerEncoder_DWid32_0_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule

