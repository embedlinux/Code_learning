
module Deserializer ( ParOut, ParValid, DecoderParClk, FIFOEmpty, FIFOFull, 
        ParOutClk, SerialIn, ReadReq, SerValid, Reset );
  output [31:0] ParOut;
  input ParOutClk, SerialIn, ReadReq, SerValid, Reset;
  output ParValid, DecoderParClk, FIFOEmpty, FIFOFull;
  wire   n152, n153, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, ParValidDecode, SerialClk,
         SerRxToDecode, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n18, n20,
         n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48,
         n50, n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76,
         n78, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151;
  wire   [31:0] FIFO_Out;
  wire   [31:0] DecodeToFIFO;

  FIFOTop_AWid5_DWid32 FIFO_U1 ( .Dout(FIFO_Out), .Din(DecodeToFIFO), .Full(
        FIFOFull), .Empty(n153), .ReadIn(n148), .WriteIn(ParValidDecode), 
        .ClkR(ParOutClk), .ClkW(n7), .Reseter(n146) );
  DesDecoder_DWid32 DesDecoder_U1 ( .ParOut(DecodeToFIFO), .ParValid(
        ParValidDecode), .ParClk(n152), .SerIn(SerRxToDecode), .SerClk(
        SerialClk), .SerValid(n147), .Reset(n146) );
  SerialRx SerialRx_U1 ( .SerClk(SerialClk), .SerData(SerRxToDecode), 
        .SerLinkIn(SerialIn), .ParClk(n7), .Reset(Reset) );
  DFCND1 \ParBuf_reg[6]  ( .D(N9), .CP(ParOutClk), .CDN(n11), .QN(n120) );
  DFCND1 \ParBuf_reg[5]  ( .D(N8), .CP(ParOutClk), .CDN(n11), .QN(n119) );
  DFCND1 \ParBuf_reg[4]  ( .D(N7), .CP(ParOutClk), .CDN(n11), .QN(n118) );
  DFCND1 \ParBuf_reg[3]  ( .D(N6), .CP(ParOutClk), .CDN(n11), .QN(n117) );
  DFCND1 \ParBuf_reg[2]  ( .D(N5), .CP(ParOutClk), .CDN(n13), .QN(n116) );
  DFCND1 \ParBuf_reg[1]  ( .D(N4), .CP(ParOutClk), .CDN(n11), .QN(n115) );
  DFCND1 \ParBuf_reg[31]  ( .D(N34), .CP(ParOutClk), .CDN(n10), .QN(n145) );
  DFCND1 \ParBuf_reg[30]  ( .D(N33), .CP(ParOutClk), .CDN(n12), .QN(n144) );
  DFCND1 \ParBuf_reg[29]  ( .D(N32), .CP(ParOutClk), .CDN(n12), .QN(n143) );
  DFCND1 \ParBuf_reg[28]  ( .D(N31), .CP(ParOutClk), .CDN(n10), .QN(n142) );
  DFCND1 \ParBuf_reg[27]  ( .D(N30), .CP(ParOutClk), .CDN(n11), .QN(n141) );
  DFCND1 \ParBuf_reg[26]  ( .D(N29), .CP(ParOutClk), .CDN(n13), .QN(n140) );
  DFCND1 \ParBuf_reg[25]  ( .D(N28), .CP(ParOutClk), .CDN(n13), .QN(n139) );
  DFCND1 \ParBuf_reg[24]  ( .D(N27), .CP(ParOutClk), .CDN(n10), .QN(n138) );
  DFCND1 \ParBuf_reg[23]  ( .D(N26), .CP(ParOutClk), .CDN(n12), .QN(n137) );
  DFCND1 \ParBuf_reg[22]  ( .D(N25), .CP(ParOutClk), .CDN(n12), .QN(n136) );
  DFCND1 \ParBuf_reg[21]  ( .D(N24), .CP(ParOutClk), .CDN(n10), .QN(n135) );
  DFCND1 \ParBuf_reg[20]  ( .D(N23), .CP(ParOutClk), .CDN(n11), .QN(n134) );
  DFCND1 \ParBuf_reg[19]  ( .D(N22), .CP(ParOutClk), .CDN(n13), .QN(n133) );
  DFCND1 \ParBuf_reg[18]  ( .D(N21), .CP(ParOutClk), .CDN(n13), .QN(n132) );
  DFCND1 \ParBuf_reg[17]  ( .D(N20), .CP(ParOutClk), .CDN(n11), .QN(n131) );
  DFCND1 \ParBuf_reg[16]  ( .D(N19), .CP(ParOutClk), .CDN(n12), .QN(n130) );
  DFCND1 \ParBuf_reg[15]  ( .D(N18), .CP(ParOutClk), .CDN(n12), .QN(n129) );
  DFCND1 \ParBuf_reg[14]  ( .D(N17), .CP(ParOutClk), .CDN(n10), .QN(n128) );
  DFCND1 \ParBuf_reg[13]  ( .D(N16), .CP(ParOutClk), .CDN(n10), .QN(n127) );
  DFCND1 \ParBuf_reg[0]  ( .D(N3), .CP(ParOutClk), .CDN(n13), .QN(n114) );
  DFCND1 \ParBuf_reg[12]  ( .D(N15), .CP(ParOutClk), .CDN(n13), .QN(n126) );
  DFCND1 \ParBuf_reg[11]  ( .D(N14), .CP(ParOutClk), .CDN(n13), .QN(n125) );
  DFCND1 \ParBuf_reg[10]  ( .D(N13), .CP(ParOutClk), .CDN(n11), .QN(n124) );
  DFCND1 \ParBuf_reg[9]  ( .D(N12), .CP(ParOutClk), .CDN(n10), .QN(n123) );
  DFCND1 \ParBuf_reg[8]  ( .D(N11), .CP(ParOutClk), .CDN(n12), .QN(n122) );
  DFCND1 \ParBuf_reg[7]  ( .D(N10), .CP(ParOutClk), .CDN(n12), .QN(n121) );
  DFCND1 ParValidr_reg ( .D(N35), .CP(ParOutClk), .CDN(n10), .QN(n113) );
  INVD1 U38 ( .I(n6), .ZN(n7) );
  INVD1 U39 ( .I(n8), .ZN(n9) );
  CKNXD16 U40 ( .I(n6), .ZN(DecoderParClk) );
  CKNXD16 U41 ( .I(n8), .ZN(FIFOEmpty) );
  CKND0 U42 ( .CLK(n152), .CN(n6) );
  CKND0 U43 ( .CLK(n153), .CN(n8) );
  INVD0 U44 ( .I(Reset), .ZN(n10) );
  INVD0 U45 ( .I(Reset), .ZN(n13) );
  INVD0 U46 ( .I(Reset), .ZN(n11) );
  INVD0 U47 ( .I(Reset), .ZN(n12) );
  CKBD0 U48 ( .CLK(n145), .C(n14) );
  CKNXD16 U49 ( .I(n14), .ZN(ParOut[31]) );
  CKBD0 U50 ( .CLK(n144), .C(n16) );
  CKNXD16 U51 ( .I(n16), .ZN(ParOut[30]) );
  CKBD0 U52 ( .CLK(n143), .C(n18) );
  CKNXD16 U53 ( .I(n18), .ZN(ParOut[29]) );
  CKBD0 U54 ( .CLK(n142), .C(n20) );
  CKNXD16 U55 ( .I(n20), .ZN(ParOut[28]) );
  CKBD0 U56 ( .CLK(n141), .C(n22) );
  CKNXD16 U57 ( .I(n22), .ZN(ParOut[27]) );
  CKBD0 U58 ( .CLK(n140), .C(n24) );
  CKNXD16 U59 ( .I(n24), .ZN(ParOut[26]) );
  CKBD0 U60 ( .CLK(n139), .C(n26) );
  CKNXD16 U61 ( .I(n26), .ZN(ParOut[25]) );
  CKBD0 U62 ( .CLK(n138), .C(n28) );
  CKNXD16 U63 ( .I(n28), .ZN(ParOut[24]) );
  CKBD0 U64 ( .CLK(n137), .C(n30) );
  CKNXD16 U65 ( .I(n30), .ZN(ParOut[23]) );
  CKBD0 U66 ( .CLK(n136), .C(n32) );
  CKNXD16 U67 ( .I(n32), .ZN(ParOut[22]) );
  CKBD0 U68 ( .CLK(n135), .C(n34) );
  CKNXD16 U69 ( .I(n34), .ZN(ParOut[21]) );
  CKBD0 U70 ( .CLK(n134), .C(n36) );
  CKNXD16 U71 ( .I(n36), .ZN(ParOut[20]) );
  CKBD0 U72 ( .CLK(n133), .C(n38) );
  CKNXD16 U73 ( .I(n38), .ZN(ParOut[19]) );
  CKBD0 U74 ( .CLK(n132), .C(n40) );
  CKNXD16 U75 ( .I(n40), .ZN(ParOut[18]) );
  CKBD0 U76 ( .CLK(n131), .C(n42) );
  CKNXD16 U77 ( .I(n42), .ZN(ParOut[17]) );
  CKBD0 U78 ( .CLK(n130), .C(n44) );
  CKNXD16 U79 ( .I(n44), .ZN(ParOut[16]) );
  CKBD0 U80 ( .CLK(n129), .C(n46) );
  CKNXD16 U81 ( .I(n46), .ZN(ParOut[15]) );
  CKBD0 U82 ( .CLK(n128), .C(n48) );
  CKNXD16 U83 ( .I(n48), .ZN(ParOut[14]) );
  CKBD0 U84 ( .CLK(n127), .C(n50) );
  CKNXD16 U85 ( .I(n50), .ZN(ParOut[13]) );
  CKBD0 U86 ( .CLK(n126), .C(n52) );
  CKNXD16 U87 ( .I(n52), .ZN(ParOut[12]) );
  CKBD0 U88 ( .CLK(n125), .C(n54) );
  CKNXD16 U89 ( .I(n54), .ZN(ParOut[11]) );
  CKBD0 U90 ( .CLK(n124), .C(n56) );
  CKNXD16 U91 ( .I(n56), .ZN(ParOut[10]) );
  CKBD0 U92 ( .CLK(n123), .C(n58) );
  CKNXD16 U93 ( .I(n58), .ZN(ParOut[9]) );
  CKBD0 U94 ( .CLK(n122), .C(n60) );
  CKNXD16 U95 ( .I(n60), .ZN(ParOut[8]) );
  CKBD0 U96 ( .CLK(n121), .C(n62) );
  CKNXD16 U97 ( .I(n62), .ZN(ParOut[7]) );
  CKBD0 U98 ( .CLK(n120), .C(n64) );
  CKNXD16 U99 ( .I(n64), .ZN(ParOut[6]) );
  CKBD0 U100 ( .CLK(n119), .C(n66) );
  CKNXD16 U101 ( .I(n66), .ZN(ParOut[5]) );
  CKBD0 U102 ( .CLK(n118), .C(n68) );
  CKNXD16 U103 ( .I(n68), .ZN(ParOut[4]) );
  CKBD0 U104 ( .CLK(n117), .C(n70) );
  CKNXD16 U105 ( .I(n70), .ZN(ParOut[3]) );
  CKBD0 U106 ( .CLK(n116), .C(n72) );
  CKNXD16 U107 ( .I(n72), .ZN(ParOut[2]) );
  CKBD0 U108 ( .CLK(n115), .C(n74) );
  CKNXD16 U109 ( .I(n74), .ZN(ParOut[1]) );
  CKBD0 U110 ( .CLK(n114), .C(n76) );
  CKNXD16 U111 ( .I(n76), .ZN(ParOut[0]) );
  CKBD0 U112 ( .CLK(n113), .C(n78) );
  CKNXD16 U113 ( .I(n78), .ZN(ParValid) );
  NR2D0 U114 ( .A1(n9), .A2(n151), .ZN(N35) );
  INVD1 U115 ( .I(n151), .ZN(n148) );
  INVD1 U116 ( .I(n151), .ZN(n149) );
  INVD1 U117 ( .I(n151), .ZN(n150) );
  BUFFD1 U118 ( .I(Reset), .Z(n146) );
  AN2D1 U119 ( .A1(FIFO_Out[0]), .A2(n150), .Z(N3) );
  AN2D1 U120 ( .A1(FIFO_Out[1]), .A2(ReadReq), .Z(N4) );
  AN2D1 U121 ( .A1(FIFO_Out[2]), .A2(ReadReq), .Z(N5) );
  AN2D1 U122 ( .A1(FIFO_Out[3]), .A2(ReadReq), .Z(N6) );
  AN2D1 U123 ( .A1(FIFO_Out[4]), .A2(ReadReq), .Z(N7) );
  AN2D1 U124 ( .A1(FIFO_Out[5]), .A2(ReadReq), .Z(N8) );
  AN2D1 U125 ( .A1(FIFO_Out[6]), .A2(ReadReq), .Z(N9) );
  AN2D1 U126 ( .A1(FIFO_Out[7]), .A2(n148), .Z(N10) );
  AN2D1 U127 ( .A1(FIFO_Out[8]), .A2(n148), .Z(N11) );
  AN2D1 U128 ( .A1(FIFO_Out[9]), .A2(n148), .Z(N12) );
  AN2D1 U129 ( .A1(FIFO_Out[10]), .A2(n148), .Z(N13) );
  AN2D1 U130 ( .A1(FIFO_Out[11]), .A2(n148), .Z(N14) );
  AN2D1 U131 ( .A1(FIFO_Out[12]), .A2(n148), .Z(N15) );
  AN2D1 U132 ( .A1(FIFO_Out[13]), .A2(n149), .Z(N16) );
  AN2D1 U133 ( .A1(FIFO_Out[14]), .A2(n149), .Z(N17) );
  AN2D1 U134 ( .A1(FIFO_Out[15]), .A2(n149), .Z(N18) );
  AN2D1 U135 ( .A1(FIFO_Out[16]), .A2(n149), .Z(N19) );
  AN2D1 U136 ( .A1(FIFO_Out[17]), .A2(n149), .Z(N20) );
  AN2D1 U137 ( .A1(FIFO_Out[18]), .A2(n149), .Z(N21) );
  AN2D1 U138 ( .A1(FIFO_Out[19]), .A2(n149), .Z(N22) );
  AN2D1 U139 ( .A1(FIFO_Out[20]), .A2(n149), .Z(N23) );
  AN2D1 U140 ( .A1(FIFO_Out[21]), .A2(n149), .Z(N24) );
  AN2D1 U141 ( .A1(FIFO_Out[22]), .A2(n149), .Z(N25) );
  AN2D1 U142 ( .A1(FIFO_Out[23]), .A2(n150), .Z(N26) );
  AN2D1 U143 ( .A1(FIFO_Out[24]), .A2(n150), .Z(N27) );
  AN2D1 U144 ( .A1(FIFO_Out[25]), .A2(n150), .Z(N28) );
  AN2D1 U145 ( .A1(FIFO_Out[26]), .A2(n150), .Z(N29) );
  AN2D1 U146 ( .A1(FIFO_Out[27]), .A2(n150), .Z(N30) );
  AN2D1 U147 ( .A1(FIFO_Out[28]), .A2(n150), .Z(N31) );
  AN2D1 U148 ( .A1(FIFO_Out[29]), .A2(n150), .Z(N32) );
  AN2D1 U149 ( .A1(FIFO_Out[30]), .A2(n150), .Z(N33) );
  AN2D1 U150 ( .A1(FIFO_Out[31]), .A2(n150), .Z(N34) );
  INVD1 U151 ( .I(ReadReq), .ZN(n151) );
  BUFFD1 U152 ( .I(SerValid), .Z(n147) );
endmodule


module FIFOTop_AWid5_DWid32 ( Dout, Din, Full, Empty, ReadIn, WriteIn, ClkR, 
        ClkW, Reseter );
  output [31:0] Dout;
  input [31:0] Din;
  input ReadIn, WriteIn, ClkR, ClkW, Reseter;
  output Full, Empty;
  wire   \*Logic1* , SM_MemReadCmd, SM_MemWriteCmd, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  wire   [4:0] SM_ReadAddr;
  wire   [4:0] SM_WriteAddr;

  FIFOStateM_AWid5 FIFO_SM1 ( .ReadAddr(SM_ReadAddr), .WriteAddr(SM_WriteAddr), 
        .EmptyFIFO(Empty), .FullFIFO(Full), .ReadCmd(SM_MemReadCmd), 
        .WriteCmd(SM_MemWriteCmd), .ReadReq(ReadIn), .WriteReq(WriteIn), 
        .ClkR(ClkR), .ClkW(ClkW), .Reset(Reseter) );
  DPMem1kx32_AWid5_DWid32 FIFO_Mem1 ( .DataO(Dout), .DataI({n33, n32, n31, n30, 
        n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, n18, n17, n16, 
        n15, n14, n13, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2}), 
        .AddrR(SM_ReadAddr), .AddrW(SM_WriteAddr), .ClkR(ClkR), .ClkW(ClkW), 
        .ChipEna(\*Logic1* ), .Read(n1), .Write(SM_MemWriteCmd), .Reset(
        Reseter) );
  BUFFD1 U2 ( .I(SM_MemReadCmd), .Z(n1) );
  BUFFD1 U3 ( .I(Din[0]), .Z(n2) );
  BUFFD1 U4 ( .I(Din[1]), .Z(n3) );
  BUFFD1 U5 ( .I(Din[2]), .Z(n4) );
  BUFFD1 U6 ( .I(Din[3]), .Z(n5) );
  BUFFD1 U7 ( .I(Din[4]), .Z(n6) );
  BUFFD1 U8 ( .I(Din[5]), .Z(n7) );
  BUFFD1 U9 ( .I(Din[6]), .Z(n8) );
  BUFFD1 U10 ( .I(Din[7]), .Z(n9) );
  BUFFD1 U11 ( .I(Din[8]), .Z(n10) );
  BUFFD1 U12 ( .I(Din[9]), .Z(n11) );
  BUFFD1 U13 ( .I(Din[10]), .Z(n12) );
  BUFFD1 U14 ( .I(Din[11]), .Z(n13) );
  BUFFD1 U15 ( .I(Din[12]), .Z(n14) );
  BUFFD1 U16 ( .I(Din[13]), .Z(n15) );
  BUFFD1 U17 ( .I(Din[14]), .Z(n16) );
  BUFFD1 U18 ( .I(Din[15]), .Z(n17) );
  BUFFD1 U19 ( .I(Din[16]), .Z(n18) );
  BUFFD1 U20 ( .I(Din[17]), .Z(n19) );
  BUFFD1 U21 ( .I(Din[18]), .Z(n20) );
  BUFFD1 U22 ( .I(Din[19]), .Z(n21) );
  BUFFD1 U23 ( .I(Din[20]), .Z(n22) );
  BUFFD1 U24 ( .I(Din[21]), .Z(n23) );
  BUFFD1 U25 ( .I(Din[22]), .Z(n24) );
  BUFFD1 U26 ( .I(Din[23]), .Z(n25) );
  BUFFD1 U27 ( .I(Din[24]), .Z(n26) );
  BUFFD1 U28 ( .I(Din[25]), .Z(n27) );
  BUFFD1 U29 ( .I(Din[26]), .Z(n28) );
  BUFFD1 U30 ( .I(Din[27]), .Z(n29) );
  BUFFD1 U31 ( .I(Din[28]), .Z(n30) );
  BUFFD1 U32 ( .I(Din[29]), .Z(n31) );
  BUFFD1 U33 ( .I(Din[30]), .Z(n32) );
  BUFFD1 U34 ( .I(Din[31]), .Z(n33) );
  TIEH U35 ( .Z(\*Logic1* ) );
endmodule


module DesDecoder_DWid32 ( ParOut, ParValid, ParClk, SerIn, SerClk, SerValid, 
        Reset );
  output [31:0] ParOut;
  input SerIn, SerClk, SerValid, Reset;
  output ParValid, ParClk;
  wire   UnLoad, N12, N44, N49, N50, N51, N52, N53, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, n2, n3, n38, n39, n40, n41, n42, n43, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n136, n137, n138, n151, n152, n153, n165, n166, n167, n168, n179,
         n180, n181, n182, n183, n184, n185, n186, n254, n255, n256, n257,
         n258, n259, n260;
  wire   [63:0] FrameSR;
  wire   [4:0] Count32;

  LHD1 SerClock_reg ( .E(N69), .D(N64), .Q(n252) );
  LHQD1 \Count32_reg[0]  ( .E(N69), .D(N65), .Q(Count32[0]) );
  LHQD1 \Count32_reg[1]  ( .E(N69), .D(N66), .Q(Count32[1]) );
  LHQD1 \Count32_reg[2]  ( .E(N69), .D(N67), .Q(Count32[2]) );
  LHQD1 \Count32_reg[3]  ( .E(N69), .D(N68), .Q(Count32[3]) );
  LHQD1 \Count32_reg[4]  ( .E(N69), .D(N70), .Q(Count32[4]) );
  LHQD1 ParClkReg_reg ( .E(N62), .D(N63), .Q(ParClk) );
  DesDecoder_DWid32_DW01_inc_0 \SerClockGen/add_170_C252_S2  ( .A(Count32), 
        .SUM({N53, N52, N51, N50, N49}) );
  DFNCND1 \FrameSR_reg[63]  ( .D(FrameSR[62]), .CPN(n122), .CDN(n114), .QN(
        n123) );
  DFNCND1 doParSync_reg ( .D(N12), .CPN(n179), .CDN(n108), .Q(n36), .QN(n2) );
  DFNCND1 \FrameSR_reg[8]  ( .D(FrameSR[7]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[8]), .QN(n178) );
  DFNCND1 \FrameSR_reg[9]  ( .D(FrameSR[8]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[9]), .QN(n177) );
  DFNCND1 \FrameSR_reg[10]  ( .D(FrameSR[9]), .CPN(n166), .CDN(n110), .Q(
        FrameSR[10]), .QN(n176) );
  DFNCND1 \FrameSR_reg[11]  ( .D(FrameSR[10]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[11]), .QN(n175) );
  DFNCND1 \FrameSR_reg[12]  ( .D(FrameSR[11]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[12]), .QN(n174) );
  DFNCND1 \FrameSR_reg[13]  ( .D(FrameSR[12]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[13]), .QN(n173) );
  DFNCND1 \FrameSR_reg[14]  ( .D(FrameSR[13]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[14]), .QN(n172) );
  DFNCND1 \FrameSR_reg[15]  ( .D(FrameSR[14]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[15]), .QN(n171) );
  DFNCND1 \FrameSR_reg[16]  ( .D(FrameSR[15]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[16]), .QN(n170) );
  DFNCND1 \FrameSR_reg[17]  ( .D(FrameSR[16]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[17]), .QN(n169) );
  DFNCND1 \FrameSR_reg[22]  ( .D(FrameSR[21]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[22]), .QN(n164) );
  DFNCND1 \FrameSR_reg[23]  ( .D(FrameSR[22]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[23]), .QN(n163) );
  DFNCND1 \FrameSR_reg[24]  ( .D(FrameSR[23]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[24]), .QN(n162) );
  DFNCND1 \FrameSR_reg[25]  ( .D(FrameSR[24]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[25]), .QN(n161) );
  DFNCND1 \FrameSR_reg[26]  ( .D(FrameSR[25]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[26]), .QN(n160) );
  DFNCND1 \FrameSR_reg[27]  ( .D(FrameSR[26]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[27]), .QN(n159) );
  DFNCND1 \FrameSR_reg[28]  ( .D(FrameSR[27]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[28]), .QN(n158) );
  DFNCND1 \FrameSR_reg[29]  ( .D(FrameSR[28]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[29]), .QN(n157) );
  DFNCND1 \FrameSR_reg[30]  ( .D(FrameSR[29]), .CPN(n153), .CDN(n112), .Q(
        FrameSR[30]), .QN(n156) );
  DFNCND1 \FrameSR_reg[31]  ( .D(FrameSR[30]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[31]), .QN(n155) );
  DFNCND1 \FrameSR_reg[32]  ( .D(FrameSR[31]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[32]), .QN(n154) );
  DFNCND1 \FrameSR_reg[36]  ( .D(FrameSR[35]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[36]), .QN(n150) );
  DFNCND1 \FrameSR_reg[37]  ( .D(FrameSR[36]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[37]), .QN(n149) );
  DFNCND1 \FrameSR_reg[38]  ( .D(FrameSR[37]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[38]), .QN(n148) );
  DFNCND1 \FrameSR_reg[39]  ( .D(FrameSR[38]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[39]), .QN(n147) );
  DFNCND1 \FrameSR_reg[40]  ( .D(FrameSR[39]), .CPN(n152), .CDN(n113), .Q(
        FrameSR[40]), .QN(n146) );
  DFNCND1 \FrameSR_reg[41]  ( .D(FrameSR[40]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[41]), .QN(n145) );
  DFNCND1 \FrameSR_reg[42]  ( .D(FrameSR[41]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[42]), .QN(n144) );
  DFNCND1 \FrameSR_reg[43]  ( .D(FrameSR[42]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[43]), .QN(n143) );
  DFNCND1 \FrameSR_reg[44]  ( .D(FrameSR[43]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[44]), .QN(n142) );
  DFNCND1 \FrameSR_reg[45]  ( .D(FrameSR[44]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[45]), .QN(n141) );
  DFNCND1 \FrameSR_reg[46]  ( .D(FrameSR[45]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[46]), .QN(n140) );
  DFNCND1 \FrameSR_reg[47]  ( .D(FrameSR[46]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[47]), .QN(n139) );
  DFNCND1 \FrameSR_reg[51]  ( .D(FrameSR[50]), .CPN(n252), .CDN(n118), .Q(
        FrameSR[51]), .QN(n135) );
  DFNCND1 \FrameSR_reg[52]  ( .D(FrameSR[51]), .CPN(n167), .CDN(n119), .Q(
        FrameSR[52]), .QN(n134) );
  DFNCND1 \FrameSR_reg[53]  ( .D(FrameSR[52]), .CPN(n180), .CDN(n118), .Q(
        FrameSR[53]), .QN(n133) );
  DFNCND1 \FrameSR_reg[54]  ( .D(FrameSR[53]), .CPN(n121), .CDN(n108), .Q(
        FrameSR[54]), .QN(n132) );
  DFNCND1 \FrameSR_reg[55]  ( .D(FrameSR[54]), .CPN(n167), .CDN(n107), .Q(
        FrameSR[55]), .QN(n131) );
  DFNCND1 \FrameSR_reg[56]  ( .D(FrameSR[55]), .CPN(n168), .CDN(n116), .Q(
        FrameSR[56]), .QN(n130) );
  DFNCND1 \FrameSR_reg[57]  ( .D(FrameSR[56]), .CPN(n167), .CDN(n253), .Q(
        FrameSR[57]), .QN(n129) );
  DFNCND1 \FrameSR_reg[58]  ( .D(FrameSR[57]), .CPN(n179), .CDN(n120), .Q(
        FrameSR[58]), .QN(n128) );
  DFNCND1 \FrameSR_reg[59]  ( .D(FrameSR[58]), .CPN(n121), .CDN(n119), .Q(
        FrameSR[59]), .QN(n127) );
  DFNCND1 \FrameSR_reg[60]  ( .D(FrameSR[59]), .CPN(n122), .CDN(n114), .Q(
        FrameSR[60]), .QN(n126) );
  DFNCND1 \FrameSR_reg[61]  ( .D(FrameSR[60]), .CPN(n252), .CDN(n114), .Q(
        FrameSR[61]), .QN(n125) );
  DFNCND1 \FrameSR_reg[62]  ( .D(FrameSR[61]), .CPN(n136), .CDN(n114), .Q(
        FrameSR[62]), .QN(n124) );
  DFNCND1 \DecodeReg_reg[31]  ( .D(n251), .CPN(n180), .CDN(n114), .QN(n4) );
  DFNCND1 \DecodeReg_reg[30]  ( .D(n250), .CPN(n121), .CDN(n114), .QN(n35) );
  DFNCND1 \DecodeReg_reg[29]  ( .D(n249), .CPN(n167), .CDN(n114), .QN(n34) );
  DFNCND1 \DecodeReg_reg[28]  ( .D(n248), .CPN(n168), .CDN(n114), .QN(n33) );
  DFNCND1 \DecodeReg_reg[27]  ( .D(n247), .CPN(n168), .CDN(n114), .QN(n32) );
  DFNCND1 \DecodeReg_reg[26]  ( .D(n246), .CPN(n179), .CDN(n115), .QN(n31) );
  DFNCND1 \DecodeReg_reg[25]  ( .D(n245), .CPN(n136), .CDN(n115), .QN(n30) );
  DFNCND1 \DecodeReg_reg[24]  ( .D(n244), .CPN(n179), .CDN(n115), .QN(n29) );
  DFNCND1 \DecodeReg_reg[23]  ( .D(n243), .CPN(n122), .CDN(n115), .QN(n28) );
  DFNCND1 \DecodeReg_reg[22]  ( .D(n242), .CPN(n252), .CDN(n115), .QN(n27) );
  DFNCND1 \DecodeReg_reg[21]  ( .D(n241), .CPN(n136), .CDN(n115), .QN(n26) );
  DFNCND1 \DecodeReg_reg[20]  ( .D(n240), .CPN(n180), .CDN(n115), .QN(n25) );
  DFNCND1 \DecodeReg_reg[19]  ( .D(n239), .CPN(n121), .CDN(n115), .QN(n24) );
  DFNCND1 \DecodeReg_reg[18]  ( .D(n238), .CPN(n168), .CDN(n115), .QN(n23) );
  DFNCND1 \DecodeReg_reg[17]  ( .D(n237), .CPN(n167), .CDN(n115), .QN(n22) );
  DFNCND1 \DecodeReg_reg[16]  ( .D(n236), .CPN(n121), .CDN(n108), .QN(n21) );
  DFNCND1 \DecodeReg_reg[15]  ( .D(n235), .CPN(n179), .CDN(n108), .QN(n20) );
  DFNCND1 \DecodeReg_reg[14]  ( .D(n234), .CPN(n122), .CDN(n107), .QN(n19) );
  DFNCND1 \DecodeReg_reg[13]  ( .D(n233), .CPN(n180), .CDN(n107), .QN(n18) );
  DFNCND1 \DecodeReg_reg[12]  ( .D(n232), .CPN(n122), .CDN(n119), .QN(n17) );
  DFNCND1 \DecodeReg_reg[11]  ( .D(n231), .CPN(n180), .CDN(n116), .QN(n16) );
  DFNCND1 \DecodeReg_reg[10]  ( .D(n230), .CPN(n167), .CDN(n253), .QN(n15) );
  DFNCND1 \DecodeReg_reg[9]  ( .D(n229), .CPN(n168), .CDN(n120), .QN(n14) );
  DFNCND1 \DecodeReg_reg[8]  ( .D(n228), .CPN(n179), .CDN(n118), .QN(n13) );
  DFNCND1 \DecodeReg_reg[7]  ( .D(n227), .CPN(n136), .CDN(n117), .QN(n12) );
  DFNCND1 \DecodeReg_reg[6]  ( .D(n226), .CPN(n252), .CDN(n119), .QN(n11) );
  DFNCND1 \DecodeReg_reg[5]  ( .D(n225), .CPN(n121), .CDN(n107), .QN(n10) );
  DFNCND1 \DecodeReg_reg[4]  ( .D(n224), .CPN(n179), .CDN(n118), .QN(n9) );
  DFNCND1 \DecodeReg_reg[3]  ( .D(n223), .CPN(n136), .CDN(n119), .QN(n8) );
  DFNCND1 \DecodeReg_reg[2]  ( .D(n222), .CPN(n122), .CDN(n116), .QN(n7) );
  DFNCND1 \DecodeReg_reg[1]  ( .D(n221), .CPN(n121), .CDN(n253), .QN(n6) );
  DFNCND1 \DecodeReg_reg[0]  ( .D(n220), .CPN(n167), .CDN(n120), .QN(n5) );
  DFNCND1 \FrameSR_reg[0]  ( .D(SerIn), .CPN(n136), .CDN(n114), .Q(FrameSR[0])
         );
  DFNCND1 \FrameSR_reg[4]  ( .D(FrameSR[3]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[4]) );
  DFNCND1 \FrameSR_reg[20]  ( .D(FrameSR[19]), .CPN(n165), .CDN(n111), .Q(
        FrameSR[20]) );
  DFNCND1 \FrameSR_reg[34]  ( .D(FrameSR[33]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[34]) );
  DFNCND1 \FrameSR_reg[49]  ( .D(FrameSR[48]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[49]) );
  DFNCND1 \FrameSR_reg[2]  ( .D(FrameSR[1]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[2]) );
  DFNCND1 \FrameSR_reg[6]  ( .D(FrameSR[5]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[6]) );
  DFNCND1 \FrameSR_reg[18]  ( .D(FrameSR[17]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[18]) );
  DFNCND1 \FrameSR_reg[33]  ( .D(FrameSR[32]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[33]) );
  DFNCND1 \FrameSR_reg[48]  ( .D(FrameSR[47]), .CPN(n151), .CDN(n113), .Q(
        FrameSR[48]) );
  DFNCND1 \FrameSR_reg[1]  ( .D(FrameSR[0]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[1]) );
  DFNCND1 \FrameSR_reg[3]  ( .D(FrameSR[2]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[3]) );
  DFNCND1 \FrameSR_reg[5]  ( .D(FrameSR[4]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[5]) );
  DFNCND1 \FrameSR_reg[7]  ( .D(FrameSR[6]), .CPN(n166), .CDN(n109), .Q(
        FrameSR[7]) );
  DFNCND1 \FrameSR_reg[21]  ( .D(FrameSR[20]), .CPN(n153), .CDN(n111), .Q(
        FrameSR[21]) );
  DFNCND1 \FrameSR_reg[35]  ( .D(FrameSR[34]), .CPN(n152), .CDN(n112), .Q(
        FrameSR[35]) );
  DFNCND1 \FrameSR_reg[50]  ( .D(FrameSR[49]), .CPN(n151), .CDN(n117), .Q(
        FrameSR[50]) );
  DFNCND1 \FrameSR_reg[19]  ( .D(FrameSR[18]), .CPN(n165), .CDN(n110), .Q(
        FrameSR[19]) );
  DFNCND1 UnLoad_reg ( .D(N44), .CPN(n168), .CDN(n118), .Q(UnLoad), .QN(n1) );
  DFNCND1 ParValidReg_reg ( .D(n187), .CPN(n137), .CDN(n116), .Q(ParValid), 
        .QN(n57) );
  DFNCND1 \ParOutReg_reg[0]  ( .D(n219), .CPN(n180), .CDN(n117), .Q(ParOut[0]), 
        .QN(n89) );
  DFNCND1 \ParOutReg_reg[1]  ( .D(n218), .CPN(n122), .CDN(n253), .Q(ParOut[1]), 
        .QN(n88) );
  DFNCND1 \ParOutReg_reg[2]  ( .D(n217), .CPN(n179), .CDN(n116), .Q(ParOut[2]), 
        .QN(n87) );
  DFNCND1 \ParOutReg_reg[3]  ( .D(n216), .CPN(n180), .CDN(n253), .Q(ParOut[3]), 
        .QN(n86) );
  DFNCND1 \ParOutReg_reg[4]  ( .D(n215), .CPN(n252), .CDN(n253), .Q(ParOut[4]), 
        .QN(n85) );
  DFNCND1 \ParOutReg_reg[5]  ( .D(n214), .CPN(n179), .CDN(n118), .Q(ParOut[5]), 
        .QN(n84) );
  DFNCND1 \ParOutReg_reg[6]  ( .D(n213), .CPN(n136), .CDN(n108), .Q(ParOut[6]), 
        .QN(n83) );
  DFNCND1 \ParOutReg_reg[7]  ( .D(n212), .CPN(n122), .CDN(n120), .Q(ParOut[7]), 
        .QN(n82) );
  DFNCND1 \ParOutReg_reg[8]  ( .D(n211), .CPN(n252), .CDN(n107), .Q(ParOut[8]), 
        .QN(n81) );
  DFNCND1 \ParOutReg_reg[9]  ( .D(n210), .CPN(n168), .CDN(n117), .Q(ParOut[9]), 
        .QN(n80) );
  DFNCND1 \ParOutReg_reg[10]  ( .D(n209), .CPN(n167), .CDN(n119), .Q(
        ParOut[10]), .QN(n79) );
  DFNCND1 \ParOutReg_reg[11]  ( .D(n208), .CPN(n180), .CDN(n116), .Q(
        ParOut[11]), .QN(n78) );
  DFNCND1 \ParOutReg_reg[12]  ( .D(n207), .CPN(n168), .CDN(n253), .Q(
        ParOut[12]), .QN(n77) );
  DFNCND1 \ParOutReg_reg[13]  ( .D(n206), .CPN(n138), .CDN(n120), .Q(
        ParOut[13]), .QN(n76) );
  DFNCND1 \ParOutReg_reg[14]  ( .D(n205), .CPN(n138), .CDN(n117), .Q(
        ParOut[14]), .QN(n75) );
  DFNCND1 \ParOutReg_reg[15]  ( .D(n204), .CPN(n138), .CDN(n118), .Q(
        ParOut[15]), .QN(n74) );
  DFNCND1 \ParOutReg_reg[16]  ( .D(n203), .CPN(n138), .CDN(n108), .Q(
        ParOut[16]), .QN(n73) );
  DFNCND1 \ParOutReg_reg[17]  ( .D(n202), .CPN(n138), .CDN(n107), .Q(
        ParOut[17]), .QN(n72) );
  DFNCND1 \ParOutReg_reg[18]  ( .D(n201), .CPN(n138), .CDN(n117), .Q(
        ParOut[18]), .QN(n71) );
  DFNCND1 \ParOutReg_reg[19]  ( .D(n200), .CPN(n138), .CDN(n117), .Q(
        ParOut[19]), .QN(n70) );
  DFNCND1 \ParOutReg_reg[20]  ( .D(n199), .CPN(n138), .CDN(n119), .Q(
        ParOut[20]), .QN(n69) );
  DFNCND1 \ParOutReg_reg[21]  ( .D(n198), .CPN(n138), .CDN(n253), .Q(
        ParOut[21]), .QN(n68) );
  DFNCND1 \ParOutReg_reg[22]  ( .D(n197), .CPN(n138), .CDN(n108), .Q(
        ParOut[22]), .QN(n67) );
  DFNCND1 \ParOutReg_reg[23]  ( .D(n196), .CPN(n137), .CDN(n120), .Q(
        ParOut[23]), .QN(n66) );
  DFNCND1 \ParOutReg_reg[24]  ( .D(n195), .CPN(n137), .CDN(n120), .Q(
        ParOut[24]), .QN(n65) );
  DFNCND1 \ParOutReg_reg[25]  ( .D(n194), .CPN(n137), .CDN(n117), .Q(
        ParOut[25]), .QN(n64) );
  DFNCND1 \ParOutReg_reg[26]  ( .D(n193), .CPN(n137), .CDN(n119), .Q(
        ParOut[26]), .QN(n63) );
  DFNCND1 \ParOutReg_reg[27]  ( .D(n192), .CPN(n137), .CDN(n118), .Q(
        ParOut[27]), .QN(n62) );
  DFNCND1 \ParOutReg_reg[28]  ( .D(n191), .CPN(n137), .CDN(n120), .Q(
        ParOut[28]), .QN(n61) );
  DFNCND1 \ParOutReg_reg[29]  ( .D(n190), .CPN(n137), .CDN(n118), .Q(
        ParOut[29]), .QN(n60) );
  DFNCND1 \ParOutReg_reg[30]  ( .D(n189), .CPN(n137), .CDN(n108), .Q(
        ParOut[30]), .QN(n59) );
  DFNCND1 \ParOutReg_reg[31]  ( .D(n188), .CPN(n137), .CDN(n116), .Q(
        ParOut[31]), .QN(n58) );
  BUFFD1 U3 ( .I(n117), .Z(n115) );
  BUFFD1 U4 ( .I(n118), .Z(n113) );
  BUFFD1 U5 ( .I(n119), .Z(n112) );
  BUFFD1 U6 ( .I(n119), .Z(n111) );
  BUFFD1 U7 ( .I(n117), .Z(n114) );
  BUFFD1 U8 ( .I(n107), .Z(n116) );
  INVD1 U9 ( .I(n186), .ZN(n181) );
  INVD1 U10 ( .I(n185), .ZN(n182) );
  INVD1 U11 ( .I(n254), .ZN(n183) );
  BUFFD1 U12 ( .I(n254), .Z(n185) );
  BUFFD1 U13 ( .I(n254), .Z(n186) );
  BUFFD1 U14 ( .I(n120), .Z(n110) );
  BUFFD1 U15 ( .I(n120), .Z(n109) );
  BUFFD1 U16 ( .I(n107), .Z(n118) );
  BUFFD1 U17 ( .I(n107), .Z(n119) );
  BUFFD1 U18 ( .I(n107), .Z(n117) );
  ND2D1 U19 ( .A1(n39), .A2(n116), .ZN(N69) );
  BUFFD1 U20 ( .I(n254), .Z(n184) );
  INVD1 U21 ( .I(N44), .ZN(n254) );
  BUFFD1 U22 ( .I(n253), .Z(n107) );
  BUFFD1 U23 ( .I(n108), .Z(n120) );
  BUFFD1 U24 ( .I(n253), .Z(n108) );
  BUFFD1 U25 ( .I(n168), .Z(n151) );
  BUFFD1 U26 ( .I(n168), .Z(n152) );
  BUFFD1 U27 ( .I(n167), .Z(n153) );
  BUFFD1 U28 ( .I(n167), .Z(n165) );
  BUFFD1 U29 ( .I(n136), .Z(n166) );
  INVD1 U30 ( .I(n260), .ZN(n256) );
  INVD1 U31 ( .I(n259), .ZN(n257) );
  INVD1 U32 ( .I(UnLoad), .ZN(n258) );
  INVD1 U33 ( .I(Reset), .ZN(n253) );
  INR2D1 U34 ( .A1(N53), .B1(n38), .ZN(N70) );
  INR2D1 U35 ( .A1(N52), .B1(n38), .ZN(N68) );
  INR2D1 U36 ( .A1(N51), .B1(n38), .ZN(N67) );
  INVD1 U37 ( .I(N50), .ZN(n40) );
  BUFFD1 U38 ( .I(n255), .Z(n259) );
  BUFFD1 U39 ( .I(n255), .Z(n260) );
  NR2D1 U40 ( .A1(n38), .A2(n40), .ZN(N66) );
  NR2D1 U41 ( .A1(n38), .A2(n41), .ZN(N65) );
  INVD1 U42 ( .I(SerValid), .ZN(n39) );
  INR2D1 U43 ( .A1(n45), .B1(n46), .ZN(N44) );
  NR2D1 U44 ( .A1(n45), .A2(n46), .ZN(N12) );
  BUFFD1 U45 ( .I(n180), .Z(n137) );
  BUFFD1 U46 ( .I(n180), .Z(n138) );
  BUFFD1 U47 ( .I(n122), .Z(n179) );
  BUFFD1 U48 ( .I(n121), .Z(n168) );
  BUFFD1 U49 ( .I(n121), .Z(n167) );
  ND3D1 U50 ( .A1(SerValid), .A2(n116), .A3(n2), .ZN(n38) );
  NR4D0 U51 ( .A1(n53), .A2(FrameSR[48]), .A3(FrameSR[50]), .A4(FrameSR[49]), 
        .ZN(n52) );
  ND3D1 U52 ( .A1(n132), .A2(n131), .A3(n133), .ZN(n53) );
  OAI21D1 U53 ( .A1(n3), .A2(n57), .B(n256), .ZN(n187) );
  OAI22D0 U54 ( .A1(n255), .A2(n58), .B1(n4), .B2(n256), .ZN(n188) );
  OAI22D0 U55 ( .A1(n255), .A2(n59), .B1(n256), .B2(n35), .ZN(n189) );
  OAI22D0 U56 ( .A1(n255), .A2(n60), .B1(n256), .B2(n34), .ZN(n190) );
  OAI22D0 U57 ( .A1(UnLoad), .A2(n61), .B1(n256), .B2(n33), .ZN(n191) );
  OAI22D0 U58 ( .A1(UnLoad), .A2(n62), .B1(n256), .B2(n32), .ZN(n192) );
  OAI22D0 U59 ( .A1(UnLoad), .A2(n63), .B1(n256), .B2(n31), .ZN(n193) );
  OAI22D0 U60 ( .A1(n255), .A2(n64), .B1(n256), .B2(n30), .ZN(n194) );
  OAI22D0 U61 ( .A1(n260), .A2(n65), .B1(n256), .B2(n29), .ZN(n195) );
  OAI22D0 U62 ( .A1(n255), .A2(n66), .B1(n256), .B2(n28), .ZN(n196) );
  OAI22D0 U63 ( .A1(n255), .A2(n67), .B1(n257), .B2(n27), .ZN(n197) );
  OAI22D0 U64 ( .A1(n259), .A2(n68), .B1(n257), .B2(n26), .ZN(n198) );
  OAI22D0 U65 ( .A1(UnLoad), .A2(n69), .B1(n257), .B2(n25), .ZN(n199) );
  OAI22D0 U66 ( .A1(n259), .A2(n70), .B1(n257), .B2(n24), .ZN(n200) );
  OAI22D0 U67 ( .A1(n259), .A2(n71), .B1(n257), .B2(n23), .ZN(n201) );
  OAI22D0 U68 ( .A1(n259), .A2(n72), .B1(n257), .B2(n22), .ZN(n202) );
  OAI22D0 U69 ( .A1(n259), .A2(n73), .B1(n257), .B2(n21), .ZN(n203) );
  OAI22D0 U70 ( .A1(n259), .A2(n74), .B1(n257), .B2(n20), .ZN(n204) );
  OAI22D0 U71 ( .A1(n259), .A2(n75), .B1(n257), .B2(n19), .ZN(n205) );
  OAI22D0 U72 ( .A1(n260), .A2(n76), .B1(n257), .B2(n18), .ZN(n206) );
  OAI22D0 U73 ( .A1(n260), .A2(n77), .B1(n258), .B2(n17), .ZN(n207) );
  OAI22D0 U74 ( .A1(n260), .A2(n78), .B1(n258), .B2(n16), .ZN(n208) );
  OAI22D0 U75 ( .A1(n260), .A2(n79), .B1(n258), .B2(n15), .ZN(n209) );
  OAI22D0 U76 ( .A1(n260), .A2(n80), .B1(n258), .B2(n14), .ZN(n210) );
  OAI22D0 U77 ( .A1(n260), .A2(n81), .B1(n258), .B2(n13), .ZN(n211) );
  OAI22D0 U78 ( .A1(n259), .A2(n82), .B1(n258), .B2(n12), .ZN(n212) );
  OAI22D0 U79 ( .A1(n255), .A2(n83), .B1(n258), .B2(n11), .ZN(n213) );
  OAI22D0 U80 ( .A1(UnLoad), .A2(n84), .B1(n258), .B2(n10), .ZN(n214) );
  OAI22D0 U81 ( .A1(n260), .A2(n85), .B1(n258), .B2(n9), .ZN(n215) );
  OAI22D0 U82 ( .A1(n255), .A2(n86), .B1(n258), .B2(n8), .ZN(n216) );
  OAI22D0 U83 ( .A1(UnLoad), .A2(n87), .B1(n1), .B2(n7), .ZN(n217) );
  OAI22D0 U84 ( .A1(UnLoad), .A2(n88), .B1(n1), .B2(n6), .ZN(n218) );
  OAI22D0 U85 ( .A1(n260), .A2(n89), .B1(n1), .B2(n5), .ZN(n219) );
  OAI22D0 U86 ( .A1(n184), .A2(n178), .B1(n181), .B2(n5), .ZN(n220) );
  OAI22D0 U87 ( .A1(n184), .A2(n177), .B1(n181), .B2(n6), .ZN(n221) );
  OAI22D0 U88 ( .A1(n184), .A2(n176), .B1(n181), .B2(n7), .ZN(n222) );
  OAI22D0 U89 ( .A1(n184), .A2(n175), .B1(n181), .B2(n8), .ZN(n223) );
  OAI22D0 U90 ( .A1(n184), .A2(n174), .B1(n181), .B2(n9), .ZN(n224) );
  OAI22D0 U91 ( .A1(n184), .A2(n173), .B1(n181), .B2(n10), .ZN(n225) );
  OAI22D0 U92 ( .A1(n185), .A2(n172), .B1(n181), .B2(n11), .ZN(n226) );
  OAI22D0 U93 ( .A1(n186), .A2(n171), .B1(n181), .B2(n12), .ZN(n227) );
  OAI22D0 U94 ( .A1(n254), .A2(n162), .B1(n181), .B2(n13), .ZN(n228) );
  OAI22D0 U95 ( .A1(n184), .A2(n161), .B1(n181), .B2(n14), .ZN(n229) );
  OAI22D0 U96 ( .A1(n254), .A2(n160), .B1(n182), .B2(n15), .ZN(n230) );
  OAI22D0 U97 ( .A1(n184), .A2(n159), .B1(n182), .B2(n16), .ZN(n231) );
  OAI22D0 U98 ( .A1(n185), .A2(n158), .B1(n182), .B2(n17), .ZN(n232) );
  OAI22D0 U99 ( .A1(n185), .A2(n157), .B1(n182), .B2(n18), .ZN(n233) );
  OAI22D0 U100 ( .A1(n185), .A2(n156), .B1(n182), .B2(n19), .ZN(n234) );
  OAI22D0 U101 ( .A1(n185), .A2(n155), .B1(n182), .B2(n20), .ZN(n235) );
  OAI22D0 U102 ( .A1(n185), .A2(n146), .B1(n182), .B2(n21), .ZN(n236) );
  OAI22D0 U103 ( .A1(n185), .A2(n145), .B1(n182), .B2(n22), .ZN(n237) );
  OAI22D0 U104 ( .A1(n186), .A2(n144), .B1(n182), .B2(n23), .ZN(n238) );
  OAI22D0 U105 ( .A1(n186), .A2(n143), .B1(n182), .B2(n24), .ZN(n239) );
  OAI22D0 U106 ( .A1(n186), .A2(n142), .B1(n183), .B2(n25), .ZN(n240) );
  OAI22D0 U107 ( .A1(n186), .A2(n141), .B1(n183), .B2(n26), .ZN(n241) );
  OAI22D0 U108 ( .A1(n186), .A2(n140), .B1(n183), .B2(n27), .ZN(n242) );
  OAI22D0 U109 ( .A1(n186), .A2(n139), .B1(n183), .B2(n28), .ZN(n243) );
  OAI22D0 U110 ( .A1(n184), .A2(n130), .B1(n183), .B2(n29), .ZN(n244) );
  OAI22D0 U111 ( .A1(n254), .A2(n129), .B1(n183), .B2(n30), .ZN(n245) );
  OAI22D0 U112 ( .A1(n185), .A2(n128), .B1(n183), .B2(n31), .ZN(n246) );
  OAI22D0 U113 ( .A1(n186), .A2(n127), .B1(n183), .B2(n32), .ZN(n247) );
  OAI22D0 U114 ( .A1(n184), .A2(n126), .B1(n183), .B2(n33), .ZN(n248) );
  OAI22D0 U115 ( .A1(n254), .A2(n125), .B1(n183), .B2(n34), .ZN(n249) );
  OAI22D0 U116 ( .A1(n254), .A2(n124), .B1(N44), .B2(n35), .ZN(n250) );
  OAI22D0 U117 ( .A1(n186), .A2(n123), .B1(N44), .B2(n4), .ZN(n251) );
  ND2D1 U118 ( .A1(n47), .A2(n48), .ZN(n46) );
  NR4D0 U119 ( .A1(FrameSR[3]), .A2(FrameSR[2]), .A3(FrameSR[1]), .A4(
        FrameSR[0]), .ZN(n47) );
  NR4D0 U120 ( .A1(FrameSR[7]), .A2(FrameSR[6]), .A3(FrameSR[5]), .A4(
        FrameSR[4]), .ZN(n48) );
  INVD1 U121 ( .I(N49), .ZN(n41) );
  OAI21D1 U122 ( .A1(n42), .A2(n39), .B(n109), .ZN(N62) );
  AOI31D0 U123 ( .A1(n41), .A2(n40), .A3(n43), .B(n36), .ZN(n42) );
  NR3D0 U124 ( .A1(N51), .A2(N53), .A3(N52), .ZN(n43) );
  AN4D1 U125 ( .A1(n49), .A2(n50), .A3(n51), .A4(n52), .Z(n45) );
  NR4D0 U126 ( .A1(n56), .A2(n134), .A3(n150), .A4(n135), .ZN(n49) );
  NR4D0 U127 ( .A1(n55), .A2(FrameSR[18]), .A3(FrameSR[21]), .A4(FrameSR[20]), 
        .ZN(n50) );
  NR4D0 U128 ( .A1(n54), .A2(FrameSR[33]), .A3(FrameSR[35]), .A4(FrameSR[34]), 
        .ZN(n51) );
  NR2D1 U129 ( .A1(ParClk), .A2(n38), .ZN(N63) );
  ND3D1 U130 ( .A1(n170), .A2(n169), .A3(FrameSR[19]), .ZN(n56) );
  ND3D1 U131 ( .A1(n148), .A2(n147), .A3(n149), .ZN(n54) );
  ND3D1 U132 ( .A1(n163), .A2(n154), .A3(n164), .ZN(n55) );
  BUFFD1 U133 ( .I(n252), .Z(n122) );
  BUFFD1 U134 ( .I(n252), .Z(n121) );
  BUFFD1 U135 ( .I(UnLoad), .Z(n255) );
  BUFFD1 U136 ( .I(n136), .Z(n180) );
  BUFFD1 U137 ( .I(n252), .Z(n136) );
  AN3D1 U138 ( .A1(SerClk), .A2(n116), .A3(SerValid), .Z(N64) );
  CKND0 U139 ( .CLK(ParClk), .CN(n3) );
endmodule


module SerialRx ( SerClk, SerData, SerLinkIn, ParClk, Reset );
  input SerLinkIn, ParClk, Reset;
  output SerClk, SerData;
  wire   n1;

  PLLTop PLL_RxU1 ( .ClockOut(SerClk), .ClockIn(n1), .Reset(Reset) );
  BUFFD0 U1 ( .I(ParClk), .Z(n1) );
  BUFFD1 U2 ( .I(SerLinkIn), .Z(SerData) );
endmodule


module FIFOStateM_AWid5 ( ReadAddr, WriteAddr, EmptyFIFO, FullFIFO, ReadCmd, 
        WriteCmd, ReadReq, WriteReq, ClkR, ClkW, Reset );
  output [4:0] ReadAddr;
  output [4:0] WriteAddr;
  input ReadReq, WriteReq, ClkR, ClkW, Reset;
  output EmptyFIFO, FullFIFO, ReadCmd, WriteCmd;
  wire   n155, StateClockRaw, StateClock, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N169, N171, N172, N173, N321, N323, N324, N325, n73, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, \add_389/carry[2] , \add_389/carry[3] ,
         \add_389/carry[4] , \add_308/carry[2] , \add_308/carry[3] ,
         \add_308/carry[4] , n3, n4, n6, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n74, n86, n88, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154;
  wire   [2:0] CurState;
  wire   [2:0] NextState;
  assign ReadAddr[0] = N169;
  assign WriteAddr[0] = N321;
  assign WriteAddr[1] = \add_389/carry[2] ;
  assign ReadAddr[1] = \add_308/carry[2] ;

  DEL005 SM_DeGlitcher1 ( .I(StateClockRaw), .Z(StateClock) );
  DFND1 FullFIFOr_reg ( .D(n93), .CPN(StateClock), .Q(n155), .QN(n76) );
  FIFOStateM_AWid5_DW01_inc_0 r151 ( .A({WriteAddr[4:2], n20, n6}), .SUM({N70, 
        N69, N68, N67, N66}) );
  FIFOStateM_AWid5_DW01_inc_1 r150 ( .A({ReadAddr[4:2], \add_308/carry[2] , 
        N169}), .SUM({N47, N46, N45, N44, N43}) );
  DFNCND1 \OldReadAr_reg[0]  ( .D(n107), .CPN(StateClock), .CDN(n22), .QN(n89)
         );
  DFNCND1 \OldWriteAr_reg[0]  ( .D(n104), .CPN(StateClock), .CDN(n21), .QN(n87) );
  DFNCND1 \OldWriteAr_reg[3]  ( .D(n97), .CPN(StateClock), .CDN(n21), .QN(n80)
         );
  DFNCND1 \OldReadAr_reg[3]  ( .D(n94), .CPN(StateClock), .CDN(n22), .QN(n77)
         );
  DFNCND1 \OldReadAr_reg[1]  ( .D(n92), .CPN(StateClock), .CDN(n22), .QN(n75)
         );
  DFNCND1 \OldWriteAr_reg[1]  ( .D(n90), .CPN(StateClock), .CDN(n22), .QN(n73)
         );
  DFNCND1 \OldWriteAr_reg[4]  ( .D(n99), .CPN(StateClock), .CDN(n21), .QN(n82)
         );
  DFNCND1 \OldWriteAr_reg[2]  ( .D(n98), .CPN(StateClock), .CDN(n21), .QN(n81)
         );
  DFNCND1 \OldReadAr_reg[4]  ( .D(n96), .CPN(StateClock), .CDN(n21), .QN(n79)
         );
  DFNCND1 \OldReadAr_reg[2]  ( .D(n95), .CPN(StateClock), .CDN(n22), .QN(n78)
         );
  DFNCND1 \NextState_reg[1]  ( .D(n102), .CPN(StateClock), .CDN(n21), .Q(
        NextState[1]), .QN(n85) );
  DFNCND1 \NextState_reg[2]  ( .D(n101), .CPN(StateClock), .CDN(n21), .Q(
        NextState[2]), .QN(n84) );
  DFNCND1 \NextState_reg[0]  ( .D(n100), .CPN(StateClock), .CDN(n21), .Q(
        NextState[0]), .QN(n83) );
  DFCNQD1 \CurState_reg[0]  ( .D(NextState[0]), .CP(StateClock), .CDN(n22), 
        .Q(CurState[0]) );
  DFCNQD1 \CurState_reg[2]  ( .D(NextState[2]), .CP(StateClock), .CDN(n22), 
        .Q(CurState[2]) );
  DFNCND1 ReadCmdr_reg ( .D(n105), .CPN(StateClock), .CDN(n21), .Q(ReadCmd) );
  DFCNQD1 \CurState_reg[1]  ( .D(NextState[1]), .CP(StateClock), .CDN(n22), 
        .Q(CurState[1]) );
  DFNCND1 WriteCmdr_reg ( .D(n103), .CPN(StateClock), .CDN(n21), .Q(WriteCmd)
         );
  EDFCNQD1 \ReadAr_reg[0]  ( .D(N48), .E(N52), .CP(StateClock), .CDN(n22), .Q(
        N169) );
  EDFCNQD1 \ReadAr_reg[1]  ( .D(N49), .E(N52), .CP(StateClock), .CDN(n106), 
        .Q(\add_308/carry[2] ) );
  EDFCNQD1 \ReadAr_reg[3]  ( .D(N51), .E(N52), .CP(StateClock), .CDN(n106), 
        .Q(ReadAddr[3]) );
  EDFCND1 \ReadAr_reg[4]  ( .D(N53), .E(N52), .CP(StateClock), .CDN(n106), .Q(
        ReadAddr[4]), .QN(n28) );
  EDFCND1 \ReadAr_reg[2]  ( .D(N50), .E(N52), .CP(StateClock), .CDN(n106), .Q(
        ReadAddr[2]), .QN(n26) );
  EDFCND1 \WriteAr_reg[4]  ( .D(N75), .E(N76), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[4]), .QN(n29) );
  EDFCND1 \WriteAr_reg[3]  ( .D(N74), .E(N76), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[3]), .QN(n32) );
  EDFCND1 \WriteAr_reg[2]  ( .D(N73), .E(N76), .CP(StateClock), .CDN(n106), 
        .Q(WriteAddr[2]), .QN(n31) );
  EDFCND1 \WriteAr_reg[1]  ( .D(N72), .E(N76), .CP(StateClock), .CDN(n106), 
        .Q(\add_389/carry[2] ), .QN(n3) );
  EDFCND1 \WriteAr_reg[0]  ( .D(N71), .E(N76), .CP(StateClock), .CDN(n106), 
        .Q(N321), .QN(n52) );
  DFND1 EmptyFIFOr_reg ( .D(n91), .CPN(StateClock), .Q(EmptyFIFO) );
  CKBD0 U3 ( .CLK(n19), .C(n4) );
  CKNXD16 U4 ( .I(n4), .ZN(FullFIFO) );
  INVD1 U5 ( .I(n52), .ZN(n6) );
  INVD1 U6 ( .I(N43), .ZN(n24) );
  INVD1 U7 ( .I(Reset), .ZN(n21) );
  INVD1 U8 ( .I(Reset), .ZN(n22) );
  INVD1 U9 ( .I(N169), .ZN(n23) );
  INVD1 U10 ( .I(\add_308/carry[2] ), .ZN(n25) );
  INVD1 U11 ( .I(ReadAddr[3]), .ZN(n27) );
  ND2D1 U12 ( .A1(CurState[1]), .A2(n109), .ZN(n34) );
  XNR2D1 U13 ( .A1(N321), .A2(n23), .ZN(n149) );
  BUFFD1 U14 ( .I(\add_389/carry[2] ), .Z(n20) );
  CKND0 U15 ( .CLK(n155), .CN(n19) );
  CKXOR2D0 U16 ( .A1(ReadAddr[4]), .A2(\add_308/carry[4] ), .Z(N173) );
  AN2D0 U17 ( .A1(ReadAddr[3]), .A2(\add_308/carry[3] ), .Z(\add_308/carry[4] ) );
  CKXOR2D0 U18 ( .A1(\add_308/carry[3] ), .A2(ReadAddr[3]), .Z(N172) );
  AN2D0 U19 ( .A1(ReadAddr[2]), .A2(\add_308/carry[2] ), .Z(\add_308/carry[3] ) );
  CKXOR2D0 U20 ( .A1(\add_308/carry[2] ), .A2(ReadAddr[2]), .Z(N171) );
  CKXOR2D0 U21 ( .A1(WriteAddr[4]), .A2(\add_389/carry[4] ), .Z(N325) );
  AN2D0 U22 ( .A1(WriteAddr[3]), .A2(\add_389/carry[3] ), .Z(
        \add_389/carry[4] ) );
  CKXOR2D0 U23 ( .A1(\add_389/carry[3] ), .A2(WriteAddr[3]), .Z(N324) );
  AN2D0 U24 ( .A1(WriteAddr[2]), .A2(n20), .Z(\add_389/carry[3] ) );
  CKXOR2D0 U25 ( .A1(n20), .A2(WriteAddr[2]), .Z(N323) );
  MUX2ND0 U26 ( .I0(n82), .I1(n29), .S(n30), .ZN(n99) );
  MUX2ND0 U27 ( .I0(n81), .I1(n31), .S(n30), .ZN(n98) );
  MUX2ND0 U28 ( .I0(n80), .I1(n32), .S(n30), .ZN(n97) );
  MUX2ND0 U29 ( .I0(n79), .I1(n28), .S(n33), .ZN(n96) );
  MUX2ND0 U30 ( .I0(n78), .I1(n26), .S(n33), .ZN(n95) );
  MUX2ND0 U31 ( .I0(n77), .I1(n27), .S(n33), .ZN(n94) );
  OAI32D0 U32 ( .A1(n34), .A2(Reset), .A3(ReadReq), .B1(n76), .B2(n35), .ZN(
        n93) );
  AOI21D0 U33 ( .A1(n36), .A2(n37), .B(Reset), .ZN(n35) );
  MUX2ND0 U34 ( .I0(n75), .I1(n25), .S(n33), .ZN(n92) );
  OAI31D0 U35 ( .A1(n37), .A2(WriteReq), .A3(Reset), .B(n38), .ZN(n91) );
  OAI21D0 U36 ( .A1(Reset), .A2(n39), .B(EmptyFIFO), .ZN(n38) );
  MUX2ND0 U37 ( .I0(n73), .I1(n3), .S(n30), .ZN(n90) );
  MUX2ND0 U38 ( .I0(n89), .I1(n23), .S(n33), .ZN(n107) );
  INR3D0 U39 ( .A1(ReadReq), .B1(n40), .B2(n41), .ZN(n33) );
  CKND0 U40 ( .CLK(Reset), .CN(n106) );
  MUX2ND0 U41 ( .I0(n42), .I1(n43), .S(n40), .ZN(n105) );
  NR2D0 U42 ( .A1(n44), .A2(n45), .ZN(n40) );
  CKND2D0 U43 ( .A1(n41), .A2(ReadReq), .ZN(n42) );
  AN3D0 U44 ( .A1(n46), .A2(n47), .A3(n48), .Z(n41) );
  NR3D0 U45 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n48) );
  CKXOR2D0 U46 ( .A1(n27), .A2(n77), .Z(n51) );
  CKXOR2D0 U47 ( .A1(n25), .A2(n75), .Z(n50) );
  CKXOR2D0 U48 ( .A1(n23), .A2(n89), .Z(n49) );
  CKXOR2D0 U49 ( .A1(n78), .A2(ReadAddr[2]), .Z(n47) );
  CKXOR2D0 U50 ( .A1(n79), .A2(ReadAddr[4]), .Z(n46) );
  MUX2ND0 U51 ( .I0(n87), .I1(n52), .S(n30), .ZN(n104) );
  NR3D0 U52 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n30) );
  MUX2ND0 U53 ( .I0(n56), .I1(n57), .S(n53), .ZN(n103) );
  NR2D0 U54 ( .A1(n44), .A2(n58), .ZN(n53) );
  CKND2D0 U55 ( .A1(n54), .A2(WriteReq), .ZN(n56) );
  AN3D0 U56 ( .A1(n59), .A2(n60), .A3(n61), .Z(n54) );
  NR3D0 U57 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n61) );
  CKXOR2D0 U58 ( .A1(n32), .A2(n80), .Z(n64) );
  CKXOR2D0 U59 ( .A1(n3), .A2(n73), .Z(n63) );
  CKXOR2D0 U60 ( .A1(n52), .A2(n87), .Z(n62) );
  CKXOR2D0 U61 ( .A1(n81), .A2(WriteAddr[2]), .Z(n60) );
  CKXOR2D0 U62 ( .A1(n82), .A2(WriteAddr[4]), .Z(n59) );
  MUX2ND0 U63 ( .I0(n65), .I1(n85), .S(n66), .ZN(n102) );
  NR2D0 U64 ( .A1(n58), .A2(n67), .ZN(n65) );
  MUX2ND0 U65 ( .I0(n68), .I1(n69), .S(CurState[1]), .ZN(n67) );
  OAI21D0 U66 ( .A1(n70), .A2(n71), .B(n72), .ZN(n69) );
  AOI31D0 U67 ( .A1(n74), .A2(n86), .A3(n88), .B(CurState[2]), .ZN(n72) );
  OAI21D0 U68 ( .A1(n88), .A2(n108), .B(n109), .ZN(n68) );
  CKND0 U69 ( .CLK(n110), .CN(n108) );
  AN3D0 U70 ( .A1(n111), .A2(n112), .A3(n113), .Z(n88) );
  NR3D0 U71 ( .A1(n114), .A2(n115), .A3(n116), .ZN(n113) );
  CKXOR2D0 U72 ( .A1(WriteAddr[3]), .A2(ReadAddr[3]), .Z(n116) );
  CKXOR2D0 U73 ( .A1(n20), .A2(\add_308/carry[2] ), .Z(n115) );
  CKXOR2D0 U74 ( .A1(N321), .A2(N169), .Z(n114) );
  CKXOR2D0 U75 ( .A1(ReadAddr[2]), .A2(n31), .Z(n112) );
  CKXOR2D0 U76 ( .A1(ReadAddr[4]), .A2(n29), .Z(n111) );
  MUX2ND0 U77 ( .I0(n117), .I1(n84), .S(n66), .ZN(n101) );
  AOI211D0 U78 ( .A1(n109), .A2(n110), .B(n45), .C(n118), .ZN(n117) );
  NR3D0 U79 ( .A1(n71), .A2(n119), .A3(n70), .ZN(n118) );
  ND3D0 U80 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n71) );
  NR3D0 U81 ( .A1(n123), .A2(n124), .A3(n125), .ZN(n122) );
  CKXOR2D0 U82 ( .A1(ReadAddr[3]), .A2(N69), .Z(n125) );
  CKXOR2D0 U83 ( .A1(\add_308/carry[2] ), .A2(N67), .Z(n124) );
  CKXOR2D0 U84 ( .A1(N169), .A2(N66), .Z(n123) );
  CKXOR2D0 U85 ( .A1(ReadAddr[2]), .A2(n126), .Z(n121) );
  CKXOR2D0 U86 ( .A1(ReadAddr[4]), .A2(n127), .Z(n120) );
  CKND0 U87 ( .CLK(n34), .CN(n45) );
  ND3D0 U88 ( .A1(n128), .A2(n129), .A3(n130), .ZN(n110) );
  NR3D0 U89 ( .A1(n131), .A2(n132), .A3(n133), .ZN(n130) );
  CKXOR2D0 U90 ( .A1(ReadAddr[3]), .A2(N324), .Z(n133) );
  CKXOR2D0 U91 ( .A1(\add_308/carry[2] ), .A2(n3), .Z(n132) );
  CKXOR2D0 U92 ( .A1(N169), .A2(N321), .Z(n131) );
  CKXOR2D0 U93 ( .A1(N323), .A2(n26), .Z(n129) );
  CKXOR2D0 U94 ( .A1(N325), .A2(n28), .Z(n128) );
  MUX2ND0 U95 ( .I0(n134), .I1(n83), .S(n66), .ZN(n100) );
  OA211D0 U96 ( .A1(n55), .A2(n37), .B(n135), .C(n136), .Z(n66) );
  AOI21D0 U97 ( .A1(CurState[0]), .A2(n119), .B(n44), .ZN(n136) );
  MUX2ND0 U98 ( .I0(CurState[2]), .I1(n36), .S(n119), .ZN(n44) );
  CKND0 U99 ( .CLK(CurState[1]), .CN(n119) );
  OAI21D0 U100 ( .A1(ReadReq), .A2(n86), .B(CurState[2]), .ZN(n135) );
  CKND0 U101 ( .CLK(WriteReq), .CN(n55) );
  AOI21D0 U102 ( .A1(CurState[1]), .A2(n137), .B(n109), .ZN(n134) );
  OAI21D0 U103 ( .A1(n39), .A2(n74), .B(n70), .ZN(n137) );
  OAI31D0 U104 ( .A1(n138), .A2(n139), .A3(n140), .B(CurState[0]), .ZN(n70) );
  CKXOR2D0 U105 ( .A1(WriteAddr[4]), .A2(N47), .Z(n140) );
  CKXOR2D0 U106 ( .A1(WriteAddr[2]), .A2(N45), .Z(n139) );
  ND3D0 U107 ( .A1(n141), .A2(n142), .A3(n143), .ZN(n138) );
  CKXOR2D0 U108 ( .A1(N321), .A2(n24), .Z(n143) );
  CKXOR2D0 U109 ( .A1(n20), .A2(n144), .Z(n142) );
  CKXOR2D0 U110 ( .A1(WriteAddr[3]), .A2(n145), .Z(n141) );
  ND3D0 U111 ( .A1(n146), .A2(n147), .A3(n148), .ZN(n74) );
  NR3D0 U112 ( .A1(n149), .A2(n150), .A3(n151), .ZN(n148) );
  CKXOR2D0 U113 ( .A1(WriteAddr[3]), .A2(N172), .Z(n151) );
  CKXOR2D0 U114 ( .A1(n20), .A2(n25), .Z(n150) );
  CKXOR2D0 U115 ( .A1(N171), .A2(n31), .Z(n147) );
  CKXOR2D0 U116 ( .A1(N173), .A2(n29), .Z(n146) );
  CKND2D0 U117 ( .A1(ClkW), .A2(ClkR), .ZN(StateClockRaw) );
  ND3D0 U118 ( .A1(n34), .A2(n37), .A3(n57), .ZN(N76) );
  OAI22D0 U119 ( .A1(n28), .A2(n34), .B1(n57), .B2(n127), .ZN(N75) );
  CKND0 U120 ( .CLK(N70), .CN(n127) );
  OAI22D0 U121 ( .A1(n27), .A2(n34), .B1(n57), .B2(n152), .ZN(N74) );
  CKND0 U122 ( .CLK(N69), .CN(n152) );
  OAI22D0 U123 ( .A1(n26), .A2(n34), .B1(n57), .B2(n126), .ZN(N73) );
  CKND0 U124 ( .CLK(N68), .CN(n126) );
  OAI22D0 U125 ( .A1(n25), .A2(n34), .B1(n57), .B2(n153), .ZN(N72) );
  CKND0 U126 ( .CLK(N67), .CN(n153) );
  OAI22D0 U127 ( .A1(n23), .A2(n34), .B1(n57), .B2(n154), .ZN(N71) );
  CKND0 U128 ( .CLK(N66), .CN(n154) );
  CKND2D0 U129 ( .A1(WriteCmd), .A2(n34), .ZN(n57) );
  CKND0 U130 ( .CLK(n36), .CN(n109) );
  CKND2D0 U131 ( .A1(CurState[2]), .A2(CurState[0]), .ZN(n36) );
  INR2D0 U132 ( .A1(N47), .B1(n43), .ZN(N53) );
  CKND2D0 U133 ( .A1(n37), .A2(n43), .ZN(N52) );
  NR2D0 U134 ( .A1(n43), .A2(n145), .ZN(N51) );
  CKND0 U135 ( .CLK(N46), .CN(n145) );
  INR2D0 U136 ( .A1(N45), .B1(n43), .ZN(N50) );
  NR2D0 U137 ( .A1(n43), .A2(n144), .ZN(N49) );
  CKND0 U138 ( .CLK(N44), .CN(n144) );
  NR2D0 U139 ( .A1(n43), .A2(n24), .ZN(N48) );
  CKND2D0 U140 ( .A1(ReadCmd), .A2(n37), .ZN(n43) );
  CKND0 U141 ( .CLK(n58), .CN(n37) );
  NR2D0 U142 ( .A1(n39), .A2(CurState[1]), .ZN(n58) );
  IND2D0 U143 ( .A1(CurState[2]), .B1(n86), .ZN(n39) );
  CKND0 U144 ( .CLK(CurState[0]), .CN(n86) );
endmodule


module DPMem1kx32_AWid5_DWid32 ( Dready, ParityErr, DataO, DataI, AddrR, AddrW, 
        ClkR, ClkW, ChipEna, Read, Write, Reset );
  output [31:0] DataO;
  input [31:0] DataI;
  input [4:0] AddrR;
  input [4:0] AddrW;
  input ClkR, ClkW, ChipEna, Read, Write, Reset;
  output Dready, ParityErr;
  wire   N44, N45, N46, N47, N48, ClockR, ClockW, Dreadyr, \Storage[31][32] ,
         \Storage[31][31] , \Storage[31][30] , \Storage[31][29] ,
         \Storage[31][28] , \Storage[31][27] , \Storage[31][26] ,
         \Storage[31][25] , \Storage[31][24] , \Storage[31][23] ,
         \Storage[31][22] , \Storage[31][21] , \Storage[31][20] ,
         \Storage[31][19] , \Storage[31][18] , \Storage[31][17] ,
         \Storage[31][16] , \Storage[31][15] , \Storage[31][14] ,
         \Storage[31][13] , \Storage[31][12] , \Storage[31][11] ,
         \Storage[31][10] , \Storage[31][9] , \Storage[31][8] ,
         \Storage[31][7] , \Storage[31][6] , \Storage[31][5] ,
         \Storage[31][4] , \Storage[31][3] , \Storage[31][2] ,
         \Storage[31][1] , \Storage[31][0] , \Storage[30][32] ,
         \Storage[30][31] , \Storage[30][30] , \Storage[30][29] ,
         \Storage[30][28] , \Storage[30][27] , \Storage[30][26] ,
         \Storage[30][25] , \Storage[30][24] , \Storage[30][23] ,
         \Storage[30][22] , \Storage[30][21] , \Storage[30][20] ,
         \Storage[30][19] , \Storage[30][18] , \Storage[30][17] ,
         \Storage[30][16] , \Storage[30][15] , \Storage[30][14] ,
         \Storage[30][13] , \Storage[30][12] , \Storage[30][11] ,
         \Storage[30][10] , \Storage[30][9] , \Storage[30][8] ,
         \Storage[30][7] , \Storage[30][6] , \Storage[30][5] ,
         \Storage[30][4] , \Storage[30][3] , \Storage[30][2] ,
         \Storage[30][1] , \Storage[30][0] , \Storage[29][32] ,
         \Storage[29][31] , \Storage[29][30] , \Storage[29][29] ,
         \Storage[29][28] , \Storage[29][27] , \Storage[29][26] ,
         \Storage[29][25] , \Storage[29][24] , \Storage[29][23] ,
         \Storage[29][22] , \Storage[29][21] , \Storage[29][20] ,
         \Storage[29][19] , \Storage[29][18] , \Storage[29][17] ,
         \Storage[29][16] , \Storage[29][15] , \Storage[29][14] ,
         \Storage[29][13] , \Storage[29][12] , \Storage[29][11] ,
         \Storage[29][10] , \Storage[29][9] , \Storage[29][8] ,
         \Storage[29][7] , \Storage[29][6] , \Storage[29][5] ,
         \Storage[29][4] , \Storage[29][3] , \Storage[29][2] ,
         \Storage[29][1] , \Storage[29][0] , \Storage[28][32] ,
         \Storage[28][31] , \Storage[28][30] , \Storage[28][29] ,
         \Storage[28][28] , \Storage[28][27] , \Storage[28][26] ,
         \Storage[28][25] , \Storage[28][24] , \Storage[28][23] ,
         \Storage[28][22] , \Storage[28][21] , \Storage[28][20] ,
         \Storage[28][19] , \Storage[28][18] , \Storage[28][17] ,
         \Storage[28][16] , \Storage[28][15] , \Storage[28][14] ,
         \Storage[28][13] , \Storage[28][12] , \Storage[28][11] ,
         \Storage[28][10] , \Storage[28][9] , \Storage[28][8] ,
         \Storage[28][7] , \Storage[28][6] , \Storage[28][5] ,
         \Storage[28][4] , \Storage[28][3] , \Storage[28][2] ,
         \Storage[28][1] , \Storage[28][0] , \Storage[27][32] ,
         \Storage[27][31] , \Storage[27][30] , \Storage[27][29] ,
         \Storage[27][28] , \Storage[27][27] , \Storage[27][26] ,
         \Storage[27][25] , \Storage[27][24] , \Storage[27][23] ,
         \Storage[27][22] , \Storage[27][21] , \Storage[27][20] ,
         \Storage[27][19] , \Storage[27][18] , \Storage[27][17] ,
         \Storage[27][16] , \Storage[27][15] , \Storage[27][14] ,
         \Storage[27][13] , \Storage[27][12] , \Storage[27][11] ,
         \Storage[27][10] , \Storage[27][9] , \Storage[27][8] ,
         \Storage[27][7] , \Storage[27][6] , \Storage[27][5] ,
         \Storage[27][4] , \Storage[27][3] , \Storage[27][2] ,
         \Storage[27][1] , \Storage[27][0] , \Storage[26][32] ,
         \Storage[26][31] , \Storage[26][30] , \Storage[26][29] ,
         \Storage[26][28] , \Storage[26][27] , \Storage[26][26] ,
         \Storage[26][25] , \Storage[26][24] , \Storage[26][23] ,
         \Storage[26][22] , \Storage[26][21] , \Storage[26][20] ,
         \Storage[26][19] , \Storage[26][18] , \Storage[26][17] ,
         \Storage[26][16] , \Storage[26][15] , \Storage[26][14] ,
         \Storage[26][13] , \Storage[26][12] , \Storage[26][11] ,
         \Storage[26][10] , \Storage[26][9] , \Storage[26][8] ,
         \Storage[26][7] , \Storage[26][6] , \Storage[26][5] ,
         \Storage[26][4] , \Storage[26][3] , \Storage[26][2] ,
         \Storage[26][1] , \Storage[26][0] , \Storage[25][32] ,
         \Storage[25][31] , \Storage[25][30] , \Storage[25][29] ,
         \Storage[25][28] , \Storage[25][27] , \Storage[25][26] ,
         \Storage[25][25] , \Storage[25][24] , \Storage[25][23] ,
         \Storage[25][22] , \Storage[25][21] , \Storage[25][20] ,
         \Storage[25][19] , \Storage[25][18] , \Storage[25][17] ,
         \Storage[25][16] , \Storage[25][15] , \Storage[25][14] ,
         \Storage[25][13] , \Storage[25][12] , \Storage[25][11] ,
         \Storage[25][10] , \Storage[25][9] , \Storage[25][8] ,
         \Storage[25][7] , \Storage[25][6] , \Storage[25][5] ,
         \Storage[25][4] , \Storage[25][3] , \Storage[25][2] ,
         \Storage[25][1] , \Storage[25][0] , \Storage[24][32] ,
         \Storage[24][31] , \Storage[24][30] , \Storage[24][29] ,
         \Storage[24][28] , \Storage[24][27] , \Storage[24][26] ,
         \Storage[24][25] , \Storage[24][24] , \Storage[24][23] ,
         \Storage[24][22] , \Storage[24][21] , \Storage[24][20] ,
         \Storage[24][19] , \Storage[24][18] , \Storage[24][17] ,
         \Storage[24][16] , \Storage[24][15] , \Storage[24][14] ,
         \Storage[24][13] , \Storage[24][12] , \Storage[24][11] ,
         \Storage[24][10] , \Storage[24][9] , \Storage[24][8] ,
         \Storage[24][7] , \Storage[24][6] , \Storage[24][5] ,
         \Storage[24][4] , \Storage[24][3] , \Storage[24][2] ,
         \Storage[24][1] , \Storage[24][0] , \Storage[23][32] ,
         \Storage[23][31] , \Storage[23][30] , \Storage[23][29] ,
         \Storage[23][28] , \Storage[23][27] , \Storage[23][26] ,
         \Storage[23][25] , \Storage[23][24] , \Storage[23][23] ,
         \Storage[23][22] , \Storage[23][21] , \Storage[23][20] ,
         \Storage[23][19] , \Storage[23][18] , \Storage[23][17] ,
         \Storage[23][16] , \Storage[23][15] , \Storage[23][14] ,
         \Storage[23][13] , \Storage[23][12] , \Storage[23][11] ,
         \Storage[23][10] , \Storage[23][9] , \Storage[23][8] ,
         \Storage[23][7] , \Storage[23][6] , \Storage[23][5] ,
         \Storage[23][4] , \Storage[23][3] , \Storage[23][2] ,
         \Storage[23][1] , \Storage[23][0] , \Storage[22][32] ,
         \Storage[22][31] , \Storage[22][30] , \Storage[22][29] ,
         \Storage[22][28] , \Storage[22][27] , \Storage[22][26] ,
         \Storage[22][25] , \Storage[22][24] , \Storage[22][23] ,
         \Storage[22][22] , \Storage[22][21] , \Storage[22][20] ,
         \Storage[22][19] , \Storage[22][18] , \Storage[22][17] ,
         \Storage[22][16] , \Storage[22][15] , \Storage[22][14] ,
         \Storage[22][13] , \Storage[22][12] , \Storage[22][11] ,
         \Storage[22][10] , \Storage[22][9] , \Storage[22][8] ,
         \Storage[22][7] , \Storage[22][6] , \Storage[22][5] ,
         \Storage[22][4] , \Storage[22][3] , \Storage[22][2] ,
         \Storage[22][1] , \Storage[22][0] , \Storage[21][32] ,
         \Storage[21][31] , \Storage[21][30] , \Storage[21][29] ,
         \Storage[21][28] , \Storage[21][27] , \Storage[21][26] ,
         \Storage[21][25] , \Storage[21][24] , \Storage[21][23] ,
         \Storage[21][22] , \Storage[21][21] , \Storage[21][20] ,
         \Storage[21][19] , \Storage[21][18] , \Storage[21][17] ,
         \Storage[21][16] , \Storage[21][15] , \Storage[21][14] ,
         \Storage[21][13] , \Storage[21][12] , \Storage[21][11] ,
         \Storage[21][10] , \Storage[21][9] , \Storage[21][8] ,
         \Storage[21][7] , \Storage[21][6] , \Storage[21][5] ,
         \Storage[21][4] , \Storage[21][3] , \Storage[21][2] ,
         \Storage[21][1] , \Storage[21][0] , \Storage[20][32] ,
         \Storage[20][31] , \Storage[20][30] , \Storage[20][29] ,
         \Storage[20][28] , \Storage[20][27] , \Storage[20][26] ,
         \Storage[20][25] , \Storage[20][24] , \Storage[20][23] ,
         \Storage[20][22] , \Storage[20][21] , \Storage[20][20] ,
         \Storage[20][19] , \Storage[20][18] , \Storage[20][17] ,
         \Storage[20][16] , \Storage[20][15] , \Storage[20][14] ,
         \Storage[20][13] , \Storage[20][12] , \Storage[20][11] ,
         \Storage[20][10] , \Storage[20][9] , \Storage[20][8] ,
         \Storage[20][7] , \Storage[20][6] , \Storage[20][5] ,
         \Storage[20][4] , \Storage[20][3] , \Storage[20][2] ,
         \Storage[20][1] , \Storage[20][0] , \Storage[19][32] ,
         \Storage[19][31] , \Storage[19][30] , \Storage[19][29] ,
         \Storage[19][28] , \Storage[19][27] , \Storage[19][26] ,
         \Storage[19][25] , \Storage[19][24] , \Storage[19][23] ,
         \Storage[19][22] , \Storage[19][21] , \Storage[19][20] ,
         \Storage[19][19] , \Storage[19][18] , \Storage[19][17] ,
         \Storage[19][16] , \Storage[19][15] , \Storage[19][14] ,
         \Storage[19][13] , \Storage[19][12] , \Storage[19][11] ,
         \Storage[19][10] , \Storage[19][9] , \Storage[19][8] ,
         \Storage[19][7] , \Storage[19][6] , \Storage[19][5] ,
         \Storage[19][4] , \Storage[19][3] , \Storage[19][2] ,
         \Storage[19][1] , \Storage[19][0] , \Storage[18][32] ,
         \Storage[18][31] , \Storage[18][30] , \Storage[18][29] ,
         \Storage[18][28] , \Storage[18][27] , \Storage[18][26] ,
         \Storage[18][25] , \Storage[18][24] , \Storage[18][23] ,
         \Storage[18][22] , \Storage[18][21] , \Storage[18][20] ,
         \Storage[18][19] , \Storage[18][18] , \Storage[18][17] ,
         \Storage[18][16] , \Storage[18][15] , \Storage[18][14] ,
         \Storage[18][13] , \Storage[18][12] , \Storage[18][11] ,
         \Storage[18][10] , \Storage[18][9] , \Storage[18][8] ,
         \Storage[18][7] , \Storage[18][6] , \Storage[18][5] ,
         \Storage[18][4] , \Storage[18][3] , \Storage[18][2] ,
         \Storage[18][1] , \Storage[18][0] , \Storage[17][32] ,
         \Storage[17][31] , \Storage[17][30] , \Storage[17][29] ,
         \Storage[17][28] , \Storage[17][27] , \Storage[17][26] ,
         \Storage[17][25] , \Storage[17][24] , \Storage[17][23] ,
         \Storage[17][22] , \Storage[17][21] , \Storage[17][20] ,
         \Storage[17][19] , \Storage[17][18] , \Storage[17][17] ,
         \Storage[17][16] , \Storage[17][15] , \Storage[17][14] ,
         \Storage[17][13] , \Storage[17][12] , \Storage[17][11] ,
         \Storage[17][10] , \Storage[17][9] , \Storage[17][8] ,
         \Storage[17][7] , \Storage[17][6] , \Storage[17][5] ,
         \Storage[17][4] , \Storage[17][3] , \Storage[17][2] ,
         \Storage[17][1] , \Storage[17][0] , \Storage[16][32] ,
         \Storage[16][31] , \Storage[16][30] , \Storage[16][29] ,
         \Storage[16][28] , \Storage[16][27] , \Storage[16][26] ,
         \Storage[16][25] , \Storage[16][24] , \Storage[16][23] ,
         \Storage[16][22] , \Storage[16][21] , \Storage[16][20] ,
         \Storage[16][19] , \Storage[16][18] , \Storage[16][17] ,
         \Storage[16][16] , \Storage[16][15] , \Storage[16][14] ,
         \Storage[16][13] , \Storage[16][12] , \Storage[16][11] ,
         \Storage[16][10] , \Storage[16][9] , \Storage[16][8] ,
         \Storage[16][7] , \Storage[16][6] , \Storage[16][5] ,
         \Storage[16][4] , \Storage[16][3] , \Storage[16][2] ,
         \Storage[16][1] , \Storage[16][0] , \Storage[15][32] ,
         \Storage[15][31] , \Storage[15][30] , \Storage[15][29] ,
         \Storage[15][28] , \Storage[15][27] , \Storage[15][26] ,
         \Storage[15][25] , \Storage[15][24] , \Storage[15][23] ,
         \Storage[15][22] , \Storage[15][21] , \Storage[15][20] ,
         \Storage[15][19] , \Storage[15][18] , \Storage[15][17] ,
         \Storage[15][16] , \Storage[15][15] , \Storage[15][14] ,
         \Storage[15][13] , \Storage[15][12] , \Storage[15][11] ,
         \Storage[15][10] , \Storage[15][9] , \Storage[15][8] ,
         \Storage[15][7] , \Storage[15][6] , \Storage[15][5] ,
         \Storage[15][4] , \Storage[15][3] , \Storage[15][2] ,
         \Storage[15][1] , \Storage[15][0] , \Storage[14][32] ,
         \Storage[14][31] , \Storage[14][30] , \Storage[14][29] ,
         \Storage[14][28] , \Storage[14][27] , \Storage[14][26] ,
         \Storage[14][25] , \Storage[14][24] , \Storage[14][23] ,
         \Storage[14][22] , \Storage[14][21] , \Storage[14][20] ,
         \Storage[14][19] , \Storage[14][18] , \Storage[14][17] ,
         \Storage[14][16] , \Storage[14][15] , \Storage[14][14] ,
         \Storage[14][13] , \Storage[14][12] , \Storage[14][11] ,
         \Storage[14][10] , \Storage[14][9] , \Storage[14][8] ,
         \Storage[14][7] , \Storage[14][6] , \Storage[14][5] ,
         \Storage[14][4] , \Storage[14][3] , \Storage[14][2] ,
         \Storage[14][1] , \Storage[14][0] , \Storage[13][32] ,
         \Storage[13][31] , \Storage[13][30] , \Storage[13][29] ,
         \Storage[13][28] , \Storage[13][27] , \Storage[13][26] ,
         \Storage[13][25] , \Storage[13][24] , \Storage[13][23] ,
         \Storage[13][22] , \Storage[13][21] , \Storage[13][20] ,
         \Storage[13][19] , \Storage[13][18] , \Storage[13][17] ,
         \Storage[13][16] , \Storage[13][15] , \Storage[13][14] ,
         \Storage[13][13] , \Storage[13][12] , \Storage[13][11] ,
         \Storage[13][10] , \Storage[13][9] , \Storage[13][8] ,
         \Storage[13][7] , \Storage[13][6] , \Storage[13][5] ,
         \Storage[13][4] , \Storage[13][3] , \Storage[13][2] ,
         \Storage[13][1] , \Storage[13][0] , \Storage[12][32] ,
         \Storage[12][31] , \Storage[12][30] , \Storage[12][29] ,
         \Storage[12][28] , \Storage[12][27] , \Storage[12][26] ,
         \Storage[12][25] , \Storage[12][24] , \Storage[12][23] ,
         \Storage[12][22] , \Storage[12][21] , \Storage[12][20] ,
         \Storage[12][19] , \Storage[12][18] , \Storage[12][17] ,
         \Storage[12][16] , \Storage[12][15] , \Storage[12][14] ,
         \Storage[12][13] , \Storage[12][12] , \Storage[12][11] ,
         \Storage[12][10] , \Storage[12][9] , \Storage[12][8] ,
         \Storage[12][7] , \Storage[12][6] , \Storage[12][5] ,
         \Storage[12][4] , \Storage[12][3] , \Storage[12][2] ,
         \Storage[12][1] , \Storage[12][0] , \Storage[11][32] ,
         \Storage[11][31] , \Storage[11][30] , \Storage[11][29] ,
         \Storage[11][28] , \Storage[11][27] , \Storage[11][26] ,
         \Storage[11][25] , \Storage[11][24] , \Storage[11][23] ,
         \Storage[11][22] , \Storage[11][21] , \Storage[11][20] ,
         \Storage[11][19] , \Storage[11][18] , \Storage[11][17] ,
         \Storage[11][16] , \Storage[11][15] , \Storage[11][14] ,
         \Storage[11][13] , \Storage[11][12] , \Storage[11][11] ,
         \Storage[11][10] , \Storage[11][9] , \Storage[11][8] ,
         \Storage[11][7] , \Storage[11][6] , \Storage[11][5] ,
         \Storage[11][4] , \Storage[11][3] , \Storage[11][2] ,
         \Storage[11][1] , \Storage[11][0] , \Storage[10][32] ,
         \Storage[10][31] , \Storage[10][30] , \Storage[10][29] ,
         \Storage[10][28] , \Storage[10][27] , \Storage[10][26] ,
         \Storage[10][25] , \Storage[10][24] , \Storage[10][23] ,
         \Storage[10][22] , \Storage[10][21] , \Storage[10][20] ,
         \Storage[10][19] , \Storage[10][18] , \Storage[10][17] ,
         \Storage[10][16] , \Storage[10][15] , \Storage[10][14] ,
         \Storage[10][13] , \Storage[10][12] , \Storage[10][11] ,
         \Storage[10][10] , \Storage[10][9] , \Storage[10][8] ,
         \Storage[10][7] , \Storage[10][6] , \Storage[10][5] ,
         \Storage[10][4] , \Storage[10][3] , \Storage[10][2] ,
         \Storage[10][1] , \Storage[10][0] , \Storage[9][32] ,
         \Storage[9][31] , \Storage[9][30] , \Storage[9][29] ,
         \Storage[9][28] , \Storage[9][27] , \Storage[9][26] ,
         \Storage[9][25] , \Storage[9][24] , \Storage[9][23] ,
         \Storage[9][22] , \Storage[9][21] , \Storage[9][20] ,
         \Storage[9][19] , \Storage[9][18] , \Storage[9][17] ,
         \Storage[9][16] , \Storage[9][15] , \Storage[9][14] ,
         \Storage[9][13] , \Storage[9][12] , \Storage[9][11] ,
         \Storage[9][10] , \Storage[9][9] , \Storage[9][8] , \Storage[9][7] ,
         \Storage[9][6] , \Storage[9][5] , \Storage[9][4] , \Storage[9][3] ,
         \Storage[9][2] , \Storage[9][1] , \Storage[9][0] , \Storage[8][32] ,
         \Storage[8][31] , \Storage[8][30] , \Storage[8][29] ,
         \Storage[8][28] , \Storage[8][27] , \Storage[8][26] ,
         \Storage[8][25] , \Storage[8][24] , \Storage[8][23] ,
         \Storage[8][22] , \Storage[8][21] , \Storage[8][20] ,
         \Storage[8][19] , \Storage[8][18] , \Storage[8][17] ,
         \Storage[8][16] , \Storage[8][15] , \Storage[8][14] ,
         \Storage[8][13] , \Storage[8][12] , \Storage[8][11] ,
         \Storage[8][10] , \Storage[8][9] , \Storage[8][8] , \Storage[8][7] ,
         \Storage[8][6] , \Storage[8][5] , \Storage[8][4] , \Storage[8][3] ,
         \Storage[8][2] , \Storage[8][1] , \Storage[8][0] , \Storage[7][32] ,
         \Storage[7][31] , \Storage[7][30] , \Storage[7][29] ,
         \Storage[7][28] , \Storage[7][27] , \Storage[7][26] ,
         \Storage[7][25] , \Storage[7][24] , \Storage[7][23] ,
         \Storage[7][22] , \Storage[7][21] , \Storage[7][20] ,
         \Storage[7][19] , \Storage[7][18] , \Storage[7][17] ,
         \Storage[7][16] , \Storage[7][15] , \Storage[7][14] ,
         \Storage[7][13] , \Storage[7][12] , \Storage[7][11] ,
         \Storage[7][10] , \Storage[7][9] , \Storage[7][8] , \Storage[7][7] ,
         \Storage[7][6] , \Storage[7][5] , \Storage[7][4] , \Storage[7][3] ,
         \Storage[7][2] , \Storage[7][1] , \Storage[7][0] , \Storage[6][32] ,
         \Storage[6][31] , \Storage[6][30] , \Storage[6][29] ,
         \Storage[6][28] , \Storage[6][27] , \Storage[6][26] ,
         \Storage[6][25] , \Storage[6][24] , \Storage[6][23] ,
         \Storage[6][22] , \Storage[6][21] , \Storage[6][20] ,
         \Storage[6][19] , \Storage[6][18] , \Storage[6][17] ,
         \Storage[6][16] , \Storage[6][15] , \Storage[6][14] ,
         \Storage[6][13] , \Storage[6][12] , \Storage[6][11] ,
         \Storage[6][10] , \Storage[6][9] , \Storage[6][8] , \Storage[6][7] ,
         \Storage[6][6] , \Storage[6][5] , \Storage[6][4] , \Storage[6][3] ,
         \Storage[6][2] , \Storage[6][1] , \Storage[6][0] , \Storage[5][32] ,
         \Storage[5][31] , \Storage[5][30] , \Storage[5][29] ,
         \Storage[5][28] , \Storage[5][27] , \Storage[5][26] ,
         \Storage[5][25] , \Storage[5][24] , \Storage[5][23] ,
         \Storage[5][22] , \Storage[5][21] , \Storage[5][20] ,
         \Storage[5][19] , \Storage[5][18] , \Storage[5][17] ,
         \Storage[5][16] , \Storage[5][15] , \Storage[5][14] ,
         \Storage[5][13] , \Storage[5][12] , \Storage[5][11] ,
         \Storage[5][10] , \Storage[5][9] , \Storage[5][8] , \Storage[5][7] ,
         \Storage[5][6] , \Storage[5][5] , \Storage[5][4] , \Storage[5][3] ,
         \Storage[5][2] , \Storage[5][1] , \Storage[5][0] , \Storage[4][32] ,
         \Storage[4][31] , \Storage[4][30] , \Storage[4][29] ,
         \Storage[4][28] , \Storage[4][27] , \Storage[4][26] ,
         \Storage[4][25] , \Storage[4][24] , \Storage[4][23] ,
         \Storage[4][22] , \Storage[4][21] , \Storage[4][20] ,
         \Storage[4][19] , \Storage[4][18] , \Storage[4][17] ,
         \Storage[4][16] , \Storage[4][15] , \Storage[4][14] ,
         \Storage[4][13] , \Storage[4][12] , \Storage[4][11] ,
         \Storage[4][10] , \Storage[4][9] , \Storage[4][8] , \Storage[4][7] ,
         \Storage[4][6] , \Storage[4][5] , \Storage[4][4] , \Storage[4][3] ,
         \Storage[4][2] , \Storage[4][1] , \Storage[4][0] , \Storage[3][32] ,
         \Storage[3][31] , \Storage[3][30] , \Storage[3][29] ,
         \Storage[3][28] , \Storage[3][27] , \Storage[3][26] ,
         \Storage[3][25] , \Storage[3][24] , \Storage[3][23] ,
         \Storage[3][22] , \Storage[3][21] , \Storage[3][20] ,
         \Storage[3][19] , \Storage[3][18] , \Storage[3][17] ,
         \Storage[3][16] , \Storage[3][15] , \Storage[3][14] ,
         \Storage[3][13] , \Storage[3][12] , \Storage[3][11] ,
         \Storage[3][10] , \Storage[3][9] , \Storage[3][8] , \Storage[3][7] ,
         \Storage[3][6] , \Storage[3][5] , \Storage[3][4] , \Storage[3][3] ,
         \Storage[3][2] , \Storage[3][1] , \Storage[3][0] , \Storage[2][32] ,
         \Storage[2][31] , \Storage[2][30] , \Storage[2][29] ,
         \Storage[2][28] , \Storage[2][27] , \Storage[2][26] ,
         \Storage[2][25] , \Storage[2][24] , \Storage[2][23] ,
         \Storage[2][22] , \Storage[2][21] , \Storage[2][20] ,
         \Storage[2][19] , \Storage[2][18] , \Storage[2][17] ,
         \Storage[2][16] , \Storage[2][15] , \Storage[2][14] ,
         \Storage[2][13] , \Storage[2][12] , \Storage[2][11] ,
         \Storage[2][10] , \Storage[2][9] , \Storage[2][8] , \Storage[2][7] ,
         \Storage[2][6] , \Storage[2][5] , \Storage[2][4] , \Storage[2][3] ,
         \Storage[2][2] , \Storage[2][1] , \Storage[2][0] , \Storage[1][32] ,
         \Storage[1][31] , \Storage[1][30] , \Storage[1][29] ,
         \Storage[1][28] , \Storage[1][27] , \Storage[1][26] ,
         \Storage[1][25] , \Storage[1][24] , \Storage[1][23] ,
         \Storage[1][22] , \Storage[1][21] , \Storage[1][20] ,
         \Storage[1][19] , \Storage[1][18] , \Storage[1][17] ,
         \Storage[1][16] , \Storage[1][15] , \Storage[1][14] ,
         \Storage[1][13] , \Storage[1][12] , \Storage[1][11] ,
         \Storage[1][10] , \Storage[1][9] , \Storage[1][8] , \Storage[1][7] ,
         \Storage[1][6] , \Storage[1][5] , \Storage[1][4] , \Storage[1][3] ,
         \Storage[1][2] , \Storage[1][1] , \Storage[1][0] , \Storage[0][32] ,
         \Storage[0][31] , \Storage[0][30] , \Storage[0][29] ,
         \Storage[0][28] , \Storage[0][27] , \Storage[0][26] ,
         \Storage[0][25] , \Storage[0][24] , \Storage[0][23] ,
         \Storage[0][22] , \Storage[0][21] , \Storage[0][20] ,
         \Storage[0][19] , \Storage[0][18] , \Storage[0][17] ,
         \Storage[0][16] , \Storage[0][15] , \Storage[0][14] ,
         \Storage[0][13] , \Storage[0][12] , \Storage[0][11] ,
         \Storage[0][10] , \Storage[0][9] , \Storage[0][8] , \Storage[0][7] ,
         \Storage[0][6] , \Storage[0][5] , \Storage[0][4] , \Storage[0][3] ,
         \Storage[0][2] , \Storage[0][1] , \Storage[0][0] , N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N85, N150, N183, N216, N249, N282, N315, N348, N381, N414,
         N447, N480, N513, N546, N579, N612, N645, N678, N711, N744, N777,
         N810, N843, N876, N909, N942, N975, N999, N1041, N1074, N1107, N1140,
         N1173, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n1, n2, n3, n4, n5, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
  wire   [31:0] DataOr;
  assign N44 = AddrR[0];
  assign N45 = AddrR[1];
  assign N46 = AddrR[2];
  assign N47 = AddrR[3];
  assign N48 = AddrR[4];

  OR2D1 U3 ( .A1(Read), .A2(Dreadyr), .Z(n107) );
  XNR4D1 U18 ( .A1(n1066), .A2(n1062), .A3(n1074), .A4(n1070), .ZN(n84) );
  XOR4D1 U19 ( .A1(n1082), .A2(n1078), .A3(n1090), .A4(n1086), .Z(n83) );
  XOR4D1 U20 ( .A1(n1050), .A2(n1046), .A3(n1058), .A4(n1054), .Z(n80) );
  XOR4D1 U21 ( .A1(n1022), .A2(n1018), .A3(n1030), .A4(n1026), .Z(n77) );
  XNR4D1 U22 ( .A1(n994), .A2(n990), .A3(n1002), .A4(n998), .ZN(n74) );
  XOR4D1 U27 ( .A1(n90), .A2(N72), .A3(n91), .A4(N75), .Z(n89) );
  XNR4D1 U28 ( .A1(N69), .A2(N68), .A3(N71), .A4(N70), .ZN(n91) );
  XNR4D1 U33 ( .A1(N51), .A2(N50), .A3(N53), .A4(N52), .ZN(n97) );
  XOR4D1 U34 ( .A1(N55), .A2(N54), .A3(N57), .A4(N56), .Z(n96) );
  XNR4D1 U35 ( .A1(N62), .A2(N61), .A3(N64), .A4(N63), .ZN(n93) );
  XNR4D1 U36 ( .A1(N80), .A2(N78), .A3(N82), .A4(N81), .ZN(n87) );
  EDFCNQD1 \Storage_reg[26][32]  ( .D(n842), .E(n734), .CP(n863), .CDN(n662), 
        .Q(\Storage[26][32] ) );
  EDFCNQD1 \Storage_reg[26][31]  ( .D(n1092), .E(n734), .CP(n863), .CDN(n662), 
        .Q(\Storage[26][31] ) );
  EDFCNQD1 \Storage_reg[26][30]  ( .D(n1088), .E(n734), .CP(n863), .CDN(n661), 
        .Q(\Storage[26][30] ) );
  EDFCNQD1 \Storage_reg[26][29]  ( .D(n1084), .E(n734), .CP(n863), .CDN(n661), 
        .Q(\Storage[26][29] ) );
  EDFCNQD1 \Storage_reg[26][28]  ( .D(n1080), .E(n734), .CP(n863), .CDN(n661), 
        .Q(\Storage[26][28] ) );
  EDFCNQD1 \Storage_reg[26][27]  ( .D(n1076), .E(n734), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][27] ) );
  EDFCNQD1 \Storage_reg[26][26]  ( .D(n1072), .E(n734), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][26] ) );
  EDFCNQD1 \Storage_reg[26][25]  ( .D(n1068), .E(n734), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][25] ) );
  EDFCNQD1 \Storage_reg[26][24]  ( .D(n1064), .E(n734), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][24] ) );
  EDFCNQD1 \Storage_reg[26][23]  ( .D(n1060), .E(n734), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][23] ) );
  EDFCNQD1 \Storage_reg[26][22]  ( .D(n1056), .E(n735), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][22] ) );
  EDFCNQD1 \Storage_reg[26][21]  ( .D(n1052), .E(n735), .CP(n864), .CDN(n661), 
        .Q(\Storage[26][21] ) );
  EDFCNQD1 \Storage_reg[26][20]  ( .D(n1048), .E(n735), .CP(n864), .CDN(n660), 
        .Q(\Storage[26][20] ) );
  EDFCNQD1 \Storage_reg[26][19]  ( .D(n1044), .E(n735), .CP(n864), .CDN(n660), 
        .Q(\Storage[26][19] ) );
  EDFCNQD1 \Storage_reg[26][18]  ( .D(n1040), .E(n735), .CP(n864), .CDN(n660), 
        .Q(\Storage[26][18] ) );
  EDFCNQD1 \Storage_reg[26][17]  ( .D(n1036), .E(n735), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][17] ) );
  EDFCNQD1 \Storage_reg[26][16]  ( .D(n1032), .E(n735), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][16] ) );
  EDFCNQD1 \Storage_reg[26][15]  ( .D(n1028), .E(n735), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][15] ) );
  EDFCNQD1 \Storage_reg[26][14]  ( .D(n1024), .E(n735), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][14] ) );
  EDFCNQD1 \Storage_reg[26][13]  ( .D(n1020), .E(n735), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][13] ) );
  EDFCNQD1 \Storage_reg[26][12]  ( .D(n1016), .E(n736), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][12] ) );
  EDFCNQD1 \Storage_reg[26][11]  ( .D(n1012), .E(n736), .CP(n865), .CDN(n660), 
        .Q(\Storage[26][11] ) );
  EDFCNQD1 \Storage_reg[26][10]  ( .D(n1008), .E(n736), .CP(n865), .CDN(n659), 
        .Q(\Storage[26][10] ) );
  EDFCNQD1 \Storage_reg[26][9]  ( .D(n1004), .E(n736), .CP(n865), .CDN(n659), 
        .Q(\Storage[26][9] ) );
  EDFCNQD1 \Storage_reg[26][8]  ( .D(n1000), .E(n736), .CP(n865), .CDN(n659), 
        .Q(\Storage[26][8] ) );
  EDFCNQD1 \Storage_reg[26][7]  ( .D(n996), .E(n736), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][7] ) );
  EDFCNQD1 \Storage_reg[26][6]  ( .D(n992), .E(n736), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][6] ) );
  EDFCNQD1 \Storage_reg[26][5]  ( .D(n988), .E(n736), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][5] ) );
  EDFCNQD1 \Storage_reg[26][4]  ( .D(n984), .E(n736), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][4] ) );
  EDFCNQD1 \Storage_reg[26][3]  ( .D(n980), .E(n736), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][3] ) );
  EDFCNQD1 \Storage_reg[26][2]  ( .D(n976), .E(N999), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][2] ) );
  EDFCNQD1 \Storage_reg[26][1]  ( .D(n972), .E(N999), .CP(n866), .CDN(n659), 
        .Q(\Storage[26][1] ) );
  EDFCNQD1 \Storage_reg[26][0]  ( .D(n968), .E(N999), .CP(n866), .CDN(n658), 
        .Q(\Storage[26][0] ) );
  EDFCNQD1 \Storage_reg[24][32]  ( .D(n842), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][32] ) );
  EDFCNQD1 \Storage_reg[24][31]  ( .D(n1092), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][31] ) );
  EDFCNQD1 \Storage_reg[24][30]  ( .D(n1088), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][30] ) );
  EDFCNQD1 \Storage_reg[24][29]  ( .D(n1084), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][29] ) );
  EDFCNQD1 \Storage_reg[24][28]  ( .D(n1080), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][28] ) );
  EDFCNQD1 \Storage_reg[24][27]  ( .D(n1076), .E(n742), .CP(n870), .CDN(n655), 
        .Q(\Storage[24][27] ) );
  EDFCNQD1 \Storage_reg[24][26]  ( .D(n1072), .E(n742), .CP(n870), .CDN(n654), 
        .Q(\Storage[24][26] ) );
  EDFCNQD1 \Storage_reg[24][25]  ( .D(n1068), .E(n742), .CP(n870), .CDN(n654), 
        .Q(\Storage[24][25] ) );
  EDFCNQD1 \Storage_reg[24][24]  ( .D(n1064), .E(n742), .CP(n870), .CDN(n654), 
        .Q(\Storage[24][24] ) );
  EDFCNQD1 \Storage_reg[24][23]  ( .D(n1060), .E(n742), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][23] ) );
  EDFCNQD1 \Storage_reg[24][22]  ( .D(n1056), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][22] ) );
  EDFCNQD1 \Storage_reg[24][21]  ( .D(n1052), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][21] ) );
  EDFCNQD1 \Storage_reg[24][20]  ( .D(n1048), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][20] ) );
  EDFCNQD1 \Storage_reg[24][19]  ( .D(n1044), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][19] ) );
  EDFCNQD1 \Storage_reg[24][18]  ( .D(n1040), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][18] ) );
  EDFCNQD1 \Storage_reg[24][17]  ( .D(n1036), .E(n743), .CP(n871), .CDN(n654), 
        .Q(\Storage[24][17] ) );
  EDFCNQD1 \Storage_reg[24][16]  ( .D(n1032), .E(n743), .CP(n871), .CDN(n653), 
        .Q(\Storage[24][16] ) );
  EDFCNQD1 \Storage_reg[24][15]  ( .D(n1028), .E(n743), .CP(n871), .CDN(n653), 
        .Q(\Storage[24][15] ) );
  EDFCNQD1 \Storage_reg[24][14]  ( .D(n1024), .E(n743), .CP(n871), .CDN(n653), 
        .Q(\Storage[24][14] ) );
  EDFCNQD1 \Storage_reg[24][13]  ( .D(n1020), .E(n743), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][13] ) );
  EDFCNQD1 \Storage_reg[24][12]  ( .D(n1016), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][12] ) );
  EDFCNQD1 \Storage_reg[24][11]  ( .D(n1012), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][11] ) );
  EDFCNQD1 \Storage_reg[24][10]  ( .D(n1008), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][10] ) );
  EDFCNQD1 \Storage_reg[24][9]  ( .D(n1004), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][9] ) );
  EDFCNQD1 \Storage_reg[24][8]  ( .D(n1000), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][8] ) );
  EDFCNQD1 \Storage_reg[24][7]  ( .D(n996), .E(n744), .CP(n872), .CDN(n653), 
        .Q(\Storage[24][7] ) );
  EDFCNQD1 \Storage_reg[24][6]  ( .D(n992), .E(n744), .CP(n872), .CDN(n652), 
        .Q(\Storage[24][6] ) );
  EDFCNQD1 \Storage_reg[24][5]  ( .D(n988), .E(n744), .CP(n872), .CDN(n652), 
        .Q(\Storage[24][5] ) );
  EDFCNQD1 \Storage_reg[24][4]  ( .D(n984), .E(n744), .CP(n872), .CDN(n652), 
        .Q(\Storage[24][4] ) );
  EDFCNQD1 \Storage_reg[24][3]  ( .D(n980), .E(n744), .CP(n873), .CDN(n652), 
        .Q(\Storage[24][3] ) );
  EDFCNQD1 \Storage_reg[24][2]  ( .D(n976), .E(N942), .CP(n873), .CDN(n652), 
        .Q(\Storage[24][2] ) );
  EDFCNQD1 \Storage_reg[24][1]  ( .D(n972), .E(N942), .CP(n873), .CDN(n652), 
        .Q(\Storage[24][1] ) );
  EDFCNQD1 \Storage_reg[24][0]  ( .D(n968), .E(N942), .CP(n873), .CDN(n652), 
        .Q(\Storage[24][0] ) );
  EDFCNQD1 \Storage_reg[30][32]  ( .D(n842), .E(n718), .CP(n850), .CDN(n675), 
        .Q(\Storage[30][32] ) );
  EDFCNQD1 \Storage_reg[30][31]  ( .D(DataI[31]), .E(n718), .CP(n850), .CDN(
        n675), .Q(\Storage[30][31] ) );
  EDFCNQD1 \Storage_reg[30][30]  ( .D(DataI[30]), .E(n718), .CP(n850), .CDN(
        n675), .Q(\Storage[30][30] ) );
  EDFCNQD1 \Storage_reg[30][29]  ( .D(DataI[29]), .E(n718), .CP(n850), .CDN(
        n675), .Q(\Storage[30][29] ) );
  EDFCNQD1 \Storage_reg[30][28]  ( .D(DataI[28]), .E(n718), .CP(n850), .CDN(
        n674), .Q(\Storage[30][28] ) );
  EDFCNQD1 \Storage_reg[30][27]  ( .D(DataI[27]), .E(n718), .CP(n850), .CDN(
        n674), .Q(\Storage[30][27] ) );
  EDFCNQD1 \Storage_reg[30][26]  ( .D(DataI[26]), .E(n718), .CP(n850), .CDN(
        n674), .Q(\Storage[30][26] ) );
  EDFCNQD1 \Storage_reg[30][25]  ( .D(DataI[25]), .E(n718), .CP(n851), .CDN(
        n674), .Q(\Storage[30][25] ) );
  EDFCNQD1 \Storage_reg[30][24]  ( .D(DataI[24]), .E(n718), .CP(n851), .CDN(
        n674), .Q(\Storage[30][24] ) );
  EDFCNQD1 \Storage_reg[30][23]  ( .D(DataI[23]), .E(n718), .CP(n851), .CDN(
        n674), .Q(\Storage[30][23] ) );
  EDFCNQD1 \Storage_reg[30][22]  ( .D(DataI[22]), .E(n719), .CP(n851), .CDN(
        n674), .Q(\Storage[30][22] ) );
  EDFCNQD1 \Storage_reg[30][21]  ( .D(DataI[21]), .E(n719), .CP(n851), .CDN(
        n674), .Q(\Storage[30][21] ) );
  EDFCNQD1 \Storage_reg[30][20]  ( .D(DataI[20]), .E(n719), .CP(n851), .CDN(
        n674), .Q(\Storage[30][20] ) );
  EDFCNQD1 \Storage_reg[30][19]  ( .D(DataI[19]), .E(n719), .CP(n851), .CDN(
        n674), .Q(\Storage[30][19] ) );
  EDFCNQD1 \Storage_reg[30][18]  ( .D(DataI[18]), .E(n719), .CP(n851), .CDN(
        n673), .Q(\Storage[30][18] ) );
  EDFCNQD1 \Storage_reg[30][17]  ( .D(DataI[17]), .E(n719), .CP(n851), .CDN(
        n673), .Q(\Storage[30][17] ) );
  EDFCNQD1 \Storage_reg[30][16]  ( .D(DataI[16]), .E(n719), .CP(n851), .CDN(
        n673), .Q(\Storage[30][16] ) );
  EDFCNQD1 \Storage_reg[30][15]  ( .D(DataI[15]), .E(n719), .CP(n852), .CDN(
        n673), .Q(\Storage[30][15] ) );
  EDFCNQD1 \Storage_reg[30][14]  ( .D(DataI[14]), .E(n719), .CP(n852), .CDN(
        n673), .Q(\Storage[30][14] ) );
  EDFCNQD1 \Storage_reg[30][13]  ( .D(DataI[13]), .E(n719), .CP(n852), .CDN(
        n673), .Q(\Storage[30][13] ) );
  EDFCNQD1 \Storage_reg[30][12]  ( .D(DataI[12]), .E(n720), .CP(n852), .CDN(
        n673), .Q(\Storage[30][12] ) );
  EDFCNQD1 \Storage_reg[30][11]  ( .D(DataI[11]), .E(n720), .CP(n852), .CDN(
        n673), .Q(\Storage[30][11] ) );
  EDFCNQD1 \Storage_reg[30][10]  ( .D(DataI[10]), .E(n720), .CP(n852), .CDN(
        n673), .Q(\Storage[30][10] ) );
  EDFCNQD1 \Storage_reg[30][9]  ( .D(DataI[9]), .E(n720), .CP(n852), .CDN(n673), .Q(\Storage[30][9] ) );
  EDFCNQD1 \Storage_reg[30][8]  ( .D(DataI[8]), .E(n720), .CP(n852), .CDN(n672), .Q(\Storage[30][8] ) );
  EDFCNQD1 \Storage_reg[30][7]  ( .D(DataI[7]), .E(n720), .CP(n852), .CDN(n672), .Q(\Storage[30][7] ) );
  EDFCNQD1 \Storage_reg[30][6]  ( .D(DataI[6]), .E(n720), .CP(n852), .CDN(n672), .Q(\Storage[30][6] ) );
  EDFCNQD1 \Storage_reg[30][5]  ( .D(DataI[5]), .E(n720), .CP(n853), .CDN(n672), .Q(\Storage[30][5] ) );
  EDFCNQD1 \Storage_reg[30][4]  ( .D(DataI[4]), .E(n720), .CP(n853), .CDN(n672), .Q(\Storage[30][4] ) );
  EDFCNQD1 \Storage_reg[30][3]  ( .D(DataI[3]), .E(n720), .CP(n853), .CDN(n672), .Q(\Storage[30][3] ) );
  EDFCNQD1 \Storage_reg[30][2]  ( .D(DataI[2]), .E(N1140), .CP(n853), .CDN(
        n672), .Q(\Storage[30][2] ) );
  EDFCNQD1 \Storage_reg[30][1]  ( .D(DataI[1]), .E(N1140), .CP(n853), .CDN(
        n672), .Q(\Storage[30][1] ) );
  EDFCNQD1 \Storage_reg[30][0]  ( .D(DataI[0]), .E(N1140), .CP(n853), .CDN(
        n672), .Q(\Storage[30][0] ) );
  EDFCNQD1 \Storage_reg[29][32]  ( .D(n842), .E(n722), .CP(n853), .CDN(n672), 
        .Q(\Storage[29][32] ) );
  EDFCNQD1 \Storage_reg[29][31]  ( .D(DataI[31]), .E(n722), .CP(n853), .CDN(
        n671), .Q(\Storage[29][31] ) );
  EDFCNQD1 \Storage_reg[29][30]  ( .D(DataI[30]), .E(n722), .CP(n853), .CDN(
        n671), .Q(\Storage[29][30] ) );
  EDFCNQD1 \Storage_reg[29][29]  ( .D(DataI[29]), .E(n722), .CP(n853), .CDN(
        n671), .Q(\Storage[29][29] ) );
  EDFCNQD1 \Storage_reg[29][28]  ( .D(DataI[28]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][28] ) );
  EDFCNQD1 \Storage_reg[29][27]  ( .D(DataI[27]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][27] ) );
  EDFCNQD1 \Storage_reg[29][26]  ( .D(DataI[26]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][26] ) );
  EDFCNQD1 \Storage_reg[29][25]  ( .D(DataI[25]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][25] ) );
  EDFCNQD1 \Storage_reg[29][24]  ( .D(DataI[24]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][24] ) );
  EDFCNQD1 \Storage_reg[29][23]  ( .D(DataI[23]), .E(n722), .CP(n854), .CDN(
        n671), .Q(\Storage[29][23] ) );
  EDFCNQD1 \Storage_reg[29][22]  ( .D(DataI[22]), .E(n723), .CP(n854), .CDN(
        n671), .Q(\Storage[29][22] ) );
  EDFCNQD1 \Storage_reg[29][21]  ( .D(DataI[21]), .E(n723), .CP(n854), .CDN(
        n670), .Q(\Storage[29][21] ) );
  EDFCNQD1 \Storage_reg[29][20]  ( .D(DataI[20]), .E(n723), .CP(n854), .CDN(
        n670), .Q(\Storage[29][20] ) );
  EDFCNQD1 \Storage_reg[29][19]  ( .D(DataI[19]), .E(n723), .CP(n854), .CDN(
        n670), .Q(\Storage[29][19] ) );
  EDFCNQD1 \Storage_reg[29][18]  ( .D(DataI[18]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][18] ) );
  EDFCNQD1 \Storage_reg[29][17]  ( .D(DataI[17]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][17] ) );
  EDFCNQD1 \Storage_reg[29][16]  ( .D(DataI[16]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][16] ) );
  EDFCNQD1 \Storage_reg[29][15]  ( .D(DataI[15]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][15] ) );
  EDFCNQD1 \Storage_reg[29][14]  ( .D(DataI[14]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][14] ) );
  EDFCNQD1 \Storage_reg[29][13]  ( .D(DataI[13]), .E(n723), .CP(n855), .CDN(
        n670), .Q(\Storage[29][13] ) );
  EDFCNQD1 \Storage_reg[29][12]  ( .D(DataI[12]), .E(n724), .CP(n855), .CDN(
        n670), .Q(\Storage[29][12] ) );
  EDFCNQD1 \Storage_reg[29][11]  ( .D(DataI[11]), .E(n724), .CP(n855), .CDN(
        n669), .Q(\Storage[29][11] ) );
  EDFCNQD1 \Storage_reg[29][10]  ( .D(DataI[10]), .E(n724), .CP(n855), .CDN(
        n669), .Q(\Storage[29][10] ) );
  EDFCNQD1 \Storage_reg[29][9]  ( .D(DataI[9]), .E(n724), .CP(n855), .CDN(n669), .Q(\Storage[29][9] ) );
  EDFCNQD1 \Storage_reg[29][8]  ( .D(DataI[8]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][8] ) );
  EDFCNQD1 \Storage_reg[29][7]  ( .D(DataI[7]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][7] ) );
  EDFCNQD1 \Storage_reg[29][6]  ( .D(DataI[6]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][6] ) );
  EDFCNQD1 \Storage_reg[29][5]  ( .D(DataI[5]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][5] ) );
  EDFCNQD1 \Storage_reg[29][4]  ( .D(DataI[4]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][4] ) );
  EDFCNQD1 \Storage_reg[29][3]  ( .D(DataI[3]), .E(n724), .CP(n856), .CDN(n669), .Q(\Storage[29][3] ) );
  EDFCNQD1 \Storage_reg[29][2]  ( .D(DataI[2]), .E(N1107), .CP(n856), .CDN(
        n669), .Q(\Storage[29][2] ) );
  EDFCNQD1 \Storage_reg[29][1]  ( .D(DataI[1]), .E(N1107), .CP(n856), .CDN(
        n668), .Q(\Storage[29][1] ) );
  EDFCNQD1 \Storage_reg[29][0]  ( .D(DataI[0]), .E(N1107), .CP(n856), .CDN(
        n668), .Q(\Storage[29][0] ) );
  EDFCNQD1 \Storage_reg[28][32]  ( .D(n842), .E(n726), .CP(n856), .CDN(n668), 
        .Q(\Storage[28][32] ) );
  EDFCNQD1 \Storage_reg[28][31]  ( .D(n1092), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][31] ) );
  EDFCNQD1 \Storage_reg[28][30]  ( .D(n1088), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][30] ) );
  EDFCNQD1 \Storage_reg[28][29]  ( .D(n1084), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][29] ) );
  EDFCNQD1 \Storage_reg[28][28]  ( .D(n1080), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][28] ) );
  EDFCNQD1 \Storage_reg[28][27]  ( .D(n1076), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][27] ) );
  EDFCNQD1 \Storage_reg[28][26]  ( .D(n1072), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][26] ) );
  EDFCNQD1 \Storage_reg[28][25]  ( .D(n1068), .E(n726), .CP(n857), .CDN(n668), 
        .Q(\Storage[28][25] ) );
  EDFCNQD1 \Storage_reg[28][24]  ( .D(n1064), .E(n726), .CP(n857), .CDN(n667), 
        .Q(\Storage[28][24] ) );
  EDFCNQD1 \Storage_reg[28][23]  ( .D(n1060), .E(n726), .CP(n857), .CDN(n667), 
        .Q(\Storage[28][23] ) );
  EDFCNQD1 \Storage_reg[28][22]  ( .D(n1056), .E(n727), .CP(n857), .CDN(n667), 
        .Q(\Storage[28][22] ) );
  EDFCNQD1 \Storage_reg[28][21]  ( .D(n1052), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][21] ) );
  EDFCNQD1 \Storage_reg[28][20]  ( .D(n1048), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][20] ) );
  EDFCNQD1 \Storage_reg[28][19]  ( .D(n1044), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][19] ) );
  EDFCNQD1 \Storage_reg[28][18]  ( .D(n1040), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][18] ) );
  EDFCNQD1 \Storage_reg[28][17]  ( .D(n1036), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][17] ) );
  EDFCNQD1 \Storage_reg[28][16]  ( .D(n1032), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][16] ) );
  EDFCNQD1 \Storage_reg[28][15]  ( .D(n1028), .E(n727), .CP(n858), .CDN(n667), 
        .Q(\Storage[28][15] ) );
  EDFCNQD1 \Storage_reg[28][14]  ( .D(n1024), .E(n727), .CP(n858), .CDN(n666), 
        .Q(\Storage[28][14] ) );
  EDFCNQD1 \Storage_reg[28][13]  ( .D(n1020), .E(n727), .CP(n858), .CDN(n666), 
        .Q(\Storage[28][13] ) );
  EDFCNQD1 \Storage_reg[28][12]  ( .D(n1016), .E(n728), .CP(n858), .CDN(n666), 
        .Q(\Storage[28][12] ) );
  EDFCNQD1 \Storage_reg[28][11]  ( .D(n1012), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][11] ) );
  EDFCNQD1 \Storage_reg[28][10]  ( .D(n1008), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][10] ) );
  EDFCNQD1 \Storage_reg[28][9]  ( .D(n1004), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][9] ) );
  EDFCNQD1 \Storage_reg[28][8]  ( .D(n1000), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][8] ) );
  EDFCNQD1 \Storage_reg[28][7]  ( .D(n996), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][7] ) );
  EDFCNQD1 \Storage_reg[28][6]  ( .D(n992), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][6] ) );
  EDFCNQD1 \Storage_reg[28][5]  ( .D(n988), .E(n728), .CP(n859), .CDN(n666), 
        .Q(\Storage[28][5] ) );
  EDFCNQD1 \Storage_reg[28][4]  ( .D(n984), .E(n728), .CP(n859), .CDN(n665), 
        .Q(\Storage[28][4] ) );
  EDFCNQD1 \Storage_reg[28][3]  ( .D(n980), .E(n728), .CP(n859), .CDN(n665), 
        .Q(\Storage[28][3] ) );
  EDFCNQD1 \Storage_reg[28][2]  ( .D(n976), .E(N1074), .CP(n859), .CDN(n665), 
        .Q(\Storage[28][2] ) );
  EDFCNQD1 \Storage_reg[28][1]  ( .D(n972), .E(N1074), .CP(n860), .CDN(n665), 
        .Q(\Storage[28][1] ) );
  EDFCNQD1 \Storage_reg[28][0]  ( .D(n968), .E(N1074), .CP(n860), .CDN(n665), 
        .Q(\Storage[28][0] ) );
  EDFCNQD1 \Storage_reg[27][32]  ( .D(n842), .E(n730), .CP(n860), .CDN(n665), 
        .Q(\Storage[27][32] ) );
  EDFCNQD1 \Storage_reg[27][31]  ( .D(n1092), .E(n730), .CP(n860), .CDN(n665), 
        .Q(\Storage[27][31] ) );
  EDFCNQD1 \Storage_reg[27][30]  ( .D(n1088), .E(n730), .CP(n860), .CDN(n665), 
        .Q(\Storage[27][30] ) );
  EDFCNQD1 \Storage_reg[27][29]  ( .D(n1084), .E(n730), .CP(n860), .CDN(n665), 
        .Q(\Storage[27][29] ) );
  EDFCNQD1 \Storage_reg[27][28]  ( .D(n1080), .E(n730), .CP(n860), .CDN(n665), 
        .Q(\Storage[27][28] ) );
  EDFCNQD1 \Storage_reg[27][27]  ( .D(n1076), .E(n730), .CP(n860), .CDN(n664), 
        .Q(\Storage[27][27] ) );
  EDFCNQD1 \Storage_reg[27][26]  ( .D(n1072), .E(n730), .CP(n860), .CDN(n664), 
        .Q(\Storage[27][26] ) );
  EDFCNQD1 \Storage_reg[27][25]  ( .D(n1068), .E(n730), .CP(n860), .CDN(n664), 
        .Q(\Storage[27][25] ) );
  EDFCNQD1 \Storage_reg[27][24]  ( .D(n1064), .E(n730), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][24] ) );
  EDFCNQD1 \Storage_reg[27][23]  ( .D(n1060), .E(n730), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][23] ) );
  EDFCNQD1 \Storage_reg[27][22]  ( .D(n1056), .E(n731), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][22] ) );
  EDFCNQD1 \Storage_reg[27][21]  ( .D(n1052), .E(n731), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][21] ) );
  EDFCNQD1 \Storage_reg[27][20]  ( .D(n1048), .E(n731), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][20] ) );
  EDFCNQD1 \Storage_reg[27][19]  ( .D(n1044), .E(n731), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][19] ) );
  EDFCNQD1 \Storage_reg[27][18]  ( .D(n1040), .E(n731), .CP(n861), .CDN(n664), 
        .Q(\Storage[27][18] ) );
  EDFCNQD1 \Storage_reg[27][17]  ( .D(n1036), .E(n731), .CP(n861), .CDN(n663), 
        .Q(\Storage[27][17] ) );
  EDFCNQD1 \Storage_reg[27][16]  ( .D(n1032), .E(n731), .CP(n861), .CDN(n663), 
        .Q(\Storage[27][16] ) );
  EDFCNQD1 \Storage_reg[27][15]  ( .D(n1028), .E(n731), .CP(n861), .CDN(n663), 
        .Q(\Storage[27][15] ) );
  EDFCNQD1 \Storage_reg[27][14]  ( .D(n1024), .E(n731), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][14] ) );
  EDFCNQD1 \Storage_reg[27][13]  ( .D(n1020), .E(n731), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][13] ) );
  EDFCNQD1 \Storage_reg[27][12]  ( .D(n1016), .E(n732), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][12] ) );
  EDFCNQD1 \Storage_reg[27][11]  ( .D(n1012), .E(n732), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][11] ) );
  EDFCNQD1 \Storage_reg[27][10]  ( .D(n1008), .E(n732), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][10] ) );
  EDFCNQD1 \Storage_reg[27][9]  ( .D(n1004), .E(n732), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][9] ) );
  EDFCNQD1 \Storage_reg[27][8]  ( .D(n1000), .E(n732), .CP(n862), .CDN(n663), 
        .Q(\Storage[27][8] ) );
  EDFCNQD1 \Storage_reg[27][7]  ( .D(n996), .E(n732), .CP(n862), .CDN(n662), 
        .Q(\Storage[27][7] ) );
  EDFCNQD1 \Storage_reg[27][6]  ( .D(n992), .E(n732), .CP(n862), .CDN(n662), 
        .Q(\Storage[27][6] ) );
  EDFCNQD1 \Storage_reg[27][5]  ( .D(n988), .E(n732), .CP(n862), .CDN(n662), 
        .Q(\Storage[27][5] ) );
  EDFCNQD1 \Storage_reg[27][4]  ( .D(n984), .E(n732), .CP(n863), .CDN(n662), 
        .Q(\Storage[27][4] ) );
  EDFCNQD1 \Storage_reg[27][3]  ( .D(n980), .E(n732), .CP(n863), .CDN(n662), 
        .Q(\Storage[27][3] ) );
  EDFCNQD1 \Storage_reg[27][2]  ( .D(n976), .E(N1041), .CP(n863), .CDN(n662), 
        .Q(\Storage[27][2] ) );
  EDFCNQD1 \Storage_reg[27][1]  ( .D(n972), .E(N1041), .CP(n863), .CDN(n662), 
        .Q(\Storage[27][1] ) );
  EDFCNQD1 \Storage_reg[27][0]  ( .D(n968), .E(N1041), .CP(n863), .CDN(n662), 
        .Q(\Storage[27][0] ) );
  EDFCNQD1 \Storage_reg[25][32]  ( .D(n842), .E(n738), .CP(n866), .CDN(n658), 
        .Q(\Storage[25][32] ) );
  EDFCNQD1 \Storage_reg[25][31]  ( .D(n1092), .E(n738), .CP(n866), .CDN(n658), 
        .Q(\Storage[25][31] ) );
  EDFCNQD1 \Storage_reg[25][30]  ( .D(n1088), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][30] ) );
  EDFCNQD1 \Storage_reg[25][29]  ( .D(n1084), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][29] ) );
  EDFCNQD1 \Storage_reg[25][28]  ( .D(n1080), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][28] ) );
  EDFCNQD1 \Storage_reg[25][27]  ( .D(n1076), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][27] ) );
  EDFCNQD1 \Storage_reg[25][26]  ( .D(n1072), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][26] ) );
  EDFCNQD1 \Storage_reg[25][25]  ( .D(n1068), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][25] ) );
  EDFCNQD1 \Storage_reg[25][24]  ( .D(n1064), .E(n738), .CP(n867), .CDN(n658), 
        .Q(\Storage[25][24] ) );
  EDFCNQD1 \Storage_reg[25][23]  ( .D(n1060), .E(n738), .CP(n867), .CDN(n657), 
        .Q(\Storage[25][23] ) );
  EDFCNQD1 \Storage_reg[25][22]  ( .D(n1056), .E(n739), .CP(n867), .CDN(n657), 
        .Q(\Storage[25][22] ) );
  EDFCNQD1 \Storage_reg[25][21]  ( .D(n1052), .E(n739), .CP(n867), .CDN(n657), 
        .Q(\Storage[25][21] ) );
  EDFCNQD1 \Storage_reg[25][20]  ( .D(n1048), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][20] ) );
  EDFCNQD1 \Storage_reg[25][19]  ( .D(n1044), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][19] ) );
  EDFCNQD1 \Storage_reg[25][18]  ( .D(n1040), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][18] ) );
  EDFCNQD1 \Storage_reg[25][17]  ( .D(n1036), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][17] ) );
  EDFCNQD1 \Storage_reg[25][16]  ( .D(n1032), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][16] ) );
  EDFCNQD1 \Storage_reg[25][15]  ( .D(n1028), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][15] ) );
  EDFCNQD1 \Storage_reg[25][14]  ( .D(n1024), .E(n739), .CP(n868), .CDN(n657), 
        .Q(\Storage[25][14] ) );
  EDFCNQD1 \Storage_reg[25][13]  ( .D(n1020), .E(n739), .CP(n868), .CDN(n656), 
        .Q(\Storage[25][13] ) );
  EDFCNQD1 \Storage_reg[25][12]  ( .D(n1016), .E(n740), .CP(n868), .CDN(n656), 
        .Q(\Storage[25][12] ) );
  EDFCNQD1 \Storage_reg[25][11]  ( .D(n1012), .E(n740), .CP(n868), .CDN(n656), 
        .Q(\Storage[25][11] ) );
  EDFCNQD1 \Storage_reg[25][10]  ( .D(n1008), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][10] ) );
  EDFCNQD1 \Storage_reg[25][9]  ( .D(n1004), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][9] ) );
  EDFCNQD1 \Storage_reg[25][8]  ( .D(n1000), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][8] ) );
  EDFCNQD1 \Storage_reg[25][7]  ( .D(n996), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][7] ) );
  EDFCNQD1 \Storage_reg[25][6]  ( .D(n992), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][6] ) );
  EDFCNQD1 \Storage_reg[25][5]  ( .D(n988), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][5] ) );
  EDFCNQD1 \Storage_reg[25][4]  ( .D(n984), .E(n740), .CP(n869), .CDN(n656), 
        .Q(\Storage[25][4] ) );
  EDFCNQD1 \Storage_reg[25][3]  ( .D(n980), .E(n740), .CP(n869), .CDN(n655), 
        .Q(\Storage[25][3] ) );
  EDFCNQD1 \Storage_reg[25][2]  ( .D(n976), .E(N975), .CP(n869), .CDN(n655), 
        .Q(\Storage[25][2] ) );
  EDFCNQD1 \Storage_reg[25][1]  ( .D(n972), .E(N975), .CP(n869), .CDN(n655), 
        .Q(\Storage[25][1] ) );
  EDFCNQD1 \Storage_reg[25][0]  ( .D(n968), .E(N975), .CP(n870), .CDN(n655), 
        .Q(\Storage[25][0] ) );
  EDFCNQD1 \Storage_reg[22][32]  ( .D(n842), .E(n750), .CP(n876), .CDN(n648), 
        .Q(\Storage[22][32] ) );
  EDFCNQD1 \Storage_reg[22][31]  ( .D(n1092), .E(n750), .CP(n876), .CDN(n648), 
        .Q(\Storage[22][31] ) );
  EDFCNQD1 \Storage_reg[22][30]  ( .D(n1088), .E(n750), .CP(n876), .CDN(n648), 
        .Q(\Storage[22][30] ) );
  EDFCNQD1 \Storage_reg[22][29]  ( .D(n1084), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][29] ) );
  EDFCNQD1 \Storage_reg[22][28]  ( .D(n1080), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][28] ) );
  EDFCNQD1 \Storage_reg[22][27]  ( .D(n1076), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][27] ) );
  EDFCNQD1 \Storage_reg[22][26]  ( .D(n1072), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][26] ) );
  EDFCNQD1 \Storage_reg[22][25]  ( .D(n1068), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][25] ) );
  EDFCNQD1 \Storage_reg[22][24]  ( .D(n1064), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][24] ) );
  EDFCNQD1 \Storage_reg[22][23]  ( .D(n1060), .E(n750), .CP(n877), .CDN(n648), 
        .Q(\Storage[22][23] ) );
  EDFCNQD1 \Storage_reg[22][22]  ( .D(n1056), .E(n751), .CP(n877), .CDN(n647), 
        .Q(\Storage[22][22] ) );
  EDFCNQD1 \Storage_reg[22][21]  ( .D(n1052), .E(n751), .CP(n877), .CDN(n647), 
        .Q(\Storage[22][21] ) );
  EDFCNQD1 \Storage_reg[22][20]  ( .D(n1048), .E(n751), .CP(n877), .CDN(n647), 
        .Q(\Storage[22][20] ) );
  EDFCNQD1 \Storage_reg[22][19]  ( .D(n1044), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][19] ) );
  EDFCNQD1 \Storage_reg[22][18]  ( .D(n1040), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][18] ) );
  EDFCNQD1 \Storage_reg[22][17]  ( .D(n1036), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][17] ) );
  EDFCNQD1 \Storage_reg[22][16]  ( .D(n1032), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][16] ) );
  EDFCNQD1 \Storage_reg[22][15]  ( .D(n1028), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][15] ) );
  EDFCNQD1 \Storage_reg[22][14]  ( .D(n1024), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][14] ) );
  EDFCNQD1 \Storage_reg[22][13]  ( .D(n1020), .E(n751), .CP(n878), .CDN(n647), 
        .Q(\Storage[22][13] ) );
  EDFCNQD1 \Storage_reg[22][12]  ( .D(n1016), .E(n752), .CP(n878), .CDN(n646), 
        .Q(\Storage[22][12] ) );
  EDFCNQD1 \Storage_reg[22][11]  ( .D(n1012), .E(n752), .CP(n878), .CDN(n646), 
        .Q(\Storage[22][11] ) );
  EDFCNQD1 \Storage_reg[22][10]  ( .D(n1008), .E(n752), .CP(n878), .CDN(n646), 
        .Q(\Storage[22][10] ) );
  EDFCNQD1 \Storage_reg[22][9]  ( .D(n1004), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][9] ) );
  EDFCNQD1 \Storage_reg[22][8]  ( .D(n1000), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][8] ) );
  EDFCNQD1 \Storage_reg[22][7]  ( .D(n996), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][7] ) );
  EDFCNQD1 \Storage_reg[22][6]  ( .D(n992), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][6] ) );
  EDFCNQD1 \Storage_reg[22][5]  ( .D(n988), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][5] ) );
  EDFCNQD1 \Storage_reg[22][4]  ( .D(n984), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][4] ) );
  EDFCNQD1 \Storage_reg[22][3]  ( .D(n980), .E(n752), .CP(n879), .CDN(n646), 
        .Q(\Storage[22][3] ) );
  EDFCNQD1 \Storage_reg[22][2]  ( .D(n976), .E(N876), .CP(n879), .CDN(n645), 
        .Q(\Storage[22][2] ) );
  EDFCNQD1 \Storage_reg[22][1]  ( .D(n972), .E(N876), .CP(n879), .CDN(n645), 
        .Q(\Storage[22][1] ) );
  EDFCNQD1 \Storage_reg[22][0]  ( .D(n968), .E(N876), .CP(n879), .CDN(n645), 
        .Q(\Storage[22][0] ) );
  EDFCNQD1 \Storage_reg[21][32]  ( .D(n843), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][32] ) );
  EDFCNQD1 \Storage_reg[21][31]  ( .D(n1092), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][31] ) );
  EDFCNQD1 \Storage_reg[21][30]  ( .D(n1088), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][30] ) );
  EDFCNQD1 \Storage_reg[21][29]  ( .D(n1084), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][29] ) );
  EDFCNQD1 \Storage_reg[21][28]  ( .D(n1080), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][28] ) );
  EDFCNQD1 \Storage_reg[21][27]  ( .D(n1076), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][27] ) );
  EDFCNQD1 \Storage_reg[21][26]  ( .D(n1072), .E(n754), .CP(n880), .CDN(n645), 
        .Q(\Storage[21][26] ) );
  EDFCNQD1 \Storage_reg[21][25]  ( .D(n1068), .E(n754), .CP(n880), .CDN(n644), 
        .Q(\Storage[21][25] ) );
  EDFCNQD1 \Storage_reg[21][24]  ( .D(n1064), .E(n754), .CP(n880), .CDN(n644), 
        .Q(\Storage[21][24] ) );
  EDFCNQD1 \Storage_reg[21][23]  ( .D(n1060), .E(n754), .CP(n880), .CDN(n644), 
        .Q(\Storage[21][23] ) );
  EDFCNQD1 \Storage_reg[21][22]  ( .D(n1056), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][22] ) );
  EDFCNQD1 \Storage_reg[21][21]  ( .D(n1052), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][21] ) );
  EDFCNQD1 \Storage_reg[21][20]  ( .D(n1048), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][20] ) );
  EDFCNQD1 \Storage_reg[21][19]  ( .D(n1044), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][19] ) );
  EDFCNQD1 \Storage_reg[21][18]  ( .D(n1040), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][18] ) );
  EDFCNQD1 \Storage_reg[21][17]  ( .D(n1036), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][17] ) );
  EDFCNQD1 \Storage_reg[21][16]  ( .D(n1032), .E(n755), .CP(n881), .CDN(n644), 
        .Q(\Storage[21][16] ) );
  EDFCNQD1 \Storage_reg[21][15]  ( .D(n1028), .E(n755), .CP(n881), .CDN(n643), 
        .Q(\Storage[21][15] ) );
  EDFCNQD1 \Storage_reg[21][14]  ( .D(n1024), .E(n755), .CP(n881), .CDN(n643), 
        .Q(\Storage[21][14] ) );
  EDFCNQD1 \Storage_reg[21][13]  ( .D(n1020), .E(n755), .CP(n881), .CDN(n643), 
        .Q(\Storage[21][13] ) );
  EDFCNQD1 \Storage_reg[21][12]  ( .D(n1016), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][12] ) );
  EDFCNQD1 \Storage_reg[21][11]  ( .D(n1012), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][11] ) );
  EDFCNQD1 \Storage_reg[21][10]  ( .D(n1008), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][10] ) );
  EDFCNQD1 \Storage_reg[21][9]  ( .D(n1004), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][9] ) );
  EDFCNQD1 \Storage_reg[21][8]  ( .D(n1000), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][8] ) );
  EDFCNQD1 \Storage_reg[21][7]  ( .D(n996), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][7] ) );
  EDFCNQD1 \Storage_reg[21][6]  ( .D(n992), .E(n756), .CP(n882), .CDN(n643), 
        .Q(\Storage[21][6] ) );
  EDFCNQD1 \Storage_reg[21][5]  ( .D(n988), .E(n756), .CP(n882), .CDN(n642), 
        .Q(\Storage[21][5] ) );
  EDFCNQD1 \Storage_reg[21][4]  ( .D(n984), .E(n756), .CP(n882), .CDN(n642), 
        .Q(\Storage[21][4] ) );
  EDFCNQD1 \Storage_reg[21][3]  ( .D(n980), .E(n756), .CP(n882), .CDN(n642), 
        .Q(\Storage[21][3] ) );
  EDFCNQD1 \Storage_reg[21][2]  ( .D(n976), .E(N843), .CP(n883), .CDN(n642), 
        .Q(\Storage[21][2] ) );
  EDFCNQD1 \Storage_reg[21][1]  ( .D(n972), .E(N843), .CP(n883), .CDN(n642), 
        .Q(\Storage[21][1] ) );
  EDFCNQD1 \Storage_reg[21][0]  ( .D(n968), .E(N843), .CP(n883), .CDN(n642), 
        .Q(\Storage[21][0] ) );
  EDFCNQD1 \Storage_reg[18][32]  ( .D(n843), .E(n766), .CP(n889), .CDN(n635), 
        .Q(\Storage[18][32] ) );
  EDFCNQD1 \Storage_reg[18][31]  ( .D(n1091), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][31] ) );
  EDFCNQD1 \Storage_reg[18][30]  ( .D(n1087), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][30] ) );
  EDFCNQD1 \Storage_reg[18][29]  ( .D(n1083), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][29] ) );
  EDFCNQD1 \Storage_reg[18][28]  ( .D(n1079), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][28] ) );
  EDFCNQD1 \Storage_reg[18][27]  ( .D(n1075), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][27] ) );
  EDFCNQD1 \Storage_reg[18][26]  ( .D(n1071), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][26] ) );
  EDFCNQD1 \Storage_reg[18][25]  ( .D(n1067), .E(n766), .CP(n890), .CDN(n635), 
        .Q(\Storage[18][25] ) );
  EDFCNQD1 \Storage_reg[18][24]  ( .D(n1063), .E(n766), .CP(n890), .CDN(n634), 
        .Q(\Storage[18][24] ) );
  EDFCNQD1 \Storage_reg[18][23]  ( .D(n1059), .E(n766), .CP(n890), .CDN(n634), 
        .Q(\Storage[18][23] ) );
  EDFCNQD1 \Storage_reg[18][22]  ( .D(n1055), .E(n767), .CP(n890), .CDN(n634), 
        .Q(\Storage[18][22] ) );
  EDFCNQD1 \Storage_reg[18][21]  ( .D(n1051), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][21] ) );
  EDFCNQD1 \Storage_reg[18][20]  ( .D(n1047), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][20] ) );
  EDFCNQD1 \Storage_reg[18][19]  ( .D(n1043), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][19] ) );
  EDFCNQD1 \Storage_reg[18][18]  ( .D(n1039), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][18] ) );
  EDFCNQD1 \Storage_reg[18][17]  ( .D(n1035), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][17] ) );
  EDFCNQD1 \Storage_reg[18][16]  ( .D(n1031), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][16] ) );
  EDFCNQD1 \Storage_reg[18][15]  ( .D(n1027), .E(n767), .CP(n891), .CDN(n634), 
        .Q(\Storage[18][15] ) );
  EDFCNQD1 \Storage_reg[18][14]  ( .D(n1023), .E(n767), .CP(n891), .CDN(n633), 
        .Q(\Storage[18][14] ) );
  EDFCNQD1 \Storage_reg[18][13]  ( .D(n1019), .E(n767), .CP(n891), .CDN(n633), 
        .Q(\Storage[18][13] ) );
  EDFCNQD1 \Storage_reg[18][12]  ( .D(n1015), .E(n768), .CP(n891), .CDN(n633), 
        .Q(\Storage[18][12] ) );
  EDFCNQD1 \Storage_reg[18][11]  ( .D(n1011), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][11] ) );
  EDFCNQD1 \Storage_reg[18][10]  ( .D(n1007), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][10] ) );
  EDFCNQD1 \Storage_reg[18][9]  ( .D(n1003), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][9] ) );
  EDFCNQD1 \Storage_reg[18][8]  ( .D(n999), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][8] ) );
  EDFCNQD1 \Storage_reg[18][7]  ( .D(n995), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][7] ) );
  EDFCNQD1 \Storage_reg[18][6]  ( .D(n991), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][6] ) );
  EDFCNQD1 \Storage_reg[18][5]  ( .D(n987), .E(n768), .CP(n892), .CDN(n633), 
        .Q(\Storage[18][5] ) );
  EDFCNQD1 \Storage_reg[18][4]  ( .D(n983), .E(n768), .CP(n892), .CDN(n632), 
        .Q(\Storage[18][4] ) );
  EDFCNQD1 \Storage_reg[18][3]  ( .D(n979), .E(n768), .CP(n892), .CDN(n632), 
        .Q(\Storage[18][3] ) );
  EDFCNQD1 \Storage_reg[18][2]  ( .D(n975), .E(N744), .CP(n892), .CDN(n632), 
        .Q(\Storage[18][2] ) );
  EDFCNQD1 \Storage_reg[18][1]  ( .D(n971), .E(N744), .CP(n893), .CDN(n632), 
        .Q(\Storage[18][1] ) );
  EDFCNQD1 \Storage_reg[18][0]  ( .D(n967), .E(N744), .CP(n893), .CDN(n632), 
        .Q(\Storage[18][0] ) );
  EDFCNQD1 \Storage_reg[17][32]  ( .D(n843), .E(n770), .CP(n893), .CDN(n632), 
        .Q(\Storage[17][32] ) );
  EDFCNQD1 \Storage_reg[17][31]  ( .D(n1091), .E(n770), .CP(n893), .CDN(n632), 
        .Q(\Storage[17][31] ) );
  EDFCNQD1 \Storage_reg[17][30]  ( .D(n1087), .E(n770), .CP(n893), .CDN(n632), 
        .Q(\Storage[17][30] ) );
  EDFCNQD1 \Storage_reg[17][29]  ( .D(n1083), .E(n770), .CP(n893), .CDN(n632), 
        .Q(\Storage[17][29] ) );
  EDFCNQD1 \Storage_reg[17][28]  ( .D(n1079), .E(n770), .CP(n893), .CDN(n632), 
        .Q(\Storage[17][28] ) );
  EDFCNQD1 \Storage_reg[17][27]  ( .D(n1075), .E(n770), .CP(n893), .CDN(n631), 
        .Q(\Storage[17][27] ) );
  EDFCNQD1 \Storage_reg[17][26]  ( .D(n1071), .E(n770), .CP(n893), .CDN(n631), 
        .Q(\Storage[17][26] ) );
  EDFCNQD1 \Storage_reg[17][25]  ( .D(n1067), .E(n770), .CP(n893), .CDN(n631), 
        .Q(\Storage[17][25] ) );
  EDFCNQD1 \Storage_reg[17][24]  ( .D(n1063), .E(n770), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][24] ) );
  EDFCNQD1 \Storage_reg[17][23]  ( .D(n1059), .E(n770), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][23] ) );
  EDFCNQD1 \Storage_reg[17][22]  ( .D(n1055), .E(n771), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][22] ) );
  EDFCNQD1 \Storage_reg[17][21]  ( .D(n1051), .E(n771), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][21] ) );
  EDFCNQD1 \Storage_reg[17][20]  ( .D(n1047), .E(n771), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][20] ) );
  EDFCNQD1 \Storage_reg[17][19]  ( .D(n1043), .E(n771), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][19] ) );
  EDFCNQD1 \Storage_reg[17][18]  ( .D(n1039), .E(n771), .CP(n894), .CDN(n631), 
        .Q(\Storage[17][18] ) );
  EDFCNQD1 \Storage_reg[17][17]  ( .D(n1035), .E(n771), .CP(n894), .CDN(n630), 
        .Q(\Storage[17][17] ) );
  EDFCNQD1 \Storage_reg[17][16]  ( .D(n1031), .E(n771), .CP(n894), .CDN(n630), 
        .Q(\Storage[17][16] ) );
  EDFCNQD1 \Storage_reg[17][15]  ( .D(n1027), .E(n771), .CP(n894), .CDN(n630), 
        .Q(\Storage[17][15] ) );
  EDFCNQD1 \Storage_reg[17][14]  ( .D(n1023), .E(n771), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][14] ) );
  EDFCNQD1 \Storage_reg[17][13]  ( .D(n1019), .E(n771), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][13] ) );
  EDFCNQD1 \Storage_reg[17][12]  ( .D(n1015), .E(n772), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][12] ) );
  EDFCNQD1 \Storage_reg[17][11]  ( .D(n1011), .E(n772), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][11] ) );
  EDFCNQD1 \Storage_reg[17][10]  ( .D(n1007), .E(n772), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][10] ) );
  EDFCNQD1 \Storage_reg[17][9]  ( .D(n1003), .E(n772), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][9] ) );
  EDFCNQD1 \Storage_reg[17][8]  ( .D(n999), .E(n772), .CP(n895), .CDN(n630), 
        .Q(\Storage[17][8] ) );
  EDFCNQD1 \Storage_reg[17][7]  ( .D(n995), .E(n772), .CP(n895), .CDN(n629), 
        .Q(\Storage[17][7] ) );
  EDFCNQD1 \Storage_reg[17][6]  ( .D(n991), .E(n772), .CP(n895), .CDN(n629), 
        .Q(\Storage[17][6] ) );
  EDFCNQD1 \Storage_reg[17][5]  ( .D(n987), .E(n772), .CP(n895), .CDN(n629), 
        .Q(\Storage[17][5] ) );
  EDFCNQD1 \Storage_reg[17][4]  ( .D(n983), .E(n772), .CP(n896), .CDN(n629), 
        .Q(\Storage[17][4] ) );
  EDFCNQD1 \Storage_reg[17][3]  ( .D(n979), .E(n772), .CP(n896), .CDN(n629), 
        .Q(\Storage[17][3] ) );
  EDFCNQD1 \Storage_reg[17][2]  ( .D(n975), .E(N711), .CP(n896), .CDN(n629), 
        .Q(\Storage[17][2] ) );
  EDFCNQD1 \Storage_reg[17][1]  ( .D(n971), .E(N711), .CP(n896), .CDN(n629), 
        .Q(\Storage[17][1] ) );
  EDFCNQD1 \Storage_reg[17][0]  ( .D(n967), .E(N711), .CP(n896), .CDN(n629), 
        .Q(\Storage[17][0] ) );
  EDFCNQD1 \Storage_reg[14][32]  ( .D(n843), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][32] ) );
  EDFCNQD1 \Storage_reg[14][31]  ( .D(n1091), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][31] ) );
  EDFCNQD1 \Storage_reg[14][30]  ( .D(n1087), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][30] ) );
  EDFCNQD1 \Storage_reg[14][29]  ( .D(n1083), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][29] ) );
  EDFCNQD1 \Storage_reg[14][28]  ( .D(n1079), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][28] ) );
  EDFCNQD1 \Storage_reg[14][27]  ( .D(n1075), .E(n782), .CP(n903), .CDN(n622), 
        .Q(\Storage[14][27] ) );
  EDFCNQD1 \Storage_reg[14][26]  ( .D(n1071), .E(n782), .CP(n903), .CDN(n621), 
        .Q(\Storage[14][26] ) );
  EDFCNQD1 \Storage_reg[14][25]  ( .D(n1067), .E(n782), .CP(n903), .CDN(n621), 
        .Q(\Storage[14][25] ) );
  EDFCNQD1 \Storage_reg[14][24]  ( .D(n1063), .E(n782), .CP(n903), .CDN(n621), 
        .Q(\Storage[14][24] ) );
  EDFCNQD1 \Storage_reg[14][23]  ( .D(n1059), .E(n782), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][23] ) );
  EDFCNQD1 \Storage_reg[14][22]  ( .D(n1055), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][22] ) );
  EDFCNQD1 \Storage_reg[14][21]  ( .D(n1051), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][21] ) );
  EDFCNQD1 \Storage_reg[14][20]  ( .D(n1047), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][20] ) );
  EDFCNQD1 \Storage_reg[14][19]  ( .D(n1043), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][19] ) );
  EDFCNQD1 \Storage_reg[14][18]  ( .D(n1039), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][18] ) );
  EDFCNQD1 \Storage_reg[14][17]  ( .D(n1035), .E(n783), .CP(n904), .CDN(n621), 
        .Q(\Storage[14][17] ) );
  EDFCNQD1 \Storage_reg[14][16]  ( .D(n1031), .E(n783), .CP(n904), .CDN(n620), 
        .Q(\Storage[14][16] ) );
  EDFCNQD1 \Storage_reg[14][15]  ( .D(n1027), .E(n783), .CP(n904), .CDN(n620), 
        .Q(\Storage[14][15] ) );
  EDFCNQD1 \Storage_reg[14][14]  ( .D(n1023), .E(n783), .CP(n904), .CDN(n620), 
        .Q(\Storage[14][14] ) );
  EDFCNQD1 \Storage_reg[14][13]  ( .D(n1019), .E(n783), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][13] ) );
  EDFCNQD1 \Storage_reg[14][12]  ( .D(n1015), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][12] ) );
  EDFCNQD1 \Storage_reg[14][11]  ( .D(n1011), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][11] ) );
  EDFCNQD1 \Storage_reg[14][10]  ( .D(n1007), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][10] ) );
  EDFCNQD1 \Storage_reg[14][9]  ( .D(n1003), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][9] ) );
  EDFCNQD1 \Storage_reg[14][8]  ( .D(n999), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][8] ) );
  EDFCNQD1 \Storage_reg[14][7]  ( .D(n995), .E(n784), .CP(n905), .CDN(n620), 
        .Q(\Storage[14][7] ) );
  EDFCNQD1 \Storage_reg[14][6]  ( .D(n991), .E(n784), .CP(n905), .CDN(n619), 
        .Q(\Storage[14][6] ) );
  EDFCNQD1 \Storage_reg[14][5]  ( .D(n987), .E(n784), .CP(n905), .CDN(n619), 
        .Q(\Storage[14][5] ) );
  EDFCNQD1 \Storage_reg[14][4]  ( .D(n983), .E(n784), .CP(n905), .CDN(n619), 
        .Q(\Storage[14][4] ) );
  EDFCNQD1 \Storage_reg[14][3]  ( .D(n979), .E(n784), .CP(n906), .CDN(n619), 
        .Q(\Storage[14][3] ) );
  EDFCNQD1 \Storage_reg[14][2]  ( .D(n975), .E(N612), .CP(n906), .CDN(n619), 
        .Q(\Storage[14][2] ) );
  EDFCNQD1 \Storage_reg[14][1]  ( .D(n971), .E(N612), .CP(n906), .CDN(n619), 
        .Q(\Storage[14][1] ) );
  EDFCNQD1 \Storage_reg[14][0]  ( .D(n967), .E(N612), .CP(n906), .CDN(n619), 
        .Q(\Storage[14][0] ) );
  EDFCNQD1 \Storage_reg[13][32]  ( .D(n843), .E(n786), .CP(n906), .CDN(n619), 
        .Q(\Storage[13][32] ) );
  EDFCNQD1 \Storage_reg[13][31]  ( .D(n1091), .E(n786), .CP(n906), .CDN(n619), 
        .Q(\Storage[13][31] ) );
  EDFCNQD1 \Storage_reg[13][30]  ( .D(n1087), .E(n786), .CP(n906), .CDN(n619), 
        .Q(\Storage[13][30] ) );
  EDFCNQD1 \Storage_reg[13][29]  ( .D(n1083), .E(n786), .CP(n906), .CDN(n618), 
        .Q(\Storage[13][29] ) );
  EDFCNQD1 \Storage_reg[13][28]  ( .D(n1079), .E(n786), .CP(n906), .CDN(n618), 
        .Q(\Storage[13][28] ) );
  EDFCNQD1 \Storage_reg[13][27]  ( .D(n1075), .E(n786), .CP(n906), .CDN(n618), 
        .Q(\Storage[13][27] ) );
  EDFCNQD1 \Storage_reg[13][26]  ( .D(n1071), .E(n786), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][26] ) );
  EDFCNQD1 \Storage_reg[13][25]  ( .D(n1067), .E(n786), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][25] ) );
  EDFCNQD1 \Storage_reg[13][24]  ( .D(n1063), .E(n786), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][24] ) );
  EDFCNQD1 \Storage_reg[13][23]  ( .D(n1059), .E(n786), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][23] ) );
  EDFCNQD1 \Storage_reg[13][22]  ( .D(n1055), .E(n787), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][22] ) );
  EDFCNQD1 \Storage_reg[13][21]  ( .D(n1051), .E(n787), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][21] ) );
  EDFCNQD1 \Storage_reg[13][20]  ( .D(n1047), .E(n787), .CP(n907), .CDN(n618), 
        .Q(\Storage[13][20] ) );
  EDFCNQD1 \Storage_reg[13][19]  ( .D(n1043), .E(n787), .CP(n907), .CDN(n617), 
        .Q(\Storage[13][19] ) );
  EDFCNQD1 \Storage_reg[13][18]  ( .D(n1039), .E(n787), .CP(n907), .CDN(n617), 
        .Q(\Storage[13][18] ) );
  EDFCNQD1 \Storage_reg[13][17]  ( .D(n1035), .E(n787), .CP(n907), .CDN(n617), 
        .Q(\Storage[13][17] ) );
  EDFCNQD1 \Storage_reg[13][16]  ( .D(n1031), .E(n787), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][16] ) );
  EDFCNQD1 \Storage_reg[13][15]  ( .D(n1027), .E(n787), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][15] ) );
  EDFCNQD1 \Storage_reg[13][14]  ( .D(n1023), .E(n787), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][14] ) );
  EDFCNQD1 \Storage_reg[13][13]  ( .D(n1019), .E(n787), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][13] ) );
  EDFCNQD1 \Storage_reg[13][12]  ( .D(n1015), .E(n788), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][12] ) );
  EDFCNQD1 \Storage_reg[13][11]  ( .D(n1011), .E(n788), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][11] ) );
  EDFCNQD1 \Storage_reg[13][10]  ( .D(n1007), .E(n788), .CP(n908), .CDN(n617), 
        .Q(\Storage[13][10] ) );
  EDFCNQD1 \Storage_reg[13][9]  ( .D(n1003), .E(n788), .CP(n908), .CDN(n616), 
        .Q(\Storage[13][9] ) );
  EDFCNQD1 \Storage_reg[13][8]  ( .D(n999), .E(n788), .CP(n908), .CDN(n616), 
        .Q(\Storage[13][8] ) );
  EDFCNQD1 \Storage_reg[13][7]  ( .D(n995), .E(n788), .CP(n908), .CDN(n616), 
        .Q(\Storage[13][7] ) );
  EDFCNQD1 \Storage_reg[13][6]  ( .D(n991), .E(n788), .CP(n918), .CDN(n616), 
        .Q(\Storage[13][6] ) );
  EDFCNQD1 \Storage_reg[13][5]  ( .D(n987), .E(n788), .CP(n934), .CDN(n616), 
        .Q(\Storage[13][5] ) );
  EDFCNQD1 \Storage_reg[13][4]  ( .D(n983), .E(n788), .CP(n933), .CDN(n616), 
        .Q(\Storage[13][4] ) );
  EDFCNQD1 \Storage_reg[13][3]  ( .D(n979), .E(n788), .CP(n932), .CDN(n616), 
        .Q(\Storage[13][3] ) );
  EDFCNQD1 \Storage_reg[13][2]  ( .D(n975), .E(N579), .CP(n931), .CDN(n616), 
        .Q(\Storage[13][2] ) );
  EDFCNQD1 \Storage_reg[13][1]  ( .D(n971), .E(N579), .CP(n930), .CDN(n616), 
        .Q(\Storage[13][1] ) );
  EDFCNQD1 \Storage_reg[13][0]  ( .D(n967), .E(N579), .CP(n929), .CDN(n616), 
        .Q(\Storage[13][0] ) );
  EDFCNQD1 \Storage_reg[10][32]  ( .D(n844), .E(n798), .CP(ClockW), .CDN(n609), 
        .Q(\Storage[10][32] ) );
  EDFCNQD1 \Storage_reg[10][31]  ( .D(n1091), .E(n798), .CP(n942), .CDN(n609), 
        .Q(\Storage[10][31] ) );
  EDFCNQD1 \Storage_reg[10][30]  ( .D(n1087), .E(n798), .CP(n955), .CDN(n609), 
        .Q(\Storage[10][30] ) );
  EDFCNQD1 \Storage_reg[10][29]  ( .D(n1083), .E(n798), .CP(n957), .CDN(n609), 
        .Q(\Storage[10][29] ) );
  EDFCNQD1 \Storage_reg[10][28]  ( .D(n1079), .E(n798), .CP(n951), .CDN(n608), 
        .Q(\Storage[10][28] ) );
  EDFCNQD1 \Storage_reg[10][27]  ( .D(n1075), .E(n798), .CP(n952), .CDN(n608), 
        .Q(\Storage[10][27] ) );
  EDFCNQD1 \Storage_reg[10][26]  ( .D(n1071), .E(n798), .CP(n953), .CDN(n608), 
        .Q(\Storage[10][26] ) );
  EDFCNQD1 \Storage_reg[10][25]  ( .D(n1067), .E(n798), .CP(n929), .CDN(n608), 
        .Q(\Storage[10][25] ) );
  EDFCNQD1 \Storage_reg[10][24]  ( .D(n1063), .E(n798), .CP(n918), .CDN(n608), 
        .Q(\Storage[10][24] ) );
  EDFCNQD1 \Storage_reg[10][23]  ( .D(n1059), .E(n798), .CP(n961), .CDN(n608), 
        .Q(\Storage[10][23] ) );
  EDFCNQD1 \Storage_reg[10][22]  ( .D(n1055), .E(n799), .CP(n940), .CDN(n608), 
        .Q(\Storage[10][22] ) );
  EDFCNQD1 \Storage_reg[10][21]  ( .D(n1051), .E(n799), .CP(n939), .CDN(n608), 
        .Q(\Storage[10][21] ) );
  EDFCNQD1 \Storage_reg[10][20]  ( .D(n1047), .E(n799), .CP(n938), .CDN(n608), 
        .Q(\Storage[10][20] ) );
  EDFCNQD1 \Storage_reg[10][19]  ( .D(n1043), .E(n799), .CP(n937), .CDN(n608), 
        .Q(\Storage[10][19] ) );
  EDFCNQD1 \Storage_reg[10][18]  ( .D(n1039), .E(n799), .CP(n936), .CDN(n607), 
        .Q(\Storage[10][18] ) );
  EDFCNQD1 \Storage_reg[10][17]  ( .D(n1035), .E(n799), .CP(n935), .CDN(n607), 
        .Q(\Storage[10][17] ) );
  EDFCNQD1 \Storage_reg[10][16]  ( .D(n1031), .E(n799), .CP(n941), .CDN(n607), 
        .Q(\Storage[10][16] ) );
  EDFCNQD1 \Storage_reg[10][15]  ( .D(n1027), .E(n799), .CP(n926), .CDN(n607), 
        .Q(\Storage[10][15] ) );
  EDFCNQD1 \Storage_reg[10][14]  ( .D(n1023), .E(n799), .CP(n919), .CDN(n607), 
        .Q(\Storage[10][14] ) );
  EDFCNQD1 \Storage_reg[10][13]  ( .D(n1019), .E(n799), .CP(n930), .CDN(n607), 
        .Q(\Storage[10][13] ) );
  EDFCNQD1 \Storage_reg[10][12]  ( .D(n1015), .E(n800), .CP(n931), .CDN(n607), 
        .Q(\Storage[10][12] ) );
  EDFCNQD1 \Storage_reg[10][11]  ( .D(n1011), .E(n800), .CP(n932), .CDN(n607), 
        .Q(\Storage[10][11] ) );
  EDFCNQD1 \Storage_reg[10][10]  ( .D(n1007), .E(n800), .CP(n933), .CDN(n607), 
        .Q(\Storage[10][10] ) );
  EDFCNQD1 \Storage_reg[10][9]  ( .D(n1003), .E(n800), .CP(n934), .CDN(n607), 
        .Q(\Storage[10][9] ) );
  EDFCNQD1 \Storage_reg[10][8]  ( .D(n999), .E(n800), .CP(n959), .CDN(n606), 
        .Q(\Storage[10][8] ) );
  EDFCNQD1 \Storage_reg[10][7]  ( .D(n995), .E(n800), .CP(n928), .CDN(n606), 
        .Q(\Storage[10][7] ) );
  EDFCNQD1 \Storage_reg[10][6]  ( .D(n991), .E(n800), .CP(n927), .CDN(n606), 
        .Q(\Storage[10][6] ) );
  EDFCNQD1 \Storage_reg[10][5]  ( .D(n987), .E(n800), .CP(n943), .CDN(n606), 
        .Q(\Storage[10][5] ) );
  EDFCNQD1 \Storage_reg[10][4]  ( .D(n983), .E(n800), .CP(n957), .CDN(n606), 
        .Q(\Storage[10][4] ) );
  EDFCNQD1 \Storage_reg[10][3]  ( .D(n979), .E(n800), .CP(n915), .CDN(n606), 
        .Q(\Storage[10][3] ) );
  EDFCNQD1 \Storage_reg[10][2]  ( .D(n975), .E(N480), .CP(n959), .CDN(n606), 
        .Q(\Storage[10][2] ) );
  EDFCNQD1 \Storage_reg[10][1]  ( .D(n971), .E(N480), .CP(n962), .CDN(n606), 
        .Q(\Storage[10][1] ) );
  EDFCNQD1 \Storage_reg[10][0]  ( .D(n967), .E(N480), .CP(n944), .CDN(n606), 
        .Q(\Storage[10][0] ) );
  EDFCNQD1 \Storage_reg[9][32]  ( .D(n844), .E(n802), .CP(n945), .CDN(n606), 
        .Q(\Storage[9][32] ) );
  EDFCNQD1 \Storage_reg[9][31]  ( .D(n1091), .E(n802), .CP(n946), .CDN(n605), 
        .Q(\Storage[9][31] ) );
  EDFCNQD1 \Storage_reg[9][30]  ( .D(n1087), .E(n802), .CP(n941), .CDN(n605), 
        .Q(\Storage[9][30] ) );
  EDFCNQD1 \Storage_reg[9][29]  ( .D(n1083), .E(n802), .CP(n942), .CDN(n605), 
        .Q(\Storage[9][29] ) );
  EDFCNQD1 \Storage_reg[9][28]  ( .D(n1079), .E(n802), .CP(n961), .CDN(n605), 
        .Q(\Storage[9][28] ) );
  EDFCNQD1 \Storage_reg[9][27]  ( .D(n1075), .E(n802), .CP(n960), .CDN(n605), 
        .Q(\Storage[9][27] ) );
  EDFCNQD1 \Storage_reg[9][26]  ( .D(n1071), .E(n802), .CP(ClockW), .CDN(n605), 
        .Q(\Storage[9][26] ) );
  EDFCNQD1 \Storage_reg[9][25]  ( .D(n1067), .E(n802), .CP(n962), .CDN(n605), 
        .Q(\Storage[9][25] ) );
  EDFCNQD1 \Storage_reg[9][24]  ( .D(n1063), .E(n802), .CP(n946), .CDN(n605), 
        .Q(\Storage[9][24] ) );
  EDFCNQD1 \Storage_reg[9][23]  ( .D(n1059), .E(n802), .CP(n945), .CDN(n605), 
        .Q(\Storage[9][23] ) );
  EDFCNQD1 \Storage_reg[9][22]  ( .D(n1055), .E(n803), .CP(n944), .CDN(n605), 
        .Q(\Storage[9][22] ) );
  EDFCNQD1 \Storage_reg[9][21]  ( .D(n1051), .E(n803), .CP(n943), .CDN(n604), 
        .Q(\Storage[9][21] ) );
  EDFCNQD1 \Storage_reg[9][20]  ( .D(n1047), .E(n803), .CP(n942), .CDN(n604), 
        .Q(\Storage[9][20] ) );
  EDFCNQD1 \Storage_reg[9][19]  ( .D(n1043), .E(n803), .CP(n941), .CDN(n604), 
        .Q(\Storage[9][19] ) );
  EDFCNQD1 \Storage_reg[9][18]  ( .D(n1039), .E(n803), .CP(n950), .CDN(n604), 
        .Q(\Storage[9][18] ) );
  EDFCNQD1 \Storage_reg[9][17]  ( .D(n1035), .E(n803), .CP(n915), .CDN(n604), 
        .Q(\Storage[9][17] ) );
  EDFCNQD1 \Storage_reg[9][16]  ( .D(n1031), .E(n803), .CP(n926), .CDN(n604), 
        .Q(\Storage[9][16] ) );
  EDFCNQD1 \Storage_reg[9][15]  ( .D(n1027), .E(n803), .CP(n914), .CDN(n604), 
        .Q(\Storage[9][15] ) );
  EDFCNQD1 \Storage_reg[9][14]  ( .D(n1023), .E(n803), .CP(n913), .CDN(n604), 
        .Q(\Storage[9][14] ) );
  EDFCNQD1 \Storage_reg[9][13]  ( .D(n1019), .E(n803), .CP(n944), .CDN(n604), 
        .Q(\Storage[9][13] ) );
  EDFCNQD1 \Storage_reg[9][12]  ( .D(n1015), .E(n804), .CP(n922), .CDN(n604), 
        .Q(\Storage[9][12] ) );
  EDFCNQD1 \Storage_reg[9][11]  ( .D(n1011), .E(n804), .CP(n940), .CDN(n603), 
        .Q(\Storage[9][11] ) );
  EDFCNQD1 \Storage_reg[9][10]  ( .D(n1007), .E(n804), .CP(n927), .CDN(n603), 
        .Q(\Storage[9][10] ) );
  EDFCNQD1 \Storage_reg[9][9]  ( .D(n1003), .E(n804), .CP(n921), .CDN(n603), 
        .Q(\Storage[9][9] ) );
  EDFCNQD1 \Storage_reg[9][8]  ( .D(n999), .E(n804), .CP(n956), .CDN(n603), 
        .Q(\Storage[9][8] ) );
  EDFCNQD1 \Storage_reg[9][7]  ( .D(n995), .E(n804), .CP(n957), .CDN(n603), 
        .Q(\Storage[9][7] ) );
  EDFCNQD1 \Storage_reg[9][6]  ( .D(n991), .E(n804), .CP(n846), .CDN(n603), 
        .Q(\Storage[9][6] ) );
  EDFCNQD1 \Storage_reg[9][5]  ( .D(n987), .E(n804), .CP(n948), .CDN(n603), 
        .Q(\Storage[9][5] ) );
  EDFCNQD1 \Storage_reg[9][4]  ( .D(n983), .E(n804), .CP(n949), .CDN(n603), 
        .Q(\Storage[9][4] ) );
  EDFCNQD1 \Storage_reg[9][3]  ( .D(n979), .E(n804), .CP(n952), .CDN(n603), 
        .Q(\Storage[9][3] ) );
  EDFCNQD1 \Storage_reg[9][2]  ( .D(n975), .E(N447), .CP(n951), .CDN(n603), 
        .Q(\Storage[9][2] ) );
  EDFCNQD1 \Storage_reg[9][1]  ( .D(n971), .E(N447), .CP(n953), .CDN(n602), 
        .Q(\Storage[9][1] ) );
  EDFCNQD1 \Storage_reg[9][0]  ( .D(n967), .E(N447), .CP(n955), .CDN(n602), 
        .Q(\Storage[9][0] ) );
  EDFCNQD1 \Storage_reg[6][32]  ( .D(n844), .E(n814), .CP(n954), .CDN(n713), 
        .Q(\Storage[6][32] ) );
  EDFCNQD1 \Storage_reg[6][31]  ( .D(n1090), .E(n814), .CP(n924), .CDN(n686), 
        .Q(\Storage[6][31] ) );
  EDFCNQD1 \Storage_reg[6][30]  ( .D(n1086), .E(n814), .CP(n951), .CDN(n710), 
        .Q(\Storage[6][30] ) );
  EDFCNQD1 \Storage_reg[6][29]  ( .D(n1082), .E(n814), .CP(n952), .CDN(n700), 
        .Q(\Storage[6][29] ) );
  EDFCNQD1 \Storage_reg[6][28]  ( .D(n1078), .E(n814), .CP(n949), .CDN(n702), 
        .Q(\Storage[6][28] ) );
  EDFCNQD1 \Storage_reg[6][27]  ( .D(n1074), .E(n814), .CP(n931), .CDN(n711), 
        .Q(\Storage[6][27] ) );
  EDFCNQD1 \Storage_reg[6][26]  ( .D(n1070), .E(n814), .CP(n935), .CDN(n712), 
        .Q(\Storage[6][26] ) );
  EDFCNQD1 \Storage_reg[6][25]  ( .D(n1066), .E(n814), .CP(n956), .CDN(n694), 
        .Q(\Storage[6][25] ) );
  EDFCNQD1 \Storage_reg[6][24]  ( .D(n1062), .E(n814), .CP(n923), .CDN(n693), 
        .Q(\Storage[6][24] ) );
  EDFCNQD1 \Storage_reg[6][23]  ( .D(n1058), .E(n814), .CP(n958), .CDN(n703), 
        .Q(\Storage[6][23] ) );
  EDFCNQD1 \Storage_reg[6][22]  ( .D(n1054), .E(n815), .CP(n932), .CDN(n704), 
        .Q(\Storage[6][22] ) );
  EDFCNQD1 \Storage_reg[6][21]  ( .D(n1050), .E(n815), .CP(n933), .CDN(n595), 
        .Q(\Storage[6][21] ) );
  EDFCNQD1 \Storage_reg[6][20]  ( .D(n1046), .E(n815), .CP(n934), .CDN(n596), 
        .Q(\Storage[6][20] ) );
  EDFCNQD1 \Storage_reg[6][19]  ( .D(n1042), .E(n815), .CP(n929), .CDN(n679), 
        .Q(\Storage[6][19] ) );
  EDFCNQD1 \Storage_reg[6][18]  ( .D(n1038), .E(n815), .CP(n930), .CDN(n708), 
        .Q(\Storage[6][18] ) );
  EDFCNQD1 \Storage_reg[6][17]  ( .D(n1034), .E(n815), .CP(n940), .CDN(n709), 
        .Q(\Storage[6][17] ) );
  EDFCNQD1 \Storage_reg[6][16]  ( .D(n1030), .E(n815), .CP(n959), .CDN(n705), 
        .Q(\Storage[6][16] ) );
  EDFCNQD1 \Storage_reg[6][15]  ( .D(n1026), .E(n815), .CP(n962), .CDN(n706), 
        .Q(\Storage[6][15] ) );
  EDFCNQD1 \Storage_reg[6][14]  ( .D(n1022), .E(n815), .CP(n946), .CDN(n707), 
        .Q(\Storage[6][14] ) );
  EDFCNQD1 \Storage_reg[6][13]  ( .D(n1018), .E(n815), .CP(n945), .CDN(n710), 
        .Q(\Storage[6][13] ) );
  EDFCNQD1 \Storage_reg[6][12]  ( .D(n1014), .E(n816), .CP(n944), .CDN(n701), 
        .Q(\Storage[6][12] ) );
  EDFCNQD1 \Storage_reg[6][11]  ( .D(n1010), .E(n816), .CP(n943), .CDN(n692), 
        .Q(\Storage[6][11] ) );
  EDFCNQD1 \Storage_reg[6][10]  ( .D(n1006), .E(n816), .CP(n942), .CDN(n680), 
        .Q(\Storage[6][10] ) );
  EDFCNQD1 \Storage_reg[6][9]  ( .D(n1002), .E(n816), .CP(n941), .CDN(n685), 
        .Q(\Storage[6][9] ) );
  EDFCNQD1 \Storage_reg[6][8]  ( .D(n998), .E(n816), .CP(n961), .CDN(n697), 
        .Q(\Storage[6][8] ) );
  EDFCNQD1 \Storage_reg[6][7]  ( .D(n994), .E(n816), .CP(n938), .CDN(n698), 
        .Q(\Storage[6][7] ) );
  EDFCNQD1 \Storage_reg[6][6]  ( .D(n990), .E(n816), .CP(n922), .CDN(n709), 
        .Q(\Storage[6][6] ) );
  EDFCNQD1 \Storage_reg[6][5]  ( .D(n986), .E(n816), .CP(n960), .CDN(n679), 
        .Q(\Storage[6][5] ) );
  EDFCNQD1 \Storage_reg[6][4]  ( .D(n982), .E(n816), .CP(n934), .CDN(n699), 
        .Q(\Storage[6][4] ) );
  EDFCNQD1 \Storage_reg[6][3]  ( .D(n978), .E(n816), .CP(n933), .CDN(n596), 
        .Q(\Storage[6][3] ) );
  EDFCNQD1 \Storage_reg[6][2]  ( .D(n974), .E(N348), .CP(n932), .CDN(n696), 
        .Q(\Storage[6][2] ) );
  EDFCNQD1 \Storage_reg[6][1]  ( .D(n970), .E(N348), .CP(n931), .CDN(n695), 
        .Q(\Storage[6][1] ) );
  EDFCNQD1 \Storage_reg[6][0]  ( .D(n966), .E(N348), .CP(n930), .CDN(n690), 
        .Q(\Storage[6][0] ) );
  EDFCNQD1 \Storage_reg[5][32]  ( .D(n844), .E(n818), .CP(n929), .CDN(n596), 
        .Q(\Storage[5][32] ) );
  EDFCNQD1 \Storage_reg[5][31]  ( .D(n1090), .E(n818), .CP(n939), .CDN(n684), 
        .Q(\Storage[5][31] ) );
  EDFCNQD1 \Storage_reg[5][30]  ( .D(n1086), .E(n818), .CP(n956), .CDN(n683), 
        .Q(\Storage[5][30] ) );
  EDFCNQD1 \Storage_reg[5][29]  ( .D(n1082), .E(n818), .CP(n960), .CDN(n682), 
        .Q(\Storage[5][29] ) );
  EDFCNQD1 \Storage_reg[5][28]  ( .D(n1078), .E(n818), .CP(n937), .CDN(n681), 
        .Q(\Storage[5][28] ) );
  EDFCNQD1 \Storage_reg[5][27]  ( .D(n1074), .E(n818), .CP(n936), .CDN(n685), 
        .Q(\Storage[5][27] ) );
  EDFCNQD1 \Storage_reg[5][26]  ( .D(n1070), .E(n818), .CP(n935), .CDN(n686), 
        .Q(\Storage[5][26] ) );
  EDFCNQD1 \Storage_reg[5][25]  ( .D(n1066), .E(n818), .CP(n928), .CDN(n688), 
        .Q(\Storage[5][25] ) );
  EDFCNQD1 \Storage_reg[5][24]  ( .D(n1062), .E(n818), .CP(n927), .CDN(n687), 
        .Q(\Storage[5][24] ) );
  EDFCNQD1 \Storage_reg[5][23]  ( .D(n1058), .E(n818), .CP(n926), .CDN(n701), 
        .Q(\Storage[5][23] ) );
  EDFCNQD1 \Storage_reg[5][22]  ( .D(n1054), .E(n819), .CP(n923), .CDN(n689), 
        .Q(\Storage[5][22] ) );
  EDFCNQD1 \Storage_reg[5][21]  ( .D(n1050), .E(n819), .CP(n958), .CDN(n693), 
        .Q(\Storage[5][21] ) );
  EDFCNQD1 \Storage_reg[5][20]  ( .D(n1046), .E(n819), .CP(n933), .CDN(n712), 
        .Q(\Storage[5][20] ) );
  EDFCNQD1 \Storage_reg[5][19]  ( .D(n1042), .E(n819), .CP(n934), .CDN(n702), 
        .Q(\Storage[5][19] ) );
  EDFCNQD1 \Storage_reg[5][18]  ( .D(n1038), .E(n819), .CP(n922), .CDN(n713), 
        .Q(\Storage[5][18] ) );
  EDFCNQD1 \Storage_reg[5][17]  ( .D(n1034), .E(n819), .CP(n846), .CDN(n687), 
        .Q(\Storage[5][17] ) );
  EDFCNQD1 \Storage_reg[5][16]  ( .D(n1030), .E(n819), .CP(n940), .CDN(n711), 
        .Q(\Storage[5][16] ) );
  EDFCNQD1 \Storage_reg[5][15]  ( .D(n1026), .E(n819), .CP(n923), .CDN(n704), 
        .Q(\Storage[5][15] ) );
  EDFCNQD1 \Storage_reg[5][14]  ( .D(n1022), .E(n819), .CP(n935), .CDN(n703), 
        .Q(\Storage[5][14] ) );
  EDFCNQD1 \Storage_reg[5][13]  ( .D(n1018), .E(n819), .CP(n961), .CDN(n707), 
        .Q(\Storage[5][13] ) );
  EDFCNQD1 \Storage_reg[5][12]  ( .D(n1014), .E(n820), .CP(n923), .CDN(n679), 
        .Q(\Storage[5][12] ) );
  EDFCNQD1 \Storage_reg[5][11]  ( .D(n1010), .E(n820), .CP(n929), .CDN(n710), 
        .Q(\Storage[5][11] ) );
  EDFCNQD1 \Storage_reg[5][10]  ( .D(n1006), .E(n820), .CP(n956), .CDN(n705), 
        .Q(\Storage[5][10] ) );
  EDFCNQD1 \Storage_reg[5][9]  ( .D(n1002), .E(n820), .CP(n946), .CDN(n595), 
        .Q(\Storage[5][9] ) );
  EDFCNQD1 \Storage_reg[5][8]  ( .D(n998), .E(n820), .CP(n954), .CDN(n695), 
        .Q(\Storage[5][8] ) );
  EDFCNQD1 \Storage_reg[5][7]  ( .D(n994), .E(n820), .CP(ClockW), .CDN(n700), 
        .Q(\Storage[5][7] ) );
  EDFCNQD1 \Storage_reg[5][6]  ( .D(n990), .E(n820), .CP(n948), .CDN(n708), 
        .Q(\Storage[5][6] ) );
  EDFCNQD1 \Storage_reg[5][5]  ( .D(n986), .E(n820), .CP(n949), .CDN(n709), 
        .Q(\Storage[5][5] ) );
  EDFCNQD1 \Storage_reg[5][4]  ( .D(n982), .E(n820), .CP(n952), .CDN(n706), 
        .Q(\Storage[5][4] ) );
  EDFCNQD1 \Storage_reg[5][3]  ( .D(n978), .E(n820), .CP(n948), .CDN(n712), 
        .Q(\Storage[5][3] ) );
  EDFCNQD1 \Storage_reg[5][2]  ( .D(n974), .E(N315), .CP(n954), .CDN(n596), 
        .Q(\Storage[5][2] ) );
  EDFCNQD1 \Storage_reg[5][1]  ( .D(n970), .E(N315), .CP(n955), .CDN(n689), 
        .Q(\Storage[5][1] ) );
  EDFCNQD1 \Storage_reg[5][0]  ( .D(n966), .E(N315), .CP(n927), .CDN(n679), 
        .Q(\Storage[5][0] ) );
  EDFCNQD1 \Storage_reg[2][32]  ( .D(n844), .E(n830), .CP(n914), .CDN(n595), 
        .Q(\Storage[2][32] ) );
  EDFCNQD1 \Storage_reg[2][31]  ( .D(n1090), .E(n830), .CP(n918), .CDN(n708), 
        .Q(\Storage[2][31] ) );
  EDFCNQD1 \Storage_reg[2][30]  ( .D(n1086), .E(n830), .CP(n949), .CDN(n688), 
        .Q(\Storage[2][30] ) );
  EDFCNQD1 \Storage_reg[2][29]  ( .D(n1082), .E(n830), .CP(n938), .CDN(n687), 
        .Q(\Storage[2][29] ) );
  EDFCNQD1 \Storage_reg[2][28]  ( .D(n1078), .E(n830), .CP(n936), .CDN(n697), 
        .Q(\Storage[2][28] ) );
  EDFCNQD1 \Storage_reg[2][27]  ( .D(n1074), .E(n830), .CP(n915), .CDN(n702), 
        .Q(\Storage[2][27] ) );
  EDFCNQD1 \Storage_reg[2][26]  ( .D(n1070), .E(n830), .CP(n920), .CDN(n713), 
        .Q(\Storage[2][26] ) );
  EDFCNQD1 \Storage_reg[2][25]  ( .D(n1066), .E(n830), .CP(n917), .CDN(n711), 
        .Q(\Storage[2][25] ) );
  EDFCNQD1 \Storage_reg[2][24]  ( .D(n1062), .E(n830), .CP(n925), .CDN(n712), 
        .Q(\Storage[2][24] ) );
  EDFCNQD1 \Storage_reg[2][23]  ( .D(n1058), .E(n830), .CP(n931), .CDN(n703), 
        .Q(\Storage[2][23] ) );
  EDFCNQD1 \Storage_reg[2][22]  ( .D(n1054), .E(n831), .CP(n937), .CDN(n680), 
        .Q(\Storage[2][22] ) );
  EDFCNQD1 \Storage_reg[2][21]  ( .D(n1050), .E(n831), .CP(n926), .CDN(n707), 
        .Q(\Storage[2][21] ) );
  EDFCNQD1 \Storage_reg[2][20]  ( .D(n1046), .E(n831), .CP(n921), .CDN(n706), 
        .Q(\Storage[2][20] ) );
  EDFCNQD1 \Storage_reg[2][19]  ( .D(n1042), .E(n831), .CP(n940), .CDN(n596), 
        .Q(\Storage[2][19] ) );
  EDFCNQD1 \Storage_reg[2][18]  ( .D(n1038), .E(n831), .CP(n944), .CDN(n679), 
        .Q(\Storage[2][18] ) );
  EDFCNQD1 \Storage_reg[2][17]  ( .D(n1034), .E(n831), .CP(n929), .CDN(n700), 
        .Q(\Storage[2][17] ) );
  EDFCNQD1 \Storage_reg[2][16]  ( .D(n1030), .E(n831), .CP(n930), .CDN(n691), 
        .Q(\Storage[2][16] ) );
  EDFCNQD1 \Storage_reg[2][15]  ( .D(n1026), .E(n831), .CP(n931), .CDN(n681), 
        .Q(\Storage[2][15] ) );
  EDFCNQD1 \Storage_reg[2][14]  ( .D(n1022), .E(n831), .CP(n935), .CDN(n678), 
        .Q(\Storage[2][14] ) );
  EDFCNQD1 \Storage_reg[2][13]  ( .D(n1018), .E(n831), .CP(n936), .CDN(n684), 
        .Q(\Storage[2][13] ) );
  EDFCNQD1 \Storage_reg[2][12]  ( .D(n1014), .E(n832), .CP(n937), .CDN(n694), 
        .Q(\Storage[2][12] ) );
  EDFCNQD1 \Storage_reg[2][11]  ( .D(n1010), .E(n832), .CP(n938), .CDN(n705), 
        .Q(\Storage[2][11] ) );
  EDFCNQD1 \Storage_reg[2][10]  ( .D(n1006), .E(n832), .CP(n939), .CDN(n697), 
        .Q(\Storage[2][10] ) );
  EDFCNQD1 \Storage_reg[2][9]  ( .D(n1002), .E(n832), .CP(n940), .CDN(n682), 
        .Q(\Storage[2][9] ) );
  EDFCNQD1 \Storage_reg[2][8]  ( .D(n998), .E(n832), .CP(n919), .CDN(n699), 
        .Q(\Storage[2][8] ) );
  EDFCNQD1 \Storage_reg[2][7]  ( .D(n994), .E(n832), .CP(n960), .CDN(n687), 
        .Q(\Storage[2][7] ) );
  EDFCNQD1 \Storage_reg[2][6]  ( .D(n990), .E(n832), .CP(n934), .CDN(n688), 
        .Q(\Storage[2][6] ) );
  EDFCNQD1 \Storage_reg[2][5]  ( .D(n986), .E(n832), .CP(n933), .CDN(n713), 
        .Q(\Storage[2][5] ) );
  EDFCNQD1 \Storage_reg[2][4]  ( .D(n982), .E(n832), .CP(n932), .CDN(n698), 
        .Q(\Storage[2][4] ) );
  EDFCNQD1 \Storage_reg[2][3]  ( .D(n978), .E(n832), .CP(n931), .CDN(n693), 
        .Q(\Storage[2][3] ) );
  EDFCNQD1 \Storage_reg[2][2]  ( .D(n974), .E(N216), .CP(n930), .CDN(n692), 
        .Q(\Storage[2][2] ) );
  EDFCNQD1 \Storage_reg[2][1]  ( .D(n970), .E(N216), .CP(n929), .CDN(n691), 
        .Q(\Storage[2][1] ) );
  EDFCNQD1 \Storage_reg[2][0]  ( .D(n966), .E(N216), .CP(n961), .CDN(n702), 
        .Q(\Storage[2][0] ) );
  EDFCNQD1 \Storage_reg[1][32]  ( .D(N85), .E(n834), .CP(n937), .CDN(n683), 
        .Q(\Storage[1][32] ) );
  EDFCNQD1 \Storage_reg[1][31]  ( .D(n1090), .E(n834), .CP(n936), .CDN(n690), 
        .Q(\Storage[1][31] ) );
  EDFCNQD1 \Storage_reg[1][30]  ( .D(n1086), .E(n834), .CP(n943), .CDN(n689), 
        .Q(\Storage[1][30] ) );
  EDFCNQD1 \Storage_reg[1][29]  ( .D(n1082), .E(n834), .CP(n942), .CDN(n685), 
        .Q(\Storage[1][29] ) );
  EDFCNQD1 \Storage_reg[1][28]  ( .D(n1078), .E(n834), .CP(n941), .CDN(n686), 
        .Q(\Storage[1][28] ) );
  EDFCNQD1 \Storage_reg[1][27]  ( .D(n1074), .E(n834), .CP(n946), .CDN(n696), 
        .Q(\Storage[1][27] ) );
  EDFCNQD1 \Storage_reg[1][26]  ( .D(n1070), .E(n834), .CP(n945), .CDN(n695), 
        .Q(\Storage[1][26] ) );
  EDFCNQD1 \Storage_reg[1][25]  ( .D(n1066), .E(n834), .CP(n944), .CDN(n708), 
        .Q(\Storage[1][25] ) );
  EDFCNQD1 \Storage_reg[1][24]  ( .D(n1062), .E(n834), .CP(n939), .CDN(n4), 
        .Q(\Storage[1][24] ) );
  EDFCNQD1 \Storage_reg[1][23]  ( .D(n1058), .E(n834), .CP(n938), .CDN(n711), 
        .Q(\Storage[1][23] ) );
  EDFCNQD1 \Storage_reg[1][22]  ( .D(n1054), .E(n835), .CP(n958), .CDN(n712), 
        .Q(\Storage[1][22] ) );
  EDFCNQD1 \Storage_reg[1][21]  ( .D(n1050), .E(n835), .CP(n918), .CDN(n704), 
        .Q(\Storage[1][21] ) );
  EDFCNQD1 \Storage_reg[1][20]  ( .D(n1046), .E(n835), .CP(n935), .CDN(n703), 
        .Q(\Storage[1][20] ) );
  EDFCNQD1 \Storage_reg[1][19]  ( .D(n1042), .E(n835), .CP(n959), .CDN(n595), 
        .Q(\Storage[1][19] ) );
  EDFCNQD1 \Storage_reg[1][18]  ( .D(n1038), .E(n835), .CP(n928), .CDN(n709), 
        .Q(\Storage[1][18] ) );
  EDFCNQD1 \Storage_reg[1][17]  ( .D(n1034), .E(n835), .CP(n927), .CDN(n701), 
        .Q(\Storage[1][17] ) );
  EDFCNQD1 \Storage_reg[1][16]  ( .D(n1030), .E(n835), .CP(n926), .CDN(n710), 
        .Q(\Storage[1][16] ) );
  EDFCNQD1 \Storage_reg[1][15]  ( .D(n1026), .E(n835), .CP(n925), .CDN(n601), 
        .Q(\Storage[1][15] ) );
  EDFCNQD1 \Storage_reg[1][14]  ( .D(n1022), .E(n835), .CP(n924), .CDN(n601), 
        .Q(\Storage[1][14] ) );
  EDFCNQD1 \Storage_reg[1][13]  ( .D(n1018), .E(n835), .CP(n923), .CDN(n601), 
        .Q(\Storage[1][13] ) );
  EDFCNQD1 \Storage_reg[1][12]  ( .D(n1014), .E(n836), .CP(n921), .CDN(n601), 
        .Q(\Storage[1][12] ) );
  EDFCNQD1 \Storage_reg[1][11]  ( .D(n1010), .E(n836), .CP(n920), .CDN(n601), 
        .Q(\Storage[1][11] ) );
  EDFCNQD1 \Storage_reg[1][10]  ( .D(n1006), .E(n836), .CP(n954), .CDN(n601), 
        .Q(\Storage[1][10] ) );
  EDFCNQD1 \Storage_reg[1][9]  ( .D(n1002), .E(n836), .CP(n916), .CDN(n601), 
        .Q(\Storage[1][9] ) );
  EDFCNQD1 \Storage_reg[1][8]  ( .D(n998), .E(n836), .CP(n915), .CDN(n601), 
        .Q(\Storage[1][8] ) );
  EDFCNQD1 \Storage_reg[1][7]  ( .D(n994), .E(n836), .CP(n914), .CDN(n601), 
        .Q(\Storage[1][7] ) );
  EDFCNQD1 \Storage_reg[1][6]  ( .D(n990), .E(n836), .CP(n913), .CDN(n601), 
        .Q(\Storage[1][6] ) );
  EDFCNQD1 \Storage_reg[1][5]  ( .D(n986), .E(n836), .CP(n958), .CDN(n600), 
        .Q(\Storage[1][5] ) );
  EDFCNQD1 \Storage_reg[1][4]  ( .D(n982), .E(n836), .CP(n925), .CDN(n600), 
        .Q(\Storage[1][4] ) );
  EDFCNQD1 \Storage_reg[1][3]  ( .D(n978), .E(n836), .CP(n922), .CDN(n600), 
        .Q(\Storage[1][3] ) );
  EDFCNQD1 \Storage_reg[1][2]  ( .D(n974), .E(N183), .CP(n948), .CDN(n600), 
        .Q(\Storage[1][2] ) );
  EDFCNQD1 \Storage_reg[1][1]  ( .D(n970), .E(N183), .CP(n952), .CDN(n600), 
        .Q(\Storage[1][1] ) );
  EDFCNQD1 \Storage_reg[1][0]  ( .D(n966), .E(N183), .CP(n941), .CDN(n600), 
        .Q(\Storage[1][0] ) );
  EDFCNQD1 \Storage_reg[0][5]  ( .D(n986), .E(n840), .CP(n937), .CDN(n597), 
        .Q(\Storage[0][5] ) );
  EDFCNQD1 \Storage_reg[0][4]  ( .D(n982), .E(n840), .CP(n945), .CDN(n597), 
        .Q(\Storage[0][4] ) );
  EDFCNQD1 \Storage_reg[0][3]  ( .D(n978), .E(n840), .CP(n950), .CDN(n597), 
        .Q(\Storage[0][3] ) );
  EDFCNQD1 \Storage_reg[0][2]  ( .D(n974), .E(N150), .CP(n958), .CDN(n597), 
        .Q(\Storage[0][2] ) );
  EDFCNQD1 \Storage_reg[0][1]  ( .D(n970), .E(N150), .CP(n947), .CDN(n597), 
        .Q(\Storage[0][1] ) );
  EDFCNQD1 \Storage_reg[0][0]  ( .D(n966), .E(N150), .CP(n932), .CDN(n597), 
        .Q(\Storage[0][0] ) );
  EDFCNQD1 \Storage_reg[23][32]  ( .D(n842), .E(n746), .CP(n873), .CDN(n652), 
        .Q(\Storage[23][32] ) );
  EDFCNQD1 \Storage_reg[23][31]  ( .D(n1092), .E(n746), .CP(n873), .CDN(n652), 
        .Q(\Storage[23][31] ) );
  EDFCNQD1 \Storage_reg[23][30]  ( .D(n1088), .E(n746), .CP(n873), .CDN(n652), 
        .Q(\Storage[23][30] ) );
  EDFCNQD1 \Storage_reg[23][29]  ( .D(n1084), .E(n746), .CP(n873), .CDN(n651), 
        .Q(\Storage[23][29] ) );
  EDFCNQD1 \Storage_reg[23][28]  ( .D(n1080), .E(n746), .CP(n873), .CDN(n651), 
        .Q(\Storage[23][28] ) );
  EDFCNQD1 \Storage_reg[23][27]  ( .D(n1076), .E(n746), .CP(n873), .CDN(n651), 
        .Q(\Storage[23][27] ) );
  EDFCNQD1 \Storage_reg[23][26]  ( .D(n1072), .E(n746), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][26] ) );
  EDFCNQD1 \Storage_reg[23][25]  ( .D(n1068), .E(n746), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][25] ) );
  EDFCNQD1 \Storage_reg[23][24]  ( .D(n1064), .E(n746), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][24] ) );
  EDFCNQD1 \Storage_reg[23][23]  ( .D(n1060), .E(n746), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][23] ) );
  EDFCNQD1 \Storage_reg[23][22]  ( .D(n1056), .E(n747), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][22] ) );
  EDFCNQD1 \Storage_reg[23][21]  ( .D(n1052), .E(n747), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][21] ) );
  EDFCNQD1 \Storage_reg[23][20]  ( .D(n1048), .E(n747), .CP(n874), .CDN(n651), 
        .Q(\Storage[23][20] ) );
  EDFCNQD1 \Storage_reg[23][19]  ( .D(n1044), .E(n747), .CP(n874), .CDN(n650), 
        .Q(\Storage[23][19] ) );
  EDFCNQD1 \Storage_reg[23][18]  ( .D(n1040), .E(n747), .CP(n874), .CDN(n650), 
        .Q(\Storage[23][18] ) );
  EDFCNQD1 \Storage_reg[23][17]  ( .D(n1036), .E(n747), .CP(n874), .CDN(n650), 
        .Q(\Storage[23][17] ) );
  EDFCNQD1 \Storage_reg[23][16]  ( .D(n1032), .E(n747), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][16] ) );
  EDFCNQD1 \Storage_reg[23][15]  ( .D(n1028), .E(n747), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][15] ) );
  EDFCNQD1 \Storage_reg[23][14]  ( .D(n1024), .E(n747), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][14] ) );
  EDFCNQD1 \Storage_reg[23][13]  ( .D(n1020), .E(n747), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][13] ) );
  EDFCNQD1 \Storage_reg[23][12]  ( .D(n1016), .E(n748), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][12] ) );
  EDFCNQD1 \Storage_reg[23][11]  ( .D(n1012), .E(n748), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][11] ) );
  EDFCNQD1 \Storage_reg[23][10]  ( .D(n1008), .E(n748), .CP(n875), .CDN(n650), 
        .Q(\Storage[23][10] ) );
  EDFCNQD1 \Storage_reg[23][9]  ( .D(n1004), .E(n748), .CP(n875), .CDN(n649), 
        .Q(\Storage[23][9] ) );
  EDFCNQD1 \Storage_reg[23][8]  ( .D(n1000), .E(n748), .CP(n875), .CDN(n649), 
        .Q(\Storage[23][8] ) );
  EDFCNQD1 \Storage_reg[23][7]  ( .D(n996), .E(n748), .CP(n875), .CDN(n649), 
        .Q(\Storage[23][7] ) );
  EDFCNQD1 \Storage_reg[23][6]  ( .D(n992), .E(n748), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][6] ) );
  EDFCNQD1 \Storage_reg[23][5]  ( .D(n988), .E(n748), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][5] ) );
  EDFCNQD1 \Storage_reg[23][4]  ( .D(n984), .E(n748), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][4] ) );
  EDFCNQD1 \Storage_reg[23][3]  ( .D(n980), .E(n748), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][3] ) );
  EDFCNQD1 \Storage_reg[23][2]  ( .D(n976), .E(N909), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][2] ) );
  EDFCNQD1 \Storage_reg[23][1]  ( .D(n972), .E(N909), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][1] ) );
  EDFCNQD1 \Storage_reg[23][0]  ( .D(n968), .E(N909), .CP(n876), .CDN(n649), 
        .Q(\Storage[23][0] ) );
  EDFCNQD1 \Storage_reg[20][32]  ( .D(n843), .E(n758), .CP(n883), .CDN(n642), 
        .Q(\Storage[20][32] ) );
  EDFCNQD1 \Storage_reg[20][31]  ( .D(n1092), .E(n758), .CP(n883), .CDN(n642), 
        .Q(\Storage[20][31] ) );
  EDFCNQD1 \Storage_reg[20][30]  ( .D(n1088), .E(n758), .CP(n883), .CDN(n642), 
        .Q(\Storage[20][30] ) );
  EDFCNQD1 \Storage_reg[20][29]  ( .D(n1084), .E(n758), .CP(n883), .CDN(n642), 
        .Q(\Storage[20][29] ) );
  EDFCNQD1 \Storage_reg[20][28]  ( .D(n1080), .E(n758), .CP(n883), .CDN(n641), 
        .Q(\Storage[20][28] ) );
  EDFCNQD1 \Storage_reg[20][27]  ( .D(n1076), .E(n758), .CP(n883), .CDN(n641), 
        .Q(\Storage[20][27] ) );
  EDFCNQD1 \Storage_reg[20][26]  ( .D(n1072), .E(n758), .CP(n883), .CDN(n641), 
        .Q(\Storage[20][26] ) );
  EDFCNQD1 \Storage_reg[20][25]  ( .D(n1068), .E(n758), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][25] ) );
  EDFCNQD1 \Storage_reg[20][24]  ( .D(n1064), .E(n758), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][24] ) );
  EDFCNQD1 \Storage_reg[20][23]  ( .D(n1060), .E(n758), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][23] ) );
  EDFCNQD1 \Storage_reg[20][22]  ( .D(n1056), .E(n759), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][22] ) );
  EDFCNQD1 \Storage_reg[20][21]  ( .D(n1052), .E(n759), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][21] ) );
  EDFCNQD1 \Storage_reg[20][20]  ( .D(n1048), .E(n759), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][20] ) );
  EDFCNQD1 \Storage_reg[20][19]  ( .D(n1044), .E(n759), .CP(n884), .CDN(n641), 
        .Q(\Storage[20][19] ) );
  EDFCNQD1 \Storage_reg[20][18]  ( .D(n1040), .E(n759), .CP(n884), .CDN(n640), 
        .Q(\Storage[20][18] ) );
  EDFCNQD1 \Storage_reg[20][17]  ( .D(n1036), .E(n759), .CP(n884), .CDN(n640), 
        .Q(\Storage[20][17] ) );
  EDFCNQD1 \Storage_reg[20][16]  ( .D(n1032), .E(n759), .CP(n884), .CDN(n640), 
        .Q(\Storage[20][16] ) );
  EDFCNQD1 \Storage_reg[20][15]  ( .D(n1028), .E(n759), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][15] ) );
  EDFCNQD1 \Storage_reg[20][14]  ( .D(n1024), .E(n759), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][14] ) );
  EDFCNQD1 \Storage_reg[20][13]  ( .D(n1020), .E(n759), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][13] ) );
  EDFCNQD1 \Storage_reg[20][12]  ( .D(n1016), .E(n760), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][12] ) );
  EDFCNQD1 \Storage_reg[20][11]  ( .D(n1012), .E(n760), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][11] ) );
  EDFCNQD1 \Storage_reg[20][10]  ( .D(n1008), .E(n760), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][10] ) );
  EDFCNQD1 \Storage_reg[20][9]  ( .D(n1004), .E(n760), .CP(n885), .CDN(n640), 
        .Q(\Storage[20][9] ) );
  EDFCNQD1 \Storage_reg[20][8]  ( .D(n1000), .E(n760), .CP(n885), .CDN(n639), 
        .Q(\Storage[20][8] ) );
  EDFCNQD1 \Storage_reg[20][7]  ( .D(n996), .E(n760), .CP(n885), .CDN(n639), 
        .Q(\Storage[20][7] ) );
  EDFCNQD1 \Storage_reg[20][6]  ( .D(n992), .E(n760), .CP(n885), .CDN(n639), 
        .Q(\Storage[20][6] ) );
  EDFCNQD1 \Storage_reg[20][5]  ( .D(n988), .E(n760), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][5] ) );
  EDFCNQD1 \Storage_reg[20][4]  ( .D(n984), .E(n760), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][4] ) );
  EDFCNQD1 \Storage_reg[20][3]  ( .D(n980), .E(n760), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][3] ) );
  EDFCNQD1 \Storage_reg[20][2]  ( .D(n976), .E(N810), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][2] ) );
  EDFCNQD1 \Storage_reg[20][1]  ( .D(n972), .E(N810), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][1] ) );
  EDFCNQD1 \Storage_reg[20][0]  ( .D(n968), .E(N810), .CP(n886), .CDN(n639), 
        .Q(\Storage[20][0] ) );
  EDFCNQD1 \Storage_reg[19][32]  ( .D(n843), .E(n762), .CP(n886), .CDN(n639), 
        .Q(\Storage[19][32] ) );
  EDFCNQD1 \Storage_reg[19][31]  ( .D(n1092), .E(n762), .CP(n886), .CDN(n638), 
        .Q(\Storage[19][31] ) );
  EDFCNQD1 \Storage_reg[19][30]  ( .D(n1088), .E(n762), .CP(n886), .CDN(n638), 
        .Q(\Storage[19][30] ) );
  EDFCNQD1 \Storage_reg[19][29]  ( .D(n1084), .E(n762), .CP(n886), .CDN(n638), 
        .Q(\Storage[19][29] ) );
  EDFCNQD1 \Storage_reg[19][28]  ( .D(n1080), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][28] ) );
  EDFCNQD1 \Storage_reg[19][27]  ( .D(n1076), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][27] ) );
  EDFCNQD1 \Storage_reg[19][26]  ( .D(n1072), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][26] ) );
  EDFCNQD1 \Storage_reg[19][25]  ( .D(n1068), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][25] ) );
  EDFCNQD1 \Storage_reg[19][24]  ( .D(n1064), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][24] ) );
  EDFCNQD1 \Storage_reg[19][23]  ( .D(n1060), .E(n762), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][23] ) );
  EDFCNQD1 \Storage_reg[19][22]  ( .D(n1056), .E(n763), .CP(n887), .CDN(n638), 
        .Q(\Storage[19][22] ) );
  EDFCNQD1 \Storage_reg[19][21]  ( .D(n1052), .E(n763), .CP(n887), .CDN(n637), 
        .Q(\Storage[19][21] ) );
  EDFCNQD1 \Storage_reg[19][20]  ( .D(n1048), .E(n763), .CP(n887), .CDN(n637), 
        .Q(\Storage[19][20] ) );
  EDFCNQD1 \Storage_reg[19][19]  ( .D(n1044), .E(n763), .CP(n887), .CDN(n637), 
        .Q(\Storage[19][19] ) );
  EDFCNQD1 \Storage_reg[19][18]  ( .D(n1040), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][18] ) );
  EDFCNQD1 \Storage_reg[19][17]  ( .D(n1036), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][17] ) );
  EDFCNQD1 \Storage_reg[19][16]  ( .D(n1032), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][16] ) );
  EDFCNQD1 \Storage_reg[19][15]  ( .D(n1028), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][15] ) );
  EDFCNQD1 \Storage_reg[19][14]  ( .D(n1024), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][14] ) );
  EDFCNQD1 \Storage_reg[19][13]  ( .D(n1020), .E(n763), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][13] ) );
  EDFCNQD1 \Storage_reg[19][12]  ( .D(n1016), .E(n764), .CP(n888), .CDN(n637), 
        .Q(\Storage[19][12] ) );
  EDFCNQD1 \Storage_reg[19][11]  ( .D(n1012), .E(n764), .CP(n888), .CDN(n636), 
        .Q(\Storage[19][11] ) );
  EDFCNQD1 \Storage_reg[19][10]  ( .D(n1008), .E(n764), .CP(n888), .CDN(n636), 
        .Q(\Storage[19][10] ) );
  EDFCNQD1 \Storage_reg[19][9]  ( .D(n1004), .E(n764), .CP(n888), .CDN(n636), 
        .Q(\Storage[19][9] ) );
  EDFCNQD1 \Storage_reg[19][8]  ( .D(n1000), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][8] ) );
  EDFCNQD1 \Storage_reg[19][7]  ( .D(n996), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][7] ) );
  EDFCNQD1 \Storage_reg[19][6]  ( .D(n992), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][6] ) );
  EDFCNQD1 \Storage_reg[19][5]  ( .D(n988), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][5] ) );
  EDFCNQD1 \Storage_reg[19][4]  ( .D(n984), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][4] ) );
  EDFCNQD1 \Storage_reg[19][3]  ( .D(n980), .E(n764), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][3] ) );
  EDFCNQD1 \Storage_reg[19][2]  ( .D(n976), .E(N777), .CP(n889), .CDN(n636), 
        .Q(\Storage[19][2] ) );
  EDFCNQD1 \Storage_reg[19][1]  ( .D(n972), .E(N777), .CP(n889), .CDN(n635), 
        .Q(\Storage[19][1] ) );
  EDFCNQD1 \Storage_reg[19][0]  ( .D(n968), .E(N777), .CP(n889), .CDN(n635), 
        .Q(\Storage[19][0] ) );
  EDFCNQD1 \Storage_reg[16][32]  ( .D(n843), .E(n774), .CP(n896), .CDN(n629), 
        .Q(\Storage[16][32] ) );
  EDFCNQD1 \Storage_reg[16][31]  ( .D(n1091), .E(n774), .CP(n896), .CDN(n629), 
        .Q(\Storage[16][31] ) );
  EDFCNQD1 \Storage_reg[16][30]  ( .D(n1087), .E(n774), .CP(n896), .CDN(n628), 
        .Q(\Storage[16][30] ) );
  EDFCNQD1 \Storage_reg[16][29]  ( .D(n1083), .E(n774), .CP(n896), .CDN(n628), 
        .Q(\Storage[16][29] ) );
  EDFCNQD1 \Storage_reg[16][28]  ( .D(n1079), .E(n774), .CP(n896), .CDN(n628), 
        .Q(\Storage[16][28] ) );
  EDFCNQD1 \Storage_reg[16][27]  ( .D(n1075), .E(n774), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][27] ) );
  EDFCNQD1 \Storage_reg[16][26]  ( .D(n1071), .E(n774), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][26] ) );
  EDFCNQD1 \Storage_reg[16][25]  ( .D(n1067), .E(n774), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][25] ) );
  EDFCNQD1 \Storage_reg[16][24]  ( .D(n1063), .E(n774), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][24] ) );
  EDFCNQD1 \Storage_reg[16][23]  ( .D(n1059), .E(n774), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][23] ) );
  EDFCNQD1 \Storage_reg[16][22]  ( .D(n1055), .E(n775), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][22] ) );
  EDFCNQD1 \Storage_reg[16][21]  ( .D(n1051), .E(n775), .CP(n897), .CDN(n628), 
        .Q(\Storage[16][21] ) );
  EDFCNQD1 \Storage_reg[16][20]  ( .D(n1047), .E(n775), .CP(n897), .CDN(n627), 
        .Q(\Storage[16][20] ) );
  EDFCNQD1 \Storage_reg[16][19]  ( .D(n1043), .E(n775), .CP(n897), .CDN(n627), 
        .Q(\Storage[16][19] ) );
  EDFCNQD1 \Storage_reg[16][18]  ( .D(n1039), .E(n775), .CP(n897), .CDN(n627), 
        .Q(\Storage[16][18] ) );
  EDFCNQD1 \Storage_reg[16][17]  ( .D(n1035), .E(n775), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][17] ) );
  EDFCNQD1 \Storage_reg[16][16]  ( .D(n1031), .E(n775), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][16] ) );
  EDFCNQD1 \Storage_reg[16][15]  ( .D(n1027), .E(n775), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][15] ) );
  EDFCNQD1 \Storage_reg[16][14]  ( .D(n1023), .E(n775), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][14] ) );
  EDFCNQD1 \Storage_reg[16][13]  ( .D(n1019), .E(n775), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][13] ) );
  EDFCNQD1 \Storage_reg[16][12]  ( .D(n1015), .E(n776), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][12] ) );
  EDFCNQD1 \Storage_reg[16][11]  ( .D(n1011), .E(n776), .CP(n898), .CDN(n627), 
        .Q(\Storage[16][11] ) );
  EDFCNQD1 \Storage_reg[16][10]  ( .D(n1007), .E(n776), .CP(n898), .CDN(n626), 
        .Q(\Storage[16][10] ) );
  EDFCNQD1 \Storage_reg[16][9]  ( .D(n1003), .E(n776), .CP(n898), .CDN(n626), 
        .Q(\Storage[16][9] ) );
  EDFCNQD1 \Storage_reg[16][8]  ( .D(n999), .E(n776), .CP(n898), .CDN(n626), 
        .Q(\Storage[16][8] ) );
  EDFCNQD1 \Storage_reg[16][7]  ( .D(n995), .E(n776), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][7] ) );
  EDFCNQD1 \Storage_reg[16][6]  ( .D(n991), .E(n776), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][6] ) );
  EDFCNQD1 \Storage_reg[16][5]  ( .D(n987), .E(n776), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][5] ) );
  EDFCNQD1 \Storage_reg[16][4]  ( .D(n983), .E(n776), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][4] ) );
  EDFCNQD1 \Storage_reg[16][3]  ( .D(n979), .E(n776), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][3] ) );
  EDFCNQD1 \Storage_reg[16][2]  ( .D(n975), .E(N678), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][2] ) );
  EDFCNQD1 \Storage_reg[16][1]  ( .D(n971), .E(N678), .CP(n899), .CDN(n626), 
        .Q(\Storage[16][1] ) );
  EDFCNQD1 \Storage_reg[16][0]  ( .D(n967), .E(N678), .CP(n899), .CDN(n625), 
        .Q(\Storage[16][0] ) );
  EDFCNQD1 \Storage_reg[15][32]  ( .D(n843), .E(n778), .CP(n899), .CDN(n625), 
        .Q(\Storage[15][32] ) );
  EDFCNQD1 \Storage_reg[15][31]  ( .D(n1091), .E(n778), .CP(n899), .CDN(n625), 
        .Q(\Storage[15][31] ) );
  EDFCNQD1 \Storage_reg[15][30]  ( .D(n1087), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][30] ) );
  EDFCNQD1 \Storage_reg[15][29]  ( .D(n1083), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][29] ) );
  EDFCNQD1 \Storage_reg[15][28]  ( .D(n1079), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][28] ) );
  EDFCNQD1 \Storage_reg[15][27]  ( .D(n1075), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][27] ) );
  EDFCNQD1 \Storage_reg[15][26]  ( .D(n1071), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][26] ) );
  EDFCNQD1 \Storage_reg[15][25]  ( .D(n1067), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][25] ) );
  EDFCNQD1 \Storage_reg[15][24]  ( .D(n1063), .E(n778), .CP(n900), .CDN(n625), 
        .Q(\Storage[15][24] ) );
  EDFCNQD1 \Storage_reg[15][23]  ( .D(n1059), .E(n778), .CP(n900), .CDN(n624), 
        .Q(\Storage[15][23] ) );
  EDFCNQD1 \Storage_reg[15][22]  ( .D(n1055), .E(n779), .CP(n900), .CDN(n624), 
        .Q(\Storage[15][22] ) );
  EDFCNQD1 \Storage_reg[15][21]  ( .D(n1051), .E(n779), .CP(n900), .CDN(n624), 
        .Q(\Storage[15][21] ) );
  EDFCNQD1 \Storage_reg[15][20]  ( .D(n1047), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][20] ) );
  EDFCNQD1 \Storage_reg[15][19]  ( .D(n1043), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][19] ) );
  EDFCNQD1 \Storage_reg[15][18]  ( .D(n1039), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][18] ) );
  EDFCNQD1 \Storage_reg[15][17]  ( .D(n1035), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][17] ) );
  EDFCNQD1 \Storage_reg[15][16]  ( .D(n1031), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][16] ) );
  EDFCNQD1 \Storage_reg[15][15]  ( .D(n1027), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][15] ) );
  EDFCNQD1 \Storage_reg[15][14]  ( .D(n1023), .E(n779), .CP(n901), .CDN(n624), 
        .Q(\Storage[15][14] ) );
  EDFCNQD1 \Storage_reg[15][13]  ( .D(n1019), .E(n779), .CP(n901), .CDN(n623), 
        .Q(\Storage[15][13] ) );
  EDFCNQD1 \Storage_reg[15][12]  ( .D(n1015), .E(n780), .CP(n901), .CDN(n623), 
        .Q(\Storage[15][12] ) );
  EDFCNQD1 \Storage_reg[15][11]  ( .D(n1011), .E(n780), .CP(n901), .CDN(n623), 
        .Q(\Storage[15][11] ) );
  EDFCNQD1 \Storage_reg[15][10]  ( .D(n1007), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][10] ) );
  EDFCNQD1 \Storage_reg[15][9]  ( .D(n1003), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][9] ) );
  EDFCNQD1 \Storage_reg[15][8]  ( .D(n999), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][8] ) );
  EDFCNQD1 \Storage_reg[15][7]  ( .D(n995), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][7] ) );
  EDFCNQD1 \Storage_reg[15][6]  ( .D(n991), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][6] ) );
  EDFCNQD1 \Storage_reg[15][5]  ( .D(n987), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][5] ) );
  EDFCNQD1 \Storage_reg[15][4]  ( .D(n983), .E(n780), .CP(n902), .CDN(n623), 
        .Q(\Storage[15][4] ) );
  EDFCNQD1 \Storage_reg[15][3]  ( .D(n979), .E(n780), .CP(n902), .CDN(n622), 
        .Q(\Storage[15][3] ) );
  EDFCNQD1 \Storage_reg[15][2]  ( .D(n975), .E(N645), .CP(n902), .CDN(n622), 
        .Q(\Storage[15][2] ) );
  EDFCNQD1 \Storage_reg[15][1]  ( .D(n971), .E(N645), .CP(n902), .CDN(n622), 
        .Q(\Storage[15][1] ) );
  EDFCNQD1 \Storage_reg[15][0]  ( .D(n967), .E(N645), .CP(n903), .CDN(n622), 
        .Q(\Storage[15][0] ) );
  EDFCNQD1 \Storage_reg[12][32]  ( .D(n843), .E(n790), .CP(n922), .CDN(n615), 
        .Q(\Storage[12][32] ) );
  EDFCNQD1 \Storage_reg[12][31]  ( .D(n1091), .E(n790), .CP(n920), .CDN(n615), 
        .Q(\Storage[12][31] ) );
  EDFCNQD1 \Storage_reg[12][30]  ( .D(n1087), .E(n790), .CP(n919), .CDN(n615), 
        .Q(\Storage[12][30] ) );
  EDFCNQD1 \Storage_reg[12][29]  ( .D(n1083), .E(n790), .CP(n925), .CDN(n615), 
        .Q(\Storage[12][29] ) );
  EDFCNQD1 \Storage_reg[12][28]  ( .D(n1079), .E(n790), .CP(n915), .CDN(n615), 
        .Q(\Storage[12][28] ) );
  EDFCNQD1 \Storage_reg[12][27]  ( .D(n1075), .E(n790), .CP(n917), .CDN(n615), 
        .Q(\Storage[12][27] ) );
  EDFCNQD1 \Storage_reg[12][26]  ( .D(n1071), .E(n790), .CP(n913), .CDN(n615), 
        .Q(\Storage[12][26] ) );
  EDFCNQD1 \Storage_reg[12][25]  ( .D(n1067), .E(n790), .CP(n940), .CDN(n615), 
        .Q(\Storage[12][25] ) );
  EDFCNQD1 \Storage_reg[12][24]  ( .D(n1063), .E(n790), .CP(n939), .CDN(n615), 
        .Q(\Storage[12][24] ) );
  EDFCNQD1 \Storage_reg[12][23]  ( .D(n1059), .E(n790), .CP(n938), .CDN(n615), 
        .Q(\Storage[12][23] ) );
  EDFCNQD1 \Storage_reg[12][22]  ( .D(n1055), .E(n791), .CP(n928), .CDN(n614), 
        .Q(\Storage[12][22] ) );
  EDFCNQD1 \Storage_reg[12][21]  ( .D(n1051), .E(n791), .CP(n927), .CDN(n614), 
        .Q(\Storage[12][21] ) );
  EDFCNQD1 \Storage_reg[12][20]  ( .D(n1047), .E(n791), .CP(n926), .CDN(n614), 
        .Q(\Storage[12][20] ) );
  EDFCNQD1 \Storage_reg[12][19]  ( .D(n1043), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][19] ) );
  EDFCNQD1 \Storage_reg[12][18]  ( .D(n1039), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][18] ) );
  EDFCNQD1 \Storage_reg[12][17]  ( .D(n1035), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][17] ) );
  EDFCNQD1 \Storage_reg[12][16]  ( .D(n1031), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][16] ) );
  EDFCNQD1 \Storage_reg[12][15]  ( .D(n1027), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][15] ) );
  EDFCNQD1 \Storage_reg[12][14]  ( .D(n1023), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][14] ) );
  EDFCNQD1 \Storage_reg[12][13]  ( .D(n1019), .E(n791), .CP(n909), .CDN(n614), 
        .Q(\Storage[12][13] ) );
  EDFCNQD1 \Storage_reg[12][12]  ( .D(n1015), .E(n792), .CP(n909), .CDN(n613), 
        .Q(\Storage[12][12] ) );
  EDFCNQD1 \Storage_reg[12][11]  ( .D(n1011), .E(n792), .CP(n909), .CDN(n613), 
        .Q(\Storage[12][11] ) );
  EDFCNQD1 \Storage_reg[12][10]  ( .D(n1007), .E(n792), .CP(n909), .CDN(n613), 
        .Q(\Storage[12][10] ) );
  EDFCNQD1 \Storage_reg[12][9]  ( .D(n1003), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][9] ) );
  EDFCNQD1 \Storage_reg[12][8]  ( .D(n999), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][8] ) );
  EDFCNQD1 \Storage_reg[12][7]  ( .D(n995), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][7] ) );
  EDFCNQD1 \Storage_reg[12][6]  ( .D(n991), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][6] ) );
  EDFCNQD1 \Storage_reg[12][5]  ( .D(n987), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][5] ) );
  EDFCNQD1 \Storage_reg[12][4]  ( .D(n983), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][4] ) );
  EDFCNQD1 \Storage_reg[12][3]  ( .D(n979), .E(n792), .CP(n910), .CDN(n613), 
        .Q(\Storage[12][3] ) );
  EDFCNQD1 \Storage_reg[12][2]  ( .D(n975), .E(N546), .CP(n910), .CDN(n612), 
        .Q(\Storage[12][2] ) );
  EDFCNQD1 \Storage_reg[12][1]  ( .D(n971), .E(N546), .CP(n910), .CDN(n612), 
        .Q(\Storage[12][1] ) );
  EDFCNQD1 \Storage_reg[12][0]  ( .D(n967), .E(N546), .CP(n910), .CDN(n612), 
        .Q(\Storage[12][0] ) );
  EDFCNQD1 \Storage_reg[11][32]  ( .D(n844), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][32] ) );
  EDFCNQD1 \Storage_reg[11][31]  ( .D(n1091), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][31] ) );
  EDFCNQD1 \Storage_reg[11][30]  ( .D(n1087), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][30] ) );
  EDFCNQD1 \Storage_reg[11][29]  ( .D(n1083), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][29] ) );
  EDFCNQD1 \Storage_reg[11][28]  ( .D(n1079), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][28] ) );
  EDFCNQD1 \Storage_reg[11][27]  ( .D(n1075), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][27] ) );
  EDFCNQD1 \Storage_reg[11][26]  ( .D(n1071), .E(n794), .CP(n911), .CDN(n612), 
        .Q(\Storage[11][26] ) );
  EDFCNQD1 \Storage_reg[11][25]  ( .D(n1067), .E(n794), .CP(n911), .CDN(n611), 
        .Q(\Storage[11][25] ) );
  EDFCNQD1 \Storage_reg[11][24]  ( .D(n1063), .E(n794), .CP(n911), .CDN(n611), 
        .Q(\Storage[11][24] ) );
  EDFCNQD1 \Storage_reg[11][23]  ( .D(n1059), .E(n794), .CP(n911), .CDN(n611), 
        .Q(\Storage[11][23] ) );
  EDFCNQD1 \Storage_reg[11][22]  ( .D(n1055), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][22] ) );
  EDFCNQD1 \Storage_reg[11][21]  ( .D(n1051), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][21] ) );
  EDFCNQD1 \Storage_reg[11][20]  ( .D(n1047), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][20] ) );
  EDFCNQD1 \Storage_reg[11][19]  ( .D(n1043), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][19] ) );
  EDFCNQD1 \Storage_reg[11][18]  ( .D(n1039), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][18] ) );
  EDFCNQD1 \Storage_reg[11][17]  ( .D(n1035), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][17] ) );
  EDFCNQD1 \Storage_reg[11][16]  ( .D(n1031), .E(n795), .CP(n912), .CDN(n611), 
        .Q(\Storage[11][16] ) );
  EDFCNQD1 \Storage_reg[11][15]  ( .D(n1027), .E(n795), .CP(n912), .CDN(n610), 
        .Q(\Storage[11][15] ) );
  EDFCNQD1 \Storage_reg[11][14]  ( .D(n1023), .E(n795), .CP(n912), .CDN(n610), 
        .Q(\Storage[11][14] ) );
  EDFCNQD1 \Storage_reg[11][13]  ( .D(n1019), .E(n795), .CP(n912), .CDN(n610), 
        .Q(\Storage[11][13] ) );
  EDFCNQD1 \Storage_reg[11][12]  ( .D(n1015), .E(n796), .CP(n950), .CDN(n610), 
        .Q(\Storage[11][12] ) );
  EDFCNQD1 \Storage_reg[11][11]  ( .D(n1011), .E(n796), .CP(n921), .CDN(n610), 
        .Q(\Storage[11][11] ) );
  EDFCNQD1 \Storage_reg[11][10]  ( .D(n1007), .E(n796), .CP(n960), .CDN(n610), 
        .Q(\Storage[11][10] ) );
  EDFCNQD1 \Storage_reg[11][9]  ( .D(n1003), .E(n796), .CP(n915), .CDN(n610), 
        .Q(\Storage[11][9] ) );
  EDFCNQD1 \Storage_reg[11][8]  ( .D(n999), .E(n796), .CP(n916), .CDN(n610), 
        .Q(\Storage[11][8] ) );
  EDFCNQD1 \Storage_reg[11][7]  ( .D(n995), .E(n796), .CP(ClockW), .CDN(n610), 
        .Q(\Storage[11][7] ) );
  EDFCNQD1 \Storage_reg[11][6]  ( .D(n991), .E(n796), .CP(n846), .CDN(n610), 
        .Q(\Storage[11][6] ) );
  EDFCNQD1 \Storage_reg[11][5]  ( .D(n987), .E(n796), .CP(n947), .CDN(n609), 
        .Q(\Storage[11][5] ) );
  EDFCNQD1 \Storage_reg[11][4]  ( .D(n983), .E(n796), .CP(n948), .CDN(n609), 
        .Q(\Storage[11][4] ) );
  EDFCNQD1 \Storage_reg[11][3]  ( .D(n979), .E(n796), .CP(n949), .CDN(n609), 
        .Q(\Storage[11][3] ) );
  EDFCNQD1 \Storage_reg[11][2]  ( .D(n975), .E(N513), .CP(n954), .CDN(n609), 
        .Q(\Storage[11][2] ) );
  EDFCNQD1 \Storage_reg[11][1]  ( .D(n971), .E(N513), .CP(n956), .CDN(n609), 
        .Q(\Storage[11][1] ) );
  EDFCNQD1 \Storage_reg[11][0]  ( .D(n967), .E(N513), .CP(n955), .CDN(n609), 
        .Q(\Storage[11][0] ) );
  EDFCNQD1 \Storage_reg[8][32]  ( .D(n844), .E(n806), .CP(n921), .CDN(n602), 
        .Q(\Storage[8][32] ) );
  EDFCNQD1 \Storage_reg[8][31]  ( .D(n1090), .E(n806), .CP(n961), .CDN(n602), 
        .Q(\Storage[8][31] ) );
  EDFCNQD1 \Storage_reg[8][30]  ( .D(n1086), .E(n806), .CP(n922), .CDN(n602), 
        .Q(\Storage[8][30] ) );
  EDFCNQD1 \Storage_reg[8][29]  ( .D(n1082), .E(n806), .CP(n962), .CDN(n602), 
        .Q(\Storage[8][29] ) );
  EDFCNQD1 \Storage_reg[8][28]  ( .D(n1078), .E(n806), .CP(ClockW), .CDN(n602), 
        .Q(\Storage[8][28] ) );
  EDFCNQD1 \Storage_reg[8][27]  ( .D(n1074), .E(n806), .CP(n941), .CDN(n602), 
        .Q(\Storage[8][27] ) );
  EDFCNQD1 \Storage_reg[8][26]  ( .D(n1070), .E(n806), .CP(n942), .CDN(n602), 
        .Q(\Storage[8][26] ) );
  EDFCNQD1 \Storage_reg[8][25]  ( .D(n1066), .E(n806), .CP(n943), .CDN(n602), 
        .Q(\Storage[8][25] ) );
  EDFCNQD1 \Storage_reg[8][24]  ( .D(n1062), .E(n806), .CP(n945), .CDN(n5), 
        .Q(\Storage[8][24] ) );
  EDFCNQD1 \Storage_reg[8][23]  ( .D(n1058), .E(n806), .CP(n946), .CDN(n706), 
        .Q(\Storage[8][23] ) );
  EDFCNQD1 \Storage_reg[8][22]  ( .D(n1054), .E(n807), .CP(n944), .CDN(n691), 
        .Q(\Storage[8][22] ) );
  EDFCNQD1 \Storage_reg[8][21]  ( .D(n1050), .E(n807), .CP(n939), .CDN(n694), 
        .Q(\Storage[8][21] ) );
  EDFCNQD1 \Storage_reg[8][20]  ( .D(n1046), .E(n807), .CP(n928), .CDN(n692), 
        .Q(\Storage[8][20] ) );
  EDFCNQD1 \Storage_reg[8][19]  ( .D(n1042), .E(n807), .CP(n960), .CDN(n693), 
        .Q(\Storage[8][19] ) );
  EDFCNQD1 \Storage_reg[8][18]  ( .D(n1038), .E(n807), .CP(n934), .CDN(n697), 
        .Q(\Storage[8][18] ) );
  EDFCNQD1 \Storage_reg[8][17]  ( .D(n1034), .E(n807), .CP(n933), .CDN(n698), 
        .Q(\Storage[8][17] ) );
  EDFCNQD1 \Storage_reg[8][16]  ( .D(n1030), .E(n807), .CP(n932), .CDN(n699), 
        .Q(\Storage[8][16] ) );
  EDFCNQD1 \Storage_reg[8][15]  ( .D(n1026), .E(n807), .CP(n929), .CDN(n701), 
        .Q(\Storage[8][15] ) );
  EDFCNQD1 \Storage_reg[8][14]  ( .D(n1022), .E(n807), .CP(n930), .CDN(n686), 
        .Q(\Storage[8][14] ) );
  EDFCNQD1 \Storage_reg[8][13]  ( .D(n1018), .E(n807), .CP(n931), .CDN(n707), 
        .Q(\Storage[8][13] ) );
  EDFCNQD1 \Storage_reg[8][12]  ( .D(n1014), .E(n808), .CP(n938), .CDN(n695), 
        .Q(\Storage[8][12] ) );
  EDFCNQD1 \Storage_reg[8][11]  ( .D(n1010), .E(n808), .CP(n920), .CDN(n696), 
        .Q(\Storage[8][11] ) );
  EDFCNQD1 \Storage_reg[8][10]  ( .D(n1006), .E(n808), .CP(n961), .CDN(n680), 
        .Q(\Storage[8][10] ) );
  EDFCNQD1 \Storage_reg[8][9]  ( .D(n1002), .E(n808), .CP(n920), .CDN(n681), 
        .Q(\Storage[8][9] ) );
  EDFCNQD1 \Storage_reg[8][8]  ( .D(n998), .E(n808), .CP(n913), .CDN(n682), 
        .Q(\Storage[8][8] ) );
  EDFCNQD1 \Storage_reg[8][7]  ( .D(n994), .E(n808), .CP(n943), .CDN(n683), 
        .Q(\Storage[8][7] ) );
  EDFCNQD1 \Storage_reg[8][6]  ( .D(n990), .E(n808), .CP(n914), .CDN(n684), 
        .Q(\Storage[8][6] ) );
  EDFCNQD1 \Storage_reg[8][5]  ( .D(n986), .E(n808), .CP(n916), .CDN(n685), 
        .Q(\Storage[8][5] ) );
  EDFCNQD1 \Storage_reg[8][4]  ( .D(n982), .E(n808), .CP(n919), .CDN(n712), 
        .Q(\Storage[8][4] ) );
  EDFCNQD1 \Storage_reg[8][3]  ( .D(n978), .E(n808), .CP(n918), .CDN(n691), 
        .Q(\Storage[8][3] ) );
  EDFCNQD1 \Storage_reg[8][2]  ( .D(n974), .E(N414), .CP(n917), .CDN(n687), 
        .Q(\Storage[8][2] ) );
  EDFCNQD1 \Storage_reg[8][1]  ( .D(n970), .E(N414), .CP(n928), .CDN(n688), 
        .Q(\Storage[8][1] ) );
  EDFCNQD1 \Storage_reg[8][0]  ( .D(n966), .E(N414), .CP(n927), .CDN(n689), 
        .Q(\Storage[8][0] ) );
  EDFCNQD1 \Storage_reg[7][32]  ( .D(n844), .E(n810), .CP(n945), .CDN(n690), 
        .Q(\Storage[7][32] ) );
  EDFCNQD1 \Storage_reg[7][31]  ( .D(n1090), .E(n810), .CP(n944), .CDN(n713), 
        .Q(\Storage[7][31] ) );
  EDFCNQD1 \Storage_reg[7][30]  ( .D(n1086), .E(n810), .CP(n943), .CDN(n689), 
        .Q(\Storage[7][30] ) );
  EDFCNQD1 \Storage_reg[7][29]  ( .D(n1082), .E(n810), .CP(n942), .CDN(n702), 
        .Q(\Storage[7][29] ) );
  EDFCNQD1 \Storage_reg[7][28]  ( .D(n1078), .E(n810), .CP(n941), .CDN(n711), 
        .Q(\Storage[7][28] ) );
  EDFCNQD1 \Storage_reg[7][27]  ( .D(n1074), .E(n810), .CP(n940), .CDN(n708), 
        .Q(\Storage[7][27] ) );
  EDFCNQD1 \Storage_reg[7][26]  ( .D(n1070), .E(n810), .CP(n939), .CDN(n679), 
        .Q(\Storage[7][26] ) );
  EDFCNQD1 \Storage_reg[7][25]  ( .D(n1066), .E(n810), .CP(n938), .CDN(n704), 
        .Q(\Storage[7][25] ) );
  EDFCNQD1 \Storage_reg[7][24]  ( .D(n1062), .E(n810), .CP(n919), .CDN(n703), 
        .Q(\Storage[7][24] ) );
  EDFCNQD1 \Storage_reg[7][23]  ( .D(n1058), .E(n810), .CP(n955), .CDN(n680), 
        .Q(\Storage[7][23] ) );
  EDFCNQD1 \Storage_reg[7][22]  ( .D(n1054), .E(n811), .CP(n928), .CDN(n701), 
        .Q(\Storage[7][22] ) );
  EDFCNQD1 \Storage_reg[7][21]  ( .D(n1050), .E(n811), .CP(n958), .CDN(n690), 
        .Q(\Storage[7][21] ) );
  EDFCNQD1 \Storage_reg[7][20]  ( .D(n1046), .E(n811), .CP(n916), .CDN(n595), 
        .Q(\Storage[7][20] ) );
  EDFCNQD1 \Storage_reg[7][19]  ( .D(n1042), .E(n811), .CP(n915), .CDN(n710), 
        .Q(\Storage[7][19] ) );
  EDFCNQD1 \Storage_reg[7][18]  ( .D(n1038), .E(n811), .CP(n914), .CDN(n709), 
        .Q(\Storage[7][18] ) );
  EDFCNQD1 \Storage_reg[7][17]  ( .D(n1034), .E(n811), .CP(n913), .CDN(n710), 
        .Q(\Storage[7][17] ) );
  EDFCNQD1 \Storage_reg[7][16]  ( .D(n1030), .E(n811), .CP(n945), .CDN(n698), 
        .Q(\Storage[7][16] ) );
  EDFCNQD1 \Storage_reg[7][15]  ( .D(n1026), .E(n811), .CP(n921), .CDN(n697), 
        .Q(\Storage[7][15] ) );
  EDFCNQD1 \Storage_reg[7][14]  ( .D(n1022), .E(n811), .CP(n947), .CDN(n692), 
        .Q(\Storage[7][14] ) );
  EDFCNQD1 \Storage_reg[7][13]  ( .D(n1018), .E(n811), .CP(n959), .CDN(n711), 
        .Q(\Storage[7][13] ) );
  EDFCNQD1 \Storage_reg[7][12]  ( .D(n1014), .E(n812), .CP(n918), .CDN(n712), 
        .Q(\Storage[7][12] ) );
  EDFCNQD1 \Storage_reg[7][11]  ( .D(n1010), .E(n812), .CP(n917), .CDN(n709), 
        .Q(\Storage[7][11] ) );
  EDFCNQD1 \Storage_reg[7][10]  ( .D(n1006), .E(n812), .CP(n920), .CDN(n704), 
        .Q(\Storage[7][10] ) );
  EDFCNQD1 \Storage_reg[7][9]  ( .D(n1002), .E(n812), .CP(n916), .CDN(n703), 
        .Q(\Storage[7][9] ) );
  EDFCNQD1 \Storage_reg[7][8]  ( .D(n998), .E(n812), .CP(n917), .CDN(n595), 
        .Q(\Storage[7][8] ) );
  EDFCNQD1 \Storage_reg[7][7]  ( .D(n994), .E(n812), .CP(n959), .CDN(n691), 
        .Q(\Storage[7][7] ) );
  EDFCNQD1 \Storage_reg[7][6]  ( .D(n990), .E(n812), .CP(n920), .CDN(n692), 
        .Q(\Storage[7][6] ) );
  EDFCNQD1 \Storage_reg[7][5]  ( .D(n986), .E(n812), .CP(n947), .CDN(n697), 
        .Q(\Storage[7][5] ) );
  EDFCNQD1 \Storage_reg[7][4]  ( .D(n982), .E(n812), .CP(n950), .CDN(n698), 
        .Q(\Storage[7][4] ) );
  EDFCNQD1 \Storage_reg[7][3]  ( .D(n978), .E(n812), .CP(n948), .CDN(n699), 
        .Q(\Storage[7][3] ) );
  EDFCNQD1 \Storage_reg[7][2]  ( .D(n974), .E(N381), .CP(n951), .CDN(n704), 
        .Q(\Storage[7][2] ) );
  EDFCNQD1 \Storage_reg[7][1]  ( .D(n970), .E(N381), .CP(n957), .CDN(n700), 
        .Q(\Storage[7][1] ) );
  EDFCNQD1 \Storage_reg[7][0]  ( .D(n966), .E(N381), .CP(n953), .CDN(n705), 
        .Q(\Storage[7][0] ) );
  EDFCNQD1 \Storage_reg[4][32]  ( .D(n844), .E(n822), .CP(n935), .CDN(n683), 
        .Q(\Storage[4][32] ) );
  EDFCNQD1 \Storage_reg[4][31]  ( .D(n1090), .E(n822), .CP(n957), .CDN(n700), 
        .Q(\Storage[4][31] ) );
  EDFCNQD1 \Storage_reg[4][30]  ( .D(n1086), .E(n822), .CP(n914), .CDN(n700), 
        .Q(\Storage[4][30] ) );
  EDFCNQD1 \Storage_reg[4][29]  ( .D(n1082), .E(n822), .CP(n925), .CDN(n713), 
        .Q(\Storage[4][29] ) );
  EDFCNQD1 \Storage_reg[4][28]  ( .D(n1078), .E(n822), .CP(n953), .CDN(n702), 
        .Q(\Storage[4][28] ) );
  EDFCNQD1 \Storage_reg[4][27]  ( .D(n1074), .E(n822), .CP(n846), .CDN(n711), 
        .Q(\Storage[4][27] ) );
  EDFCNQD1 \Storage_reg[4][26]  ( .D(n1070), .E(n822), .CP(n951), .CDN(n708), 
        .Q(\Storage[4][26] ) );
  EDFCNQD1 \Storage_reg[4][25]  ( .D(n1066), .E(n822), .CP(n947), .CDN(n685), 
        .Q(\Storage[4][25] ) );
  EDFCNQD1 \Storage_reg[4][24]  ( .D(n1062), .E(n822), .CP(n950), .CDN(n693), 
        .Q(\Storage[4][24] ) );
  EDFCNQD1 \Storage_reg[4][23]  ( .D(n1058), .E(n822), .CP(n923), .CDN(n690), 
        .Q(\Storage[4][23] ) );
  EDFCNQD1 \Storage_reg[4][22]  ( .D(n1054), .E(n823), .CP(n916), .CDN(n596), 
        .Q(\Storage[4][22] ) );
  EDFCNQD1 \Storage_reg[4][21]  ( .D(n1050), .E(n823), .CP(n918), .CDN(n704), 
        .Q(\Storage[4][21] ) );
  EDFCNQD1 \Storage_reg[4][20]  ( .D(n1046), .E(n823), .CP(n962), .CDN(n703), 
        .Q(\Storage[4][20] ) );
  EDFCNQD1 \Storage_reg[4][19]  ( .D(n1042), .E(n823), .CP(n959), .CDN(n595), 
        .Q(\Storage[4][19] ) );
  EDFCNQD1 \Storage_reg[4][18]  ( .D(n1038), .E(n823), .CP(n928), .CDN(n710), 
        .Q(\Storage[4][18] ) );
  EDFCNQD1 \Storage_reg[4][17]  ( .D(n1034), .E(n823), .CP(n927), .CDN(n709), 
        .Q(\Storage[4][17] ) );
  EDFCNQD1 \Storage_reg[4][16]  ( .D(n1030), .E(n823), .CP(n926), .CDN(n684), 
        .Q(\Storage[4][16] ) );
  EDFCNQD1 \Storage_reg[4][15]  ( .D(n1026), .E(n823), .CP(n925), .CDN(n686), 
        .Q(\Storage[4][15] ) );
  EDFCNQD1 \Storage_reg[4][14]  ( .D(n1022), .E(n823), .CP(n924), .CDN(n707), 
        .Q(\Storage[4][14] ) );
  EDFCNQD1 \Storage_reg[4][13]  ( .D(n1018), .E(n823), .CP(n920), .CDN(n706), 
        .Q(\Storage[4][13] ) );
  EDFCNQD1 \Storage_reg[4][12]  ( .D(n1014), .E(n824), .CP(n913), .CDN(n705), 
        .Q(\Storage[4][12] ) );
  EDFCNQD1 \Storage_reg[4][11]  ( .D(n1010), .E(n824), .CP(n916), .CDN(n694), 
        .Q(\Storage[4][11] ) );
  EDFCNQD1 \Storage_reg[4][10]  ( .D(n1006), .E(n824), .CP(n915), .CDN(n682), 
        .Q(\Storage[4][10] ) );
  EDFCNQD1 \Storage_reg[4][9]  ( .D(n1002), .E(n824), .CP(n914), .CDN(n701), 
        .Q(\Storage[4][9] ) );
  EDFCNQD1 \Storage_reg[4][8]  ( .D(n998), .E(n824), .CP(n913), .CDN(n694), 
        .Q(\Storage[4][8] ) );
  EDFCNQD1 \Storage_reg[4][7]  ( .D(n994), .E(n824), .CP(n962), .CDN(n679), 
        .Q(\Storage[4][7] ) );
  EDFCNQD1 \Storage_reg[4][6]  ( .D(n990), .E(n824), .CP(n924), .CDN(n684), 
        .Q(\Storage[4][6] ) );
  EDFCNQD1 \Storage_reg[4][5]  ( .D(n986), .E(n824), .CP(n922), .CDN(n687), 
        .Q(\Storage[4][5] ) );
  EDFCNQD1 \Storage_reg[4][4]  ( .D(n982), .E(n824), .CP(n921), .CDN(n700), 
        .Q(\Storage[4][4] ) );
  EDFCNQD1 \Storage_reg[4][3]  ( .D(n978), .E(n824), .CP(n936), .CDN(n688), 
        .Q(\Storage[4][3] ) );
  EDFCNQD1 \Storage_reg[4][2]  ( .D(n974), .E(N282), .CP(n923), .CDN(n695), 
        .Q(\Storage[4][2] ) );
  EDFCNQD1 \Storage_reg[4][1]  ( .D(n970), .E(N282), .CP(n919), .CDN(n696), 
        .Q(\Storage[4][1] ) );
  EDFCNQD1 \Storage_reg[4][0]  ( .D(n966), .E(N282), .CP(n918), .CDN(n680), 
        .Q(\Storage[4][0] ) );
  EDFCNQD1 \Storage_reg[3][32]  ( .D(n844), .E(n826), .CP(n917), .CDN(n681), 
        .Q(\Storage[3][32] ) );
  EDFCNQD1 \Storage_reg[3][31]  ( .D(n1090), .E(n826), .CP(n958), .CDN(n682), 
        .Q(\Storage[3][31] ) );
  EDFCNQD1 \Storage_reg[3][30]  ( .D(n1086), .E(n826), .CP(ClockW), .CDN(n683), 
        .Q(\Storage[3][30] ) );
  EDFCNQD1 \Storage_reg[3][29]  ( .D(n1082), .E(n826), .CP(n939), .CDN(n696), 
        .Q(\Storage[3][29] ) );
  EDFCNQD1 \Storage_reg[3][28]  ( .D(n1078), .E(n826), .CP(n924), .CDN(n705), 
        .Q(\Storage[3][28] ) );
  EDFCNQD1 \Storage_reg[3][27]  ( .D(n1074), .E(n826), .CP(n930), .CDN(n701), 
        .Q(\Storage[3][27] ) );
  EDFCNQD1 \Storage_reg[3][26]  ( .D(n1070), .E(n826), .CP(n913), .CDN(n708), 
        .Q(\Storage[3][26] ) );
  EDFCNQD1 \Storage_reg[3][25]  ( .D(n1066), .E(n826), .CP(n925), .CDN(n707), 
        .Q(\Storage[3][25] ) );
  EDFCNQD1 \Storage_reg[3][24]  ( .D(n1062), .E(n826), .CP(n937), .CDN(n706), 
        .Q(\Storage[3][24] ) );
  EDFCNQD1 \Storage_reg[3][23]  ( .D(n1058), .E(n826), .CP(n922), .CDN(n705), 
        .Q(\Storage[3][23] ) );
  EDFCNQD1 \Storage_reg[3][22]  ( .D(n1054), .E(n827), .CP(n946), .CDN(n596), 
        .Q(\Storage[3][22] ) );
  EDFCNQD1 \Storage_reg[3][21]  ( .D(n1050), .E(n827), .CP(n921), .CDN(n679), 
        .Q(\Storage[3][21] ) );
  EDFCNQD1 \Storage_reg[3][20]  ( .D(n1046), .E(n827), .CP(n919), .CDN(n700), 
        .Q(\Storage[3][20] ) );
  EDFCNQD1 \Storage_reg[3][19]  ( .D(n1042), .E(n827), .CP(n936), .CDN(n695), 
        .Q(\Storage[3][19] ) );
  EDFCNQD1 \Storage_reg[3][18]  ( .D(n1038), .E(n827), .CP(n924), .CDN(n707), 
        .Q(\Storage[3][18] ) );
  EDFCNQD1 \Storage_reg[3][17]  ( .D(n1034), .E(n827), .CP(ClockW), .CDN(n691), 
        .Q(\Storage[3][17] ) );
  EDFCNQD1 \Storage_reg[3][16]  ( .D(n1030), .E(n827), .CP(n952), .CDN(n681), 
        .Q(\Storage[3][16] ) );
  EDFCNQD1 \Storage_reg[3][15]  ( .D(n1026), .E(n827), .CP(n924), .CDN(n678), 
        .Q(\Storage[3][15] ) );
  EDFCNQD1 \Storage_reg[3][14]  ( .D(n1022), .E(n827), .CP(n957), .CDN(n706), 
        .Q(\Storage[3][14] ) );
  EDFCNQD1 \Storage_reg[3][13]  ( .D(n1018), .E(n827), .CP(n953), .CDN(n692), 
        .Q(\Storage[3][13] ) );
  EDFCNQD1 \Storage_reg[3][12]  ( .D(n1014), .E(n828), .CP(n955), .CDN(n693), 
        .Q(\Storage[3][12] ) );
  EDFCNQD1 \Storage_reg[3][11]  ( .D(n1010), .E(n828), .CP(n956), .CDN(n694), 
        .Q(\Storage[3][11] ) );
  EDFCNQD1 \Storage_reg[3][10]  ( .D(n1006), .E(n828), .CP(n954), .CDN(n698), 
        .Q(\Storage[3][10] ) );
  EDFCNQD1 \Storage_reg[3][9]  ( .D(n1002), .E(n828), .CP(n953), .CDN(n685), 
        .Q(\Storage[3][9] ) );
  EDFCNQD1 \Storage_reg[3][8]  ( .D(n998), .E(n828), .CP(n846), .CDN(n696), 
        .Q(\Storage[3][8] ) );
  EDFCNQD1 \Storage_reg[3][7]  ( .D(n994), .E(n828), .CP(n951), .CDN(n682), 
        .Q(\Storage[3][7] ) );
  EDFCNQD1 \Storage_reg[3][6]  ( .D(n990), .E(n828), .CP(n950), .CDN(n699), 
        .Q(\Storage[3][6] ) );
  EDFCNQD1 \Storage_reg[3][5]  ( .D(n986), .E(n828), .CP(n948), .CDN(n680), 
        .Q(\Storage[3][5] ) );
  EDFCNQD1 \Storage_reg[3][4]  ( .D(n982), .E(n828), .CP(n947), .CDN(n684), 
        .Q(\Storage[3][4] ) );
  EDFCNQD1 \Storage_reg[3][3]  ( .D(n978), .E(n828), .CP(n926), .CDN(n683), 
        .Q(\Storage[3][3] ) );
  EDFCNQD1 \Storage_reg[3][2]  ( .D(n974), .E(N249), .CP(n950), .CDN(n689), 
        .Q(\Storage[3][2] ) );
  EDFCNQD1 \Storage_reg[3][1]  ( .D(n970), .E(N249), .CP(n962), .CDN(n690), 
        .Q(\Storage[3][1] ) );
  EDFCNQD1 \Storage_reg[3][0]  ( .D(n966), .E(N249), .CP(n917), .CDN(n686), 
        .Q(\Storage[3][0] ) );
  EDFCNQD1 \Storage_reg[0][32]  ( .D(N85), .E(n838), .CP(n943), .CDN(n600), 
        .Q(\Storage[0][32] ) );
  EDFCNQD1 \Storage_reg[0][31]  ( .D(n1090), .E(n838), .CP(n962), .CDN(n600), 
        .Q(\Storage[0][31] ) );
  EDFCNQD1 \Storage_reg[0][30]  ( .D(n1086), .E(n838), .CP(n946), .CDN(n600), 
        .Q(\Storage[0][30] ) );
  EDFCNQD1 \Storage_reg[0][29]  ( .D(n1082), .E(n838), .CP(n919), .CDN(n600), 
        .Q(\Storage[0][29] ) );
  EDFCNQD1 \Storage_reg[0][28]  ( .D(n1078), .E(n838), .CP(ClockW), .CDN(n599), 
        .Q(\Storage[0][28] ) );
  EDFCNQD1 \Storage_reg[0][27]  ( .D(n1074), .E(n838), .CP(n846), .CDN(n599), 
        .Q(\Storage[0][27] ) );
  EDFCNQD1 \Storage_reg[0][26]  ( .D(n1070), .E(n838), .CP(n947), .CDN(n599), 
        .Q(\Storage[0][26] ) );
  EDFCNQD1 \Storage_reg[0][25]  ( .D(n1066), .E(n838), .CP(n951), .CDN(n599), 
        .Q(\Storage[0][25] ) );
  EDFCNQD1 \Storage_reg[0][24]  ( .D(n1062), .E(n838), .CP(n949), .CDN(n599), 
        .Q(\Storage[0][24] ) );
  EDFCNQD1 \Storage_reg[0][23]  ( .D(n1058), .E(n838), .CP(n952), .CDN(n599), 
        .Q(\Storage[0][23] ) );
  EDFCNQD1 \Storage_reg[0][22]  ( .D(n1054), .E(n839), .CP(n957), .CDN(n599), 
        .Q(\Storage[0][22] ) );
  EDFCNQD1 \Storage_reg[0][21]  ( .D(n1050), .E(n839), .CP(n915), .CDN(n599), 
        .Q(\Storage[0][21] ) );
  EDFCNQD1 \Storage_reg[0][20]  ( .D(n1046), .E(n839), .CP(n955), .CDN(n599), 
        .Q(\Storage[0][20] ) );
  EDFCNQD1 \Storage_reg[0][19]  ( .D(n1042), .E(n839), .CP(n956), .CDN(n599), 
        .Q(\Storage[0][19] ) );
  EDFCNQD1 \Storage_reg[0][18]  ( .D(n1038), .E(n839), .CP(n917), .CDN(n598), 
        .Q(\Storage[0][18] ) );
  EDFCNQD1 \Storage_reg[0][17]  ( .D(n1034), .E(n839), .CP(n953), .CDN(n598), 
        .Q(\Storage[0][17] ) );
  EDFCNQD1 \Storage_reg[0][16]  ( .D(n1030), .E(n839), .CP(n954), .CDN(n598), 
        .Q(\Storage[0][16] ) );
  EDFCNQD1 \Storage_reg[0][15]  ( .D(n1026), .E(n839), .CP(n932), .CDN(n598), 
        .Q(\Storage[0][15] ) );
  EDFCNQD1 \Storage_reg[0][14]  ( .D(n1022), .E(n839), .CP(n942), .CDN(n598), 
        .Q(\Storage[0][14] ) );
  EDFCNQD1 \Storage_reg[0][13]  ( .D(n1018), .E(n839), .CP(n925), .CDN(n598), 
        .Q(\Storage[0][13] ) );
  EDFCNQD1 \Storage_reg[0][12]  ( .D(n1014), .E(n840), .CP(n959), .CDN(n598), 
        .Q(\Storage[0][12] ) );
  EDFCNQD1 \Storage_reg[0][11]  ( .D(n1010), .E(n840), .CP(n960), .CDN(n598), 
        .Q(\Storage[0][11] ) );
  EDFCNQD1 \Storage_reg[0][10]  ( .D(n1006), .E(n840), .CP(n961), .CDN(n598), 
        .Q(\Storage[0][10] ) );
  EDFCNQD1 \Storage_reg[0][9]  ( .D(n1002), .E(n840), .CP(n937), .CDN(n598), 
        .Q(\Storage[0][9] ) );
  EDFCNQD1 \Storage_reg[0][8]  ( .D(n998), .E(n840), .CP(n958), .CDN(n597), 
        .Q(\Storage[0][8] ) );
  EDFCNQD1 \Storage_reg[0][7]  ( .D(n994), .E(n840), .CP(n934), .CDN(n597), 
        .Q(\Storage[0][7] ) );
  EDFCNQD1 \Storage_reg[0][6]  ( .D(n990), .E(n840), .CP(n933), .CDN(n597), 
        .Q(\Storage[0][6] ) );
  EDFCNQD1 \Storage_reg[31][32]  ( .D(n842), .E(n714), .CP(n847), .CDN(n678), 
        .Q(\Storage[31][32] ) );
  EDFCNQD1 \Storage_reg[31][31]  ( .D(DataI[31]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][31] ) );
  EDFCNQD1 \Storage_reg[31][30]  ( .D(DataI[30]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][30] ) );
  EDFCNQD1 \Storage_reg[31][29]  ( .D(DataI[29]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][29] ) );
  EDFCNQD1 \Storage_reg[31][28]  ( .D(DataI[28]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][28] ) );
  EDFCNQD1 \Storage_reg[31][27]  ( .D(DataI[27]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][27] ) );
  EDFCNQD1 \Storage_reg[31][26]  ( .D(DataI[26]), .E(n714), .CP(n847), .CDN(
        n678), .Q(\Storage[31][26] ) );
  EDFCNQD1 \Storage_reg[31][25]  ( .D(DataI[25]), .E(n714), .CP(n847), .CDN(
        n677), .Q(\Storage[31][25] ) );
  EDFCNQD1 \Storage_reg[31][24]  ( .D(DataI[24]), .E(n714), .CP(n847), .CDN(
        n677), .Q(\Storage[31][24] ) );
  EDFCNQD1 \Storage_reg[31][23]  ( .D(DataI[23]), .E(n714), .CP(n847), .CDN(
        n677), .Q(\Storage[31][23] ) );
  EDFCNQD1 \Storage_reg[31][22]  ( .D(DataI[22]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][22] ) );
  EDFCNQD1 \Storage_reg[31][21]  ( .D(DataI[21]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][21] ) );
  EDFCNQD1 \Storage_reg[31][20]  ( .D(DataI[20]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][20] ) );
  EDFCNQD1 \Storage_reg[31][19]  ( .D(DataI[19]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][19] ) );
  EDFCNQD1 \Storage_reg[31][18]  ( .D(DataI[18]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][18] ) );
  EDFCNQD1 \Storage_reg[31][17]  ( .D(DataI[17]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][17] ) );
  EDFCNQD1 \Storage_reg[31][16]  ( .D(DataI[16]), .E(n715), .CP(n848), .CDN(
        n677), .Q(\Storage[31][16] ) );
  EDFCNQD1 \Storage_reg[31][15]  ( .D(DataI[15]), .E(n715), .CP(n848), .CDN(
        n676), .Q(\Storage[31][15] ) );
  EDFCNQD1 \Storage_reg[31][14]  ( .D(DataI[14]), .E(n715), .CP(n848), .CDN(
        n676), .Q(\Storage[31][14] ) );
  EDFCNQD1 \Storage_reg[31][13]  ( .D(DataI[13]), .E(n715), .CP(n848), .CDN(
        n676), .Q(\Storage[31][13] ) );
  EDFCNQD1 \Storage_reg[31][12]  ( .D(DataI[12]), .E(n716), .CP(n849), .CDN(
        n676), .Q(\Storage[31][12] ) );
  EDFCNQD1 \Storage_reg[31][11]  ( .D(DataI[11]), .E(n716), .CP(n849), .CDN(
        n676), .Q(\Storage[31][11] ) );
  EDFCNQD1 \Storage_reg[31][10]  ( .D(DataI[10]), .E(n716), .CP(n849), .CDN(
        n676), .Q(\Storage[31][10] ) );
  EDFCNQD1 \Storage_reg[31][9]  ( .D(DataI[9]), .E(n716), .CP(n849), .CDN(n676), .Q(\Storage[31][9] ) );
  EDFCNQD1 \Storage_reg[31][8]  ( .D(DataI[8]), .E(n716), .CP(n849), .CDN(n676), .Q(\Storage[31][8] ) );
  EDFCNQD1 \Storage_reg[31][7]  ( .D(DataI[7]), .E(n716), .CP(n849), .CDN(n676), .Q(\Storage[31][7] ) );
  EDFCNQD1 \Storage_reg[31][6]  ( .D(DataI[6]), .E(n716), .CP(n849), .CDN(n676), .Q(\Storage[31][6] ) );
  EDFCNQD1 \Storage_reg[31][5]  ( .D(DataI[5]), .E(n716), .CP(n849), .CDN(n675), .Q(\Storage[31][5] ) );
  EDFCNQD1 \Storage_reg[31][4]  ( .D(DataI[4]), .E(n716), .CP(n849), .CDN(n675), .Q(\Storage[31][4] ) );
  EDFCNQD1 \Storage_reg[31][3]  ( .D(DataI[3]), .E(n716), .CP(n849), .CDN(n675), .Q(\Storage[31][3] ) );
  EDFCNQD1 \Storage_reg[31][2]  ( .D(DataI[2]), .E(N1173), .CP(n850), .CDN(
        n675), .Q(\Storage[31][2] ) );
  EDFCNQD1 \Storage_reg[31][1]  ( .D(DataI[1]), .E(N1173), .CP(n850), .CDN(
        n675), .Q(\Storage[31][1] ) );
  EDFCNQD1 \Storage_reg[31][0]  ( .D(DataI[0]), .E(N1173), .CP(n850), .CDN(
        n675), .Q(\Storage[31][0] ) );
  DFCNQD1 Dreadyr_reg ( .D(n107), .CP(ClockR), .CDN(n597), .Q(Dreadyr) );
  BUFTD0 \DataO_tri[0]  ( .I(DataOr[0]), .OE(ChipEna), .Z(DataO[0]) );
  BUFTD0 \DataO_tri[1]  ( .I(DataOr[1]), .OE(ChipEna), .Z(DataO[1]) );
  BUFTD0 \DataO_tri[2]  ( .I(DataOr[2]), .OE(ChipEna), .Z(DataO[2]) );
  BUFTD0 \DataO_tri[3]  ( .I(DataOr[3]), .OE(ChipEna), .Z(DataO[3]) );
  BUFTD0 \DataO_tri[4]  ( .I(DataOr[4]), .OE(ChipEna), .Z(DataO[4]) );
  BUFTD0 \DataO_tri[5]  ( .I(DataOr[5]), .OE(ChipEna), .Z(DataO[5]) );
  BUFTD0 \DataO_tri[6]  ( .I(DataOr[6]), .OE(ChipEna), .Z(DataO[6]) );
  BUFTD0 \DataO_tri[7]  ( .I(DataOr[7]), .OE(ChipEna), .Z(DataO[7]) );
  BUFTD0 \DataO_tri[8]  ( .I(DataOr[8]), .OE(ChipEna), .Z(DataO[8]) );
  BUFTD0 \DataO_tri[9]  ( .I(DataOr[9]), .OE(ChipEna), .Z(DataO[9]) );
  BUFTD0 \DataO_tri[10]  ( .I(DataOr[10]), .OE(ChipEna), .Z(DataO[10]) );
  BUFTD0 \DataO_tri[11]  ( .I(DataOr[11]), .OE(ChipEna), .Z(DataO[11]) );
  BUFTD0 \DataO_tri[12]  ( .I(DataOr[12]), .OE(ChipEna), .Z(DataO[12]) );
  BUFTD0 \DataO_tri[13]  ( .I(DataOr[13]), .OE(ChipEna), .Z(DataO[13]) );
  BUFTD0 \DataO_tri[14]  ( .I(DataOr[14]), .OE(ChipEna), .Z(DataO[14]) );
  BUFTD0 \DataO_tri[15]  ( .I(DataOr[15]), .OE(ChipEna), .Z(DataO[15]) );
  BUFTD0 \DataO_tri[16]  ( .I(DataOr[16]), .OE(ChipEna), .Z(DataO[16]) );
  BUFTD0 \DataO_tri[17]  ( .I(DataOr[17]), .OE(ChipEna), .Z(DataO[17]) );
  BUFTD0 \DataO_tri[18]  ( .I(DataOr[18]), .OE(ChipEna), .Z(DataO[18]) );
  BUFTD0 \DataO_tri[19]  ( .I(DataOr[19]), .OE(ChipEna), .Z(DataO[19]) );
  BUFTD0 \DataO_tri[20]  ( .I(DataOr[20]), .OE(ChipEna), .Z(DataO[20]) );
  BUFTD0 \DataO_tri[21]  ( .I(DataOr[21]), .OE(ChipEna), .Z(DataO[21]) );
  BUFTD0 \DataO_tri[22]  ( .I(DataOr[22]), .OE(ChipEna), .Z(DataO[22]) );
  BUFTD0 \DataO_tri[23]  ( .I(DataOr[23]), .OE(ChipEna), .Z(DataO[23]) );
  BUFTD0 \DataO_tri[24]  ( .I(DataOr[24]), .OE(ChipEna), .Z(DataO[24]) );
  BUFTD0 \DataO_tri[25]  ( .I(DataOr[25]), .OE(ChipEna), .Z(DataO[25]) );
  BUFTD0 \DataO_tri[26]  ( .I(DataOr[26]), .OE(ChipEna), .Z(DataO[26]) );
  BUFTD0 \DataO_tri[27]  ( .I(DataOr[27]), .OE(ChipEna), .Z(DataO[27]) );
  BUFTD0 \DataO_tri[28]  ( .I(DataOr[28]), .OE(ChipEna), .Z(DataO[28]) );
  BUFTD0 \DataO_tri[29]  ( .I(DataOr[29]), .OE(ChipEna), .Z(DataO[29]) );
  BUFTD0 \DataO_tri[30]  ( .I(DataOr[30]), .OE(ChipEna), .Z(DataO[30]) );
  BUFTD0 \DataO_tri[31]  ( .I(DataOr[31]), .OE(ChipEna), .Z(DataO[31]) );
  EDFCND1 \DataOr_reg[29]  ( .D(N53), .E(n1), .CP(ClockR), .CDN(n701), .Q(
        DataOr[29]) );
  EDFCND1 \DataOr_reg[28]  ( .D(N54), .E(Read), .CP(ClockR), .CDN(n708), .Q(
        DataOr[28]) );
  EDFCND1 \DataOr_reg[25]  ( .D(N57), .E(n1), .CP(ClockR), .CDN(n709), .Q(
        DataOr[25]) );
  EDFCND1 \DataOr_reg[22]  ( .D(N60), .E(Read), .CP(ClockR), .CDN(n5), .Q(
        DataOr[22]) );
  EDFCND1 \DataOr_reg[21]  ( .D(N61), .E(Read), .CP(ClockR), .CDN(n688), .Q(
        DataOr[21]) );
  EDFCND1 \DataOr_reg[18]  ( .D(N64), .E(n3), .CP(ClockR), .CDN(n4), .Q(
        DataOr[18]) );
  EDFCND1 \DataOr_reg[17]  ( .D(N65), .E(n2), .CP(ClockR), .CDN(n4), .Q(
        DataOr[17]) );
  EDFCND1 \DataOr_reg[15]  ( .D(N67), .E(n3), .CP(ClockR), .CDN(n5), .Q(
        DataOr[15]) );
  EDFCND1 \DataOr_reg[14]  ( .D(N68), .E(n2), .CP(ClockR), .CDN(n5), .Q(
        DataOr[14]) );
  EDFCND1 \DataOr_reg[11]  ( .D(N71), .E(n1), .CP(ClockR), .CDN(n4), .Q(
        DataOr[11]) );
  EDFCND1 \DataOr_reg[10]  ( .D(N72), .E(n3), .CP(ClockR), .CDN(n596), .Q(
        DataOr[10]) );
  EDFCND1 \DataOr_reg[9]  ( .D(N73), .E(n2), .CP(ClockR), .CDN(n710), .Q(
        DataOr[9]) );
  EDFCND1 \DataOr_reg[5]  ( .D(N77), .E(n1), .CP(ClockR), .CDN(n707), .Q(
        DataOr[5]) );
  EDFCND1 \DataOr_reg[4]  ( .D(N78), .E(Read), .CP(ClockR), .CDN(n700), .Q(
        DataOr[4]) );
  EDFCND1 \DataOr_reg[3]  ( .D(N79), .E(Read), .CP(ClockR), .CDN(n596), .Q(
        DataOr[3]) );
  EDFCND1 \DataOr_reg[0]  ( .D(N82), .E(Read), .CP(ClockR), .CDN(n4), .Q(
        DataOr[0]) );
  EDFCND1 \DataOr_reg[24]  ( .D(N58), .E(n3), .CP(ClockR), .CDN(n5), .Q(
        DataOr[24]) );
  EDFCND1 \DataOr_reg[23]  ( .D(N59), .E(n1), .CP(ClockR), .CDN(n4), .Q(
        DataOr[23]) );
  EDFCND1 \DataOr_reg[16]  ( .D(N66), .E(n2), .CP(ClockR), .CDN(n704), .Q(
        DataOr[16]) );
  EDFCND1 \DataOr_reg[8]  ( .D(N74), .E(n3), .CP(ClockR), .CDN(n4), .Q(
        DataOr[8]) );
  EDFCND1 \DataOr_reg[6]  ( .D(N76), .E(n1), .CP(ClockR), .CDN(n4), .Q(
        DataOr[6]) );
  EDFCND1 \DataOr_reg[31]  ( .D(N51), .E(n2), .CP(ClockR), .CDN(n5), .Q(
        DataOr[31]) );
  EDFCND1 \DataOr_reg[30]  ( .D(N52), .E(n3), .CP(ClockR), .CDN(n705), .Q(
        DataOr[30]) );
  EDFCND1 \DataOr_reg[27]  ( .D(N55), .E(n1), .CP(ClockR), .CDN(n679), .Q(
        DataOr[27]) );
  EDFCND1 \DataOr_reg[26]  ( .D(N56), .E(n2), .CP(ClockR), .CDN(n703), .Q(
        DataOr[26]) );
  EDFCND1 \DataOr_reg[20]  ( .D(N62), .E(n3), .CP(ClockR), .CDN(n595), .Q(
        DataOr[20]) );
  EDFCND1 \DataOr_reg[19]  ( .D(N63), .E(n1), .CP(ClockR), .CDN(n5), .Q(
        DataOr[19]) );
  EDFCND1 \DataOr_reg[13]  ( .D(N69), .E(n2), .CP(ClockR), .CDN(n4), .Q(
        DataOr[13]) );
  EDFCND1 \DataOr_reg[12]  ( .D(N70), .E(n3), .CP(ClockR), .CDN(n4), .Q(
        DataOr[12]) );
  EDFCND1 \DataOr_reg[7]  ( .D(N75), .E(n2), .CP(ClockR), .CDN(n5), .Q(
        DataOr[7]) );
  EDFCND1 \DataOr_reg[2]  ( .D(N80), .E(n1), .CP(ClockR), .CDN(n706), .Q(
        DataOr[2]) );
  EDFCND1 \DataOr_reg[1]  ( .D(N81), .E(n3), .CP(ClockR), .CDN(n699), .Q(
        DataOr[1]) );
  EDFCND1 Parityr_reg ( .D(N83), .E(n2), .CP(ClockR), .CDN(n5), .Q(ParityErr)
         );
  BUFFD0 U4 ( .I(Read), .Z(n3) );
  BUFFD0 U5 ( .I(Read), .Z(n2) );
  BUFFD0 U6 ( .I(Read), .Z(n1) );
  INVD0 U7 ( .I(Reset), .ZN(n4) );
  INVD0 U8 ( .I(Reset), .ZN(n5) );
  CKAN2D0 U9 ( .A1(ChipEna), .A2(Dreadyr), .Z(Dready) );
  BUFFD1 U10 ( .I(n698), .Z(n602) );
  BUFFD1 U11 ( .I(n698), .Z(n603) );
  BUFFD1 U12 ( .I(n698), .Z(n604) );
  BUFFD1 U13 ( .I(n698), .Z(n605) );
  BUFFD1 U14 ( .I(n697), .Z(n606) );
  BUFFD1 U15 ( .I(n697), .Z(n607) );
  BUFFD1 U16 ( .I(n697), .Z(n608) );
  BUFFD1 U17 ( .I(n697), .Z(n609) );
  BUFFD1 U23 ( .I(n696), .Z(n610) );
  BUFFD1 U24 ( .I(n696), .Z(n611) );
  BUFFD1 U25 ( .I(n696), .Z(n612) );
  BUFFD1 U26 ( .I(n696), .Z(n613) );
  BUFFD1 U29 ( .I(n695), .Z(n614) );
  BUFFD1 U30 ( .I(n695), .Z(n615) );
  BUFFD1 U31 ( .I(n695), .Z(n616) );
  BUFFD1 U32 ( .I(n695), .Z(n617) );
  BUFFD1 U37 ( .I(n694), .Z(n618) );
  BUFFD1 U38 ( .I(n694), .Z(n619) );
  BUFFD1 U39 ( .I(n694), .Z(n620) );
  BUFFD1 U40 ( .I(n694), .Z(n621) );
  BUFFD1 U41 ( .I(n693), .Z(n622) );
  BUFFD1 U42 ( .I(n693), .Z(n623) );
  BUFFD1 U43 ( .I(n693), .Z(n624) );
  BUFFD1 U44 ( .I(n693), .Z(n625) );
  BUFFD1 U45 ( .I(n692), .Z(n626) );
  BUFFD1 U46 ( .I(n692), .Z(n627) );
  BUFFD1 U47 ( .I(n692), .Z(n628) );
  BUFFD1 U48 ( .I(n692), .Z(n629) );
  BUFFD1 U49 ( .I(n691), .Z(n630) );
  BUFFD1 U50 ( .I(n691), .Z(n631) );
  BUFFD1 U51 ( .I(n691), .Z(n632) );
  BUFFD1 U52 ( .I(n691), .Z(n633) );
  BUFFD1 U53 ( .I(n690), .Z(n634) );
  BUFFD1 U54 ( .I(n690), .Z(n635) );
  BUFFD1 U55 ( .I(n690), .Z(n636) );
  BUFFD1 U56 ( .I(n690), .Z(n637) );
  BUFFD1 U57 ( .I(n689), .Z(n638) );
  BUFFD1 U58 ( .I(n689), .Z(n639) );
  BUFFD1 U59 ( .I(n689), .Z(n640) );
  BUFFD1 U60 ( .I(n689), .Z(n641) );
  BUFFD1 U61 ( .I(n688), .Z(n642) );
  BUFFD1 U62 ( .I(n688), .Z(n643) );
  BUFFD1 U63 ( .I(n688), .Z(n644) );
  BUFFD1 U64 ( .I(n688), .Z(n645) );
  BUFFD1 U65 ( .I(n687), .Z(n646) );
  BUFFD1 U66 ( .I(n687), .Z(n647) );
  BUFFD1 U67 ( .I(n687), .Z(n648) );
  BUFFD1 U68 ( .I(n687), .Z(n649) );
  BUFFD1 U69 ( .I(n686), .Z(n650) );
  BUFFD1 U70 ( .I(n686), .Z(n651) );
  BUFFD1 U71 ( .I(n686), .Z(n652) );
  BUFFD1 U72 ( .I(n686), .Z(n653) );
  BUFFD1 U73 ( .I(n685), .Z(n654) );
  BUFFD1 U74 ( .I(n685), .Z(n655) );
  BUFFD1 U75 ( .I(n685), .Z(n656) );
  BUFFD1 U76 ( .I(n685), .Z(n657) );
  BUFFD1 U77 ( .I(n684), .Z(n658) );
  BUFFD1 U78 ( .I(n684), .Z(n659) );
  BUFFD1 U79 ( .I(n684), .Z(n660) );
  BUFFD1 U80 ( .I(n684), .Z(n661) );
  BUFFD1 U81 ( .I(n683), .Z(n662) );
  BUFFD1 U82 ( .I(n683), .Z(n663) );
  BUFFD1 U83 ( .I(n683), .Z(n664) );
  BUFFD1 U84 ( .I(n683), .Z(n665) );
  BUFFD1 U85 ( .I(n682), .Z(n666) );
  BUFFD1 U86 ( .I(n682), .Z(n667) );
  BUFFD1 U87 ( .I(n682), .Z(n668) );
  BUFFD1 U88 ( .I(n682), .Z(n669) );
  BUFFD1 U89 ( .I(n681), .Z(n670) );
  BUFFD1 U90 ( .I(n681), .Z(n671) );
  BUFFD1 U91 ( .I(n681), .Z(n672) );
  BUFFD1 U92 ( .I(n681), .Z(n673) );
  BUFFD1 U93 ( .I(n680), .Z(n674) );
  BUFFD1 U94 ( .I(n680), .Z(n675) );
  BUFFD1 U95 ( .I(n680), .Z(n676) );
  BUFFD1 U96 ( .I(n680), .Z(n677) );
  BUFFD1 U97 ( .I(n679), .Z(n678) );
  BUFFD1 U98 ( .I(n570), .Z(n581) );
  BUFFD1 U99 ( .I(n570), .Z(n582) );
  BUFFD1 U100 ( .I(n569), .Z(n583) );
  BUFFD1 U101 ( .I(n569), .Z(n584) );
  BUFFD1 U102 ( .I(n569), .Z(n585) );
  BUFFD1 U103 ( .I(n568), .Z(n586) );
  BUFFD1 U104 ( .I(n568), .Z(n587) );
  BUFFD1 U105 ( .I(n568), .Z(n588) );
  BUFFD1 U106 ( .I(n567), .Z(n589) );
  BUFFD1 U107 ( .I(n567), .Z(n590) );
  BUFFD1 U108 ( .I(n567), .Z(n591) );
  BUFFD1 U109 ( .I(n566), .Z(n592) );
  BUFFD1 U110 ( .I(n566), .Z(n593) );
  BUFFD1 U111 ( .I(n566), .Z(n594) );
  BUFFD1 U112 ( .I(n570), .Z(n580) );
  BUFFD1 U113 ( .I(n571), .Z(n579) );
  BUFFD1 U114 ( .I(n571), .Z(n578) );
  BUFFD1 U115 ( .I(n571), .Z(n577) );
  BUFFD1 U116 ( .I(n565), .Z(n576) );
  BUFFD1 U117 ( .I(n562), .Z(n575) );
  BUFFD1 U118 ( .I(n536), .Z(n560) );
  BUFFD1 U119 ( .I(n536), .Z(n561) );
  BUFFD1 U120 ( .I(n536), .Z(n559) );
  BUFFD1 U121 ( .I(n520), .Z(n530) );
  BUFFD1 U122 ( .I(n519), .Z(n531) );
  BUFFD1 U123 ( .I(n519), .Z(n532) );
  BUFFD1 U124 ( .I(n537), .Z(n558) );
  BUFFD1 U125 ( .I(n520), .Z(n529) );
  BUFFD1 U126 ( .I(n540), .Z(n551) );
  BUFFD1 U127 ( .I(n572), .Z(n574) );
  BUFFD1 U128 ( .I(n540), .Z(n552) );
  BUFFD1 U129 ( .I(n539), .Z(n553) );
  BUFFD1 U130 ( .I(n539), .Z(n554) );
  BUFFD1 U131 ( .I(n539), .Z(n555) );
  BUFFD1 U132 ( .I(n537), .Z(n556) );
  BUFFD1 U133 ( .I(n537), .Z(n557) );
  BUFFD1 U134 ( .I(n535), .Z(n546) );
  BUFFD1 U135 ( .I(n541), .Z(n547) );
  BUFFD1 U136 ( .I(n541), .Z(n548) );
  BUFFD1 U137 ( .I(n541), .Z(n549) );
  BUFFD1 U138 ( .I(n540), .Z(n550) );
  BUFFD1 U139 ( .I(n520), .Z(n528) );
  BUFFD1 U140 ( .I(n522), .Z(n527) );
  BUFFD1 U141 ( .I(n520), .Z(n526) );
  BUFFD1 U142 ( .I(n521), .Z(n525) );
  BUFFD1 U143 ( .I(n521), .Z(n524) );
  BUFFD1 U144 ( .I(n542), .Z(n545) );
  BUFFD1 U145 ( .I(n542), .Z(n544) );
  BUFFD1 U146 ( .I(n562), .Z(n573) );
  BUFFD1 U147 ( .I(n542), .Z(n543) );
  BUFFD1 U148 ( .I(n522), .Z(n523) );
  BUFFD1 U149 ( .I(n699), .Z(n598) );
  BUFFD1 U150 ( .I(n699), .Z(n599) );
  BUFFD1 U151 ( .I(n699), .Z(n600) );
  BUFFD1 U152 ( .I(n699), .Z(n601) );
  BUFFD1 U153 ( .I(n913), .Z(n912) );
  BUFFD1 U154 ( .I(n913), .Z(n911) );
  BUFFD1 U155 ( .I(n914), .Z(n910) );
  BUFFD1 U156 ( .I(n914), .Z(n909) );
  BUFFD1 U157 ( .I(n916), .Z(n908) );
  BUFFD1 U158 ( .I(n916), .Z(n907) );
  BUFFD1 U159 ( .I(n917), .Z(n906) );
  BUFFD1 U160 ( .I(n917), .Z(n905) );
  BUFFD1 U161 ( .I(n918), .Z(n904) );
  BUFFD1 U162 ( .I(n918), .Z(n903) );
  BUFFD1 U163 ( .I(n919), .Z(n902) );
  BUFFD1 U164 ( .I(n919), .Z(n901) );
  BUFFD1 U165 ( .I(n920), .Z(n900) );
  BUFFD1 U166 ( .I(n920), .Z(n899) );
  BUFFD1 U167 ( .I(n921), .Z(n898) );
  BUFFD1 U168 ( .I(n921), .Z(n897) );
  BUFFD1 U169 ( .I(n922), .Z(n896) );
  BUFFD1 U170 ( .I(n922), .Z(n895) );
  BUFFD1 U171 ( .I(n923), .Z(n894) );
  BUFFD1 U172 ( .I(n923), .Z(n893) );
  BUFFD1 U173 ( .I(n924), .Z(n892) );
  BUFFD1 U174 ( .I(n924), .Z(n891) );
  BUFFD1 U175 ( .I(n925), .Z(n890) );
  BUFFD1 U176 ( .I(n925), .Z(n889) );
  BUFFD1 U177 ( .I(n926), .Z(n888) );
  BUFFD1 U178 ( .I(n926), .Z(n887) );
  BUFFD1 U179 ( .I(n927), .Z(n886) );
  BUFFD1 U180 ( .I(n927), .Z(n885) );
  BUFFD1 U181 ( .I(n928), .Z(n884) );
  BUFFD1 U182 ( .I(n928), .Z(n883) );
  BUFFD1 U183 ( .I(n929), .Z(n882) );
  BUFFD1 U184 ( .I(n929), .Z(n881) );
  BUFFD1 U185 ( .I(n930), .Z(n880) );
  BUFFD1 U186 ( .I(n930), .Z(n879) );
  BUFFD1 U187 ( .I(n931), .Z(n878) );
  BUFFD1 U188 ( .I(n931), .Z(n877) );
  BUFFD1 U189 ( .I(n932), .Z(n876) );
  BUFFD1 U190 ( .I(n932), .Z(n875) );
  BUFFD1 U191 ( .I(n933), .Z(n874) );
  BUFFD1 U192 ( .I(n933), .Z(n873) );
  BUFFD1 U193 ( .I(n934), .Z(n872) );
  BUFFD1 U194 ( .I(n934), .Z(n871) );
  BUFFD1 U195 ( .I(n935), .Z(n870) );
  BUFFD1 U196 ( .I(n935), .Z(n869) );
  BUFFD1 U197 ( .I(n936), .Z(n868) );
  BUFFD1 U198 ( .I(n936), .Z(n867) );
  BUFFD1 U199 ( .I(n937), .Z(n866) );
  BUFFD1 U200 ( .I(n937), .Z(n865) );
  BUFFD1 U201 ( .I(n938), .Z(n864) );
  BUFFD1 U202 ( .I(n938), .Z(n863) );
  BUFFD1 U203 ( .I(n939), .Z(n862) );
  BUFFD1 U204 ( .I(n939), .Z(n861) );
  BUFFD1 U205 ( .I(n940), .Z(n860) );
  BUFFD1 U206 ( .I(n940), .Z(n859) );
  BUFFD1 U207 ( .I(n941), .Z(n858) );
  BUFFD1 U208 ( .I(n941), .Z(n857) );
  BUFFD1 U209 ( .I(n942), .Z(n856) );
  BUFFD1 U210 ( .I(n942), .Z(n855) );
  BUFFD1 U211 ( .I(n943), .Z(n854) );
  BUFFD1 U212 ( .I(n943), .Z(n853) );
  BUFFD1 U213 ( .I(n944), .Z(n852) );
  BUFFD1 U214 ( .I(n944), .Z(n851) );
  BUFFD1 U215 ( .I(n945), .Z(n850) );
  BUFFD1 U216 ( .I(n945), .Z(n849) );
  BUFFD1 U217 ( .I(n946), .Z(n848) );
  BUFFD1 U218 ( .I(n946), .Z(n847) );
  BUFFD1 U219 ( .I(n713), .Z(n698) );
  BUFFD1 U220 ( .I(n702), .Z(n697) );
  BUFFD1 U221 ( .I(n702), .Z(n696) );
  BUFFD1 U222 ( .I(n702), .Z(n695) );
  BUFFD1 U223 ( .I(n703), .Z(n694) );
  BUFFD1 U224 ( .I(n703), .Z(n693) );
  BUFFD1 U225 ( .I(n704), .Z(n692) );
  BUFFD1 U226 ( .I(n704), .Z(n691) );
  BUFFD1 U227 ( .I(n705), .Z(n690) );
  BUFFD1 U228 ( .I(n705), .Z(n689) );
  BUFFD1 U229 ( .I(n706), .Z(n688) );
  BUFFD1 U230 ( .I(n706), .Z(n687) );
  BUFFD1 U231 ( .I(n707), .Z(n686) );
  BUFFD1 U232 ( .I(n707), .Z(n685) );
  BUFFD1 U233 ( .I(n708), .Z(n684) );
  BUFFD1 U234 ( .I(n708), .Z(n683) );
  BUFFD1 U235 ( .I(n709), .Z(n682) );
  BUFFD1 U236 ( .I(n709), .Z(n681) );
  BUFFD1 U237 ( .I(n710), .Z(n680) );
  BUFFD1 U238 ( .I(n710), .Z(n679) );
  INVD1 U239 ( .I(n845), .ZN(n844) );
  INVD1 U240 ( .I(n845), .ZN(n843) );
  INVD1 U241 ( .I(n845), .ZN(n842) );
  BUFFD1 U242 ( .I(n534), .Z(n539) );
  BUFFD1 U243 ( .I(n535), .Z(n538) );
  BUFFD1 U244 ( .I(n535), .Z(n537) );
  BUFFD1 U245 ( .I(n535), .Z(n536) );
  BUFFD1 U246 ( .I(n534), .Z(n541) );
  BUFFD1 U247 ( .I(n534), .Z(n540) );
  BUFFD1 U248 ( .I(N46), .Z(n521) );
  BUFFD1 U249 ( .I(n562), .Z(n572) );
  BUFFD1 U250 ( .I(n564), .Z(n569) );
  BUFFD1 U251 ( .I(n564), .Z(n568) );
  BUFFD1 U252 ( .I(n565), .Z(n567) );
  BUFFD1 U253 ( .I(n565), .Z(n566) );
  BUFFD1 U254 ( .I(n563), .Z(n570) );
  BUFFD1 U255 ( .I(n563), .Z(n571) );
  BUFFD1 U256 ( .I(n533), .Z(n520) );
  BUFFD1 U257 ( .I(n515), .Z(n518) );
  BUFFD1 U258 ( .I(n515), .Z(n517) );
  BUFFD1 U259 ( .I(n534), .Z(n542) );
  BUFFD1 U260 ( .I(N46), .Z(n522) );
  BUFFD1 U261 ( .I(n533), .Z(n519) );
  BUFFD1 U262 ( .I(n515), .Z(n516) );
  INVD1 U263 ( .I(n510), .ZN(n511) );
  INVD1 U264 ( .I(n510), .ZN(n512) );
  BUFFD1 U265 ( .I(n700), .Z(n597) );
  BUFFD1 U266 ( .I(n701), .Z(n700) );
  INVD1 U267 ( .I(N85), .ZN(n845) );
  BUFFD1 U268 ( .I(n713), .Z(n702) );
  BUFFD1 U269 ( .I(n713), .Z(n703) );
  BUFFD1 U270 ( .I(n713), .Z(n704) );
  BUFFD1 U271 ( .I(n712), .Z(n705) );
  BUFFD1 U272 ( .I(n712), .Z(n706) );
  BUFFD1 U273 ( .I(n712), .Z(n707) );
  BUFFD1 U274 ( .I(n711), .Z(n708) );
  BUFFD1 U275 ( .I(n711), .Z(n709) );
  BUFFD1 U276 ( .I(n711), .Z(n710) );
  BUFFD1 U277 ( .I(n846), .Z(n913) );
  BUFFD1 U278 ( .I(n957), .Z(n914) );
  BUFFD1 U279 ( .I(n957), .Z(n915) );
  BUFFD1 U280 ( .I(n957), .Z(n916) );
  BUFFD1 U281 ( .I(n956), .Z(n917) );
  BUFFD1 U282 ( .I(n956), .Z(n918) );
  BUFFD1 U283 ( .I(n956), .Z(n919) );
  BUFFD1 U284 ( .I(n955), .Z(n920) );
  BUFFD1 U285 ( .I(n955), .Z(n921) );
  BUFFD1 U286 ( .I(n955), .Z(n922) );
  BUFFD1 U287 ( .I(n954), .Z(n923) );
  BUFFD1 U288 ( .I(n954), .Z(n924) );
  BUFFD1 U289 ( .I(n954), .Z(n925) );
  BUFFD1 U290 ( .I(n953), .Z(n926) );
  BUFFD1 U291 ( .I(n953), .Z(n927) );
  BUFFD1 U292 ( .I(n953), .Z(n928) );
  BUFFD1 U293 ( .I(n952), .Z(n929) );
  BUFFD1 U294 ( .I(n952), .Z(n930) );
  BUFFD1 U295 ( .I(n952), .Z(n931) );
  BUFFD1 U296 ( .I(n951), .Z(n932) );
  BUFFD1 U297 ( .I(n951), .Z(n933) );
  BUFFD1 U298 ( .I(n951), .Z(n934) );
  BUFFD1 U299 ( .I(n950), .Z(n935) );
  BUFFD1 U300 ( .I(n950), .Z(n936) );
  BUFFD1 U301 ( .I(n950), .Z(n937) );
  BUFFD1 U302 ( .I(n949), .Z(n938) );
  BUFFD1 U303 ( .I(n949), .Z(n939) );
  BUFFD1 U304 ( .I(n949), .Z(n940) );
  BUFFD1 U305 ( .I(n948), .Z(n941) );
  BUFFD1 U306 ( .I(n948), .Z(n942) );
  BUFFD1 U307 ( .I(n948), .Z(n943) );
  BUFFD1 U308 ( .I(n947), .Z(n944) );
  BUFFD1 U309 ( .I(n947), .Z(n945) );
  BUFFD1 U310 ( .I(n947), .Z(n946) );
  BUFFD1 U311 ( .I(n701), .Z(n699) );
  BUFFD1 U312 ( .I(n964), .Z(n513) );
  BUFFD1 U313 ( .I(n964), .Z(n514) );
  BUFFD1 U314 ( .I(n964), .Z(n515) );
  BUFFD1 U315 ( .I(n963), .Z(n535) );
  BUFFD1 U316 ( .I(n963), .Z(n534) );
  BUFFD1 U317 ( .I(N44), .Z(n562) );
  BUFFD1 U318 ( .I(N44), .Z(n564) );
  BUFFD1 U319 ( .I(N44), .Z(n565) );
  BUFFD1 U320 ( .I(N44), .Z(n563) );
  BUFFD1 U321 ( .I(N46), .Z(n533) );
  XOR3D1 U322 ( .A1(n80), .A2(n1006), .A3(n81), .Z(n79) );
  XOR3D1 U323 ( .A1(n1042), .A2(n1038), .A3(n82), .Z(n81) );
  XOR3D1 U324 ( .A1(n83), .A2(n1034), .A3(n84), .Z(n82) );
  XOR3D1 U325 ( .A1(n986), .A2(n982), .A3(n76), .Z(n75) );
  XOR3D1 U326 ( .A1(n77), .A2(n978), .A3(n78), .Z(n76) );
  XOR3D1 U327 ( .A1(n1014), .A2(n1010), .A3(n79), .Z(n78) );
  XOR3D1 U328 ( .A1(n974), .A2(n970), .A3(n73), .Z(N85) );
  XOR3D1 U329 ( .A1(n966), .A2(n74), .A3(n75), .Z(n73) );
  BUFFD1 U330 ( .I(n681), .Z(n701) );
  BUFFD1 U331 ( .I(n596), .Z(n713) );
  BUFFD1 U332 ( .I(n595), .Z(n712) );
  BUFFD1 U333 ( .I(n595), .Z(n711) );
  BUFFD1 U334 ( .I(n936), .Z(n957) );
  BUFFD1 U335 ( .I(n958), .Z(n956) );
  BUFFD1 U336 ( .I(n958), .Z(n955) );
  BUFFD1 U337 ( .I(n959), .Z(n954) );
  BUFFD1 U338 ( .I(n959), .Z(n953) );
  BUFFD1 U339 ( .I(n960), .Z(n952) );
  BUFFD1 U340 ( .I(n960), .Z(n951) );
  BUFFD1 U341 ( .I(n961), .Z(n950) );
  BUFFD1 U342 ( .I(n961), .Z(n949) );
  BUFFD1 U343 ( .I(n962), .Z(n948) );
  BUFFD1 U344 ( .I(n962), .Z(n947) );
  INVD1 U345 ( .I(n765), .ZN(n764) );
  INVD1 U346 ( .I(n765), .ZN(n763) );
  INVD1 U347 ( .I(n765), .ZN(n762) );
  INVD1 U348 ( .I(n761), .ZN(n760) );
  INVD1 U349 ( .I(n761), .ZN(n759) );
  INVD1 U350 ( .I(n761), .ZN(n758) );
  INVD1 U351 ( .I(n757), .ZN(n756) );
  INVD1 U352 ( .I(n757), .ZN(n755) );
  INVD1 U353 ( .I(n757), .ZN(n754) );
  INVD1 U354 ( .I(n753), .ZN(n752) );
  INVD1 U355 ( .I(n753), .ZN(n751) );
  INVD1 U356 ( .I(n753), .ZN(n750) );
  INVD1 U357 ( .I(n749), .ZN(n748) );
  INVD1 U358 ( .I(n749), .ZN(n747) );
  INVD1 U359 ( .I(n749), .ZN(n746) );
  INVD1 U360 ( .I(n745), .ZN(n744) );
  INVD1 U361 ( .I(n745), .ZN(n743) );
  INVD1 U362 ( .I(n745), .ZN(n742) );
  INVD1 U363 ( .I(n741), .ZN(n740) );
  INVD1 U364 ( .I(n741), .ZN(n739) );
  INVD1 U365 ( .I(n741), .ZN(n738) );
  INVD1 U366 ( .I(n737), .ZN(n736) );
  INVD1 U367 ( .I(n737), .ZN(n735) );
  INVD1 U368 ( .I(n737), .ZN(n734) );
  INVD1 U369 ( .I(n733), .ZN(n732) );
  INVD1 U370 ( .I(n733), .ZN(n731) );
  INVD1 U371 ( .I(n733), .ZN(n730) );
  INVD1 U372 ( .I(n729), .ZN(n728) );
  INVD1 U373 ( .I(n729), .ZN(n727) );
  INVD1 U374 ( .I(n729), .ZN(n726) );
  INVD1 U375 ( .I(n725), .ZN(n724) );
  INVD1 U376 ( .I(n725), .ZN(n723) );
  INVD1 U377 ( .I(n725), .ZN(n722) );
  INVD1 U378 ( .I(n721), .ZN(n720) );
  INVD1 U379 ( .I(n721), .ZN(n719) );
  INVD1 U380 ( .I(n721), .ZN(n718) );
  INVD1 U381 ( .I(n717), .ZN(n716) );
  INVD1 U382 ( .I(n717), .ZN(n715) );
  INVD1 U383 ( .I(n717), .ZN(n714) );
  INVD1 U384 ( .I(n841), .ZN(n840) );
  INVD1 U385 ( .I(n841), .ZN(n839) );
  INVD1 U386 ( .I(n841), .ZN(n838) );
  INVD1 U387 ( .I(n837), .ZN(n836) );
  INVD1 U388 ( .I(n837), .ZN(n835) );
  INVD1 U389 ( .I(n837), .ZN(n834) );
  INVD1 U390 ( .I(n833), .ZN(n832) );
  INVD1 U391 ( .I(n833), .ZN(n831) );
  INVD1 U392 ( .I(n833), .ZN(n830) );
  INVD1 U393 ( .I(n829), .ZN(n828) );
  INVD1 U394 ( .I(n829), .ZN(n827) );
  INVD1 U395 ( .I(n829), .ZN(n826) );
  INVD1 U396 ( .I(n825), .ZN(n824) );
  INVD1 U397 ( .I(n825), .ZN(n823) );
  INVD1 U398 ( .I(n825), .ZN(n822) );
  INVD1 U399 ( .I(n821), .ZN(n820) );
  INVD1 U400 ( .I(n821), .ZN(n819) );
  INVD1 U401 ( .I(n821), .ZN(n818) );
  INVD1 U402 ( .I(n817), .ZN(n816) );
  INVD1 U403 ( .I(n817), .ZN(n815) );
  INVD1 U404 ( .I(n817), .ZN(n814) );
  INVD1 U405 ( .I(n813), .ZN(n812) );
  INVD1 U406 ( .I(n813), .ZN(n811) );
  INVD1 U407 ( .I(n813), .ZN(n810) );
  INVD1 U408 ( .I(n809), .ZN(n808) );
  INVD1 U409 ( .I(n809), .ZN(n807) );
  INVD1 U410 ( .I(n809), .ZN(n806) );
  INVD1 U411 ( .I(n805), .ZN(n804) );
  INVD1 U412 ( .I(n805), .ZN(n803) );
  INVD1 U413 ( .I(n805), .ZN(n802) );
  INVD1 U414 ( .I(n801), .ZN(n800) );
  INVD1 U415 ( .I(n801), .ZN(n799) );
  INVD1 U416 ( .I(n801), .ZN(n798) );
  INVD1 U417 ( .I(n797), .ZN(n796) );
  INVD1 U418 ( .I(n797), .ZN(n795) );
  INVD1 U419 ( .I(n797), .ZN(n794) );
  INVD1 U420 ( .I(n793), .ZN(n792) );
  INVD1 U421 ( .I(n793), .ZN(n791) );
  INVD1 U422 ( .I(n793), .ZN(n790) );
  INVD1 U423 ( .I(n789), .ZN(n788) );
  INVD1 U424 ( .I(n789), .ZN(n787) );
  INVD1 U425 ( .I(n789), .ZN(n786) );
  INVD1 U426 ( .I(n785), .ZN(n784) );
  INVD1 U427 ( .I(n785), .ZN(n783) );
  INVD1 U428 ( .I(n785), .ZN(n782) );
  INVD1 U429 ( .I(n781), .ZN(n780) );
  INVD1 U430 ( .I(n781), .ZN(n779) );
  INVD1 U431 ( .I(n781), .ZN(n778) );
  INVD1 U432 ( .I(n777), .ZN(n776) );
  INVD1 U433 ( .I(n777), .ZN(n775) );
  INVD1 U434 ( .I(n777), .ZN(n774) );
  INVD1 U435 ( .I(n773), .ZN(n772) );
  INVD1 U436 ( .I(n773), .ZN(n771) );
  INVD1 U437 ( .I(n773), .ZN(n770) );
  INVD1 U438 ( .I(n769), .ZN(n768) );
  INVD1 U439 ( .I(n769), .ZN(n767) );
  INVD1 U440 ( .I(n769), .ZN(n766) );
  XOR3D1 U441 ( .A1(N60), .A2(N59), .A3(n95), .Z(n94) );
  XOR3D1 U442 ( .A1(n96), .A2(N58), .A3(n97), .Z(n95) );
  XOR3D1 U443 ( .A1(N79), .A2(N74), .A3(n86), .Z(N83) );
  XOR3D1 U444 ( .A1(N73), .A2(n87), .A3(n88), .Z(n86) );
  XOR3D1 U445 ( .A1(N77), .A2(N76), .A3(n89), .Z(n88) );
  XOR3D1 U446 ( .A1(N67), .A2(N66), .A3(n92), .Z(n90) );
  XOR3D1 U447 ( .A1(N65), .A2(n93), .A3(n94), .Z(n92) );
  BUFFD1 U448 ( .I(N45), .Z(n963) );
  BUFFD1 U449 ( .I(N47), .Z(n964) );
  INVD1 U450 ( .I(n965), .ZN(n510) );
  BUFFD1 U451 ( .I(N48), .Z(n965) );
  INVD1 U452 ( .I(N150), .ZN(n841) );
  INVD1 U453 ( .I(N183), .ZN(n837) );
  INVD1 U454 ( .I(N216), .ZN(n833) );
  INVD1 U455 ( .I(N249), .ZN(n829) );
  INVD1 U456 ( .I(N282), .ZN(n825) );
  INVD1 U457 ( .I(N315), .ZN(n821) );
  INVD1 U458 ( .I(N348), .ZN(n817) );
  INVD1 U459 ( .I(N381), .ZN(n813) );
  INVD1 U460 ( .I(N414), .ZN(n809) );
  INVD1 U461 ( .I(N447), .ZN(n805) );
  INVD1 U462 ( .I(N480), .ZN(n801) );
  INVD1 U463 ( .I(N513), .ZN(n797) );
  INVD1 U464 ( .I(N546), .ZN(n793) );
  INVD1 U465 ( .I(N579), .ZN(n789) );
  INVD1 U466 ( .I(N612), .ZN(n785) );
  INVD1 U467 ( .I(N645), .ZN(n781) );
  INVD1 U468 ( .I(N678), .ZN(n777) );
  INVD1 U469 ( .I(N711), .ZN(n773) );
  INVD1 U470 ( .I(N744), .ZN(n769) );
  INVD1 U471 ( .I(N777), .ZN(n765) );
  INVD1 U472 ( .I(N810), .ZN(n761) );
  INVD1 U473 ( .I(N843), .ZN(n757) );
  INVD1 U474 ( .I(N876), .ZN(n753) );
  INVD1 U475 ( .I(N909), .ZN(n749) );
  INVD1 U476 ( .I(N942), .ZN(n745) );
  INVD1 U477 ( .I(N975), .ZN(n741) );
  INVD1 U478 ( .I(N999), .ZN(n737) );
  INVD1 U479 ( .I(N1041), .ZN(n733) );
  INVD1 U480 ( .I(N1074), .ZN(n729) );
  INVD1 U481 ( .I(N1107), .ZN(n725) );
  INVD1 U482 ( .I(N1140), .ZN(n721) );
  INVD1 U483 ( .I(N1173), .ZN(n717) );
  BUFFD1 U484 ( .I(n5), .Z(n596) );
  BUFFD1 U485 ( .I(n702), .Z(n595) );
  BUFFD1 U486 ( .I(n960), .Z(n958) );
  BUFFD1 U487 ( .I(n949), .Z(n959) );
  BUFFD1 U488 ( .I(n846), .Z(n960) );
  BUFFD1 U489 ( .I(n846), .Z(n961) );
  BUFFD1 U490 ( .I(n846), .Z(n962) );
  INVD1 U491 ( .I(n997), .ZN(n994) );
  INVD1 U492 ( .I(n1001), .ZN(n998) );
  INVD1 U493 ( .I(n1025), .ZN(n1022) );
  INVD1 U494 ( .I(n1029), .ZN(n1026) );
  INVD1 U495 ( .I(n1053), .ZN(n1050) );
  INVD1 U496 ( .I(n1057), .ZN(n1054) );
  INVD1 U497 ( .I(n1069), .ZN(n1066) );
  INVD1 U498 ( .I(n1073), .ZN(n1070) );
  INVD1 U499 ( .I(n1085), .ZN(n1082) );
  INVD1 U500 ( .I(n1089), .ZN(n1086) );
  INVD1 U501 ( .I(n973), .ZN(n970) );
  INVD1 U502 ( .I(n981), .ZN(n978) );
  INVD1 U503 ( .I(n985), .ZN(n982) );
  INVD1 U504 ( .I(n1009), .ZN(n1006) );
  INVD1 U505 ( .I(n1013), .ZN(n1010) );
  INVD1 U506 ( .I(n1037), .ZN(n1034) );
  INVD1 U507 ( .I(n1041), .ZN(n1038) );
  INVD1 U508 ( .I(n993), .ZN(n990) );
  INVD1 U509 ( .I(n1005), .ZN(n1002) );
  INVD1 U510 ( .I(n1021), .ZN(n1018) );
  INVD1 U511 ( .I(n1033), .ZN(n1030) );
  INVD1 U512 ( .I(n1049), .ZN(n1046) );
  INVD1 U513 ( .I(n1061), .ZN(n1058) );
  INVD1 U514 ( .I(n1065), .ZN(n1062) );
  INVD1 U515 ( .I(n1077), .ZN(n1074) );
  INVD1 U516 ( .I(n1081), .ZN(n1078) );
  INVD1 U517 ( .I(n1093), .ZN(n1090) );
  INVD1 U518 ( .I(n969), .ZN(n966) );
  INVD1 U519 ( .I(n977), .ZN(n974) );
  INVD1 U520 ( .I(n989), .ZN(n986) );
  INVD1 U521 ( .I(n1017), .ZN(n1014) );
  INVD1 U522 ( .I(n1045), .ZN(n1042) );
  INVD1 U523 ( .I(n969), .ZN(n967) );
  INVD1 U524 ( .I(n973), .ZN(n971) );
  INVD1 U525 ( .I(n977), .ZN(n975) );
  INVD1 U526 ( .I(n981), .ZN(n979) );
  INVD1 U527 ( .I(n985), .ZN(n983) );
  INVD1 U528 ( .I(n989), .ZN(n987) );
  INVD1 U529 ( .I(n993), .ZN(n991) );
  INVD1 U530 ( .I(n997), .ZN(n995) );
  INVD1 U531 ( .I(n1001), .ZN(n999) );
  INVD1 U532 ( .I(n1005), .ZN(n1003) );
  INVD1 U533 ( .I(n1009), .ZN(n1007) );
  INVD1 U534 ( .I(n1013), .ZN(n1011) );
  INVD1 U535 ( .I(n1017), .ZN(n1015) );
  INVD1 U536 ( .I(n1021), .ZN(n1019) );
  INVD1 U537 ( .I(n1025), .ZN(n1023) );
  INVD1 U538 ( .I(n1029), .ZN(n1027) );
  INVD1 U539 ( .I(n1033), .ZN(n1031) );
  INVD1 U540 ( .I(n1037), .ZN(n1035) );
  INVD1 U541 ( .I(n1041), .ZN(n1039) );
  INVD1 U542 ( .I(n1045), .ZN(n1043) );
  INVD1 U543 ( .I(n1049), .ZN(n1047) );
  INVD1 U544 ( .I(n1053), .ZN(n1051) );
  INVD1 U545 ( .I(n1057), .ZN(n1055) );
  INVD1 U546 ( .I(n1061), .ZN(n1059) );
  INVD1 U547 ( .I(n1065), .ZN(n1063) );
  INVD1 U548 ( .I(n1069), .ZN(n1067) );
  INVD1 U549 ( .I(n1073), .ZN(n1071) );
  INVD1 U550 ( .I(n1077), .ZN(n1075) );
  INVD1 U551 ( .I(n1081), .ZN(n1079) );
  INVD1 U552 ( .I(n1085), .ZN(n1083) );
  INVD1 U553 ( .I(n1089), .ZN(n1087) );
  INVD1 U554 ( .I(n1093), .ZN(n1091) );
  INVD1 U555 ( .I(n969), .ZN(n968) );
  INVD1 U556 ( .I(n973), .ZN(n972) );
  INVD1 U557 ( .I(n977), .ZN(n976) );
  INVD1 U558 ( .I(n981), .ZN(n980) );
  INVD1 U559 ( .I(n985), .ZN(n984) );
  INVD1 U560 ( .I(n989), .ZN(n988) );
  INVD1 U561 ( .I(n993), .ZN(n992) );
  INVD1 U562 ( .I(n997), .ZN(n996) );
  INVD1 U563 ( .I(n1001), .ZN(n1000) );
  INVD1 U564 ( .I(n1005), .ZN(n1004) );
  INVD1 U565 ( .I(n1009), .ZN(n1008) );
  INVD1 U566 ( .I(n1013), .ZN(n1012) );
  INVD1 U567 ( .I(n1017), .ZN(n1016) );
  INVD1 U568 ( .I(n1021), .ZN(n1020) );
  INVD1 U569 ( .I(n1025), .ZN(n1024) );
  INVD1 U570 ( .I(n1029), .ZN(n1028) );
  INVD1 U571 ( .I(n1033), .ZN(n1032) );
  INVD1 U572 ( .I(n1037), .ZN(n1036) );
  INVD1 U573 ( .I(n1041), .ZN(n1040) );
  INVD1 U574 ( .I(n1045), .ZN(n1044) );
  INVD1 U575 ( .I(n1049), .ZN(n1048) );
  INVD1 U576 ( .I(n1053), .ZN(n1052) );
  INVD1 U577 ( .I(n1057), .ZN(n1056) );
  INVD1 U578 ( .I(n1061), .ZN(n1060) );
  INVD1 U579 ( .I(n1065), .ZN(n1064) );
  INVD1 U580 ( .I(n1069), .ZN(n1068) );
  INVD1 U581 ( .I(n1073), .ZN(n1072) );
  INVD1 U582 ( .I(n1077), .ZN(n1076) );
  INVD1 U583 ( .I(n1081), .ZN(n1080) );
  INVD1 U584 ( .I(n1085), .ZN(n1084) );
  INVD1 U585 ( .I(n1089), .ZN(n1088) );
  INVD1 U586 ( .I(n1093), .ZN(n1092) );
  ND3D1 U587 ( .A1(n106), .A2(n105), .A3(n104), .ZN(n69) );
  ND3D1 U588 ( .A1(n104), .A2(n105), .A3(AddrW[1]), .ZN(n67) );
  INVD1 U589 ( .I(AddrW[1]), .ZN(n106) );
  INVD1 U590 ( .I(DataI[0]), .ZN(n969) );
  INVD1 U591 ( .I(DataI[1]), .ZN(n973) );
  INVD1 U592 ( .I(DataI[2]), .ZN(n977) );
  INVD1 U593 ( .I(DataI[3]), .ZN(n981) );
  INVD1 U594 ( .I(DataI[4]), .ZN(n985) );
  INVD1 U595 ( .I(DataI[5]), .ZN(n989) );
  INVD1 U596 ( .I(DataI[10]), .ZN(n1009) );
  INVD1 U597 ( .I(DataI[11]), .ZN(n1013) );
  INVD1 U598 ( .I(DataI[12]), .ZN(n1017) );
  INVD1 U599 ( .I(DataI[17]), .ZN(n1037) );
  INVD1 U600 ( .I(DataI[18]), .ZN(n1041) );
  INVD1 U601 ( .I(DataI[19]), .ZN(n1045) );
  INVD1 U602 ( .I(DataI[6]), .ZN(n993) );
  INVD1 U603 ( .I(DataI[7]), .ZN(n997) );
  INVD1 U604 ( .I(DataI[8]), .ZN(n1001) );
  INVD1 U605 ( .I(DataI[9]), .ZN(n1005) );
  INVD1 U606 ( .I(DataI[13]), .ZN(n1021) );
  INVD1 U607 ( .I(DataI[14]), .ZN(n1025) );
  INVD1 U608 ( .I(DataI[15]), .ZN(n1029) );
  INVD1 U609 ( .I(DataI[16]), .ZN(n1033) );
  INVD1 U610 ( .I(DataI[20]), .ZN(n1049) );
  INVD1 U611 ( .I(DataI[21]), .ZN(n1053) );
  INVD1 U612 ( .I(DataI[22]), .ZN(n1057) );
  INVD1 U613 ( .I(DataI[23]), .ZN(n1061) );
  INVD1 U614 ( .I(DataI[24]), .ZN(n1065) );
  INVD1 U615 ( .I(DataI[25]), .ZN(n1069) );
  INVD1 U616 ( .I(DataI[26]), .ZN(n1073) );
  INVD1 U617 ( .I(DataI[27]), .ZN(n1077) );
  INVD1 U618 ( .I(DataI[28]), .ZN(n1081) );
  INVD1 U619 ( .I(DataI[29]), .ZN(n1085) );
  INVD1 U620 ( .I(DataI[30]), .ZN(n1089) );
  INVD1 U621 ( .I(DataI[31]), .ZN(n1093) );
  BUFFD1 U622 ( .I(ClockW), .Z(n846) );
  NR2D1 U623 ( .A1(n70), .A2(n99), .ZN(N777) );
  NR2D1 U624 ( .A1(n70), .A2(n98), .ZN(N810) );
  NR2D1 U625 ( .A1(n70), .A2(n85), .ZN(N843) );
  NR2D1 U626 ( .A1(n70), .A2(n72), .ZN(N876) );
  NR2D1 U627 ( .A1(n70), .A2(n71), .ZN(N909) );
  NR2D1 U628 ( .A1(n66), .A2(n69), .ZN(N942) );
  NR2D1 U629 ( .A1(n66), .A2(n68), .ZN(N975) );
  NR2D1 U630 ( .A1(n66), .A2(n67), .ZN(N999) );
  NR2D1 U631 ( .A1(n66), .A2(n99), .ZN(N1041) );
  NR2D1 U632 ( .A1(n66), .A2(n98), .ZN(N1074) );
  NR2D1 U633 ( .A1(n66), .A2(n85), .ZN(N1107) );
  NR2D1 U634 ( .A1(n66), .A2(n72), .ZN(N1140) );
  NR2D1 U635 ( .A1(n66), .A2(n71), .ZN(N1173) );
  NR2D1 U636 ( .A1(n69), .A2(n103), .ZN(N150) );
  NR2D1 U637 ( .A1(n68), .A2(n103), .ZN(N183) );
  NR2D1 U638 ( .A1(n67), .A2(n103), .ZN(N216) );
  NR2D1 U639 ( .A1(n99), .A2(n103), .ZN(N249) );
  NR2D1 U640 ( .A1(n98), .A2(n103), .ZN(N282) );
  NR2D1 U641 ( .A1(n85), .A2(n103), .ZN(N315) );
  NR2D1 U642 ( .A1(n72), .A2(n103), .ZN(N348) );
  NR2D1 U643 ( .A1(n71), .A2(n103), .ZN(N381) );
  NR2D1 U644 ( .A1(n69), .A2(n101), .ZN(N414) );
  NR2D1 U645 ( .A1(n68), .A2(n101), .ZN(N447) );
  NR2D1 U646 ( .A1(n67), .A2(n101), .ZN(N480) );
  NR2D1 U647 ( .A1(n99), .A2(n101), .ZN(N513) );
  NR2D1 U648 ( .A1(n98), .A2(n101), .ZN(N546) );
  NR2D1 U649 ( .A1(n85), .A2(n101), .ZN(N579) );
  NR2D1 U650 ( .A1(n72), .A2(n101), .ZN(N612) );
  NR2D1 U651 ( .A1(n71), .A2(n101), .ZN(N645) );
  NR2D1 U652 ( .A1(n69), .A2(n70), .ZN(N678) );
  NR2D1 U653 ( .A1(n68), .A2(n70), .ZN(N711) );
  NR2D1 U654 ( .A1(n67), .A2(n70), .ZN(N744) );
  MUX4ND0 U655 ( .I0(\Storage[28][32] ), .I1(\Storage[29][32] ), .I2(
        \Storage[30][32] ), .I3(\Storage[31][32] ), .S0(n576), .S1(n543), .ZN(
        n500) );
  MUX4ND0 U656 ( .I0(\Storage[28][0] ), .I1(\Storage[29][0] ), .I2(
        \Storage[30][0] ), .I3(\Storage[31][0] ), .S0(n576), .S1(n543), .ZN(
        n42) );
  MUX4ND0 U657 ( .I0(\Storage[28][1] ), .I1(\Storage[29][1] ), .I2(
        \Storage[30][1] ), .I3(\Storage[31][1] ), .S0(n569), .S1(n963), .ZN(
        n55) );
  MUX4ND0 U658 ( .I0(\Storage[28][2] ), .I1(\Storage[29][2] ), .I2(
        \Storage[30][2] ), .I3(\Storage[31][2] ), .S0(n573), .S1(n535), .ZN(
        n110) );
  MUX4ND0 U659 ( .I0(\Storage[28][3] ), .I1(\Storage[29][3] ), .I2(
        \Storage[30][3] ), .I3(\Storage[31][3] ), .S0(n567), .S1(n540), .ZN(
        n123) );
  MUX4ND0 U660 ( .I0(\Storage[28][4] ), .I1(\Storage[29][4] ), .I2(
        \Storage[30][4] ), .I3(\Storage[31][4] ), .S0(n572), .S1(n543), .ZN(
        n136) );
  MUX4ND0 U661 ( .I0(\Storage[28][5] ), .I1(\Storage[29][5] ), .I2(
        \Storage[30][5] ), .I3(\Storage[31][5] ), .S0(n568), .S1(n543), .ZN(
        n149) );
  MUX4ND0 U662 ( .I0(\Storage[28][6] ), .I1(\Storage[29][6] ), .I2(
        \Storage[30][6] ), .I3(\Storage[31][6] ), .S0(n567), .S1(n963), .ZN(
        n162) );
  MUX4ND0 U663 ( .I0(\Storage[28][7] ), .I1(\Storage[29][7] ), .I2(
        \Storage[30][7] ), .I3(\Storage[31][7] ), .S0(n568), .S1(n543), .ZN(
        n175) );
  MUX4ND0 U664 ( .I0(\Storage[28][8] ), .I1(\Storage[29][8] ), .I2(
        \Storage[30][8] ), .I3(\Storage[31][8] ), .S0(n572), .S1(n540), .ZN(
        n188) );
  MUX4ND0 U665 ( .I0(\Storage[28][9] ), .I1(\Storage[29][9] ), .I2(
        \Storage[30][9] ), .I3(\Storage[31][9] ), .S0(n573), .S1(n545), .ZN(
        n201) );
  MUX4ND0 U666 ( .I0(\Storage[28][10] ), .I1(\Storage[29][10] ), .I2(
        \Storage[30][10] ), .I3(\Storage[31][10] ), .S0(n564), .S1(n545), .ZN(
        n214) );
  MUX4ND0 U667 ( .I0(\Storage[28][11] ), .I1(\Storage[29][11] ), .I2(
        \Storage[30][11] ), .I3(\Storage[31][11] ), .S0(n566), .S1(n545), .ZN(
        n227) );
  MUX4ND0 U668 ( .I0(\Storage[28][12] ), .I1(\Storage[29][12] ), .I2(
        \Storage[30][12] ), .I3(\Storage[31][12] ), .S0(n568), .S1(n545), .ZN(
        n240) );
  MUX4ND0 U669 ( .I0(\Storage[28][13] ), .I1(\Storage[29][13] ), .I2(
        \Storage[30][13] ), .I3(\Storage[31][13] ), .S0(n567), .S1(n545), .ZN(
        n253) );
  MUX4ND0 U670 ( .I0(\Storage[28][14] ), .I1(\Storage[29][14] ), .I2(
        \Storage[30][14] ), .I3(\Storage[31][14] ), .S0(n570), .S1(n545), .ZN(
        n266) );
  MUX4ND0 U671 ( .I0(\Storage[28][15] ), .I1(\Storage[29][15] ), .I2(
        \Storage[30][15] ), .I3(\Storage[31][15] ), .S0(n568), .S1(n545), .ZN(
        n279) );
  MUX4ND0 U672 ( .I0(\Storage[28][16] ), .I1(\Storage[29][16] ), .I2(
        \Storage[30][16] ), .I3(\Storage[31][16] ), .S0(n567), .S1(n545), .ZN(
        n292) );
  MUX4ND0 U673 ( .I0(\Storage[28][17] ), .I1(\Storage[29][17] ), .I2(
        \Storage[30][17] ), .I3(\Storage[31][17] ), .S0(n566), .S1(n545), .ZN(
        n305) );
  MUX4ND0 U674 ( .I0(\Storage[28][18] ), .I1(\Storage[29][18] ), .I2(
        \Storage[30][18] ), .I3(\Storage[31][18] ), .S0(n570), .S1(n545), .ZN(
        n318) );
  MUX4ND0 U675 ( .I0(\Storage[28][19] ), .I1(\Storage[29][19] ), .I2(
        \Storage[30][19] ), .I3(\Storage[31][19] ), .S0(n568), .S1(n544), .ZN(
        n331) );
  MUX4ND0 U676 ( .I0(\Storage[28][20] ), .I1(\Storage[29][20] ), .I2(
        \Storage[30][20] ), .I3(\Storage[31][20] ), .S0(n573), .S1(n544), .ZN(
        n344) );
  MUX4ND0 U677 ( .I0(\Storage[28][21] ), .I1(\Storage[29][21] ), .I2(
        \Storage[30][21] ), .I3(\Storage[31][21] ), .S0(n572), .S1(n544), .ZN(
        n357) );
  MUX4ND0 U678 ( .I0(\Storage[28][22] ), .I1(\Storage[29][22] ), .I2(
        \Storage[30][22] ), .I3(\Storage[31][22] ), .S0(n575), .S1(n544), .ZN(
        n370) );
  MUX4ND0 U679 ( .I0(\Storage[28][23] ), .I1(\Storage[29][23] ), .I2(
        \Storage[30][23] ), .I3(\Storage[31][23] ), .S0(n575), .S1(n544), .ZN(
        n383) );
  MUX4ND0 U680 ( .I0(\Storage[28][24] ), .I1(\Storage[29][24] ), .I2(
        \Storage[30][24] ), .I3(\Storage[31][24] ), .S0(n575), .S1(n544), .ZN(
        n396) );
  MUX4ND0 U681 ( .I0(\Storage[28][25] ), .I1(\Storage[29][25] ), .I2(
        \Storage[30][25] ), .I3(\Storage[31][25] ), .S0(n575), .S1(n544), .ZN(
        n409) );
  MUX4ND0 U682 ( .I0(\Storage[28][26] ), .I1(\Storage[29][26] ), .I2(
        \Storage[30][26] ), .I3(\Storage[31][26] ), .S0(n575), .S1(n544), .ZN(
        n422) );
  MUX4ND0 U683 ( .I0(\Storage[28][27] ), .I1(\Storage[29][27] ), .I2(
        \Storage[30][27] ), .I3(\Storage[31][27] ), .S0(n575), .S1(n544), .ZN(
        n435) );
  MUX4ND0 U684 ( .I0(\Storage[28][28] ), .I1(\Storage[29][28] ), .I2(
        \Storage[30][28] ), .I3(\Storage[31][28] ), .S0(n575), .S1(n544), .ZN(
        n448) );
  MUX4ND0 U685 ( .I0(\Storage[28][29] ), .I1(\Storage[29][29] ), .I2(
        \Storage[30][29] ), .I3(\Storage[31][29] ), .S0(n575), .S1(n543), .ZN(
        n461) );
  MUX4ND0 U686 ( .I0(\Storage[28][30] ), .I1(\Storage[29][30] ), .I2(
        \Storage[30][30] ), .I3(\Storage[31][30] ), .S0(n575), .S1(n543), .ZN(
        n474) );
  MUX4ND0 U687 ( .I0(\Storage[28][31] ), .I1(\Storage[29][31] ), .I2(
        \Storage[30][31] ), .I3(\Storage[31][31] ), .S0(n575), .S1(n543), .ZN(
        n487) );
  MUX4D0 U688 ( .I0(\Storage[20][32] ), .I1(\Storage[21][32] ), .I2(
        \Storage[22][32] ), .I3(\Storage[23][32] ), .S0(n576), .S1(n550), .Z(
        n501) );
  MUX4D0 U689 ( .I0(\Storage[20][0] ), .I1(\Storage[21][0] ), .I2(
        \Storage[22][0] ), .I3(\Storage[23][0] ), .S0(n587), .S1(n558), .Z(n43) );
  MUX4D0 U690 ( .I0(\Storage[20][1] ), .I1(\Storage[21][1] ), .I2(
        \Storage[22][1] ), .I3(\Storage[23][1] ), .S0(n580), .S1(n551), .Z(n56) );
  MUX4D0 U691 ( .I0(\Storage[20][2] ), .I1(\Storage[21][2] ), .I2(
        \Storage[22][2] ), .I3(\Storage[23][2] ), .S0(n581), .S1(n552), .Z(
        n111) );
  MUX4D0 U692 ( .I0(\Storage[20][4] ), .I1(\Storage[21][4] ), .I2(
        \Storage[22][4] ), .I3(\Storage[23][4] ), .S0(n582), .S1(n553), .Z(
        n137) );
  MUX4D0 U693 ( .I0(\Storage[20][5] ), .I1(\Storage[21][5] ), .I2(
        \Storage[22][5] ), .I3(\Storage[23][5] ), .S0(n583), .S1(n554), .Z(
        n150) );
  MUX4D0 U694 ( .I0(\Storage[20][6] ), .I1(\Storage[21][6] ), .I2(
        \Storage[22][6] ), .I3(\Storage[23][6] ), .S0(n583), .S1(n554), .Z(
        n163) );
  MUX4D0 U695 ( .I0(\Storage[20][7] ), .I1(\Storage[21][7] ), .I2(
        \Storage[22][7] ), .I3(\Storage[23][7] ), .S0(n584), .S1(n555), .Z(
        n176) );
  MUX4D0 U696 ( .I0(\Storage[20][9] ), .I1(\Storage[21][9] ), .I2(
        \Storage[22][9] ), .I3(\Storage[23][9] ), .S0(n585), .S1(n536), .Z(
        n202) );
  MUX4D0 U697 ( .I0(\Storage[20][10] ), .I1(\Storage[21][10] ), .I2(
        \Storage[22][10] ), .I3(\Storage[23][10] ), .S0(n586), .S1(n538), .Z(
        n215) );
  MUX4D0 U698 ( .I0(\Storage[20][11] ), .I1(\Storage[21][11] ), .I2(
        \Storage[22][11] ), .I3(\Storage[23][11] ), .S0(n586), .S1(n534), .Z(
        n228) );
  MUX4D0 U699 ( .I0(\Storage[20][12] ), .I1(\Storage[21][12] ), .I2(
        \Storage[22][12] ), .I3(\Storage[23][12] ), .S0(n587), .S1(n534), .Z(
        n241) );
  MUX4D0 U700 ( .I0(\Storage[20][13] ), .I1(\Storage[21][13] ), .I2(
        \Storage[22][13] ), .I3(\Storage[23][13] ), .S0(n587), .S1(n556), .Z(
        n254) );
  MUX4D0 U701 ( .I0(\Storage[20][14] ), .I1(\Storage[21][14] ), .I2(
        \Storage[22][14] ), .I3(\Storage[23][14] ), .S0(n588), .S1(n556), .Z(
        n267) );
  MUX4D0 U702 ( .I0(\Storage[20][15] ), .I1(\Storage[21][15] ), .I2(
        \Storage[22][15] ), .I3(\Storage[23][15] ), .S0(n589), .S1(n557), .Z(
        n280) );
  MUX4D0 U703 ( .I0(\Storage[20][16] ), .I1(\Storage[21][16] ), .I2(
        \Storage[22][16] ), .I3(\Storage[23][16] ), .S0(n589), .S1(n557), .Z(
        n293) );
  MUX4D0 U704 ( .I0(\Storage[20][17] ), .I1(\Storage[21][17] ), .I2(
        \Storage[22][17] ), .I3(\Storage[23][17] ), .S0(n590), .S1(n557), .Z(
        n306) );
  MUX4D0 U705 ( .I0(\Storage[20][18] ), .I1(\Storage[21][18] ), .I2(
        \Storage[22][18] ), .I3(\Storage[23][18] ), .S0(n590), .S1(n537), .Z(
        n319) );
  MUX4D0 U706 ( .I0(\Storage[20][19] ), .I1(\Storage[21][19] ), .I2(
        \Storage[22][19] ), .I3(\Storage[23][19] ), .S0(n591), .S1(n536), .Z(
        n332) );
  MUX4D0 U707 ( .I0(\Storage[20][20] ), .I1(\Storage[21][20] ), .I2(
        \Storage[22][20] ), .I3(\Storage[23][20] ), .S0(n592), .S1(n963), .Z(
        n345) );
  MUX4D0 U708 ( .I0(\Storage[20][21] ), .I1(\Storage[21][21] ), .I2(
        \Storage[22][21] ), .I3(\Storage[23][21] ), .S0(n592), .S1(N45), .Z(
        n358) );
  MUX4D0 U709 ( .I0(\Storage[20][22] ), .I1(\Storage[21][22] ), .I2(
        \Storage[22][22] ), .I3(\Storage[23][22] ), .S0(n593), .S1(n543), .Z(
        n371) );
  MUX4D0 U710 ( .I0(\Storage[20][23] ), .I1(\Storage[21][23] ), .I2(
        \Storage[22][23] ), .I3(\Storage[23][23] ), .S0(n593), .S1(n539), .Z(
        n384) );
  MUX4D0 U711 ( .I0(\Storage[20][24] ), .I1(\Storage[21][24] ), .I2(
        \Storage[22][24] ), .I3(\Storage[23][24] ), .S0(n594), .S1(n539), .Z(
        n397) );
  MUX4D0 U712 ( .I0(\Storage[20][25] ), .I1(\Storage[21][25] ), .I2(
        \Storage[22][25] ), .I3(\Storage[23][25] ), .S0(n579), .S1(n546), .Z(
        n410) );
  MUX4D0 U713 ( .I0(\Storage[20][26] ), .I1(\Storage[21][26] ), .I2(
        \Storage[22][26] ), .I3(\Storage[23][26] ), .S0(n579), .S1(n546), .Z(
        n423) );
  MUX4D0 U714 ( .I0(\Storage[20][27] ), .I1(\Storage[21][27] ), .I2(
        \Storage[22][27] ), .I3(\Storage[23][27] ), .S0(n578), .S1(n547), .Z(
        n436) );
  MUX4D0 U715 ( .I0(\Storage[20][28] ), .I1(\Storage[21][28] ), .I2(
        \Storage[22][28] ), .I3(\Storage[23][28] ), .S0(n578), .S1(n548), .Z(
        n449) );
  MUX4D0 U716 ( .I0(\Storage[20][29] ), .I1(\Storage[21][29] ), .I2(
        \Storage[22][29] ), .I3(\Storage[23][29] ), .S0(n577), .S1(n548), .Z(
        n462) );
  MUX4D0 U717 ( .I0(\Storage[20][30] ), .I1(\Storage[21][30] ), .I2(
        \Storage[22][30] ), .I3(\Storage[23][30] ), .S0(n564), .S1(n549), .Z(
        n475) );
  MUX4D0 U718 ( .I0(\Storage[20][31] ), .I1(\Storage[21][31] ), .I2(
        \Storage[22][31] ), .I3(\Storage[23][31] ), .S0(n572), .S1(n549), .Z(
        n488) );
  MUX4D0 U719 ( .I0(\Storage[12][32] ), .I1(\Storage[13][32] ), .I2(
        \Storage[14][32] ), .I3(\Storage[15][32] ), .S0(n576), .S1(n550), .Z(
        n503) );
  MUX4D0 U720 ( .I0(\Storage[4][32] ), .I1(\Storage[5][32] ), .I2(
        \Storage[6][32] ), .I3(\Storage[7][32] ), .S0(n576), .S1(n550), .Z(
        n505) );
  MUX4D0 U721 ( .I0(\Storage[12][0] ), .I1(\Storage[13][0] ), .I2(
        \Storage[14][0] ), .I3(\Storage[15][0] ), .S0(n580), .S1(n551), .Z(n45) );
  MUX4D0 U722 ( .I0(\Storage[4][0] ), .I1(\Storage[5][0] ), .I2(
        \Storage[6][0] ), .I3(\Storage[7][0] ), .S0(n580), .S1(n551), .Z(n47)
         );
  MUX4D0 U723 ( .I0(\Storage[12][1] ), .I1(\Storage[13][1] ), .I2(
        \Storage[14][1] ), .I3(\Storage[15][1] ), .S0(n580), .S1(n551), .Z(n58) );
  MUX4D0 U724 ( .I0(\Storage[4][1] ), .I1(\Storage[5][1] ), .I2(
        \Storage[6][1] ), .I3(\Storage[7][1] ), .S0(n581), .S1(n552), .Z(n60)
         );
  MUX4D0 U725 ( .I0(\Storage[12][2] ), .I1(\Storage[13][2] ), .I2(
        \Storage[14][2] ), .I3(\Storage[15][2] ), .S0(n581), .S1(n552), .Z(
        n113) );
  MUX4D0 U726 ( .I0(\Storage[4][2] ), .I1(\Storage[5][2] ), .I2(
        \Storage[6][2] ), .I3(\Storage[7][2] ), .S0(n581), .S1(n552), .Z(n115)
         );
  MUX4D0 U727 ( .I0(\Storage[12][4] ), .I1(\Storage[13][4] ), .I2(
        \Storage[14][4] ), .I3(\Storage[15][4] ), .S0(n582), .S1(n553), .Z(
        n139) );
  MUX4D0 U728 ( .I0(\Storage[4][4] ), .I1(\Storage[5][4] ), .I2(
        \Storage[6][4] ), .I3(\Storage[7][4] ), .S0(n582), .S1(n553), .Z(n141)
         );
  MUX4D0 U729 ( .I0(\Storage[12][5] ), .I1(\Storage[13][5] ), .I2(
        \Storage[14][5] ), .I3(\Storage[15][5] ), .S0(n583), .S1(n554), .Z(
        n152) );
  MUX4D0 U730 ( .I0(\Storage[4][5] ), .I1(\Storage[5][5] ), .I2(
        \Storage[6][5] ), .I3(\Storage[7][5] ), .S0(n583), .S1(n554), .Z(n154)
         );
  MUX4D0 U731 ( .I0(\Storage[12][6] ), .I1(\Storage[13][6] ), .I2(
        \Storage[14][6] ), .I3(\Storage[15][6] ), .S0(n583), .S1(n554), .Z(
        n165) );
  MUX4D0 U732 ( .I0(\Storage[4][6] ), .I1(\Storage[5][6] ), .I2(
        \Storage[6][6] ), .I3(\Storage[7][6] ), .S0(n584), .S1(n555), .Z(n167)
         );
  MUX4D0 U733 ( .I0(\Storage[12][7] ), .I1(\Storage[13][7] ), .I2(
        \Storage[14][7] ), .I3(\Storage[15][7] ), .S0(n584), .S1(n555), .Z(
        n178) );
  MUX4D0 U734 ( .I0(\Storage[4][7] ), .I1(\Storage[5][7] ), .I2(
        \Storage[6][7] ), .I3(\Storage[7][7] ), .S0(n584), .S1(n555), .Z(n180)
         );
  MUX4D0 U735 ( .I0(\Storage[12][9] ), .I1(\Storage[13][9] ), .I2(
        \Storage[14][9] ), .I3(\Storage[15][9] ), .S0(n585), .S1(n546), .Z(
        n204) );
  MUX4D0 U736 ( .I0(\Storage[4][9] ), .I1(\Storage[5][9] ), .I2(
        \Storage[6][9] ), .I3(\Storage[7][9] ), .S0(n585), .S1(n537), .Z(n206)
         );
  MUX4D0 U737 ( .I0(\Storage[12][10] ), .I1(\Storage[13][10] ), .I2(
        \Storage[14][10] ), .I3(\Storage[15][10] ), .S0(n586), .S1(n963), .Z(
        n217) );
  MUX4D0 U738 ( .I0(\Storage[4][10] ), .I1(\Storage[5][10] ), .I2(
        \Storage[6][10] ), .I3(\Storage[7][10] ), .S0(n586), .S1(n535), .Z(
        n219) );
  MUX4D0 U739 ( .I0(\Storage[12][11] ), .I1(\Storage[13][11] ), .I2(
        \Storage[14][11] ), .I3(\Storage[15][11] ), .S0(n586), .S1(n535), .Z(
        n230) );
  MUX4D0 U740 ( .I0(\Storage[4][11] ), .I1(\Storage[5][11] ), .I2(
        \Storage[6][11] ), .I3(\Storage[7][11] ), .S0(n587), .S1(n540), .Z(
        n232) );
  MUX4D0 U741 ( .I0(\Storage[12][12] ), .I1(\Storage[13][12] ), .I2(
        \Storage[14][12] ), .I3(\Storage[15][12] ), .S0(n587), .S1(n542), .Z(
        n243) );
  MUX4D0 U742 ( .I0(\Storage[4][12] ), .I1(\Storage[5][12] ), .I2(
        \Storage[6][12] ), .I3(\Storage[7][12] ), .S0(n587), .S1(n537), .Z(
        n245) );
  MUX4D0 U743 ( .I0(\Storage[12][13] ), .I1(\Storage[13][13] ), .I2(
        \Storage[14][13] ), .I3(\Storage[15][13] ), .S0(n588), .S1(n541), .Z(
        n256) );
  MUX4D0 U744 ( .I0(\Storage[4][13] ), .I1(\Storage[5][13] ), .I2(
        \Storage[6][13] ), .I3(\Storage[7][13] ), .S0(n588), .S1(n557), .Z(
        n258) );
  MUX4D0 U745 ( .I0(\Storage[12][14] ), .I1(\Storage[13][14] ), .I2(
        \Storage[14][14] ), .I3(\Storage[15][14] ), .S0(n588), .S1(n556), .Z(
        n269) );
  MUX4D0 U746 ( .I0(\Storage[4][14] ), .I1(\Storage[5][14] ), .I2(
        \Storage[6][14] ), .I3(\Storage[7][14] ), .S0(n588), .S1(n556), .Z(
        n271) );
  MUX4D0 U747 ( .I0(\Storage[12][15] ), .I1(\Storage[13][15] ), .I2(
        \Storage[14][15] ), .I3(\Storage[15][15] ), .S0(n589), .S1(n557), .Z(
        n282) );
  MUX4D0 U748 ( .I0(\Storage[4][15] ), .I1(\Storage[5][15] ), .I2(
        \Storage[6][15] ), .I3(\Storage[7][15] ), .S0(n589), .S1(n557), .Z(
        n284) );
  MUX4D0 U749 ( .I0(\Storage[12][16] ), .I1(\Storage[13][16] ), .I2(
        \Storage[14][16] ), .I3(\Storage[15][16] ), .S0(n589), .S1(n558), .Z(
        n295) );
  MUX4D0 U750 ( .I0(\Storage[4][16] ), .I1(\Storage[5][16] ), .I2(
        \Storage[6][16] ), .I3(\Storage[7][16] ), .S0(n590), .S1(n558), .Z(
        n297) );
  MUX4D0 U751 ( .I0(\Storage[12][17] ), .I1(\Storage[13][17] ), .I2(
        \Storage[14][17] ), .I3(\Storage[15][17] ), .S0(n590), .S1(n557), .Z(
        n308) );
  MUX4D0 U752 ( .I0(\Storage[4][17] ), .I1(\Storage[5][17] ), .I2(
        \Storage[6][17] ), .I3(\Storage[7][17] ), .S0(n590), .S1(n538), .Z(
        n310) );
  MUX4D0 U753 ( .I0(\Storage[12][18] ), .I1(\Storage[13][18] ), .I2(
        \Storage[14][18] ), .I3(\Storage[15][18] ), .S0(n591), .S1(n963), .Z(
        n321) );
  MUX4D0 U754 ( .I0(\Storage[4][18] ), .I1(\Storage[5][18] ), .I2(
        \Storage[6][18] ), .I3(\Storage[7][18] ), .S0(n591), .S1(n537), .Z(
        n323) );
  MUX4D0 U755 ( .I0(\Storage[12][19] ), .I1(\Storage[13][19] ), .I2(
        \Storage[14][19] ), .I3(\Storage[15][19] ), .S0(n591), .S1(n542), .Z(
        n334) );
  MUX4D0 U756 ( .I0(\Storage[4][19] ), .I1(\Storage[5][19] ), .I2(
        \Storage[6][19] ), .I3(\Storage[7][19] ), .S0(n591), .S1(n540), .Z(
        n336) );
  MUX4D0 U757 ( .I0(\Storage[12][20] ), .I1(\Storage[13][20] ), .I2(
        \Storage[14][20] ), .I3(\Storage[15][20] ), .S0(n592), .S1(n536), .Z(
        n347) );
  MUX4D0 U758 ( .I0(\Storage[4][20] ), .I1(\Storage[5][20] ), .I2(
        \Storage[6][20] ), .I3(\Storage[7][20] ), .S0(n592), .S1(n540), .Z(
        n349) );
  MUX4D0 U759 ( .I0(\Storage[12][21] ), .I1(\Storage[13][21] ), .I2(
        \Storage[14][21] ), .I3(\Storage[15][21] ), .S0(n592), .S1(n539), .Z(
        n360) );
  MUX4D0 U760 ( .I0(\Storage[4][21] ), .I1(\Storage[5][21] ), .I2(
        \Storage[6][21] ), .I3(\Storage[7][21] ), .S0(n593), .S1(n539), .Z(
        n362) );
  MUX4D0 U761 ( .I0(\Storage[12][22] ), .I1(\Storage[13][22] ), .I2(
        \Storage[14][22] ), .I3(\Storage[15][22] ), .S0(n593), .S1(n543), .Z(
        n373) );
  MUX4D0 U762 ( .I0(\Storage[4][22] ), .I1(\Storage[5][22] ), .I2(
        \Storage[6][22] ), .I3(\Storage[7][22] ), .S0(n593), .S1(n536), .Z(
        n375) );
  MUX4D0 U763 ( .I0(\Storage[12][23] ), .I1(\Storage[13][23] ), .I2(
        \Storage[14][23] ), .I3(\Storage[15][23] ), .S0(n594), .S1(n539), .Z(
        n386) );
  MUX4D0 U764 ( .I0(\Storage[4][23] ), .I1(\Storage[5][23] ), .I2(
        \Storage[6][23] ), .I3(\Storage[7][23] ), .S0(n594), .S1(n539), .Z(
        n388) );
  MUX4D0 U765 ( .I0(\Storage[12][24] ), .I1(\Storage[13][24] ), .I2(
        \Storage[14][24] ), .I3(\Storage[15][24] ), .S0(n594), .S1(n539), .Z(
        n399) );
  MUX4D0 U766 ( .I0(\Storage[4][24] ), .I1(\Storage[5][24] ), .I2(
        \Storage[6][24] ), .I3(\Storage[7][24] ), .S0(n580), .S1(n546), .Z(
        n401) );
  MUX4D0 U767 ( .I0(\Storage[12][25] ), .I1(\Storage[13][25] ), .I2(
        \Storage[14][25] ), .I3(\Storage[15][25] ), .S0(n579), .S1(n546), .Z(
        n412) );
  MUX4D0 U768 ( .I0(\Storage[4][25] ), .I1(\Storage[5][25] ), .I2(
        \Storage[6][25] ), .I3(\Storage[7][25] ), .S0(n579), .S1(n546), .Z(
        n414) );
  MUX4D0 U769 ( .I0(\Storage[12][26] ), .I1(\Storage[13][26] ), .I2(
        \Storage[14][26] ), .I3(\Storage[15][26] ), .S0(n579), .S1(n547), .Z(
        n425) );
  MUX4D0 U770 ( .I0(\Storage[4][26] ), .I1(\Storage[5][26] ), .I2(
        \Storage[6][26] ), .I3(\Storage[7][26] ), .S0(n578), .S1(n547), .Z(
        n427) );
  MUX4D0 U771 ( .I0(\Storage[12][27] ), .I1(\Storage[13][27] ), .I2(
        \Storage[14][27] ), .I3(\Storage[15][27] ), .S0(n578), .S1(n547), .Z(
        n438) );
  MUX4D0 U772 ( .I0(\Storage[4][27] ), .I1(\Storage[5][27] ), .I2(
        \Storage[6][27] ), .I3(\Storage[7][27] ), .S0(n578), .S1(n547), .Z(
        n440) );
  MUX4D0 U773 ( .I0(\Storage[12][28] ), .I1(\Storage[13][28] ), .I2(
        \Storage[14][28] ), .I3(\Storage[15][28] ), .S0(n577), .S1(n548), .Z(
        n451) );
  MUX4D0 U774 ( .I0(\Storage[4][28] ), .I1(\Storage[5][28] ), .I2(
        \Storage[6][28] ), .I3(\Storage[7][28] ), .S0(n577), .S1(n548), .Z(
        n453) );
  MUX4D0 U775 ( .I0(\Storage[12][29] ), .I1(\Storage[13][29] ), .I2(
        \Storage[14][29] ), .I3(\Storage[15][29] ), .S0(n577), .S1(n548), .Z(
        n464) );
  MUX4D0 U776 ( .I0(\Storage[4][29] ), .I1(\Storage[5][29] ), .I2(
        \Storage[6][29] ), .I3(\Storage[7][29] ), .S0(n577), .S1(n549), .Z(
        n466) );
  MUX4D0 U777 ( .I0(\Storage[12][30] ), .I1(\Storage[13][30] ), .I2(
        \Storage[14][30] ), .I3(\Storage[15][30] ), .S0(n572), .S1(n549), .Z(
        n477) );
  MUX4D0 U778 ( .I0(\Storage[4][30] ), .I1(\Storage[5][30] ), .I2(
        \Storage[6][30] ), .I3(\Storage[7][30] ), .S0(n564), .S1(n549), .Z(
        n479) );
  MUX4D0 U779 ( .I0(\Storage[12][31] ), .I1(\Storage[13][31] ), .I2(
        \Storage[14][31] ), .I3(\Storage[15][31] ), .S0(n564), .S1(n550), .Z(
        n490) );
  MUX4D0 U780 ( .I0(\Storage[4][31] ), .I1(\Storage[5][31] ), .I2(
        \Storage[6][31] ), .I3(\Storage[7][31] ), .S0(n576), .S1(n550), .Z(
        n492) );
  MUX4D0 U781 ( .I0(\Storage[16][32] ), .I1(\Storage[17][32] ), .I2(
        \Storage[18][32] ), .I3(\Storage[19][32] ), .S0(n576), .S1(n550), .Z(
        n502) );
  MUX4D0 U782 ( .I0(\Storage[16][0] ), .I1(\Storage[17][0] ), .I2(
        \Storage[18][0] ), .I3(\Storage[19][0] ), .S0(n594), .S1(n551), .Z(n44) );
  MUX4D0 U783 ( .I0(\Storage[16][1] ), .I1(\Storage[17][1] ), .I2(
        \Storage[18][1] ), .I3(\Storage[19][1] ), .S0(n580), .S1(n551), .Z(n57) );
  MUX4D0 U784 ( .I0(\Storage[16][2] ), .I1(\Storage[17][2] ), .I2(
        \Storage[18][2] ), .I3(\Storage[19][2] ), .S0(n581), .S1(n552), .Z(
        n112) );
  MUX4D0 U785 ( .I0(\Storage[16][4] ), .I1(\Storage[17][4] ), .I2(
        \Storage[18][4] ), .I3(\Storage[19][4] ), .S0(n582), .S1(n553), .Z(
        n138) );
  MUX4D0 U786 ( .I0(\Storage[16][5] ), .I1(\Storage[17][5] ), .I2(
        \Storage[18][5] ), .I3(\Storage[19][5] ), .S0(n583), .S1(n554), .Z(
        n151) );
  MUX4D0 U787 ( .I0(\Storage[16][6] ), .I1(\Storage[17][6] ), .I2(
        \Storage[18][6] ), .I3(\Storage[19][6] ), .S0(n583), .S1(n554), .Z(
        n164) );
  MUX4D0 U788 ( .I0(\Storage[16][7] ), .I1(\Storage[17][7] ), .I2(
        \Storage[18][7] ), .I3(\Storage[19][7] ), .S0(n584), .S1(n555), .Z(
        n177) );
  MUX4D0 U789 ( .I0(\Storage[16][9] ), .I1(\Storage[17][9] ), .I2(
        \Storage[18][9] ), .I3(\Storage[19][9] ), .S0(n585), .S1(n542), .Z(
        n203) );
  MUX4D0 U790 ( .I0(\Storage[16][10] ), .I1(\Storage[17][10] ), .I2(
        \Storage[18][10] ), .I3(\Storage[19][10] ), .S0(n586), .S1(n534), .Z(
        n216) );
  MUX4D0 U791 ( .I0(\Storage[16][11] ), .I1(\Storage[17][11] ), .I2(
        \Storage[18][11] ), .I3(\Storage[19][11] ), .S0(n586), .S1(n542), .Z(
        n229) );
  MUX4D0 U792 ( .I0(\Storage[16][12] ), .I1(\Storage[17][12] ), .I2(
        \Storage[18][12] ), .I3(\Storage[19][12] ), .S0(n587), .S1(n534), .Z(
        n242) );
  MUX4D0 U793 ( .I0(\Storage[16][13] ), .I1(\Storage[17][13] ), .I2(
        \Storage[18][13] ), .I3(\Storage[19][13] ), .S0(n588), .S1(n556), .Z(
        n255) );
  MUX4D0 U794 ( .I0(\Storage[16][14] ), .I1(\Storage[17][14] ), .I2(
        \Storage[18][14] ), .I3(\Storage[19][14] ), .S0(n588), .S1(n537), .Z(
        n268) );
  MUX4D0 U795 ( .I0(\Storage[16][15] ), .I1(\Storage[17][15] ), .I2(
        \Storage[18][15] ), .I3(\Storage[19][15] ), .S0(n589), .S1(n556), .Z(
        n281) );
  MUX4D0 U796 ( .I0(\Storage[16][16] ), .I1(\Storage[17][16] ), .I2(
        \Storage[18][16] ), .I3(\Storage[19][16] ), .S0(n589), .S1(n558), .Z(
        n294) );
  MUX4D0 U797 ( .I0(\Storage[16][17] ), .I1(\Storage[17][17] ), .I2(
        \Storage[18][17] ), .I3(\Storage[19][17] ), .S0(n590), .S1(n558), .Z(
        n307) );
  MUX4D0 U798 ( .I0(\Storage[16][18] ), .I1(\Storage[17][18] ), .I2(
        \Storage[18][18] ), .I3(\Storage[19][18] ), .S0(n591), .S1(N45), .Z(
        n320) );
  MUX4D0 U799 ( .I0(\Storage[16][19] ), .I1(\Storage[17][19] ), .I2(
        \Storage[18][19] ), .I3(\Storage[19][19] ), .S0(n591), .S1(n963), .Z(
        n333) );
  MUX4D0 U800 ( .I0(\Storage[16][20] ), .I1(\Storage[17][20] ), .I2(
        \Storage[18][20] ), .I3(\Storage[19][20] ), .S0(n592), .S1(n535), .Z(
        n346) );
  MUX4D0 U801 ( .I0(\Storage[16][21] ), .I1(\Storage[17][21] ), .I2(
        \Storage[18][21] ), .I3(\Storage[19][21] ), .S0(n592), .S1(n540), .Z(
        n359) );
  MUX4D0 U802 ( .I0(\Storage[16][22] ), .I1(\Storage[17][22] ), .I2(
        \Storage[18][22] ), .I3(\Storage[19][22] ), .S0(n593), .S1(n542), .Z(
        n372) );
  MUX4D0 U803 ( .I0(\Storage[16][23] ), .I1(\Storage[17][23] ), .I2(
        \Storage[18][23] ), .I3(\Storage[19][23] ), .S0(n594), .S1(n538), .Z(
        n385) );
  MUX4D0 U804 ( .I0(\Storage[16][24] ), .I1(\Storage[17][24] ), .I2(
        \Storage[18][24] ), .I3(\Storage[19][24] ), .S0(n594), .S1(n538), .Z(
        n398) );
  MUX4D0 U805 ( .I0(\Storage[16][25] ), .I1(\Storage[17][25] ), .I2(
        \Storage[18][25] ), .I3(\Storage[19][25] ), .S0(n579), .S1(n546), .Z(
        n411) );
  MUX4D0 U806 ( .I0(\Storage[16][26] ), .I1(\Storage[17][26] ), .I2(
        \Storage[18][26] ), .I3(\Storage[19][26] ), .S0(n579), .S1(n547), .Z(
        n424) );
  MUX4D0 U807 ( .I0(\Storage[16][27] ), .I1(\Storage[17][27] ), .I2(
        \Storage[18][27] ), .I3(\Storage[19][27] ), .S0(n578), .S1(n547), .Z(
        n437) );
  MUX4D0 U808 ( .I0(\Storage[16][28] ), .I1(\Storage[17][28] ), .I2(
        \Storage[18][28] ), .I3(\Storage[19][28] ), .S0(n578), .S1(n548), .Z(
        n450) );
  MUX4D0 U809 ( .I0(\Storage[16][29] ), .I1(\Storage[17][29] ), .I2(
        \Storage[18][29] ), .I3(\Storage[19][29] ), .S0(n577), .S1(n548), .Z(
        n463) );
  MUX4D0 U810 ( .I0(\Storage[16][30] ), .I1(\Storage[17][30] ), .I2(
        \Storage[18][30] ), .I3(\Storage[19][30] ), .S0(n572), .S1(n549), .Z(
        n476) );
  MUX4D0 U811 ( .I0(\Storage[16][31] ), .I1(\Storage[17][31] ), .I2(
        \Storage[18][31] ), .I3(\Storage[19][31] ), .S0(n564), .S1(n550), .Z(
        n489) );
  MUX4D0 U812 ( .I0(\Storage[8][32] ), .I1(\Storage[9][32] ), .I2(
        \Storage[10][32] ), .I3(\Storage[11][32] ), .S0(n576), .S1(n550), .Z(
        n504) );
  MUX4D0 U813 ( .I0(\Storage[0][32] ), .I1(\Storage[1][32] ), .I2(
        \Storage[2][32] ), .I3(\Storage[3][32] ), .S0(n576), .S1(n551), .Z(
        n506) );
  MUX4D0 U814 ( .I0(\Storage[8][0] ), .I1(\Storage[9][0] ), .I2(
        \Storage[10][0] ), .I3(\Storage[11][0] ), .S0(n580), .S1(n551), .Z(n46) );
  MUX4D0 U815 ( .I0(\Storage[0][0] ), .I1(\Storage[1][0] ), .I2(
        \Storage[2][0] ), .I3(\Storage[3][0] ), .S0(n580), .S1(n551), .Z(n48)
         );
  MUX4D0 U816 ( .I0(\Storage[8][1] ), .I1(\Storage[9][1] ), .I2(
        \Storage[10][1] ), .I3(\Storage[11][1] ), .S0(n580), .S1(n551), .Z(n59) );
  MUX4D0 U817 ( .I0(\Storage[0][1] ), .I1(\Storage[1][1] ), .I2(
        \Storage[2][1] ), .I3(\Storage[3][1] ), .S0(n581), .S1(n552), .Z(n61)
         );
  MUX4D0 U818 ( .I0(\Storage[8][2] ), .I1(\Storage[9][2] ), .I2(
        \Storage[10][2] ), .I3(\Storage[11][2] ), .S0(n581), .S1(n552), .Z(
        n114) );
  MUX4D0 U819 ( .I0(\Storage[0][2] ), .I1(\Storage[1][2] ), .I2(
        \Storage[2][2] ), .I3(\Storage[3][2] ), .S0(n581), .S1(n552), .Z(n116)
         );
  MUX4D0 U820 ( .I0(\Storage[8][4] ), .I1(\Storage[9][4] ), .I2(
        \Storage[10][4] ), .I3(\Storage[11][4] ), .S0(n582), .S1(n553), .Z(
        n140) );
  MUX4D0 U821 ( .I0(\Storage[0][4] ), .I1(\Storage[1][4] ), .I2(
        \Storage[2][4] ), .I3(\Storage[3][4] ), .S0(n582), .S1(n553), .Z(n142)
         );
  MUX4D0 U822 ( .I0(\Storage[8][5] ), .I1(\Storage[9][5] ), .I2(
        \Storage[10][5] ), .I3(\Storage[11][5] ), .S0(n583), .S1(n554), .Z(
        n153) );
  MUX4D0 U823 ( .I0(\Storage[0][5] ), .I1(\Storage[1][5] ), .I2(
        \Storage[2][5] ), .I3(\Storage[3][5] ), .S0(n583), .S1(n554), .Z(n155)
         );
  MUX4D0 U824 ( .I0(\Storage[8][6] ), .I1(\Storage[9][6] ), .I2(
        \Storage[10][6] ), .I3(\Storage[11][6] ), .S0(n583), .S1(n554), .Z(
        n166) );
  MUX4D0 U825 ( .I0(\Storage[0][6] ), .I1(\Storage[1][6] ), .I2(
        \Storage[2][6] ), .I3(\Storage[3][6] ), .S0(n584), .S1(n555), .Z(n168)
         );
  MUX4D0 U826 ( .I0(\Storage[8][7] ), .I1(\Storage[9][7] ), .I2(
        \Storage[10][7] ), .I3(\Storage[11][7] ), .S0(n584), .S1(n555), .Z(
        n179) );
  MUX4D0 U827 ( .I0(\Storage[0][7] ), .I1(\Storage[1][7] ), .I2(
        \Storage[2][7] ), .I3(\Storage[3][7] ), .S0(n584), .S1(n555), .Z(n181)
         );
  MUX4D0 U828 ( .I0(\Storage[8][9] ), .I1(\Storage[9][9] ), .I2(
        \Storage[10][9] ), .I3(\Storage[11][9] ), .S0(n585), .S1(n541), .Z(
        n205) );
  MUX4D0 U829 ( .I0(\Storage[0][9] ), .I1(\Storage[1][9] ), .I2(
        \Storage[2][9] ), .I3(\Storage[3][9] ), .S0(n585), .S1(n536), .Z(n207)
         );
  MUX4D0 U830 ( .I0(\Storage[8][10] ), .I1(\Storage[9][10] ), .I2(
        \Storage[10][10] ), .I3(\Storage[11][10] ), .S0(n586), .S1(n963), .Z(
        n218) );
  MUX4D0 U831 ( .I0(\Storage[0][10] ), .I1(\Storage[1][10] ), .I2(
        \Storage[2][10] ), .I3(\Storage[3][10] ), .S0(n586), .S1(n536), .Z(
        n220) );
  MUX4D0 U832 ( .I0(\Storage[8][11] ), .I1(\Storage[9][11] ), .I2(
        \Storage[10][11] ), .I3(\Storage[11][11] ), .S0(n586), .S1(n541), .Z(
        n231) );
  MUX4D0 U833 ( .I0(\Storage[0][11] ), .I1(\Storage[1][11] ), .I2(
        \Storage[2][11] ), .I3(\Storage[3][11] ), .S0(n587), .S1(n536), .Z(
        n233) );
  MUX4D0 U834 ( .I0(\Storage[8][12] ), .I1(\Storage[9][12] ), .I2(
        \Storage[10][12] ), .I3(\Storage[11][12] ), .S0(n587), .S1(n535), .Z(
        n244) );
  MUX4D0 U835 ( .I0(\Storage[0][12] ), .I1(\Storage[1][12] ), .I2(
        \Storage[2][12] ), .I3(\Storage[3][12] ), .S0(n587), .S1(n556), .Z(
        n246) );
  MUX4D0 U836 ( .I0(\Storage[8][13] ), .I1(\Storage[9][13] ), .I2(
        \Storage[10][13] ), .I3(\Storage[11][13] ), .S0(n588), .S1(n556), .Z(
        n257) );
  MUX4D0 U837 ( .I0(\Storage[0][13] ), .I1(\Storage[1][13] ), .I2(
        \Storage[2][13] ), .I3(\Storage[3][13] ), .S0(n588), .S1(n556), .Z(
        n259) );
  MUX4D0 U838 ( .I0(\Storage[8][14] ), .I1(\Storage[9][14] ), .I2(
        \Storage[10][14] ), .I3(\Storage[11][14] ), .S0(n588), .S1(n557), .Z(
        n270) );
  MUX4D0 U839 ( .I0(\Storage[0][14] ), .I1(\Storage[1][14] ), .I2(
        \Storage[2][14] ), .I3(\Storage[3][14] ), .S0(n589), .S1(n557), .Z(
        n272) );
  MUX4D0 U840 ( .I0(\Storage[8][15] ), .I1(\Storage[9][15] ), .I2(
        \Storage[10][15] ), .I3(\Storage[11][15] ), .S0(n589), .S1(n557), .Z(
        n283) );
  MUX4D0 U841 ( .I0(\Storage[0][15] ), .I1(\Storage[1][15] ), .I2(
        \Storage[2][15] ), .I3(\Storage[3][15] ), .S0(n589), .S1(n558), .Z(
        n285) );
  MUX4D0 U842 ( .I0(\Storage[8][16] ), .I1(\Storage[9][16] ), .I2(
        \Storage[10][16] ), .I3(\Storage[11][16] ), .S0(n590), .S1(n556), .Z(
        n296) );
  MUX4D0 U843 ( .I0(\Storage[0][16] ), .I1(\Storage[1][16] ), .I2(
        \Storage[2][16] ), .I3(\Storage[3][16] ), .S0(n590), .S1(n558), .Z(
        n298) );
  MUX4D0 U844 ( .I0(\Storage[8][17] ), .I1(\Storage[9][17] ), .I2(
        \Storage[10][17] ), .I3(\Storage[11][17] ), .S0(n590), .S1(n538), .Z(
        n309) );
  MUX4D0 U845 ( .I0(\Storage[0][17] ), .I1(\Storage[1][17] ), .I2(
        \Storage[2][17] ), .I3(\Storage[3][17] ), .S0(n590), .S1(n963), .Z(
        n311) );
  MUX4D0 U846 ( .I0(\Storage[8][18] ), .I1(\Storage[9][18] ), .I2(
        \Storage[10][18] ), .I3(\Storage[11][18] ), .S0(n591), .S1(n541), .Z(
        n322) );
  MUX4D0 U847 ( .I0(\Storage[0][18] ), .I1(\Storage[1][18] ), .I2(
        \Storage[2][18] ), .I3(\Storage[3][18] ), .S0(n591), .S1(n540), .Z(
        n324) );
  MUX4D0 U848 ( .I0(\Storage[8][19] ), .I1(\Storage[9][19] ), .I2(
        \Storage[10][19] ), .I3(\Storage[11][19] ), .S0(n591), .S1(n534), .Z(
        n335) );
  MUX4D0 U849 ( .I0(\Storage[0][19] ), .I1(\Storage[1][19] ), .I2(
        \Storage[2][19] ), .I3(\Storage[3][19] ), .S0(n592), .S1(n541), .Z(
        n337) );
  MUX4D0 U850 ( .I0(\Storage[8][20] ), .I1(\Storage[9][20] ), .I2(
        \Storage[10][20] ), .I3(\Storage[11][20] ), .S0(n592), .S1(n535), .Z(
        n348) );
  MUX4D0 U851 ( .I0(\Storage[0][20] ), .I1(\Storage[1][20] ), .I2(
        \Storage[2][20] ), .I3(\Storage[3][20] ), .S0(n592), .S1(n537), .Z(
        n350) );
  MUX4D0 U852 ( .I0(\Storage[8][21] ), .I1(\Storage[9][21] ), .I2(
        \Storage[10][21] ), .I3(\Storage[11][21] ), .S0(n593), .S1(n538), .Z(
        n361) );
  MUX4D0 U853 ( .I0(\Storage[0][21] ), .I1(\Storage[1][21] ), .I2(
        \Storage[2][21] ), .I3(\Storage[3][21] ), .S0(n593), .S1(n538), .Z(
        n363) );
  MUX4D0 U854 ( .I0(\Storage[8][22] ), .I1(\Storage[9][22] ), .I2(
        \Storage[10][22] ), .I3(\Storage[11][22] ), .S0(n593), .S1(n537), .Z(
        n374) );
  MUX4D0 U855 ( .I0(\Storage[0][22] ), .I1(\Storage[1][22] ), .I2(
        \Storage[2][22] ), .I3(\Storage[3][22] ), .S0(n593), .S1(n534), .Z(
        n376) );
  MUX4D0 U856 ( .I0(\Storage[8][23] ), .I1(\Storage[9][23] ), .I2(
        \Storage[10][23] ), .I3(\Storage[11][23] ), .S0(n594), .S1(n538), .Z(
        n387) );
  MUX4D0 U857 ( .I0(\Storage[0][23] ), .I1(\Storage[1][23] ), .I2(
        \Storage[2][23] ), .I3(\Storage[3][23] ), .S0(n594), .S1(n538), .Z(
        n389) );
  MUX4D0 U858 ( .I0(\Storage[8][24] ), .I1(\Storage[9][24] ), .I2(
        \Storage[10][24] ), .I3(\Storage[11][24] ), .S0(n594), .S1(n538), .Z(
        n400) );
  MUX4D0 U859 ( .I0(\Storage[0][24] ), .I1(\Storage[1][24] ), .I2(
        \Storage[2][24] ), .I3(\Storage[3][24] ), .S0(n580), .S1(n546), .Z(
        n402) );
  MUX4D0 U860 ( .I0(\Storage[8][25] ), .I1(\Storage[9][25] ), .I2(
        \Storage[10][25] ), .I3(\Storage[11][25] ), .S0(n579), .S1(n546), .Z(
        n413) );
  MUX4D0 U861 ( .I0(\Storage[0][25] ), .I1(\Storage[1][25] ), .I2(
        \Storage[2][25] ), .I3(\Storage[3][25] ), .S0(n579), .S1(n546), .Z(
        n415) );
  MUX4D0 U862 ( .I0(\Storage[8][26] ), .I1(\Storage[9][26] ), .I2(
        \Storage[10][26] ), .I3(\Storage[11][26] ), .S0(n579), .S1(n547), .Z(
        n426) );
  MUX4D0 U863 ( .I0(\Storage[0][26] ), .I1(\Storage[1][26] ), .I2(
        \Storage[2][26] ), .I3(\Storage[3][26] ), .S0(n578), .S1(n547), .Z(
        n428) );
  MUX4D0 U864 ( .I0(\Storage[8][27] ), .I1(\Storage[9][27] ), .I2(
        \Storage[10][27] ), .I3(\Storage[11][27] ), .S0(n578), .S1(n547), .Z(
        n439) );
  MUX4D0 U865 ( .I0(\Storage[0][27] ), .I1(\Storage[1][27] ), .I2(
        \Storage[2][27] ), .I3(\Storage[3][27] ), .S0(n578), .S1(n548), .Z(
        n441) );
  MUX4D0 U866 ( .I0(\Storage[8][28] ), .I1(\Storage[9][28] ), .I2(
        \Storage[10][28] ), .I3(\Storage[11][28] ), .S0(n577), .S1(n548), .Z(
        n452) );
  MUX4D0 U867 ( .I0(\Storage[0][28] ), .I1(\Storage[1][28] ), .I2(
        \Storage[2][28] ), .I3(\Storage[3][28] ), .S0(n577), .S1(n548), .Z(
        n454) );
  MUX4D0 U868 ( .I0(\Storage[8][29] ), .I1(\Storage[9][29] ), .I2(
        \Storage[10][29] ), .I3(\Storage[11][29] ), .S0(n577), .S1(n549), .Z(
        n465) );
  MUX4D0 U869 ( .I0(\Storage[0][29] ), .I1(\Storage[1][29] ), .I2(
        \Storage[2][29] ), .I3(\Storage[3][29] ), .S0(n577), .S1(n549), .Z(
        n467) );
  MUX4D0 U870 ( .I0(\Storage[8][30] ), .I1(\Storage[9][30] ), .I2(
        \Storage[10][30] ), .I3(\Storage[11][30] ), .S0(n564), .S1(n549), .Z(
        n478) );
  MUX4D0 U871 ( .I0(\Storage[0][30] ), .I1(\Storage[1][30] ), .I2(
        \Storage[2][30] ), .I3(\Storage[3][30] ), .S0(n564), .S1(n549), .Z(
        n480) );
  MUX4D0 U872 ( .I0(\Storage[8][31] ), .I1(\Storage[9][31] ), .I2(
        \Storage[10][31] ), .I3(\Storage[11][31] ), .S0(n572), .S1(n550), .Z(
        n491) );
  MUX4D0 U873 ( .I0(\Storage[0][31] ), .I1(\Storage[1][31] ), .I2(
        \Storage[2][31] ), .I3(\Storage[3][31] ), .S0(n576), .S1(n550), .Z(
        n493) );
  MUX4D0 U874 ( .I0(\Storage[20][3] ), .I1(\Storage[21][3] ), .I2(
        \Storage[22][3] ), .I3(\Storage[23][3] ), .S0(n581), .S1(n552), .Z(
        n124) );
  MUX4D0 U875 ( .I0(\Storage[20][8] ), .I1(\Storage[21][8] ), .I2(
        \Storage[22][8] ), .I3(\Storage[23][8] ), .S0(n584), .S1(n555), .Z(
        n189) );
  MUX4D0 U876 ( .I0(\Storage[12][3] ), .I1(\Storage[13][3] ), .I2(
        \Storage[14][3] ), .I3(\Storage[15][3] ), .S0(n582), .S1(n553), .Z(
        n126) );
  MUX4D0 U877 ( .I0(\Storage[4][3] ), .I1(\Storage[5][3] ), .I2(
        \Storage[6][3] ), .I3(\Storage[7][3] ), .S0(n582), .S1(n553), .Z(n128)
         );
  MUX4D0 U878 ( .I0(\Storage[12][8] ), .I1(\Storage[13][8] ), .I2(
        \Storage[14][8] ), .I3(\Storage[15][8] ), .S0(n585), .S1(n542), .Z(
        n191) );
  MUX4D0 U879 ( .I0(\Storage[4][8] ), .I1(\Storage[5][8] ), .I2(
        \Storage[6][8] ), .I3(\Storage[7][8] ), .S0(n585), .S1(n542), .Z(n193)
         );
  MUX4D0 U880 ( .I0(\Storage[16][3] ), .I1(\Storage[17][3] ), .I2(
        \Storage[18][3] ), .I3(\Storage[19][3] ), .S0(n581), .S1(n552), .Z(
        n125) );
  MUX4D0 U881 ( .I0(\Storage[16][8] ), .I1(\Storage[17][8] ), .I2(
        \Storage[18][8] ), .I3(\Storage[19][8] ), .S0(n584), .S1(n555), .Z(
        n190) );
  MUX4D0 U882 ( .I0(\Storage[8][3] ), .I1(\Storage[9][3] ), .I2(
        \Storage[10][3] ), .I3(\Storage[11][3] ), .S0(n582), .S1(n553), .Z(
        n127) );
  MUX4D0 U883 ( .I0(\Storage[0][3] ), .I1(\Storage[1][3] ), .I2(
        \Storage[2][3] ), .I3(\Storage[3][3] ), .S0(n582), .S1(n553), .Z(n129)
         );
  MUX4D0 U884 ( .I0(\Storage[8][8] ), .I1(\Storage[9][8] ), .I2(
        \Storage[10][8] ), .I3(\Storage[11][8] ), .S0(n585), .S1(n541), .Z(
        n192) );
  MUX4D0 U885 ( .I0(\Storage[0][8] ), .I1(\Storage[1][8] ), .I2(
        \Storage[2][8] ), .I3(\Storage[3][8] ), .S0(n585), .S1(n541), .Z(n194)
         );
  ND3D1 U886 ( .A1(n100), .A2(n102), .A3(Write), .ZN(n103) );
  ND3D1 U887 ( .A1(AddrW[3]), .A2(n102), .A3(Write), .ZN(n101) );
  ND3D1 U888 ( .A1(AddrW[4]), .A2(n100), .A3(Write), .ZN(n70) );
  ND3D1 U889 ( .A1(AddrW[4]), .A2(AddrW[3]), .A3(Write), .ZN(n66) );
  ND3D1 U890 ( .A1(AddrW[0]), .A2(n106), .A3(AddrW[2]), .ZN(n85) );
  ND3D1 U891 ( .A1(AddrW[0]), .A2(AddrW[1]), .A3(AddrW[2]), .ZN(n71) );
  ND3D1 U892 ( .A1(AddrW[1]), .A2(n105), .A3(AddrW[0]), .ZN(n99) );
  ND3D1 U893 ( .A1(n106), .A2(n105), .A3(AddrW[0]), .ZN(n68) );
  ND3D1 U894 ( .A1(n104), .A2(n106), .A3(AddrW[2]), .ZN(n98) );
  ND3D1 U895 ( .A1(AddrW[1]), .A2(n104), .A3(AddrW[2]), .ZN(n72) );
  CKAN2D0 U896 ( .A1(ClkW), .A2(ChipEna), .Z(ClockW) );
  INVD1 U897 ( .I(AddrW[0]), .ZN(n104) );
  INVD1 U898 ( .I(AddrW[2]), .ZN(n105) );
  INVD1 U899 ( .I(AddrW[3]), .ZN(n100) );
  INVD1 U900 ( .I(AddrW[4]), .ZN(n102) );
  AN2D1 U901 ( .A1(ClkR), .A2(ChipEna), .Z(ClockR) );
  MUX3ND0 U902 ( .I0(n40), .I1(n41), .I2(n42), .S0(n558), .S1(n523), .ZN(n39)
         );
  MUX3ND0 U903 ( .I0(n49), .I1(n50), .I2(n51), .S0(n964), .S1(n965), .ZN(N82)
         );
  MUX3ND0 U904 ( .I0(n53), .I1(n54), .I2(n55), .S0(n561), .S1(n523), .ZN(n52)
         );
  MUX3ND0 U905 ( .I0(n62), .I1(n63), .I2(n64), .S0(n515), .S1(n965), .ZN(N81)
         );
  MUX3ND0 U906 ( .I0(n108), .I1(n109), .I2(n110), .S0(n561), .S1(n519), .ZN(
        n65) );
  MUX3ND0 U907 ( .I0(n117), .I1(n118), .I2(n119), .S0(n964), .S1(n965), .ZN(
        N80) );
  MUX3ND0 U908 ( .I0(n121), .I1(n122), .I2(n123), .S0(n560), .S1(n533), .ZN(
        n120) );
  MUX3ND0 U909 ( .I0(n130), .I1(n131), .I2(n132), .S0(n515), .S1(n511), .ZN(
        N79) );
  MUX3ND0 U910 ( .I0(n134), .I1(n135), .I2(n136), .S0(n561), .S1(n533), .ZN(
        n133) );
  MUX3ND0 U911 ( .I0(n143), .I1(n144), .I2(n145), .S0(n964), .S1(n511), .ZN(
        N78) );
  MUX3ND0 U912 ( .I0(n147), .I1(n148), .I2(n149), .S0(n559), .S1(N46), .ZN(
        n146) );
  MUX3ND0 U913 ( .I0(n156), .I1(n157), .I2(n158), .S0(n515), .S1(n511), .ZN(
        N77) );
  MUX3ND0 U914 ( .I0(n160), .I1(n161), .I2(n162), .S0(n559), .S1(n521), .ZN(
        n159) );
  MUX3ND0 U915 ( .I0(n169), .I1(n170), .I2(n171), .S0(n515), .S1(n511), .ZN(
        N76) );
  MUX3ND0 U916 ( .I0(n173), .I1(n174), .I2(n175), .S0(n559), .S1(n522), .ZN(
        n172) );
  MUX3ND0 U917 ( .I0(n182), .I1(n183), .I2(n184), .S0(n513), .S1(n511), .ZN(
        N75) );
  MUX3ND0 U918 ( .I0(n186), .I1(n187), .I2(n188), .S0(n559), .S1(n521), .ZN(
        n185) );
  MUX3ND0 U919 ( .I0(n195), .I1(n196), .I2(n197), .S0(n515), .S1(n511), .ZN(
        N74) );
  MUX3ND0 U920 ( .I0(n199), .I1(n200), .I2(n201), .S0(n559), .S1(n533), .ZN(
        n198) );
  MUX3ND0 U921 ( .I0(n208), .I1(n209), .I2(n210), .S0(n515), .S1(n511), .ZN(
        N73) );
  MUX3ND0 U922 ( .I0(n212), .I1(n213), .I2(n214), .S0(n560), .S1(n521), .ZN(
        n211) );
  MUX3ND0 U923 ( .I0(n221), .I1(n222), .I2(n223), .S0(n964), .S1(n511), .ZN(
        N72) );
  MUX3ND0 U924 ( .I0(n225), .I1(n226), .I2(n227), .S0(n560), .S1(n522), .ZN(
        n224) );
  MUX3ND0 U925 ( .I0(n234), .I1(n235), .I2(n236), .S0(n515), .S1(n511), .ZN(
        N71) );
  MUX3ND0 U926 ( .I0(n238), .I1(n239), .I2(n240), .S0(n560), .S1(n522), .ZN(
        n237) );
  MUX3ND0 U927 ( .I0(n247), .I1(n248), .I2(n249), .S0(N47), .S1(n511), .ZN(N70) );
  MUX3ND0 U928 ( .I0(n251), .I1(n252), .I2(n253), .S0(n561), .S1(n520), .ZN(
        n250) );
  MUX3ND0 U929 ( .I0(n260), .I1(n261), .I2(n262), .S0(n964), .S1(n965), .ZN(
        N69) );
  MUX3ND0 U930 ( .I0(n264), .I1(n265), .I2(n266), .S0(n559), .S1(n520), .ZN(
        n263) );
  MUX3ND0 U931 ( .I0(n273), .I1(n274), .I2(n275), .S0(N47), .S1(n965), .ZN(N68) );
  MUX3ND0 U932 ( .I0(n277), .I1(n278), .I2(n279), .S0(n560), .S1(n522), .ZN(
        n276) );
  MUX3ND0 U933 ( .I0(n286), .I1(n287), .I2(n288), .S0(n964), .S1(n965), .ZN(
        N67) );
  MUX3ND0 U934 ( .I0(n290), .I1(n291), .I2(n292), .S0(n560), .S1(n522), .ZN(
        n289) );
  MUX3ND0 U935 ( .I0(n299), .I1(n300), .I2(n301), .S0(n964), .S1(n965), .ZN(
        N66) );
  MUX3ND0 U936 ( .I0(n303), .I1(n304), .I2(n305), .S0(n561), .S1(n522), .ZN(
        n302) );
  MUX3ND0 U937 ( .I0(n312), .I1(n313), .I2(n314), .S0(n516), .S1(N48), .ZN(N65) );
  MUX3ND0 U938 ( .I0(n316), .I1(n317), .I2(n318), .S0(n561), .S1(n520), .ZN(
        n315) );
  MUX3ND0 U939 ( .I0(n325), .I1(n326), .I2(n327), .S0(n516), .S1(N48), .ZN(N64) );
  MUX3ND0 U940 ( .I0(n329), .I1(n330), .I2(n331), .S0(n561), .S1(n522), .ZN(
        n328) );
  MUX3ND0 U941 ( .I0(n338), .I1(n339), .I2(n340), .S0(n514), .S1(n965), .ZN(
        N63) );
  MUX3ND0 U942 ( .I0(n342), .I1(n343), .I2(n344), .S0(n561), .S1(n520), .ZN(
        n341) );
  MUX3ND0 U943 ( .I0(n351), .I1(n352), .I2(n353), .S0(n514), .S1(n965), .ZN(
        N62) );
  MUX3ND0 U944 ( .I0(n355), .I1(n356), .I2(n357), .S0(n561), .S1(n522), .ZN(
        n354) );
  MUX3ND0 U945 ( .I0(n364), .I1(n365), .I2(n366), .S0(n514), .S1(N48), .ZN(N61) );
  MUX3ND0 U946 ( .I0(n368), .I1(n369), .I2(n370), .S0(n560), .S1(n533), .ZN(
        n367) );
  MUX3ND0 U947 ( .I0(n377), .I1(n378), .I2(n379), .S0(n516), .S1(N48), .ZN(N60) );
  MUX3ND0 U948 ( .I0(n381), .I1(n382), .I2(n383), .S0(n560), .S1(n533), .ZN(
        n380) );
  MUX3ND0 U949 ( .I0(n390), .I1(n391), .I2(n392), .S0(n514), .S1(n512), .ZN(
        N59) );
  MUX3ND0 U950 ( .I0(n394), .I1(n395), .I2(n396), .S0(n559), .S1(n521), .ZN(
        n393) );
  MUX3ND0 U951 ( .I0(n403), .I1(n404), .I2(n405), .S0(n514), .S1(n512), .ZN(
        N58) );
  MUX3ND0 U952 ( .I0(n407), .I1(n408), .I2(n409), .S0(n559), .S1(n521), .ZN(
        n406) );
  MUX3ND0 U953 ( .I0(n416), .I1(n417), .I2(n418), .S0(n514), .S1(n512), .ZN(
        N57) );
  MUX3ND0 U954 ( .I0(n420), .I1(n421), .I2(n422), .S0(n558), .S1(n521), .ZN(
        n419) );
  MUX3ND0 U955 ( .I0(n429), .I1(n430), .I2(n431), .S0(n514), .S1(n512), .ZN(
        N56) );
  MUX3ND0 U956 ( .I0(n433), .I1(n434), .I2(n435), .S0(n558), .S1(n521), .ZN(
        n432) );
  MUX3ND0 U957 ( .I0(n442), .I1(n443), .I2(n444), .S0(n514), .S1(n512), .ZN(
        N55) );
  MUX3ND0 U958 ( .I0(n446), .I1(n447), .I2(n448), .S0(n560), .S1(n519), .ZN(
        n445) );
  MUX3ND0 U959 ( .I0(n455), .I1(n456), .I2(n457), .S0(n514), .S1(n512), .ZN(
        N54) );
  MUX3ND0 U960 ( .I0(n459), .I1(n460), .I2(n461), .S0(n559), .S1(n533), .ZN(
        n458) );
  MUX3ND0 U961 ( .I0(n468), .I1(n469), .I2(n470), .S0(n514), .S1(n512), .ZN(
        N53) );
  MUX3ND0 U962 ( .I0(n472), .I1(n473), .I2(n474), .S0(n561), .S1(n521), .ZN(
        n471) );
  MUX3ND0 U963 ( .I0(n481), .I1(n482), .I2(n483), .S0(n513), .S1(n512), .ZN(
        N52) );
  MUX3ND0 U964 ( .I0(n485), .I1(n486), .I2(n487), .S0(n559), .S1(n533), .ZN(
        n484) );
  MUX3ND0 U965 ( .I0(n494), .I1(n495), .I2(n496), .S0(n513), .S1(n512), .ZN(
        N51) );
  MUX3ND0 U966 ( .I0(n498), .I1(n499), .I2(n500), .S0(n560), .S1(n524), .ZN(
        n497) );
  MUX3ND0 U967 ( .I0(n507), .I1(n508), .I2(n509), .S0(n513), .S1(n512), .ZN(
        N50) );
  MUX2ND0 U968 ( .I0(\Storage[26][0] ), .I1(\Storage[27][0] ), .S(n573), .ZN(
        n41) );
  MUX2ND0 U969 ( .I0(\Storage[24][0] ), .I1(\Storage[25][0] ), .S(n573), .ZN(
        n40) );
  MUX3ND0 U970 ( .I0(n44), .I1(n43), .I2(n39), .S0(n532), .S1(n513), .ZN(n51)
         );
  MUX2ND0 U971 ( .I0(n46), .I1(n45), .S(n529), .ZN(n50) );
  MUX2ND0 U972 ( .I0(n48), .I1(n47), .S(n528), .ZN(n49) );
  MUX2ND0 U973 ( .I0(\Storage[26][1] ), .I1(\Storage[27][1] ), .S(n566), .ZN(
        n54) );
  MUX2ND0 U974 ( .I0(\Storage[24][1] ), .I1(\Storage[25][1] ), .S(n570), .ZN(
        n53) );
  MUX3ND0 U975 ( .I0(n57), .I1(n56), .I2(n52), .S0(n532), .S1(n513), .ZN(n64)
         );
  MUX2ND0 U976 ( .I0(n59), .I1(n58), .S(n527), .ZN(n63) );
  MUX2ND0 U977 ( .I0(n61), .I1(n60), .S(n529), .ZN(n62) );
  MUX2ND0 U978 ( .I0(\Storage[26][2] ), .I1(\Storage[27][2] ), .S(n566), .ZN(
        n109) );
  MUX2ND0 U979 ( .I0(\Storage[24][2] ), .I1(\Storage[25][2] ), .S(n570), .ZN(
        n108) );
  MUX3ND0 U980 ( .I0(n112), .I1(n111), .I2(n65), .S0(n532), .S1(n513), .ZN(
        n119) );
  MUX2ND0 U981 ( .I0(n114), .I1(n113), .S(n529), .ZN(n118) );
  MUX2ND0 U982 ( .I0(n116), .I1(n115), .S(n529), .ZN(n117) );
  MUX2ND0 U983 ( .I0(\Storage[26][3] ), .I1(\Storage[27][3] ), .S(n562), .ZN(
        n122) );
  MUX2ND0 U984 ( .I0(\Storage[24][3] ), .I1(\Storage[25][3] ), .S(n565), .ZN(
        n121) );
  MUX3ND0 U985 ( .I0(n125), .I1(n124), .I2(n120), .S0(n531), .S1(n516), .ZN(
        n132) );
  MUX2ND0 U986 ( .I0(n127), .I1(n126), .S(n529), .ZN(n131) );
  MUX2ND0 U987 ( .I0(n129), .I1(n128), .S(n528), .ZN(n130) );
  MUX2ND0 U988 ( .I0(\Storage[26][4] ), .I1(\Storage[27][4] ), .S(n566), .ZN(
        n135) );
  MUX2ND0 U989 ( .I0(\Storage[24][4] ), .I1(\Storage[25][4] ), .S(n562), .ZN(
        n134) );
  MUX3ND0 U990 ( .I0(n138), .I1(n137), .I2(n133), .S0(n531), .S1(n513), .ZN(
        n145) );
  MUX2ND0 U991 ( .I0(n140), .I1(n139), .S(n529), .ZN(n144) );
  MUX2ND0 U992 ( .I0(n142), .I1(n141), .S(n529), .ZN(n143) );
  MUX2ND0 U993 ( .I0(\Storage[26][5] ), .I1(\Storage[27][5] ), .S(n571), .ZN(
        n148) );
  MUX2ND0 U994 ( .I0(\Storage[24][5] ), .I1(\Storage[25][5] ), .S(n563), .ZN(
        n147) );
  MUX3ND0 U995 ( .I0(n151), .I1(n150), .I2(n146), .S0(n531), .S1(n513), .ZN(
        n158) );
  MUX2ND0 U996 ( .I0(n153), .I1(n152), .S(n528), .ZN(n157) );
  MUX2ND0 U997 ( .I0(n155), .I1(n154), .S(n528), .ZN(n156) );
  MUX2ND0 U998 ( .I0(\Storage[26][6] ), .I1(\Storage[27][6] ), .S(n574), .ZN(
        n161) );
  MUX2ND0 U999 ( .I0(\Storage[24][6] ), .I1(\Storage[25][6] ), .S(n574), .ZN(
        n160) );
  MUX3ND0 U1000 ( .I0(n164), .I1(n163), .I2(n159), .S0(n530), .S1(n513), .ZN(
        n171) );
  MUX2ND0 U1001 ( .I0(n166), .I1(n165), .S(n528), .ZN(n170) );
  MUX2ND0 U1002 ( .I0(n168), .I1(n167), .S(n528), .ZN(n169) );
  MUX2ND0 U1003 ( .I0(\Storage[26][7] ), .I1(\Storage[27][7] ), .S(n574), .ZN(
        n174) );
  MUX2ND0 U1004 ( .I0(\Storage[24][7] ), .I1(\Storage[25][7] ), .S(n569), .ZN(
        n173) );
  MUX3ND0 U1005 ( .I0(n177), .I1(n176), .I2(n172), .S0(n530), .S1(n518), .ZN(
        n184) );
  MUX2ND0 U1006 ( .I0(n179), .I1(n178), .S(n528), .ZN(n183) );
  MUX2ND0 U1007 ( .I0(n181), .I1(n180), .S(n528), .ZN(n182) );
  MUX2ND0 U1008 ( .I0(\Storage[26][8] ), .I1(\Storage[27][8] ), .S(n568), .ZN(
        n187) );
  MUX2ND0 U1009 ( .I0(\Storage[24][8] ), .I1(\Storage[25][8] ), .S(n568), .ZN(
        n186) );
  MUX3ND0 U1010 ( .I0(n190), .I1(n189), .I2(n185), .S0(n532), .S1(n518), .ZN(
        n197) );
  MUX2ND0 U1011 ( .I0(n192), .I1(n191), .S(n528), .ZN(n196) );
  MUX2ND0 U1012 ( .I0(n194), .I1(n193), .S(n528), .ZN(n195) );
  MUX2ND0 U1013 ( .I0(\Storage[26][9] ), .I1(\Storage[27][9] ), .S(n569), .ZN(
        n200) );
  MUX2ND0 U1014 ( .I0(\Storage[24][9] ), .I1(\Storage[25][9] ), .S(n569), .ZN(
        n199) );
  MUX3ND0 U1015 ( .I0(n203), .I1(n202), .I2(n198), .S0(n531), .S1(n518), .ZN(
        n210) );
  MUX2ND0 U1016 ( .I0(n205), .I1(n204), .S(n527), .ZN(n209) );
  MUX2ND0 U1017 ( .I0(n207), .I1(n206), .S(n527), .ZN(n208) );
  MUX2ND0 U1018 ( .I0(\Storage[26][10] ), .I1(\Storage[27][10] ), .S(n569), 
        .ZN(n213) );
  MUX2ND0 U1019 ( .I0(\Storage[24][10] ), .I1(\Storage[25][10] ), .S(n574), 
        .ZN(n212) );
  MUX3ND0 U1020 ( .I0(n216), .I1(n215), .I2(n211), .S0(n529), .S1(n518), .ZN(
        n223) );
  MUX2ND0 U1021 ( .I0(n218), .I1(n217), .S(n527), .ZN(n222) );
  MUX2ND0 U1022 ( .I0(n220), .I1(n219), .S(n527), .ZN(n221) );
  MUX2ND0 U1023 ( .I0(\Storage[26][11] ), .I1(\Storage[27][11] ), .S(n574), 
        .ZN(n226) );
  MUX2ND0 U1024 ( .I0(\Storage[24][11] ), .I1(\Storage[25][11] ), .S(n569), 
        .ZN(n225) );
  MUX3ND0 U1025 ( .I0(n229), .I1(n228), .I2(n224), .S0(n529), .S1(n518), .ZN(
        n236) );
  MUX2ND0 U1026 ( .I0(n231), .I1(n230), .S(n527), .ZN(n235) );
  MUX2ND0 U1027 ( .I0(n233), .I1(n232), .S(n527), .ZN(n234) );
  MUX2ND0 U1028 ( .I0(\Storage[26][12] ), .I1(\Storage[27][12] ), .S(n569), 
        .ZN(n239) );
  MUX2ND0 U1029 ( .I0(\Storage[24][12] ), .I1(\Storage[25][12] ), .S(n574), 
        .ZN(n238) );
  MUX3ND0 U1030 ( .I0(n242), .I1(n241), .I2(n237), .S0(n530), .S1(n518), .ZN(
        n249) );
  MUX2ND0 U1031 ( .I0(n244), .I1(n243), .S(n527), .ZN(n248) );
  MUX2ND0 U1032 ( .I0(n246), .I1(n245), .S(n527), .ZN(n247) );
  MUX2ND0 U1033 ( .I0(\Storage[26][13] ), .I1(\Storage[27][13] ), .S(n574), 
        .ZN(n252) );
  MUX2ND0 U1034 ( .I0(\Storage[24][13] ), .I1(\Storage[25][13] ), .S(n574), 
        .ZN(n251) );
  MUX3ND0 U1035 ( .I0(n255), .I1(n254), .I2(n250), .S0(n531), .S1(n518), .ZN(
        n262) );
  MUX2ND0 U1036 ( .I0(n257), .I1(n256), .S(n523), .ZN(n261) );
  MUX2ND0 U1037 ( .I0(n259), .I1(n258), .S(n523), .ZN(n260) );
  MUX2ND0 U1038 ( .I0(\Storage[26][14] ), .I1(\Storage[27][14] ), .S(n574), 
        .ZN(n265) );
  MUX2ND0 U1039 ( .I0(\Storage[24][14] ), .I1(\Storage[25][14] ), .S(n563), 
        .ZN(n264) );
  MUX3ND0 U1040 ( .I0(n268), .I1(n267), .I2(n263), .S0(n530), .S1(n518), .ZN(
        n275) );
  MUX2ND0 U1041 ( .I0(n270), .I1(n269), .S(n523), .ZN(n274) );
  MUX2ND0 U1042 ( .I0(n272), .I1(n271), .S(n523), .ZN(n273) );
  MUX2ND0 U1043 ( .I0(\Storage[26][15] ), .I1(\Storage[27][15] ), .S(n563), 
        .ZN(n278) );
  MUX2ND0 U1044 ( .I0(\Storage[24][15] ), .I1(\Storage[25][15] ), .S(n574), 
        .ZN(n277) );
  MUX3ND0 U1045 ( .I0(n281), .I1(n280), .I2(n276), .S0(n530), .S1(n518), .ZN(
        n288) );
  MUX2ND0 U1046 ( .I0(n283), .I1(n282), .S(n520), .ZN(n287) );
  MUX2ND0 U1047 ( .I0(n285), .I1(n284), .S(n520), .ZN(n286) );
  MUX2ND0 U1048 ( .I0(\Storage[26][16] ), .I1(\Storage[27][16] ), .S(n563), 
        .ZN(n291) );
  MUX2ND0 U1049 ( .I0(\Storage[24][16] ), .I1(\Storage[25][16] ), .S(n563), 
        .ZN(n290) );
  MUX3ND0 U1050 ( .I0(n294), .I1(n293), .I2(n289), .S0(n530), .S1(n518), .ZN(
        n301) );
  MUX2ND0 U1051 ( .I0(n296), .I1(n295), .S(n523), .ZN(n300) );
  MUX2ND0 U1052 ( .I0(n298), .I1(n297), .S(n523), .ZN(n299) );
  MUX2ND0 U1053 ( .I0(\Storage[26][17] ), .I1(\Storage[27][17] ), .S(n571), 
        .ZN(n304) );
  MUX2ND0 U1054 ( .I0(\Storage[24][17] ), .I1(\Storage[25][17] ), .S(n566), 
        .ZN(n303) );
  MUX3ND0 U1055 ( .I0(n307), .I1(n306), .I2(n302), .S0(n530), .S1(n517), .ZN(
        n314) );
  MUX2ND0 U1056 ( .I0(n309), .I1(n308), .S(n523), .ZN(n313) );
  MUX2ND0 U1057 ( .I0(n311), .I1(n310), .S(n523), .ZN(n312) );
  MUX2ND0 U1058 ( .I0(\Storage[26][18] ), .I1(\Storage[27][18] ), .S(n562), 
        .ZN(n317) );
  MUX2ND0 U1059 ( .I0(\Storage[24][18] ), .I1(\Storage[25][18] ), .S(n571), 
        .ZN(n316) );
  MUX3ND0 U1060 ( .I0(n320), .I1(n319), .I2(n315), .S0(n530), .S1(n517), .ZN(
        n327) );
  MUX2ND0 U1061 ( .I0(n322), .I1(n321), .S(n526), .ZN(n326) );
  MUX2ND0 U1062 ( .I0(n324), .I1(n323), .S(n526), .ZN(n325) );
  MUX2ND0 U1063 ( .I0(\Storage[26][19] ), .I1(\Storage[27][19] ), .S(n563), 
        .ZN(n330) );
  MUX2ND0 U1064 ( .I0(\Storage[24][19] ), .I1(\Storage[25][19] ), .S(n572), 
        .ZN(n329) );
  MUX3ND0 U1065 ( .I0(n333), .I1(n332), .I2(n328), .S0(n529), .S1(n517), .ZN(
        n340) );
  MUX2ND0 U1066 ( .I0(n335), .I1(n334), .S(n526), .ZN(n339) );
  MUX2ND0 U1067 ( .I0(n337), .I1(n336), .S(n526), .ZN(n338) );
  MUX2ND0 U1068 ( .I0(\Storage[26][20] ), .I1(\Storage[27][20] ), .S(n562), 
        .ZN(n343) );
  MUX2ND0 U1069 ( .I0(\Storage[24][20] ), .I1(\Storage[25][20] ), .S(n572), 
        .ZN(n342) );
  MUX3ND0 U1070 ( .I0(n346), .I1(n345), .I2(n341), .S0(n531), .S1(n517), .ZN(
        n353) );
  MUX2ND0 U1071 ( .I0(n348), .I1(n347), .S(n526), .ZN(n352) );
  MUX2ND0 U1072 ( .I0(n350), .I1(n349), .S(n526), .ZN(n351) );
  MUX2ND0 U1073 ( .I0(\Storage[26][21] ), .I1(\Storage[27][21] ), .S(n565), 
        .ZN(n356) );
  MUX2ND0 U1074 ( .I0(\Storage[24][21] ), .I1(\Storage[25][21] ), .S(n567), 
        .ZN(n355) );
  MUX3ND0 U1075 ( .I0(n359), .I1(n358), .I2(n354), .S0(n530), .S1(n517), .ZN(
        n366) );
  MUX2ND0 U1076 ( .I0(n361), .I1(n360), .S(n526), .ZN(n365) );
  MUX2ND0 U1077 ( .I0(n363), .I1(n362), .S(n526), .ZN(n364) );
  MUX2ND0 U1078 ( .I0(\Storage[26][22] ), .I1(\Storage[27][22] ), .S(n563), 
        .ZN(n369) );
  MUX2ND0 U1079 ( .I0(\Storage[24][22] ), .I1(\Storage[25][22] ), .S(n567), 
        .ZN(n368) );
  MUX3ND0 U1080 ( .I0(n372), .I1(n371), .I2(n367), .S0(n532), .S1(n517), .ZN(
        n379) );
  MUX2ND0 U1081 ( .I0(n374), .I1(n373), .S(n526), .ZN(n378) );
  MUX2ND0 U1082 ( .I0(n376), .I1(n375), .S(n526), .ZN(n377) );
  MUX2ND0 U1083 ( .I0(\Storage[26][23] ), .I1(\Storage[27][23] ), .S(n566), 
        .ZN(n382) );
  MUX2ND0 U1084 ( .I0(\Storage[24][23] ), .I1(\Storage[25][23] ), .S(n562), 
        .ZN(n381) );
  MUX3ND0 U1085 ( .I0(n385), .I1(n384), .I2(n380), .S0(n530), .S1(n517), .ZN(
        n392) );
  MUX2ND0 U1086 ( .I0(n387), .I1(n386), .S(n525), .ZN(n391) );
  MUX2ND0 U1087 ( .I0(n389), .I1(n388), .S(n525), .ZN(n390) );
  MUX2ND0 U1088 ( .I0(\Storage[26][24] ), .I1(\Storage[27][24] ), .S(n570), 
        .ZN(n395) );
  MUX2ND0 U1089 ( .I0(\Storage[24][24] ), .I1(\Storage[25][24] ), .S(n567), 
        .ZN(n394) );
  MUX3ND0 U1090 ( .I0(n398), .I1(n397), .I2(n393), .S0(n531), .S1(n517), .ZN(
        n405) );
  MUX2ND0 U1091 ( .I0(n400), .I1(n399), .S(n525), .ZN(n404) );
  MUX2ND0 U1092 ( .I0(n402), .I1(n401), .S(n525), .ZN(n403) );
  MUX2ND0 U1093 ( .I0(\Storage[26][25] ), .I1(\Storage[27][25] ), .S(n565), 
        .ZN(n408) );
  MUX2ND0 U1094 ( .I0(\Storage[24][25] ), .I1(\Storage[25][25] ), .S(n565), 
        .ZN(n407) );
  MUX3ND0 U1095 ( .I0(n411), .I1(n410), .I2(n406), .S0(n531), .S1(n517), .ZN(
        n418) );
  MUX2ND0 U1096 ( .I0(n413), .I1(n412), .S(n525), .ZN(n417) );
  MUX2ND0 U1097 ( .I0(n415), .I1(n414), .S(n525), .ZN(n416) );
  MUX2ND0 U1098 ( .I0(\Storage[26][26] ), .I1(\Storage[27][26] ), .S(n562), 
        .ZN(n421) );
  MUX2ND0 U1099 ( .I0(\Storage[24][26] ), .I1(\Storage[25][26] ), .S(n565), 
        .ZN(n420) );
  MUX3ND0 U1100 ( .I0(n424), .I1(n423), .I2(n419), .S0(n531), .S1(n517), .ZN(
        n431) );
  MUX2ND0 U1101 ( .I0(n426), .I1(n425), .S(n525), .ZN(n430) );
  MUX2ND0 U1102 ( .I0(n428), .I1(n427), .S(n525), .ZN(n429) );
  MUX2ND0 U1103 ( .I0(\Storage[26][27] ), .I1(\Storage[27][27] ), .S(n565), 
        .ZN(n434) );
  MUX2ND0 U1104 ( .I0(\Storage[24][27] ), .I1(\Storage[25][27] ), .S(n570), 
        .ZN(n433) );
  MUX3ND0 U1105 ( .I0(n437), .I1(n436), .I2(n432), .S0(n531), .S1(n516), .ZN(
        n444) );
  MUX2ND0 U1106 ( .I0(n439), .I1(n438), .S(n525), .ZN(n443) );
  MUX2ND0 U1107 ( .I0(n441), .I1(n440), .S(n525), .ZN(n442) );
  MUX2ND0 U1108 ( .I0(\Storage[26][28] ), .I1(\Storage[27][28] ), .S(n570), 
        .ZN(n447) );
  MUX2ND0 U1109 ( .I0(\Storage[24][28] ), .I1(\Storage[25][28] ), .S(n563), 
        .ZN(n446) );
  MUX3ND0 U1110 ( .I0(n450), .I1(n449), .I2(n445), .S0(n532), .S1(n516), .ZN(
        n457) );
  MUX2ND0 U1111 ( .I0(n452), .I1(n451), .S(n524), .ZN(n456) );
  MUX2ND0 U1112 ( .I0(n454), .I1(n453), .S(n524), .ZN(n455) );
  MUX2ND0 U1113 ( .I0(\Storage[26][29] ), .I1(\Storage[27][29] ), .S(n565), 
        .ZN(n460) );
  MUX2ND0 U1114 ( .I0(\Storage[24][29] ), .I1(\Storage[25][29] ), .S(n562), 
        .ZN(n459) );
  MUX3ND0 U1115 ( .I0(n463), .I1(n462), .I2(n458), .S0(n532), .S1(n516), .ZN(
        n470) );
  MUX2ND0 U1116 ( .I0(n465), .I1(n464), .S(n524), .ZN(n469) );
  MUX2ND0 U1117 ( .I0(n467), .I1(n466), .S(n524), .ZN(n468) );
  MUX2ND0 U1118 ( .I0(\Storage[26][30] ), .I1(\Storage[27][30] ), .S(n573), 
        .ZN(n473) );
  MUX2ND0 U1119 ( .I0(\Storage[24][30] ), .I1(\Storage[25][30] ), .S(n573), 
        .ZN(n472) );
  MUX3ND0 U1120 ( .I0(n476), .I1(n475), .I2(n471), .S0(n532), .S1(n516), .ZN(
        n483) );
  MUX2ND0 U1121 ( .I0(n478), .I1(n477), .S(n524), .ZN(n482) );
  MUX2ND0 U1122 ( .I0(n480), .I1(n479), .S(n524), .ZN(n481) );
  MUX2ND0 U1123 ( .I0(\Storage[26][31] ), .I1(\Storage[27][31] ), .S(n573), 
        .ZN(n486) );
  MUX2ND0 U1124 ( .I0(\Storage[24][31] ), .I1(\Storage[25][31] ), .S(n573), 
        .ZN(n485) );
  MUX3ND0 U1125 ( .I0(n489), .I1(n488), .I2(n484), .S0(n532), .S1(n516), .ZN(
        n496) );
  MUX2ND0 U1126 ( .I0(n491), .I1(n490), .S(n524), .ZN(n495) );
  MUX2ND0 U1127 ( .I0(n493), .I1(n492), .S(n524), .ZN(n494) );
  MUX2ND0 U1128 ( .I0(\Storage[26][32] ), .I1(\Storage[27][32] ), .S(n573), 
        .ZN(n499) );
  MUX2ND0 U1129 ( .I0(\Storage[24][32] ), .I1(\Storage[25][32] ), .S(n564), 
        .ZN(n498) );
  MUX3ND0 U1130 ( .I0(n502), .I1(n501), .I2(n497), .S0(n532), .S1(n516), .ZN(
        n509) );
  MUX2ND0 U1131 ( .I0(n504), .I1(n503), .S(n524), .ZN(n508) );
  MUX2ND0 U1132 ( .I0(n506), .I1(n505), .S(n527), .ZN(n507) );
endmodule


module PLLTop ( ClockOut, ClockIn, Reset );
  input ClockIn, Reset;
  output ClockOut;
  wire   SampleWire, CtrCarry;
  wire   [1:0] AdjFreq;

  DEL005 SampleDelay1 ( .I(ClockIn), .Z(SampleWire) );
  ClockComparator Comp1 ( .AdjustFreq(AdjFreq), .ClockIn(ClockIn), 
        .CounterClock(CtrCarry), .Reset(Reset) );
  VFO VFO1 ( .ClockOut(ClockOut), .AdjustFreq(AdjFreq), .Sample(SampleWire), 
        .Reset(Reset) );
  MultiCounter MCntr1 ( .CarryOut(CtrCarry), .Clock(ClockOut), .Reset(Reset)
         );
endmodule


module ClockComparator ( AdjustFreq, ClockIn, CounterClock, Reset );
  output [1:0] AdjustFreq;
  input ClockIn, CounterClock, Reset;
  wire   ZeroCounters, N5, N6, N7, N8, N9, N19, N20, n2, n3, n4, n5, n6, n7;
  wire   [1:0] ClockInN;
  wire   [1:0] CounterClockN;

  MOAI22D1 U5 ( .A1(N8), .A2(n4), .B1(n5), .B2(ClockInN[1]), .ZN(N20) );
  MOAI22D1 U8 ( .A1(CounterClockN[1]), .A2(n6), .B1(n5), .B2(N9), .ZN(N19) );
  DFSNQD1 ZeroCounters_reg ( .D(N9), .CP(ClockIn), .SDN(n3), .Q(ZeroCounters)
         );
  DFCND1 \ClockInN_reg[1]  ( .D(N6), .CP(ClockIn), .CDN(n2), .Q(ClockInN[1]), 
        .QN(n7) );
  DFCND1 \ClockInN_reg[0]  ( .D(N5), .CP(ClockIn), .CDN(n2), .Q(ClockInN[0]), 
        .QN(N5) );
  DFCND1 \CounterClockN_reg[0]  ( .D(N7), .CP(CounterClock), .CDN(n2), .Q(
        CounterClockN[0]), .QN(N7) );
  DFSNQD1 \AdjustFreq_reg[0]  ( .D(N19), .CP(CounterClock), .SDN(n3), .Q(
        AdjustFreq[0]) );
  DFCNQD1 \CounterClockN_reg[1]  ( .D(N8), .CP(CounterClock), .CDN(n2), .Q(
        CounterClockN[1]) );
  DFCNQD1 \AdjustFreq_reg[1]  ( .D(N20), .CP(CounterClock), .CDN(n3), .Q(
        AdjustFreq[1]) );
  INVD1 U3 ( .I(Reset), .ZN(n3) );
  INVD1 U4 ( .I(ZeroCounters), .ZN(n2) );
  AOI21D1 U6 ( .A1(ClockInN[0]), .A2(n5), .B(N9), .ZN(n4) );
  NR2D1 U7 ( .A1(N7), .A2(N6), .ZN(n6) );
  ND2D1 U9 ( .A1(CounterClockN[1]), .A2(CounterClockN[0]), .ZN(n5) );
  NR2D1 U10 ( .A1(n7), .A2(N5), .ZN(N9) );
  XOR2D1 U11 ( .A1(N5), .A2(n7), .Z(N6) );
  XNR2D1 U12 ( .A1(N7), .A2(CounterClockN[1]), .ZN(N8) );
endmodule


module VFO ( ClockOut, AdjustFreq, Sample, Reset );
  input [1:0] AdjustFreq;
  input Sample, Reset;
  output ClockOut;
  wire   FastClock, N9, N10, N11, N12, N13, N14, N16, N17, N18, N19, N20, N21,
         N27, N28, N29, N30, N31, N32, N35, N36, N37, N38, N39, N40, N49, N51,
         N54, N55, n17, n18, n19, n20, n21, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32;
  wire   [5:0] WireD;
  wire   [5:0] FastDivvy;
  wire   [5:0] DivideFactor;

  DEL005 \DelayLine[0].Delay83ps  ( .I(WireD[0]), .Z(WireD[1]) );
  DEL005 \DelayLine[1].Delay83ps  ( .I(WireD[1]), .Z(WireD[2]) );
  DEL005 \DelayLine[2].Delay83ps  ( .I(WireD[2]), .Z(WireD[3]) );
  DEL005 \DelayLine[3].Delay83ps  ( .I(WireD[3]), .Z(WireD[4]) );
  DEL005 \DelayLine[4].Delay83ps  ( .I(WireD[4]), .Z(WireD[5]) );
  VFO_DW01_dec_0 \Sampler/sub_183  ( .A(DivideFactor), .SUM({N40, N39, N38, 
        N37, N36, N35}) );
  VFO_DW01_inc_0 \Sampler/add_180  ( .A(DivideFactor), .SUM({N32, N31, N30, 
        N29, N28, N27}) );
  VFO_DW01_inc_1 \ClockOutGen/add_161  ( .A(FastDivvy), .SUM({N14, N13, N12, 
        N11, N10, N9}) );
  DFCNQD1 ClockOutReg_reg ( .D(n17), .CP(FastClock), .CDN(n2), .Q(ClockOut) );
  DFCNQD1 \FastDivvy_reg[5]  ( .D(N21), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[5]) );
  DFCNQD1 \FastDivvy_reg[2]  ( .D(N18), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[2]) );
  DFCNQD1 \FastDivvy_reg[0]  ( .D(N16), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[0]) );
  DFCNQD1 \FastDivvy_reg[1]  ( .D(N17), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[1]) );
  DFCNQD1 \FastDivvy_reg[4]  ( .D(N20), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[4]) );
  DFCNQD1 \FastDivvy_reg[3]  ( .D(N19), .CP(FastClock), .CDN(n2), .Q(
        FastDivvy[3]) );
  EDFCND1 \DivideFactor_reg[3]  ( .D(N51), .E(N54), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[3]), .QN(n22) );
  EDFCND1 \DivideFactor_reg[2]  ( .D(N49), .E(N54), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[2]) );
  EDFCND1 \DivideFactor_reg[5]  ( .D(N55), .E(N54), .CP(Sample), .CDN(n20), 
        .Q(DivideFactor[5]), .QN(n14) );
  DFSND1 \DivideFactor_reg[4]  ( .D(n19), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[4]), .QN(n13) );
  DFSND1 \DivideFactor_reg[1]  ( .D(n18), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[1]), .QN(n23) );
  DFSND1 \DivideFactor_reg[0]  ( .D(n21), .CP(Sample), .SDN(n20), .Q(
        DivideFactor[0]), .QN(n31) );
  BUFFD1 U3 ( .I(n20), .Z(n2) );
  INVD1 U4 ( .I(Reset), .ZN(n20) );
  AO222D0 U5 ( .A1(N35), .A2(n3), .B1(N27), .B2(n4), .C1(DivideFactor[0]), 
        .C2(n5), .Z(n21) );
  AO222D0 U6 ( .A1(N39), .A2(n3), .B1(N31), .B2(n4), .C1(DivideFactor[4]), 
        .C2(n5), .Z(n19) );
  AO222D0 U7 ( .A1(N36), .A2(n3), .B1(N28), .B2(n4), .C1(DivideFactor[1]), 
        .C2(n5), .Z(n18) );
  CKND0 U8 ( .CLK(N54), .CN(n5) );
  AN2D0 U9 ( .A1(n6), .A2(n7), .Z(n4) );
  AN2D0 U10 ( .A1(n8), .A2(n9), .Z(n3) );
  CKXOR2D0 U11 ( .A1(ClockOut), .A2(n10), .Z(n17) );
  AO22D0 U12 ( .A1(N40), .A2(n8), .B1(N32), .B2(n6), .Z(N55) );
  MUX2ND0 U13 ( .I0(n11), .I1(n12), .S(AdjustFreq[0]), .ZN(N54) );
  CKND2D0 U14 ( .A1(AdjustFreq[1]), .A2(n9), .ZN(n12) );
  ND3D0 U15 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n9) );
  ND3D0 U16 ( .A1(DivideFactor[2]), .A2(DivideFactor[1]), .A3(DivideFactor[3]), 
        .ZN(n15) );
  IND2D0 U17 ( .A1(AdjustFreq[1]), .B1(n7), .ZN(n11) );
  ND3D0 U18 ( .A1(DivideFactor[5]), .A2(DivideFactor[4]), .A3(n16), .ZN(n7) );
  INR3D0 U19 ( .A1(DivideFactor[2]), .B1(n22), .B2(n23), .ZN(n16) );
  AO22D0 U20 ( .A1(N38), .A2(n8), .B1(N30), .B2(n6), .Z(N51) );
  AO22D0 U21 ( .A1(N37), .A2(n8), .B1(N29), .B2(n6), .Z(N49) );
  NR2D0 U22 ( .A1(AdjustFreq[0]), .A2(AdjustFreq[1]), .ZN(n6) );
  AN2D0 U23 ( .A1(AdjustFreq[1]), .A2(AdjustFreq[0]), .Z(n8) );
  INR2D0 U24 ( .A1(N14), .B1(n10), .ZN(N21) );
  INR2D0 U25 ( .A1(N13), .B1(n10), .ZN(N20) );
  INR2D0 U26 ( .A1(N12), .B1(n10), .ZN(N19) );
  INR2D0 U27 ( .A1(N11), .B1(n10), .ZN(N18) );
  INR2D0 U28 ( .A1(N10), .B1(n10), .ZN(N17) );
  INR2D0 U29 ( .A1(N9), .B1(n10), .ZN(N16) );
  OA21D0 U30 ( .A1(FastDivvy[5]), .A2(n14), .B(n24), .Z(n10) );
  IOA22D0 U31 ( .B1(n25), .B2(n26), .A1(n14), .A2(FastDivvy[5]), .ZN(n24) );
  AOI221D0 U32 ( .A1(FastDivvy[4]), .A2(n13), .B1(FastDivvy[3]), .B2(n22), .C(
        n27), .ZN(n26) );
  AOI221D0 U33 ( .A1(DivideFactor[3]), .A2(n28), .B1(DivideFactor[2]), .B2(n29), .C(n30), .ZN(n27) );
  IAO21D0 U34 ( .A1(n29), .A2(DivideFactor[2]), .B(FastDivvy[2]), .ZN(n30) );
  OAI32D0 U35 ( .A1(n31), .A2(FastDivvy[0]), .A3(n32), .B1(FastDivvy[1]), .B2(
        n23), .ZN(n29) );
  AN2D0 U36 ( .A1(FastDivvy[1]), .A2(n23), .Z(n32) );
  CKND0 U37 ( .CLK(FastDivvy[3]), .CN(n28) );
  NR2D0 U38 ( .A1(FastDivvy[4]), .A2(n13), .ZN(n25) );
  CKND0 U39 ( .CLK(WireD[0]), .CN(FastClock) );
  CKND2D0 U40 ( .A1(WireD[5]), .A2(n20), .ZN(WireD[0]) );
endmodule


module MultiCounter ( CarryOut, Clock, Reset );
  input Clock, Reset;
  output CarryOut;
  wire   N1, N2, N3, N4, N5, n1;
  wire   [3:0] Ctr;

  MultiCounter_DW01_inc_0 add_16 ( .A({CarryOut, Ctr}), .SUM({N5, N4, N3, N2, 
        N1}) );
  DFCNQD1 \Ctr_reg[1]  ( .D(N2), .CP(Clock), .CDN(n1), .Q(Ctr[1]) );
  DFCNQD1 \Ctr_reg[2]  ( .D(N3), .CP(Clock), .CDN(n1), .Q(Ctr[2]) );
  DFCNQD1 \Ctr_reg[3]  ( .D(N4), .CP(Clock), .CDN(n1), .Q(Ctr[3]) );
  DFCNQD1 \Ctr_reg[0]  ( .D(N1), .CP(Clock), .CDN(n1), .Q(Ctr[0]) );
  DFCNQD1 \Ctr_reg[4]  ( .D(N5), .CP(Clock), .CDN(n1), .Q(CarryOut) );
  INVD1 U3 ( .I(Reset), .ZN(n1) );
endmodule


module MultiCounter_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_dec_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   n1, n2, n3, n4, n5;

  CKXOR2D0 U1 ( .A1(A[5]), .A2(n1), .Z(SUM[5]) );
  NR2D0 U2 ( .A1(A[4]), .A2(n2), .ZN(n1) );
  XNR2D0 U3 ( .A1(n2), .A2(A[4]), .ZN(SUM[4]) );
  OAI21D0 U4 ( .A1(n3), .A2(n4), .B(n2), .ZN(SUM[3]) );
  CKND2D0 U5 ( .A1(n3), .A2(n4), .ZN(n2) );
  CKND0 U6 ( .CLK(A[3]), .CN(n4) );
  AO21D0 U7 ( .A1(n5), .A2(A[2]), .B(n3), .Z(SUM[2]) );
  NR2D0 U8 ( .A1(n5), .A2(A[2]), .ZN(n3) );
  IOA21D0 U9 ( .A1(A[0]), .A2(A[1]), .B(n5), .ZN(SUM[1]) );
  IND2D0 U10 ( .A1(A[1]), .B1(SUM[0]), .ZN(n5) );
  CKND0 U11 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module VFO_DW01_inc_1 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  CKXOR2D0 U1 ( .A1(\carry[5] ), .A2(A[5]), .Z(SUM[5]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module DesDecoder_DWid32_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  CKXOR2D0 U1 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
  CKND0 U2 ( .CLK(A[0]), .CN(SUM[0]) );
endmodule


module FIFOStateM_AWid5_DW01_inc_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   \carry[4] , \carry[3] , \carry[2] ;

  HA1D0 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA1D0 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  HA1D0 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  INVD1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  CKXOR2D0 U2 ( .A1(\carry[4] ), .A2(A[4]), .Z(SUM[4]) );
endmodule

