library verilog;
use verilog.vl_types.all;
entity ir_decode_tb is
end ir_decode_tb;
