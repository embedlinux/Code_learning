library verilog;
use verilog.vl_types.all;
entity key_led_top_tb is
end key_led_top_tb;
